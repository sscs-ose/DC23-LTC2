** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/resistor/resistor-test.sch

.include /home/designer/.volare/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_statistical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical

**.subckt resistor-test out vin vin
*.opin out
*.iopin vin
*.iopin vin
vin vin GND 4
x1 vin GND out GND resistor
**** begin user architecture code

.control
dc vin 0 3.3 0.01
plot V(vin) V(out)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  resistor.sym # of pins=4
** sym_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/resistor/resistor.sym
** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/resistor/resistor.sch
.subckt resistor VDD BULK OUT VSS
*.iopin OUT1
*.iopin VSS
*.iopin VDD
*.iopin B
*.iopin OUT2
XR1 OUT1 VDD B ppolyf_u r_width=1e-6 r_length=200e-6 m=1
XR2 VSS OUT2 B ppolyf_u r_width=1e-6 r_length=120e-6 m=1
XR3 B B B ppolyf_u r_width=1e-6 r_length=20e-6 m=1
XR4 B B B ppolyf_u r_width=1e-6 r_length=20e-6 m=1
.ends

.GLOBAL GND
.end

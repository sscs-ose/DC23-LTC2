* Extracted by KLayout with GF180MCU LVS runset on : 03/02/2024 16:18

.SUBCKT waffle_1984 S G D
M$1 S G D S pfet_03v3 L=0.5U W=8689.92U AS=5051.0418P AD=5049.1178P
+ PS=17554.32U PD=17507.92U
.ENDS waffle_1984

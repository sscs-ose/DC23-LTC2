* NGSPICE file created from inv_sample.ext - technology: gf180mcuD

.subckt pfet a_n92_0# a_94_0# a_28_312# w_n230_n138#
X0 a_94_0# a_28_312# a_n92_0# w_n230_n138# pfet_03v3 ad=0.819p pd=3.82u as=0.819p ps=3.82u w=1.26u l=0.28u
.ends

.subckt nfet$1 a_n84_n2# a_216_n2# a_30_n132# a_94_0#
X0 a_94_0# a_30_n132# a_n84_n2# a_216_n2# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
.ends

.subckt inv_sample vdd vss out in
Xpfet_0 out vdd in vdd pfet
Xnfet$1_0 out vss in vss nfet$1
.ends


* NGSPICE file created from sar.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VNW VPW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 VDD Q CLK VSS D VNW VPW VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X1 Q a_2304_115# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 a_2304_115# a_2011_527# VSS VSUBS nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X3 a_1004_159# D a_836_159# VSUBS nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.187p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X5 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.166p pd=1.28u as=0.179p ps=1.36u w=0.36u l=0.5u
X6 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.4f pd=0.64u as=0.166p ps=1.28u w=0.36u l=0.5u
X7 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.179p pd=1.36u as=0.104p ps=0.94u w=0.36u l=0.5u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
X9 VSS a_1376_115# a_1328_159# VSUBS nfet_06v0 ad=0.264p pd=1.82u as=43.2f ps=0.6u w=0.36u l=0.6u
X10 a_2011_527# a_448_472# a_1376_115# VSUBS nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X11 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
X12 Q a_2304_115# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=0.5u
X13 a_1376_115# a_1004_159# VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.264p ps=1.82u w=0.36u l=0.6u
X14 VSS a_2304_115# a_2256_159# VSUBS nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X15 a_836_159# a_36_151# VSS VSUBS nfet_06v0 ad=43.2f pd=0.6u as=0.158p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X17 a_2256_159# a_36_151# a_2011_527# VSUBS nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X18 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=54f pd=0.66u as=0.455p ps=3.25u w=0.36u l=0.5u
X19 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.2f pd=0.6u as=0.187p ps=1.4u w=0.36u l=0.5u
X20 a_1328_159# a_448_472# a_1004_159# VSUBS nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X21 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.104p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X22 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X23 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VNW VPW VSUBS
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.146p pd=1.46u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VSUBS nfet_06v0 ad=98.4f pd=1.06u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=98.4f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.439p pd=1.94u as=0.348p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.146p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.476p pd=2u as=0.439p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.348p pd=1.79u as=0.537p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.197p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VSUBS nfet_06v0 ad=0.197p pd=1.3u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.476p ps=2u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 ZN A2 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.497p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.497p pd=3.14u as=0.294p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 Z VSS VDD I VNW VPW VSUBS
X0 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u
X1 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.361p ps=2.52u w=0.82u l=0.5u
X3 a_224_552# I VSS VSUBS nfet_06v0 ad=0.266p pd=2.09u as=0.266p ps=2.09u w=0.605u l=0.6u
X4 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X6 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.2p pd=1.79u as=0.118p ps=0.975u w=0.455u l=0.6u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X8 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.118p pd=0.975u as=0.2p ps=1.79u w=0.455u l=0.6u
X9 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.254p ps=1.44u w=0.82u l=0.5u
X10 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 VSS Z I VDD VNW VPW VSUBS
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.494p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VSUBS nfet_06v0 ad=0.291p pd=1.53u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_68# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X4 Z a_36_68# VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.291p ps=1.53u w=0.82u l=0.6u
X5 VDD I a_36_68# VNW pfet_06v0 ad=0.494p pd=2.03u as=0.537p ps=3.32u w=1.22u l=0.5u
X6 VSS a_36_68# Z VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 VDD a_36_68# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A3 A4 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 ZN A2 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.406p pd=1.81u as=0.22p ps=1.37u w=0.845u l=0.5u
X2 ZN A3 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.372p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A3 a_36_68# VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 VSS A4 a_244_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X5 a_1468_68# A4 VSS VSUBS nfet_06v0 ad=0.152p pd=1.19u as=0.213p ps=1.34u w=0.82u l=0.6u
X6 VDD A4 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X7 a_1866_68# A2 a_1662_68# VSUBS nfet_06v0 ad=0.152p pd=1.19u as=0.172p ps=1.24u w=0.82u l=0.6u
X8 ZN A4 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X9 ZN A1 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.406p ps=1.81u w=0.845u l=0.5u
X10 a_3276_68# A1 ZN VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.416p ps=1.9u w=0.82u l=0.6u
X11 a_652_68# A4 VSS VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 a_36_68# A3 a_652_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X13 VDD A2 ZN VNW pfet_06v0 ad=0.372p pd=2.57u as=0.22p ps=1.37u w=0.845u l=0.5u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X15 VSS A4 a_1060_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X16 ZN A3 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X17 a_2372_68# A1 ZN VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.416p ps=1.9u w=0.82u l=0.6u
X18 a_36_68# A2 a_2372_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X19 ZN A1 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.406p ps=1.81u w=0.845u l=0.5u
X20 a_1060_68# A3 a_36_68# VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X21 VDD A2 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X22 VDD A4 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X23 ZN A2 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X24 ZN A1 a_2780_68# VSUBS nfet_06v0 ad=0.416p pd=1.9u as=0.131p ps=1.14u w=0.82u l=0.6u
X25 a_2780_68# A2 a_36_68# VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X26 ZN A4 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X27 VDD A1 ZN VNW pfet_06v0 ad=0.406p pd=1.81u as=0.22p ps=1.37u w=0.845u l=0.5u
X28 a_36_68# A2 a_3276_68# VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X29 VDD A3 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X30 a_1662_68# A3 a_1468_68# VSUBS nfet_06v0 ad=0.172p pd=1.24u as=0.152p ps=1.19u w=0.82u l=0.6u
X31 ZN A1 a_1866_68# VSUBS nfet_06v0 ad=0.416p pd=1.9u as=0.152p ps=1.19u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VNW VPW VSUBS
X0 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VNW VPW VSUBS
X0 VSS B a_36_68# VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.497p pd=3.14u as=0.425p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.598p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.425p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.409p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VSUBS nfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.409p pd=1.89u as=0.537p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VSUBS nfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.348p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VSUBS nfet_06v0 ad=0.205p pd=1.81u as=0.121p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VSUBS nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VSUBS nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.348p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VSUBS nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VSUBS nfet_06v0 ad=0.121p pd=0.985u as=0.205p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VNW VPW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 B C VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 a_692_68# B a_36_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# A2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.598p ps=3.42u w=1.22u l=0.5u
X3 VDD B ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.402p ps=1.94u w=0.985u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.402p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.443p pd=2.87u as=0.256p ps=1.5u w=0.985u l=0.5u
X6 VSS C a_692_68# VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 a_36_68# A1 ZN VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.409p pd=1.89u as=0.348p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VSUBS nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VSUBS nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.409p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VSUBS nfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.6u
X7 ZN A2 VSS VSUBS nfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 VDD VSS Z I VNW VPW VSUBS
X0 VSS I a_224_552# VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X1 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X3 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X4 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.361p ps=2.52u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X10 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X11 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X12 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X13 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X14 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X15 VSS I a_224_552# VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X16 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X17 a_224_552# I VSS VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X18 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X19 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X20 VDD I a_224_552# VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X21 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X22 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X23 VSS I a_224_552# VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X24 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X25 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X26 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X27 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X28 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.254p ps=1.44u w=0.82u l=0.5u
X29 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X30 a_224_552# I VSS VSUBS nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X31 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X32 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X33 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X34 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.213p pd=1.85u as=0.126p ps=1u w=0.485u l=0.6u
X35 VDD I a_224_552# VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X36 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X37 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X38 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X39 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X40 a_224_552# I VSS VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X41 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.213p ps=1.85u w=0.485u l=0.6u
X42 VDD I a_224_552# VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X43 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X44 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X45 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A3 A4 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X1 a_1213_472# A2 a_943_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.518p ps=2.07u w=1.22u l=0.5u
X2 VSS A2 ZN VSUBS nfet_06v0 ad=0.158p pd=1.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X3 a_943_472# A3 a_683_472# VNW pfet_06v0 ad=0.518p pd=2.07u as=0.488p ps=2.02u w=1.22u l=0.5u
X4 VSS A1 ZN VSUBS nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X5 a_1661_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.409p ps=1.89u w=1.22u l=0.5u
X6 VSS A4 ZN VSUBS nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X7 a_57_472# A2 a_1661_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X9 VDD A4 a_245_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.348p ps=1.79u w=1.22u l=0.5u
X10 ZN A2 VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
X12 a_245_472# A3 a_57_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.537p ps=3.32u w=1.22u l=0.5u
X13 ZN A3 VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
X14 ZN A1 a_1213_472# VNW pfet_06v0 ad=0.409p pd=1.89u as=0.348p ps=1.79u w=1.22u l=0.5u
X15 a_683_472# A4 VDD VNW pfet_06v0 ad=0.488p pd=2.02u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VNW VPW VSUBS
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.449p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VSUBS nfet_06v0 ad=0.151p pd=1.18u as=0.158p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VSUBS nfet_06v0 ad=0.213p pd=1.85u as=0.126p ps=1u w=0.485u l=0.6u
X5 Z a_36_160# VSS VSUBS nfet_06v0 ad=0.126p pd=1u as=0.151p ps=1.18u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 a_244_68# A2 VSS VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VSUBS nfet_06v0 ad=0.257p pd=1.56u as=0.131p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.535p pd=3.31u as=0.45p ps=1.96u w=1.22u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.45p pd=1.96u as=0.316p ps=1.74u w=1.22u l=0.5u
X5 VSS B ZN VSUBS nfet_06v0 ad=0.224p pd=1.9u as=0.257p ps=1.56u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 Z VSS VDD I VNW VPW VSUBS
X0 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.112p pd=0.95u as=0.189p ps=1.74u w=0.43u l=0.6u
X1 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X2 VDD a_224_552# Z VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X3 a_224_552# I VDD VNW pfet_06v0 ad=0.295p pd=1.54u as=0.361p ps=2.52u w=0.82u l=0.5u
X4 VDD I a_224_552# VNW pfet_06v0 ad=0.213p pd=1.34u as=0.295p ps=1.54u w=0.82u l=0.5u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X7 VSS I a_224_552# VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.295p pd=1.54u as=0.213p ps=1.34u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X10 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.189p pd=1.74u as=0.112p ps=0.95u w=0.43u l=0.6u
X11 Z a_224_552# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X12 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X13 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X14 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X15 Z a_224_552# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X16 VDD I a_224_552# VNW pfet_06v0 ad=0.367p pd=1.92u as=0.295p ps=1.54u w=0.82u l=0.5u
X17 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.439p ps=1.94u w=1.22u l=0.5u
X18 a_224_552# I VSS VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X19 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X20 Z a_224_552# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X21 a_224_552# I VSS VSUBS nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X22 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VNW VPW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.211p pd=1.84u as=0.211p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VNW VPW VSUBS
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.361p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VSUBS nfet_06v0 ad=0.2p pd=1.79u as=0.118p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.118p pd=0.975u as=0.234p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.254p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VSUBS nfet_06v0 ad=0.514p pd=2.91u as=0.266p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VSUBS nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 Z I VDD VSS VNW VPW VSUBS
X0 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 VDD a_224_472# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 a_224_472# I VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 VDD I a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X7 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 VSS a_224_472# Z VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X9 a_224_472# I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X10 VSS I a_224_472# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X11 Z a_224_472# VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 VDD ZN I VSS VNW VPW VSUBS
X0 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.125p pd=1u as=0.211p ps=1.84u w=0.48u l=0.6u
X2 VDD I ZN VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 ZN I VSS VSUBS nfet_06v0 ad=0.211p pd=1.84u as=0.125p ps=1u w=0.48u l=0.6u
X4 ZN I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X5 VSS I ZN VSUBS nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW VSUBS
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.401p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.401p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VSUBS nfet_06v0 ad=0.218p pd=1.87u as=0.153p ps=1.19u w=0.495u l=0.6u
X3 VSS I a_36_113# VSUBS nfet_06v0 ad=0.153p pd=1.19u as=0.158p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VNW VPW VSUBS
X0 ZN I VSS VSUBS nfet_06v0 ad=0.125p pd=1u as=0.211p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VSUBS nfet_06v0 ad=0.211p pd=1.84u as=0.125p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A3 VDD VSS Z A1 A2 VNW VPW VSUBS
X0 a_224_604# A1 a_36_88# VNW pfet_06v0 ad=0.174p pd=1.18u as=0.246p ps=2u w=0.56u l=0.5u
X1 a_36_88# A2 VSS VSUBS nfet_06v0 ad=0.14p pd=1.1u as=0.104p ps=0.92u w=0.4u l=0.6u
X2 Z a_36_88# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.389p ps=2.02u w=1.22u l=0.5u
X3 VSS A1 a_36_88# VSUBS nfet_06v0 ad=0.104p pd=0.92u as=0.176p ps=1.68u w=0.4u l=0.6u
X4 a_448_604# A2 a_224_604# VNW pfet_06v0 ad=0.224p pd=1.36u as=0.174p ps=1.18u w=0.56u l=0.5u
X5 VSS A3 a_36_88# VSUBS nfet_06v0 ad=0.224p pd=1.52u as=0.14p ps=1.1u w=0.4u l=0.6u
X6 VDD A3 a_448_604# VNW pfet_06v0 ad=0.389p pd=2.02u as=0.224p ps=1.36u w=0.56u l=0.5u
X7 Z a_36_88# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.224p ps=1.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 VSS ZN I VDD VNW VPW VSUBS
X0 ZN I VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 ZN I VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 VDD I ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.439p ps=1.94u w=1.22u l=0.5u
X4 VSS I ZN VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 ZN I VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.537p ps=3.32u w=1.22u l=0.5u
X6 VSS I ZN VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 VDD I ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X1 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.456p pd=1.96u as=0.486p ps=2.02u w=1.22u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.486p ps=2.02u w=1.22u l=0.5u
X6 VSS A3 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.535p pd=3.31u as=0.456p ps=1.96u w=1.22u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X10 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.346p ps=1.78u w=1.22u l=0.5u
X12 VSS A4 ZN VSUBS nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.02u as=0.377p ps=1.83u w=1.22u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X16 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346p pd=1.78u as=0.535p ps=3.31u w=1.22u l=0.5u
X18 VSS A4 ZN VSUBS nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X20 VSS A2 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.377p ps=1.83u w=1.22u l=0.5u
X26 VSS A1 ZN VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.02u as=0.377p ps=1.83u w=1.22u l=0.5u
X28 ZN A2 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VSUBS nfet_06v0 ad=0.158p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X31 ZN A1 VSS VSUBS nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 ZN A1 a_455_68# VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.172p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.433p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VSUBS nfet_06v0 ad=0.172p pd=1.24u as=0.131p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 VDD VSS Z A1 A2 VNW VPW VSUBS
X0 a_728_472# a_56_604# VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.4p ps=2.12u w=1.22u l=0.5u
X1 Z A1 a_728_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X2 VSS A1 a_56_604# VSUBS nfet_06v0 ad=0.218p pd=1.52u as=93.6f ps=0.88u w=0.36u l=0.6u
X3 a_728_472# A2 Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X4 Z a_56_604# VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X5 VSS A2 a_952_68# VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X6 a_244_604# A2 a_56_604# VNW pfet_06v0 ad=0.146p pd=1.08u as=0.246p ps=2u w=0.56u l=0.5u
X7 a_56_604# A2 VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
X8 a_952_68# A1 Z VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X9 VDD A1 a_244_604# VNW pfet_06v0 ad=0.4p pd=2.12u as=0.146p ps=1.08u w=0.56u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D VDD VSS CLK Q VNW VPW VSUBS
X0 VSS a_2304_115# Q VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X2 Q a_2304_115# VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 a_2304_115# a_2011_527# VSS VSUBS nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X4 a_1004_159# D a_836_159# VSUBS nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.187p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.166p pd=1.28u as=0.179p ps=1.36u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.4f pd=0.64u as=0.166p ps=1.28u w=0.36u l=0.5u
X8 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.179p pd=1.36u as=0.104p ps=0.94u w=0.36u l=0.5u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
X10 VDD a_2304_115# Q VNW pfet_06v0 ad=0.854p pd=3.84u as=0.317p ps=1.74u w=1.22u l=0.5u
X11 VSS a_1376_115# a_1328_159# VSUBS nfet_06v0 ad=0.264p pd=1.82u as=43.2f ps=0.6u w=0.36u l=0.6u
X12 a_2011_527# a_448_472# a_1376_115# VSUBS nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
X14 Q a_2304_115# VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X15 a_1376_115# a_1004_159# VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.264p ps=1.82u w=0.36u l=0.6u
X16 VSS a_2304_115# a_2256_159# VSUBS nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X17 a_836_159# a_36_151# VSS VSUBS nfet_06v0 ad=43.2f pd=0.6u as=0.158p ps=1.6u w=0.36u l=0.6u
X18 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X19 a_2256_159# a_36_151# a_2011_527# VSUBS nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X20 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=54f pd=0.66u as=0.455p ps=3.25u w=0.36u l=0.5u
X21 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.2f pd=0.6u as=0.187p ps=1.4u w=0.36u l=0.5u
X22 a_1328_159# a_448_472# a_1004_159# VSUBS nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X23 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.104p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X24 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X25 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D Q VDD VSS CLK VNW VPW VSUBS
X0 VSS CLK a_36_151# VSUBS nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X1 VDD a_2011_527# a_2304_115# VNW pfet_06v0 ad=0.386p pd=1.92u as=0.246p ps=1.46u w=0.945u l=0.5u
X2 a_1004_159# D a_836_159# VSUBS nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X3 VSS a_2304_115# Q VSUBS nfet_06v0 ad=0.359p pd=2.51u as=0.212p ps=1.34u w=0.815u l=0.6u
X4 a_2304_115# a_2011_527# VSS VSUBS nfet_06v0 ad=0.212p pd=1.34u as=0.233p ps=1.55u w=0.815u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.187p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.166p pd=1.28u as=0.179p ps=1.36u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.4f pd=0.64u as=0.166p ps=1.28u w=0.36u l=0.5u
X8 Q a_2304_115# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.386p ps=1.92u w=1.22u l=0.5u
X9 VSS a_2304_115# Q VSUBS nfet_06v0 ad=0.212p pd=1.34u as=0.212p ps=1.34u w=0.815u l=0.6u
X10 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.179p pd=1.36u as=0.104p ps=0.94u w=0.36u l=0.5u
X11 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
X12 VDD a_2304_115# Q VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X13 VSS a_1376_115# a_1328_159# VSUBS nfet_06v0 ad=0.264p pd=1.82u as=43.2f ps=0.6u w=0.36u l=0.6u
X14 a_2011_527# a_448_472# a_1376_115# VSUBS nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X15 Q a_2304_115# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X16 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
X17 Q a_2304_115# VSS VSUBS nfet_06v0 ad=0.212p pd=1.34u as=0.212p ps=1.34u w=0.815u l=0.6u
X18 a_1376_115# a_1004_159# VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.264p ps=1.82u w=0.36u l=0.6u
X19 VSS a_2304_115# a_2256_159# VSUBS nfet_06v0 ad=0.233p pd=1.55u as=43.2f ps=0.6u w=0.36u l=0.6u
X20 Q a_2304_115# VSS VSUBS nfet_06v0 ad=0.212p pd=1.34u as=0.261p ps=1.45u w=0.815u l=0.6u
X21 a_836_159# a_36_151# VSS VSUBS nfet_06v0 ad=43.2f pd=0.6u as=0.158p ps=1.6u w=0.36u l=0.6u
X22 a_448_472# a_36_151# VSS VSUBS nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X23 a_2256_159# a_36_151# a_2011_527# VSUBS nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X24 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=54f pd=0.66u as=0.455p ps=3.25u w=0.36u l=0.5u
X25 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.2f pd=0.6u as=0.187p ps=1.4u w=0.36u l=0.5u
X26 VDD a_2304_115# Q VNW pfet_06v0 ad=0.537p pd=3.32u as=0.439p ps=1.94u w=1.22u l=0.5u
X27 a_1328_159# a_448_472# a_1004_159# VSUBS nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X28 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.104p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X29 VSS a_2011_527# a_2304_115# VSUBS nfet_06v0 ad=0.261p pd=1.45u as=0.212p ps=1.34u w=0.815u l=0.6u
X30 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.262p pd=1.68u as=50.4f ps=0.64u w=0.36u l=0.5u
X31 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.246p pd=1.46u as=0.262p ps=1.68u w=0.945u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 VSS ZN I VDD VNW VPW VSUBS
X0 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 ZN I VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 ZN I VSS VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.537p ps=3.32u w=1.22u l=0.5u
X4 VSS I ZN VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VDD I ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VNW VPW VSUBS
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.229p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.387p pd=2.08u as=0.147p ps=1.09u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VSUBS nfet_06v0 ad=0.229p pd=1.58u as=93.6f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.387p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VSUBS nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VNW VPW VSUBS
X0 ZN A1 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VSUBS nfet_06v0 ad=0.172p pd=1.24u as=0.131p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.172p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VSUBS nfet_06v0 ad=0.115p pd=1.1u as=0.361p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.433p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VSUBS nfet_06v0 ad=0.131p pd=1.14u as=0.115p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VSUBS nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VNW VPW VSUBS
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VSUBS nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
.ends

.subckt sar_logic EOC VDD VSS clk comp dbot[0] dbot[10] dbot[11] dbot[1] dbot[2] dbot[3]
+ dbot[4] dbot[5] dbot[6] dbot[7] dbot[8] dbot[9] dtop[0] dtop[10] dtop[11] dtop[1]
+ dtop[2] dtop[3] dtop[4] dtop[5] dtop[6] dtop[7] dtop[8] dtop[9] rst
XFILLER_0_18_18 VDD VSS VDD FILLER_0_18_18/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_200_ VDD net27 clknet_2_3__leaf_clk VSS _025_ VDD _200_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_131_ _032_ VDD VSS _033_ net34 net11 VDD _131_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_114_ VDD VSS _004_ net28 _078_ VDD _114_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput7 dbot[1] VSS VDD net7 VDD output7/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput20 VSS dtop[2] net20 VDD VDD output20/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_130_ _059_ net32 VDD VSS _032_ net33 _058_ VDD _130_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_19_62 VDD VSS VDD FILLER_0_19_62/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_113_ VDD _077_ _071_ _078_ net4 VSS VDD _113_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput10 VSS dbot[4] net10 VDD VDD output10/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput21 VSS dtop[3] net21 VDD VDD output21/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput8 VSS dbot[2] net8 VDD VDD output8/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_19_138 VDD VSS VDD FILLER_0_19_138/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_189_ VDD net5 clknet_2_3__leaf_clk VSS _014_ VDD _189_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_112_ VDD VSS _077_ _062_ _071_ VDD _112_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput22 VSS dtop[4] net22 VDD VDD output22/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput11 VSS dbot[5] net11 VDD VDD output11/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput9 dbot[3] VSS VDD net9 VDD output9/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_188_ VDD net15 clknet_2_3__leaf_clk VSS _013_ VDD _188_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_111_ VDD VSS _076_ net32 net34 VDD _111_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput23 VSS dtop[5] net23 VDD VDD output23/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput12 VSS dbot[6] net12 VDD VDD output12/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_187_ VDD net14 clknet_2_2__leaf_clk VSS _012_ VDD _187_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_110_ net31 VDD VSS _075_ net33 current_bit\[1\] VDD _110_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_18_2 VDD VSS VDD FILLER_0_18_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput24 VSS dtop[6] net24 VDD VDD output24/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput13 VSS dbot[7] net13 VDD VDD output13/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_2 VDD VSS VDD FILLER_0_7_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_186_ VDD net13 clknet_2_0__leaf_clk VSS _011_ VDD _186_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_169_ _054_ net30 VDD VSS _025_ _059_ _080_ VDD _169_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput14 dbot[8] VSS VDD net14 VDD output14/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput25 dtop[7] VSS VDD net25 VDD output25/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_1_136 VDD VSS VDD FILLER_0_1_136/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_185_ VDD net12 clknet_2_0__leaf_clk VSS _010_ VDD _185_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_168_ VDD VSS _054_ net27 _040_ VDD _168_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_099_ VDD VSS _067_ net33 current_bit\[1\] VDD _099_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput15 VSS dbot[9] net15 VDD VDD output15/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput26 dtop[8] VSS VDD net26 VDD output26/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_184_ VDD net11 clknet_2_0__leaf_clk VSS _009_ VDD _184_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_138 VDD VSS VDD FILLER_0_12_138/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_167_ _053_ net30 VDD VSS _024_ net1 _074_ VDD _167_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_098_ VDD VSS _066_ _057_ _058_ VDD _098_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xoutput16 VSS dtop[0] net16 VDD VDD output16/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_16_2 VDD VSS VDD FILLER_0_16_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput27 dtop[9] VSS VDD net27 VDD output27/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xclkbuf_0_clk VDD VSS clknet_0_clk clk VDD clkbuf_0_clk/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_2 VDD VSS VDD FILLER_0_5_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_183_ VDD net10 clknet_2_3__leaf_clk VSS _008_ VDD _183_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_166_ VDD VSS _053_ net26 _074_ VDD _166_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_097_ VDD VSS _065_ _057_ _058_ VDD _097_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_149_ _062_ _067_ VDD VSS _045_ _059_ net32 VDD _149_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xoutput17 VSS dtop[10] net17 VDD VDD output17/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xfanout30 net30 VSS VDD current_state VDD fanout30/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_2_0__f_clk VDD VSS clknet_2_0__leaf_clk clknet_0_clk VDD clkbuf_2_0__f_clk/VPW
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_182_ VDD net9 clknet_2_1__leaf_clk VSS _007_ VDD _182_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_096_ VDD VSS _000_ net33 net28 VDD _096_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_148_ _064_ VDD VSS _044_ _066_ _073_ VDD _148_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_165_ _052_ net28 VDD VSS _023_ net34 _036_ VDD _165_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput18 VSS dtop[11] net18 VDD VDD output18/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xfanout31 net31 VSS VDD current_bit\[3\] VDD fanout31/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_181_ VDD net8 clknet_2_1__leaf_clk VSS _006_ VDD _181_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_095_ VDD VSS net6 _064_ VDD _095_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_164_ VDD VSS _052_ net25 _036_ VDD _164_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput19 dtop[1] VSS VDD net19 VDD output19/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_147_ _043_ net29 VDD VSS _014_ _062_ _042_ VDD _147_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_4_138 VDD VSS VDD FILLER_0_4_138/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_180_ VDD net7 clknet_2_3__leaf_clk VSS _005_ VDD _180_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout32 net32 current_bit\[2\] VDD VSS VDD fanout32/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_3_2 VDD VSS VDD FILLER_0_3_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_18 VDD VSS VDD FILLER_0_16_18/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_094_ VDD VSS net21 _063_ VDD _094_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_163_ _051_ net28 VDD VSS _022_ net34 _034_ VDD _163_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_129_ _030_ net29 VDD VSS _008_ _062_ _029_ VDD _129_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_146_ VDD VSS _043_ net5 _042_ VDD _146_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_18 VDD VSS VDD FILLER_0_19_18/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout33 net33 current_bit\[0\] VDD VSS VDD fanout33/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_162_ VDD VSS _051_ net24 _034_ VDD _162_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_093_ VDD _062_ net34 VSS VDD _093_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
Xinput1 VSS net1 comp VDD VDD input1/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_145_ net31 _060_ VDD VSS _042_ _057_ current_bit\[1\] VDD _145_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_1_18 VDD VSS VDD FILLER_0_1_18/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_128_ VDD VSS _031_ _062_ _029_ VDD _128_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout34 net34 VSS VDD net1 VDD fanout34/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_092_ VDD VSS net16 _061_ VDD _092_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput2 VSS net2 rst VDD VDD input2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_161_ _050_ net28 VDD VSS _021_ net34 _032_ VDD _161_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_144_ _041_ net29 VDD VSS _013_ _062_ _040_ VDD _144_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_127_ VDD VSS _030_ net10 _029_ VDD _127_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_143_ VDD VSS _041_ net15 _040_ VDD _143_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_091_ VDD VSS net32 _060_ VDD _091_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_160_ VDD VSS _050_ net23 _032_ VDD _160_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_2 VDD VSS VDD FILLER_0_1_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_126_ VDD VSS _029_ current_bit\[2\] _075_ VDD _126_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_109_ _072_ VDD VSS _003_ net3 _071_ VDD _109_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
Xclkbuf_2_1__f_clk VDD VSS clknet_2_1__leaf_clk clknet_0_clk VDD clkbuf_2_1__f_clk/VPW
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_090_ VSS _059_ net31 VDD VDD _090_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_142_ net31 _060_ VDD VSS _040_ current_bit\[0\] _058_ VDD _142_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_2_31 VDD VSS VDD FILLER_0_2_31/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_125_ VDD net29 _086_ _007_ _085_ VSS VDD _125_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_108_ VDD VSS _074_ net31 _068_ VDD _108_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_141_ VDD net28 _039_ _012_ _038_ VSS VDD _141_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_124_ net34 _067_ VDD VSS _086_ net31 net32 VDD _124_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_2_54 VDD VSS VDD FILLER_0_2_54/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_107_ VDD VSS _073_ _059_ net32 VDD _107_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_2 VDD VSS VDD FILLER_0_10_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_10 VDD VSS VDD FILLER_0_5_10/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_140_ net14 VDD VSS _039_ net31 _068_ VDD _140_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_106_ VDD VSS _072_ _059_ _068_ VDD _106_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_123_ net9 VDD VSS _085_ _066_ _070_ VDD _123_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout28 net28 VSS VDD net30 VDD fanout28/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_199_ VDD net26 clknet_2_2__leaf_clk VSS _024_ VDD _199_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_122_ _084_ net29 VDD VSS _006_ _062_ _082_ VDD _122_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_105_ net31 current_bit\[2\] VDD VSS _071_ net33 current_bit\[1\] VDD _105_/VPW VSS
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_0_138 VDD VSS VDD FILLER_0_0_138/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout29 net29 VSS VDD net30 VDD fanout29/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_198_ VDD net25 clknet_2_0__leaf_clk VSS _023_ VDD _198_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_121_ VDD VSS _084_ net8 _082_ VDD _121_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_104_ VDD VSS _070_ net31 net32 VDD _104_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_11_16 VDD VSS VDD FILLER_0_11_16/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_120_ _076_ VDD VSS _083_ _057_ current_bit\[1\] VDD _120_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_197_ VDD net24 clknet_2_0__leaf_clk VSS _022_ VDD _197_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_2 VDD VSS VDD FILLER_0_19_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_103_ VDD VSS _002_ net28 _069_ VDD _103_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_2 VDD VSS VDD FILLER_0_8_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_196_ VDD net23 clknet_2_0__leaf_clk VSS _021_ VDD _196_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_179_ VDD net4 clknet_2_2__leaf_clk VSS _004_ VDD _179_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_2_2__f_clk VDD VSS clknet_2_2__leaf_clk clknet_0_clk VDD clkbuf_2_2__f_clk/VPW
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_102_ VDD VSS _069_ net32 _065_ VDD _102_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_195_ VDD net22 clknet_2_3__leaf_clk VSS _020_ VDD _195_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_101_ current_bit\[2\] VDD VSS _068_ net33 current_bit\[1\] VDD _101_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_178_ VDD current_bit\[3\] clknet_2_2__leaf_clk VSS _003_ VDD _178_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_194_ VDD net21 clknet_2_1__leaf_clk VSS _019_ VDD _194_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_177_ _002_ VDD VSS clknet_2_3__leaf_clk current_bit\[2\] VDD _177_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_100_ _067_ VDD VSS _001_ net28 _065_ VDD _100_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_2 VDD VSS VDD FILLER_0_17_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_193_ VDD net20 clknet_2_1__leaf_clk VSS _018_ VDD _193_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_159_ VDD net30 _049_ _020_ _031_ VSS VDD _159_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_176_ _001_ current_bit\[1\] VDD VSS clknet_2_1__leaf_clk VDD _176_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_192_ VDD net19 clknet_2_3__leaf_clk VSS _017_ VDD _192_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_175_ VDD current_bit\[0\] clknet_2_2__leaf_clk VSS _000_ VDD _175_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_31 VDD VSS VDD FILLER_0_12_31/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_96 VDD VSS VDD FILLER_0_18_96/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_158_ net22 VDD VSS _049_ current_bit\[2\] _075_ VDD _158_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_089_ VSS _058_ current_bit\[1\] VDD VDD _089_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_191_ VDD net16 clknet_2_2__leaf_clk VSS _016_ VDD _191_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_174_ net2 VDD VSS _028_ net30 _071_ VDD _174_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_088_ VDD VSS net28 net3 VDD _088_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_157_ _048_ VDD VSS _019_ net3 _086_ VDD _157_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_173_ VDD net29 _056_ _027_ _045_ VSS VDD _173_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_2 VDD VSS VDD FILLER_0_4_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_190_ VDD net6 clknet_2_1__leaf_clk VSS _015_ VDD _190_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_087_ VSS _057_ net33 VDD VDD _087_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_156_ _063_ VDD VSS _048_ _066_ _070_ VDD _156_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_2_3__f_clk VDD VSS clknet_2_3__leaf_clk clknet_0_clk VDD clkbuf_2_3__f_clk/VPW
+ VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_139_ VDD VSS _038_ net34 _074_ VDD _139_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_172_ net18 VDD VSS _056_ _066_ _073_ VDD _172_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_155_ _047_ net29 VDD VSS _018_ current_bit\[3\] _083_ VDD _155_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_138_ VDD VSS _011_ net3 _037_ VDD _138_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_171_ _055_ net29 VDD VSS _026_ _059_ _083_ VDD _171_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_154_ VDD VSS _047_ net20 _082_ VDD _154_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_137_ _036_ VDD VSS _037_ net34 net13 VDD _137_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_2 VDD VSS VDD FILLER_0_13_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_170_ VDD VSS _055_ net17 _042_ VDD _170_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_153_ _046_ net29 VDD VSS _017_ net31 _080_ VDD _153_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_136_ _059_ net32 VDD VSS _036_ net33 current_bit\[1\] VDD _136_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_119_ _070_ VDD VSS _082_ _057_ current_bit\[1\] VDD _119_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_152_ VDD VSS _046_ net19 _079_ VDD _152_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_118_ _081_ net29 VDD VSS _005_ _062_ _079_ VDD _118_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_36 VDD VSS VDD FILLER_0_0_36/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_135_ VDD VSS _010_ net3 _035_ VDD _135_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput3 VSS EOC net3 VDD VDD output3/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_151_ _077_ net28 VDD VSS _016_ _061_ _071_ VDD _151_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_203_ VDD current_state clknet_2_2__leaf_clk VSS _028_ VDD _203_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_134_ _034_ VDD VSS _035_ net34 net12 VDD _134_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_80 VDD VSS VDD FILLER_0_19_80/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_117_ VDD VSS _081_ net7 _079_ VDD _117_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_8 VDD VSS VDD FILLER_0_15_8/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput4 VSS dbot[0] net4 VDD VDD output4/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_0_2 VDD VSS VDD FILLER_0_0_2/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_150_ _045_ VDD VSS _015_ net3 _044_ VDD _150_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_133_ _059_ net32 VDD VSS _034_ _057_ current_bit\[1\] VDD _133_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_202_ VDD net18 clknet_2_0__leaf_clk VSS _027_ VDD _202_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_116_ _076_ VDD VSS _080_ net33 _058_ VDD _116_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput5 VSS dbot[10] net5 VDD VDD output5/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_201_ VDD net17 clknet_2_1__leaf_clk VSS _026_ VDD _201_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_132_ VDD VSS _009_ net3 _033_ VDD _132_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_10_51 VDD VSS VDD FILLER_0_10_51/VPW VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_115_ _070_ VDD VSS _079_ net33 _058_ VDD _115_/VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xoutput6 VSS dbot[11] net6 VDD VDD output6/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
.ends


** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/waffle_1984/waffle_1984-test.sch

.include /home/designer/.volare/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_statistical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice bjt_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical

**.subckt waffle_1984-test
XM2 D G S B pfet_03v3 L=0.5u W=4.38u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1984
**** begin user architecture code


.param v_max=3.3
.param t_on=10n
.param t_total=20n




vg g 0 0
vd d 0 0
vs s 0 6
vb b 0 6
*XDUT0 S G D1   waffle_1984
.control
save all
dc vd 0 6 0.01 vg 0 6 1
write waffle_1984-test.raw
.endc



*.include waffle_1984-noprefix.spice

.include /home/designer/.volare/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/smbb000149.ngspice typical

**** end user architecture code
**.ends
.end

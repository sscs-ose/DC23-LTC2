** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/test/bjt/bjt.sch
.subckt bjt C E G
*.PININFO C:B E:B G:B
Q1 E G C pnp_05p00x05p00 m=1
.ends
.end

* NGSPICE file created from TOP_CHILE_LDO_pex.ext - technology: gf180mcuD

.subckt TOP_CHILE_LDO_pex ref out vdd vss iref
X0 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X3 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X4 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X5 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X6 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X7 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X8 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X9 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X10 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X11 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X12 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X13 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X14 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X15 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X16 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X17 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X18 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X19 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X20 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X21 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X22 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X23 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X24 vdd vdd vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.366214n ps=0.01721 w=25u l=1u
X25 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X26 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X27 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X28 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X29 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X30 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X31 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X32 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X33 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X34 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X35 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X36 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X37 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X38 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X39 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X40 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X41 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X42 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X43 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X44 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X45 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X46 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X47 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X48 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X49 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X50 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X51 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X52 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X53 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X54 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X55 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X56 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X57 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X58 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X59 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X60 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X61 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X62 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X63 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X64 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X65 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X66 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X67 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X68 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X69 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X70 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X71 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X72 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X73 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X74 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X75 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X76 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X77 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X78 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X79 a_206772_74418# iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X80 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X81 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X82 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X83 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X84 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X85 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X86 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X87 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X88 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X89 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X90 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X91 a_210297_77537# ldo_0.ota_0.vin_p a_206772_74418# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X92 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X93 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X94 a_194221_76595# a_194821_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X95 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X96 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X97 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X98 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X99 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X100 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X101 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X102 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X103 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X104 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X105 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X106 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X107 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X108 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X109 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X110 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X111 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X112 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X113 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X114 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X115 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X116 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X117 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X118 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X119 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X120 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X121 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=3.2335p pd=9.38u as=3.8988p ps=13.77u w=4.38u l=0.5u
X122 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X123 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X124 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X125 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X126 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X127 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X128 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X129 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X130 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X131 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X132 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X133 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X134 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X135 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X136 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X137 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X138 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X139 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X140 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X141 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X142 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X143 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X144 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X145 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X146 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X147 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X148 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X149 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X150 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X151 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X152 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X153 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X154 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X155 vss iref ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X156 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X157 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X158 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X159 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X160 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X161 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X162 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X163 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X164 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X165 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X166 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X167 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X168 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X169 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X170 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X171 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X172 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X173 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X174 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X175 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X176 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X177 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X178 a_189421_76595# a_188821_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X179 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X180 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X181 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X182 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X183 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X184 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X185 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X186 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X187 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X188 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X189 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X190 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X191 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X192 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X193 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X194 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X195 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X196 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X197 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X198 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X199 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X200 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X201 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X202 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X203 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X204 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X205 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X206 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X207 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X208 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X209 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X210 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X211 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X212 a_191821_76595# a_190021_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X213 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X214 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X215 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X216 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X217 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X218 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X219 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X220 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X221 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X222 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X223 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X224 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X225 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X226 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X227 ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X228 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X229 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X230 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X231 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X232 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X233 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X234 a_210297_77537# a_209689_77537# vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X235 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X236 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X237 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=2.6079p pd=9.38u as=4.814p ps=13.61u w=4.38u l=0.5u
X238 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X239 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X240 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X241 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X242 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X243 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X244 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X245 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X246 vss vss vss ppolyf_u_1k r_width=1u r_length=5u
X247 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X248 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X249 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X250 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X251 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X252 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X253 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X254 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X255 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X256 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X257 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X258 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X259 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X260 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X261 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X262 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X263 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X264 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X265 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X266 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X267 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X268 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X269 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X270 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X271 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X272 ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X273 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X274 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X275 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X276 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X277 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X278 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X279 vdd a_210297_77537# ldo_0.ota_0.vout vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X280 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X281 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X282 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X283 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X284 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X285 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X286 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X287 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X288 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X289 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X290 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X291 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X292 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X293 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X294 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X295 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X296 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X297 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X298 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X299 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X300 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X301 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X302 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X303 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X304 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X305 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X306 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X307 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X308 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X309 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X310 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X311 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X312 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X313 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X314 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X315 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X316 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X317 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X318 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X319 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X320 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X321 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X322 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X323 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X324 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X325 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X326 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X327 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X328 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X329 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X330 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X331 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X332 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X333 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X334 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X335 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X336 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X337 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X338 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X339 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X340 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X341 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X342 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X343 vss iref iref vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X344 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X345 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X346 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X347 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X348 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X349 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X350 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X351 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X352 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X353 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X354 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X355 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X356 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X357 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X358 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X359 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X360 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X361 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X362 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X363 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X364 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X365 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X366 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X367 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X368 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X369 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X370 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X371 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X372 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X373 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X374 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X375 ldo_0.ota_0.vin_p a_194821_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X376 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X377 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X378 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X379 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X380 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X381 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X382 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X383 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X384 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X385 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X386 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X387 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X388 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X389 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X390 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X391 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X392 vss vss a_206772_74418# vss nfet_03v3 ad=3.05p pd=11.219999u as=1.3p ps=5.52u w=5u l=1u
X393 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X394 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X395 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X396 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X397 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X398 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X399 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X400 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X401 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X402 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X403 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X404 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X405 a_206772_74418# ref a_209689_77537# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X406 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X407 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X408 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X409 ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X410 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X411 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X412 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X413 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X414 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X415 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X416 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X417 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X418 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X419 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X420 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X421 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X422 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X423 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X424 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X425 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X426 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X427 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X428 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X429 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X430 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X431 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X432 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X433 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X434 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X435 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X436 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X437 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X438 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X439 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X440 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X441 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X442 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X443 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X444 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X445 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X446 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X447 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X448 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X449 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X450 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X451 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X452 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X453 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X454 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X455 ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X456 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X457 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X458 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X459 vdd a_210297_77537# ldo_0.ota_0.vout vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X460 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X461 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X462 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X463 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X464 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X465 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X466 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X467 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X468 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X469 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X470 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X471 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X472 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X473 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X474 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X475 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X476 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X477 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X478 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X479 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X480 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X481 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X482 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X483 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X484 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X485 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X486 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X487 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X488 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X489 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X490 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X491 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X492 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X493 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X494 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X495 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X496 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X497 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X498 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X499 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X500 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X501 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X502 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X503 a_193621_76595# a_193021_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X504 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X505 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X506 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X507 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X508 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X509 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X510 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X511 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X512 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X513 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X514 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X515 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X516 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X517 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X518 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X519 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X520 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X521 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X522 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X523 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X524 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X525 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X526 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X527 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X528 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X529 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X530 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X531 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X532 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X533 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X534 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X535 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X536 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X537 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X538 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X539 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X540 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X541 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X542 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X543 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X544 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X545 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X546 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X547 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X548 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X549 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X550 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X551 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X552 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X553 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X554 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X555 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X556 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X557 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X558 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X559 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X560 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X561 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X562 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X563 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X564 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X565 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X566 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X567 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X568 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X569 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X570 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X571 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X572 a_209689_77537# a_209689_77537# vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X573 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X574 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X575 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X576 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X577 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X578 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X579 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X580 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X581 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X582 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X583 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X584 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X585 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X586 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X587 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X588 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X589 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X590 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X591 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X592 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X593 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X594 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X595 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X596 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X597 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X598 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X599 vss vss vss ppolyf_u_1k r_width=1u r_length=20u
X600 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X601 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X602 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X603 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X604 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X605 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X606 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X607 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X608 ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X609 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X610 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X611 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X612 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X613 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X614 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X615 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X616 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X617 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X618 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X619 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X620 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X621 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X622 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X623 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X624 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X625 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X626 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X627 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X628 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X629 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X630 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X631 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X632 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X633 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X634 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X635 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X636 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X637 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X638 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X639 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X640 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X641 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X642 a_189421_76595# a_190621_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X643 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X644 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X645 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X646 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X647 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X648 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X649 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X650 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X651 vss vss vss ppolyf_u_1k r_width=1u r_length=20u
X652 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X653 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X654 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X655 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X656 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X657 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X658 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X659 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X660 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X661 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X662 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X663 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X664 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X665 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X666 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X667 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X668 a_211573_72398# a_212701_72398# vss ppolyf_u_1k r_width=1u r_length=5u
X669 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X670 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X671 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X672 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X673 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X674 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X675 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X676 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X677 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X678 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X679 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X680 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X681 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X682 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X683 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X684 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X685 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X686 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X687 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X688 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X689 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X690 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X691 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X692 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X693 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X694 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X695 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X696 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X697 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X698 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X699 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X700 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X701 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X702 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X703 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X704 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X705 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X706 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X707 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X708 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X709 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X710 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X711 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X712 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X713 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X714 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X715 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X716 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X717 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X718 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X719 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X720 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X721 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X722 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X723 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X724 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X725 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X726 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X727 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X728 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X729 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X730 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X731 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X732 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X733 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X734 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X735 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X736 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X737 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X738 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X739 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X740 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X741 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X742 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X743 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X744 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X745 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X746 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X747 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X748 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X749 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X750 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X751 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X752 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X753 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X754 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X755 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X756 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X757 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X758 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X759 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X760 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X761 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X762 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X763 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X764 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X765 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X766 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X767 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X768 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X769 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X770 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X771 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X772 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X773 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X774 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X775 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X776 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X777 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X778 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X779 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X780 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X781 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X782 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X783 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X784 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X785 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=33.475p ps=0.14433m w=2.5u l=1u
X786 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X787 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X788 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X789 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X790 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X791 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X792 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X793 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X794 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X795 a_193621_76595# a_195421_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X796 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X797 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X798 a_206772_74418# vss vss vss nfet_03v3 ad=1.3p pd=5.52u as=3.075p ps=11.23u w=5u l=1u
X799 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X800 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X801 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X802 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X803 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X804 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X805 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X806 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X807 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X808 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X809 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X810 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X811 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X812 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X813 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X814 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X815 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X816 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X817 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X818 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X819 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X820 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X821 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X822 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X823 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X824 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X825 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X826 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X827 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X828 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X829 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X830 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X831 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X832 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X833 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X834 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X835 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X836 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X837 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=0 ps=0 w=2.5u l=1u
X838 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X839 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X840 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X841 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X842 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X843 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X844 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X845 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X846 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X847 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X848 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X849 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X850 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X851 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X852 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X853 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X854 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X855 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X856 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X857 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X858 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X859 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X860 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X861 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X862 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X863 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X864 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X865 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X866 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X867 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X868 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X869 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X870 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X871 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X872 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X873 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=2.6079p pd=9.38u as=4.814p ps=13.61u w=4.38u l=0.5u
X874 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X875 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X876 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X877 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X878 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X879 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X880 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X881 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X882 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X883 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X884 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X885 iref iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X886 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X887 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X888 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X889 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X890 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X891 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X892 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X893 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X894 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X895 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X896 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X897 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X898 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X899 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X900 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X901 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X902 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X903 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X904 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X905 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X906 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X907 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X908 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X909 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X910 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X911 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X912 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X913 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X914 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X915 a_191821_76595# a_192421_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X916 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X917 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X918 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X919 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X920 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X921 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X922 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X923 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X924 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X925 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X926 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X927 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X928 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X929 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X930 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X931 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X932 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X933 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X934 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X935 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X936 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X937 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X938 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X939 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X940 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X941 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X942 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X943 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X944 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X945 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X946 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X947 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X948 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X949 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X950 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X951 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X952 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X953 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X954 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X955 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X956 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X957 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X958 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X959 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X960 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X961 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X962 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X963 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X964 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X965 a_211573_72398# a_210297_77537# vss ppolyf_u_1k r_width=1u r_length=5u
X966 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=2.6079p ps=9.38u w=4.38u l=0.5u
X967 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X968 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X969 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X970 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X971 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X972 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X973 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X974 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X975 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X976 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X977 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X978 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X979 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X980 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X981 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X982 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X983 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X984 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X985 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X986 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X987 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X988 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X989 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X990 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X991 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X992 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X993 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X994 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X995 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X996 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X997 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X998 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X999 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1000 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1001 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=2.6079p ps=9.38u w=4.38u l=0.5u
X1002 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1003 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1004 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1005 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1006 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1007 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1008 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1009 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1010 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1011 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1012 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1013 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1014 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1015 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1016 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1017 ldo_0.ota_0.vout a_210297_77537# vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X1018 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1019 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1020 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1021 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1022 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1023 vdd vdd vdd vdd pfet_03v3 ad=3.25p pd=11.299999u as=0 ps=0 w=5u l=1u
X1024 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1025 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1026 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1027 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1028 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1029 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1030 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1031 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1032 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1033 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1034 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1035 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1036 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1037 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1038 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1039 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1040 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1041 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1042 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1043 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1044 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1045 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1046 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1047 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1048 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1049 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1050 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1051 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1052 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1053 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1054 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1055 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1056 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1057 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1058 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1059 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1060 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=0 ps=0 w=2.5u l=1u
X1061 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1062 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1063 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1064 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1065 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1066 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1067 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1068 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1069 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1070 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1071 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1072 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1073 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1074 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1075 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1076 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1077 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1078 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1079 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1080 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1081 a_196021_76595# a_197221_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1082 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1083 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1084 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1085 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1086 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1087 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1088 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1089 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1090 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1091 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1092 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1093 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1094 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1095 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1096 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1097 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1098 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1099 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1100 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1101 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1102 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1103 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1104 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1105 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1106 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1107 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1108 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1109 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1110 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1111 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1112 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1113 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1114 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1115 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1116 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1117 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1118 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1119 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1120 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1121 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1122 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1123 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1124 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1125 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1126 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1127 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1128 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1129 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1130 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1131 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1132 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1133 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1134 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1135 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1136 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1137 vss iref ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1138 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1139 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1140 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1141 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1142 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1143 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1144 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1145 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1146 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1147 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1148 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1149 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1150 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1151 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1152 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1153 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1154 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1155 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1156 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1157 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1158 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1159 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1160 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1161 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1162 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1163 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1164 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1165 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1166 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1167 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1168 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1169 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1170 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1171 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1172 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1173 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1174 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1175 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1176 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1177 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1178 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1179 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1180 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1181 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1182 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1183 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1184 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1185 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1186 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1187 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1188 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1189 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1190 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1191 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1192 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1193 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1194 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1195 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1196 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1197 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1198 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1199 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1200 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1201 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1202 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1203 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1204 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1205 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1206 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1207 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1208 a_194221_76595# a_192421_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1209 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1210 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1211 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1212 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1213 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1214 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1215 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1216 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1217 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1218 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1219 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1220 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1221 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1222 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1223 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1224 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1225 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=3.2335p ps=9.38u w=4.38u l=0.5u
X1226 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1227 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1228 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1229 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1230 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1231 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1232 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1233 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1234 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1235 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1236 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1237 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1238 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1239 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1240 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1241 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1242 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1243 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1244 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1245 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1246 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1247 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1248 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1249 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1250 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1251 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1252 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1253 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1254 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1255 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1256 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1257 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1258 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1259 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1260 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1261 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1262 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1263 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1264 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1265 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1266 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1267 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1268 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1269 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1270 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1271 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1272 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1273 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1274 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1275 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1276 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1277 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1278 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1279 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1280 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1281 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1282 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1283 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1284 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1285 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1286 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1287 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1288 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1289 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1290 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1291 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1292 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1293 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1294 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1295 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1296 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1297 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1298 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1299 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1300 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1301 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1302 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1303 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1304 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1305 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1306 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1307 vdd vdd vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=0 ps=0 w=5u l=1u
X1308 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1309 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1310 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1311 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1312 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1313 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1314 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1315 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1316 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1317 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1318 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1319 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1320 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1321 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1322 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1323 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1324 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1325 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1326 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1327 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1328 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1329 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1330 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1331 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1332 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1333 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1334 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1335 vss iref ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1336 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1337 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1338 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1339 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1340 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1341 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1342 a_191221_76595# a_190621_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1343 ldo_0.ota_0.vout a_210297_77537# vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X1344 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1345 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1346 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1347 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1348 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1349 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1350 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1351 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1352 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1353 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1354 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1355 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1356 a_206772_74418# ldo_0.ota_0.vin_p a_210297_77537# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1357 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1358 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1359 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1360 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1361 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1362 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1363 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1364 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1365 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1366 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1367 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1368 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1369 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1370 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1371 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1372 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1373 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1374 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1375 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1376 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1377 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1378 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1379 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1380 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1381 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1382 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1383 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1384 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1385 vss vss vss ppolyf_u_1k r_width=1u r_length=5u
X1386 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1387 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1388 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1389 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1390 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1391 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1392 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1393 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1394 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1395 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1396 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1397 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1398 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1399 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1400 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1401 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1402 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1403 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1404 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1405 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1406 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1407 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1408 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1409 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1410 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1411 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1412 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1413 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1414 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1415 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1416 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1417 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1418 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1419 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1420 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1421 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1422 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1423 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1424 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1425 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1426 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1427 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1428 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1429 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1430 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1431 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1432 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1433 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1434 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1435 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1436 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1437 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1438 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1439 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1440 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1441 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1442 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1443 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1444 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1445 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1446 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1447 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1448 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1449 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1450 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1451 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1452 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1453 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1454 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1455 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1456 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1457 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1458 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1459 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1460 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1461 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1462 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1463 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1464 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1465 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1466 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1467 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1468 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1469 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1470 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1471 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1472 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1473 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1474 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1475 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1476 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1477 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1478 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1479 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1480 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1481 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1482 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1483 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1484 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1485 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1486 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1487 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1488 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1489 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1490 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1491 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=3.2335p pd=9.38u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1492 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1493 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1494 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1495 a_196021_76595# a_195421_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1496 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1497 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1498 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1499 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1500 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1501 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1502 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1503 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1504 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1505 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1506 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1507 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1508 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1509 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1510 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1511 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1512 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1513 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1514 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1515 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1516 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1517 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1518 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1519 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1520 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1521 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1522 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1523 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1524 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1525 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1526 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1527 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1528 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1529 out a_188821_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1530 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1531 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1532 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1533 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1534 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1535 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1536 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1537 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1538 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1539 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1540 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1541 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1542 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1543 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1544 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1545 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1546 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1547 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1548 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1549 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1550 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1551 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1552 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1553 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1554 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1555 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1556 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1557 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1558 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1559 vss iref a_206772_74418# vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1560 vdd a_209689_77537# a_209689_77537# vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1561 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1562 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1563 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1564 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1565 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1566 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1567 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1568 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1569 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1570 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1571 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1572 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1573 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1574 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1575 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1576 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1577 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1578 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1579 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1580 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1581 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1582 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1583 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1584 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1585 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1586 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1587 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1588 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1589 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1590 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1591 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1592 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1593 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1594 ldo_0.ota_0.vout a_212701_72398# cap_mim_2f0_m4m5_noshield c_width=22u c_length=22u
X1595 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1596 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1597 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1598 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1599 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1600 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1601 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1602 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1603 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1604 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1605 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1606 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1607 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1608 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1609 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1610 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1611 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1612 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1613 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1614 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1615 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1616 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1617 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1618 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1619 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1620 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1621 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1622 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1623 a_191221_76595# a_193021_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1624 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1625 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1626 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1627 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1628 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1629 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1630 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1631 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1632 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1633 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1634 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1635 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1636 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1637 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1638 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1639 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1640 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1641 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1642 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1643 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1644 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1645 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1646 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1647 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1648 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1649 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1650 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1651 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1652 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1653 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1654 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1655 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1656 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1657 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1658 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1659 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1660 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=0 ps=0 w=2.5u l=1u
X1661 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1662 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1663 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1664 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1665 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1666 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1667 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1668 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1669 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1670 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1671 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1672 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1673 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1674 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1675 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1676 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1677 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1678 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1679 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1680 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1681 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1682 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1683 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1684 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1685 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1686 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1687 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1688 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1689 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1690 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1691 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1692 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1693 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1694 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1695 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1696 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1697 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1698 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1699 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1700 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1701 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1702 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1703 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1704 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1705 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1706 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1707 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1708 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1709 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1710 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1711 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1712 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1713 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1714 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1715 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1716 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1717 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1718 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1719 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1720 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1721 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1722 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1723 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1724 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1725 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1726 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1727 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1728 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1729 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1730 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1731 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1732 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1733 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1734 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1735 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1736 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1737 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1738 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1739 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1740 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1741 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1742 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1743 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1744 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1745 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1746 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1747 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1748 vdd a_209689_77537# a_210297_77537# vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1749 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1750 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1751 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1752 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1753 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1754 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1755 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1756 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1757 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1758 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1759 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1760 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1761 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1762 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1763 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1764 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1765 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1766 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1767 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1768 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1769 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1770 vss a_190021_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1771 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1772 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1773 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1774 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1775 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1776 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1777 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1778 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1779 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1780 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1781 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1782 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1783 vss iref ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1784 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1785 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1786 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1787 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1788 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1789 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1790 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1791 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1792 vdd vdd vdd vdd pfet_03v3 ad=16.25p pd=51.3u as=0 ps=0 w=25u l=1u
X1793 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1794 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1795 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1796 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1797 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1798 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1799 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1800 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1801 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1802 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1803 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1804 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1805 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1806 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1807 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1808 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1809 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1810 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1811 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1812 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1813 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1814 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1815 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1816 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1817 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1818 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1819 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1820 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1821 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1822 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1823 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1824 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1825 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1826 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1827 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1828 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1829 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1830 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1831 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1832 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1833 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1834 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1835 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1836 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1837 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1838 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1839 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1840 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1841 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1842 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1843 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1844 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1845 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1846 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1847 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1848 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1849 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1850 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1851 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1852 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1853 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1854 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1855 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1856 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1857 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1858 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1859 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1860 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1861 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1862 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1863 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1864 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1865 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1866 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1867 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1868 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1869 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1870 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1871 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1872 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1873 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1874 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1875 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1876 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1877 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1878 a_209689_77537# ref a_206772_74418# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1879 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1880 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1881 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1882 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1883 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1884 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1885 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1886 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1887 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1888 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1889 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1890 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1891 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1892 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1893 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1894 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1895 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1896 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1897 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1898 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1899 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1900 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=3.2335p ps=9.38u w=4.38u l=0.5u
X1901 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1902 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1903 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1904 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1905 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1906 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1907 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1908 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1909 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1910 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1911 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1912 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1913 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1914 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1915 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1916 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1917 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1918 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1919 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1920 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1921 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1922 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1923 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1924 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1925 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1926 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1927 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1928 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1929 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1930 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1931 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1932 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1933 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1934 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1935 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1936 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1937 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1938 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1939 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1940 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1941 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1942 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1943 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1944 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1945 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1946 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1947 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1948 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1949 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1950 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1951 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1952 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1953 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1954 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1955 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1956 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1957 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1958 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1959 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1960 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1961 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1962 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1963 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1964 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1965 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1966 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1967 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1968 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1969 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1970 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1971 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1972 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1973 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1974 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1975 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1976 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1977 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1978 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1979 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1980 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1981 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1982 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1983 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1984 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1985 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1986 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1987 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1988 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1989 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1990 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1991 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1992 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1993 ldo_0.ota_0.vin_p a_197221_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1994 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1995 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1996 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1997 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1998 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1999 vss iref ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X2000 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2001 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2002 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2003 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2004 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2005 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2006 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2007 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X2008 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2009 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2010 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2011 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2012 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2013 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2014 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2015 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2016 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2017 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2018 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2019 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2020 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2021 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2022 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2023 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2024 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2025 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X2026 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2027 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2028 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2029 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2030 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2031 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2032 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2033 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2034 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2035 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X2036 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2037 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2038 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2039 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X2040 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2041 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2042 out ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2043 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2044 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2045 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2046 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2047 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2048 vdd ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
C0 out a_189421_76595# 0.120238f
C1 vdd a_210297_77537# 9.19771f
C2 a_191221_76595# a_189421_76595# 0.14109f
C3 a_206772_74418# a_209689_77537# 0.250752f
C4 a_191221_76595# a_191821_76595# 0.802011f
C5 a_206772_74418# ldo_0.ota_0.vin_p 1.25837f
C6 vdd iref 12.6709f
C7 vdd ldo_0.ota_0.vout 1.77298p
C8 a_206772_74418# vdd 1.60493f
C9 a_210297_77537# ldo_0.ota_0.vout 2.87172f
C10 a_195421_72467# a_194821_72467# 0.864964f
C11 vdd out 2.35078p
C12 a_206772_74418# a_210297_77537# 0.514834f
C13 a_192421_72467# a_190021_72467# 0.14109f
C14 iref ldo_0.ota_0.vout 1.74891f
C15 vdd a_188821_72467# 0.121652f
C16 a_209689_77537# ref 1.11601f
C17 a_206772_74418# iref 0.340145f
C18 a_212701_72398# vdd 0.511061f
C19 a_196021_76595# a_193621_76595# 0.14109f
C20 out ldo_0.ota_0.vout 1.31128p
C21 a_192421_72467# a_193021_72467# 0.864964f
C22 a_212701_72398# a_210297_77537# 0.332743f
C23 a_192421_72467# a_194821_72467# 0.14109f
C24 vdd ref 8.751969f
C25 a_188821_72467# a_190021_72467# 0.120932f
C26 a_190621_72467# a_190021_72467# 0.864964f
C27 a_212701_72398# iref 0.423537f
C28 a_194221_76595# a_193621_76595# 0.802011f
C29 a_212701_72398# ldo_0.ota_0.vout 2.74789f
C30 a_194821_72467# a_197221_72467# 0.120932f
C31 a_196021_76595# ldo_0.ota_0.vin_p 0.592967f
C32 ref iref 0.300994f
C33 a_209689_77537# ldo_0.ota_0.vin_p 0.412413f
C34 a_206772_74418# ref 2.52489f
C35 a_209689_77537# vdd 3.29537f
C36 m1_197211_77525# ldo_0.ota_0.vin_p 0.10346f
C37 a_209689_77537# a_210297_77537# 0.91529f
C38 a_210297_77537# ldo_0.ota_0.vin_p 1.11127f
C39 a_191221_76595# a_193621_76595# 0.14109f
C40 iref vss 18.8374f
C41 ref vss 10.4156f
C42 out vss 0.147504p
C43 vdd vss 25.2192p
C44 m1_198411_71393# vss 0.237793f $ **FLOATING
C45 m1_196611_71393# vss 0.193159f $ **FLOATING
C46 m1_194811_71393# vss 0.192608f $ **FLOATING
C47 m1_194211_71393# vss 0.193159f $ **FLOATING
C48 m1_192411_71393# vss 0.192608f $ **FLOATING
C49 m1_191811_71393# vss 0.193159f $ **FLOATING
C50 m1_190011_71393# vss 0.192608f $ **FLOATING
C51 m1_188211_71393# vss 0.217848f $ **FLOATING
C52 m1_198411_71793# vss 0.269211f $ **FLOATING
C53 m1_188211_71793# vss 0.248714f $ **FLOATING
C54 m1_198411_77125# vss 0.31235f $ **FLOATING
C55 m1_188211_77125# vss 0.270516f $ **FLOATING
C56 m1_198411_77525# vss 0.262201f $ **FLOATING
C57 m1_197211_77525# vss 0.195149f $ **FLOATING
C58 m1_196011_77525# vss 0.205536f $ **FLOATING
C59 m1_195411_77525# vss 0.205536f $ **FLOATING
C60 m1_193611_77525# vss 0.205536f $ **FLOATING
C61 m1_193011_77525# vss 0.205536f $ **FLOATING
C62 m1_191211_77525# vss 0.205536f $ **FLOATING
C63 m1_190611_77525# vss 0.269682f $ **FLOATING
C64 m1_189411_77525# vss 0.267473f $ **FLOATING
C65 m1_188211_77525# vss 0.227432f $ **FLOATING
C66 a_212701_72398# vss 3.08142f
C67 a_211573_72398# vss 1.30871f
C68 a_197221_72467# vss 1.84846f
C69 a_196021_76595# vss 2.16629f
C70 a_195421_72467# vss 1.55755f
C71 a_194821_72467# vss 1.94527f
C72 a_194221_76595# vss 1.80662f
C73 a_193621_76595# vss 2.46883f
C74 a_193021_72467# vss 1.56132f
C75 a_192421_72467# vss 1.93093f
C76 a_191821_76595# vss 1.81178f
C77 a_191221_76595# vss 2.46883f
C78 a_190621_72467# vss 1.55755f
C79 a_190021_72467# vss 1.94527f
C80 a_189421_76595# vss 2.67953f
C81 a_188821_72467# vss 1.81856f
C82 a_210297_77537# vss 3.7114f
C83 a_209689_77537# vss 1.53708f
C84 a_206772_74418# vss 5.20193f
C85 ldo_0.ota_0.vin_p vss 12.9019f
C86 ldo_0.ota_0.vout vss 0.129471p
.ends


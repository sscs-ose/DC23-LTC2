* Extracted by KLayout with GF180MCU LVS runset on : 30/12/2023 05:58

.SUBCKT resistor_core IN1 IN2 gf180mcu_gnd
R$1 IN1 IN2 gf180mcu_gnd 7000 ppolyf_u L=20U W=1U
.ENDS resistor_core

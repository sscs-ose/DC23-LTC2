* Extracted by KLayout with GF180MCU LVS runset on : 24/12/2023 04:22

* cell resistor_core
* pin A,B,BULK
* pin gf180mcu_gnd
.SUBCKT resistor_core A|B|BULK gf180mcu_gnd
* device instance $1 r0 *1 9.505,0.36 ppolyf_u
R$1 A|B|BULK A|B|BULK gf180mcu_gnd 7000 ppolyf_u L=20U W=1U
.ENDS resistor_core

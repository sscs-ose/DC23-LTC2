** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/test/resistor_core/resistor_core.sch
.subckt resistor_core IN2 IN1 B
*.PININFO IN2:B IN1:B B:B
R2 IN2 IN1 B ppolyf_u W=1e-6 L=20e-6 m=1
.ends
.end

** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/test/waffle_1984/waffle_1984.sch
**.subckt waffle_1984 S G D
*.iopin S
*.iopin G
*.iopin D
XM1 D G S S pfet_03v3 L=0.5u W=4.38u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1860
**.ends
.end

* Extracted by KLayout with GF180MCU LVS runset on : 27/12/2023 05:25

* cell pmos
* pin S
* pin D
* pin G
.SUBCKT pmos S D G
* device instance $1 r0 *1 0.35,0.5 pfet_03v3
M$1 S G D S pfet_03v3 L=0.7U W=5U AS=1.69P AD=1.69P PS=9.38U PD=9.38U
.ENDS pmos

** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/resistor/resistor.sch
**.subckt resistor OUT1 VSS VDD B OUT2
*.iopin OUT1
*.iopin VSS
*.iopin VDD
*.iopin B
*.iopin OUT2
XR1 OUT1 VDD B ppolyf_u r_width=1e-6 r_length=200e-6 m=1
XR2 VSS OUT2 B ppolyf_u r_width=1e-6 r_length=120e-6 m=1
XR3 B B B ppolyf_u r_width=1e-6 r_length=20e-6 m=1
XR4 B B B ppolyf_u r_width=1e-6 r_length=20e-6 m=1
**.ends
.end

** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/ldo/ldo-full-test.sch

.include /home/designer/.volare/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_statistical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical

**.subckt ldo-full-test out
*.iopin out
I1 GND net1 3u
V1 ref GND 1.25
XM1 out op_out vin vin pfet_03v3 L=0.3u W=10u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=800
XR1 net2 out GND ppolyf_u_2k r_width=1e-6 r_length=164e-6 m=1
XR2 GND pos GND ppolyf_u_2k r_width=1e-6 r_length=100e-6 m=1
v4 net2 pos 0
X1 op_out GND vin net3 ref net1 ota-ldo
vt net3 pos 0
**** begin user architecture code

.param R=66
R10 out 0 {R}
IL out 0 PWL(0 0.1m 10u 0.1m 20u 10m 30u 10m)
*CL out 0 10p

Vs vin 0 PULSE(5 5 50u 20u 1u 100u 100u)

.nodeset v(out)=0
.nodeset v(x1.pos)=0

*TRANSIENT
.control
save all
tran 1ns 200us
let gds =
print ic
plot gds
plot v(out) v(ref) v(pos) v(vin)
*plot v(op_out)
*plot v(out)
*plot i(out)
*plot i(v3)*v(vin)
.endc



*SUPPLY SWEEP
.control
dc Vs 4 0 -0.01
plot v(out) v(ref) v(vin)
*plot v(x1.op_out)
*plot i(v.x1.v4)
.endc

*Stability_Analysis (openloop)
.control
alter Vs AC=0
alter Vt AC =1
ac dec 100 1 1G
plot vdb(out)
let phase_val = 180/PI*cph(out)
plot phase_val
meas ac pm FIND phase_val WHEN vdb(out)=0
*plot (180/pi)*vp(out)
*let gm0=
*let Zout=(1.5)/(gm0*v(op_out))
*let Zout2=v(out)/gm0
*plot vdb(Zout2)
*wrdata /foss/designs/LDO_Design/data/data_PSRR.dat vdb(out)
.endc

*PSRR_Analysis
.control
alter Vs AC =1
alter Vt AC=0
ac dec 100 1 1G
plot vdb(out)
let phase_val = 180/PI*cph(out)
plot phase_val
*plot (180/pi)*vp(out)
*let gm0=
*let Zout=(1.5)/(gm0*v(op_out))
*let Zout2=v(out)/gm0
*plot vdb(Zout2)
*wrdata /foss/designs/LDO_Design/data/data_PSRR.dat vdb(out)
.endc


**Load_Transient
.control
alter IL 50u
alter R10 3600k
tran 0.1u 100u
meas TRAN V_ldo_100u FIND v(out) AT=5u
meas TRAN V_ldo_10m FIND v(out) AT=100u
let load_reg= V_ldo_100u-V_ldo_10m
let load_current =(-1*i(Vs)-131.8e-6)
print load_reg
plot load_current v(out)-3.3
.endc



.control
alter R10 36k
alter  0 0 10u 0 20u 0 30u 0 ]
alter  3.3 50u 1u 1u 10u 100u]
alter IL 0
tran 0.1u 100u
plot v(vin) v(out)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  ota-ldo.sym # of pins=6
** sym_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/ota-ldo/ota-ldo.sym
** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/ota-ldo/ota-ldo.sch
.subckt ota-ldo out agnd avdd pos neg vb
*.iopin vb
*.iopin avdd
*.iopin agnd
*.ipin neg
*.ipin pos
*.opin out
XC2 net2 net4 cap_mim_2f0fF c_width=50e-6 c_length=50e-6 m=1
XM1 net1 neg net3 agnd nfet_03v3 L=0.5u W=9u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 net1 avdd avdd pfet_03v3 L=1.5u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net2 pos net3 agnd nfet_03v3 L=0.5u W=9u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net2 net1 avdd avdd pfet_03v3 L=1.5u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 net3 vb agnd agnd nfet_03v3 L=0.7u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 vb vb agnd agnd nfet_03v3 L=0.7u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 out net2 avdd avdd pfet_03v3 L=0.5u W=35u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 out vb agnd agnd nfet_03v3 L=0.7u W=36.3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
R1 net4 out 10k m=1
.ends

.GLOBAL GND
.end

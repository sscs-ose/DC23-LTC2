* Extracted by KLayout with GF180MCU LVS runset on : 27/12/2023 05:24

* cell resistor_core
* pin A
* pin B
.SUBCKT resistor_core A B
* device instance $1 r0 *1 9.505,0.36 ppolyf_u
R$1 A B B 7000 ppolyf_u L=20U W=1U
.ENDS resistor_core

* NGSPICE file created from open_ldo_pex.ext - technology: gf180mcuD

.subckt open_ldo_pex out vin_p feedback ref iref vdd vss
X0 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X2 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X3 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X4 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X5 a_29974_15620# out vss ppolyf_u_1k r_width=1u r_length=20u
X6 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X7 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X8 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X9 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X10 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X11 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X12 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X13 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X14 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X15 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X16 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X17 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X18 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X19 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=33.475p ps=0.14433m w=2.5u l=1u
X20 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X21 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X22 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X23 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X24 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X25 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X26 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X27 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X28 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X29 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X30 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X31 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X32 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X33 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X34 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X35 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X36 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X37 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X38 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X39 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X40 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X41 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X42 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X43 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X44 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X45 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X46 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X47 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X48 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X49 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X50 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X51 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X52 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X53 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X54 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X55 vdd ota_0.vout out vdd pfet_03v3 ad=3.2335p pd=9.38u as=3.8988p ps=13.77u w=4.38u l=0.5u
X56 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X57 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X58 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X59 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X60 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X61 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X62 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X63 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X64 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X65 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X66 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X67 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X68 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X69 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X70 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X71 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X72 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X73 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X74 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X75 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X76 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X77 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X78 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X79 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X80 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X81 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X82 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X83 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X84 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X85 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X86 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X87 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X88 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X89 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X90 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X91 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X92 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X93 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X94 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X95 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X96 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X97 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X98 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X99 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X100 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X101 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X102 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X103 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X104 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X105 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X106 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X107 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X108 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X109 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X110 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X111 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X112 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X113 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X114 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X115 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X116 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X117 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X118 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X119 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X120 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X121 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X122 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X123 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X124 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X125 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X126 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X127 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X128 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X129 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X130 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X131 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X132 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X133 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X134 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X135 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X136 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X137 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X138 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X139 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X140 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X141 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X142 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X143 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X144 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X145 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X146 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X147 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X148 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X149 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X150 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X151 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X152 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X153 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X154 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X155 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X156 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X157 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X158 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X159 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X160 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X161 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X162 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X163 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X164 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X165 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X166 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X167 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X168 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X169 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X170 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X171 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X172 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X173 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X174 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X175 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X176 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X177 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X178 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X179 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X180 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X181 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X182 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X183 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X184 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X185 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X186 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X187 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X188 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X189 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X190 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X191 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X192 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X193 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X194 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X195 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X196 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X197 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X198 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X199 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X200 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X201 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X202 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X203 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X204 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X205 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X206 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X207 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X208 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X209 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X210 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X211 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X212 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X213 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X214 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X215 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X216 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X217 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X218 a_29974_9020# a_34102_7820# vss ppolyf_u_1k r_width=1u r_length=20u
X219 vdd a_34724_n8101# a_34724_n8101# vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X220 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X221 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X222 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X223 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X224 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X225 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X226 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X227 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X228 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X229 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X230 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X231 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X232 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X233 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X234 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X235 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X236 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X237 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X238 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X239 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X240 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X241 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X242 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X243 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X244 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X245 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X246 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X247 ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X248 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X249 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X250 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X251 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X252 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X253 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X254 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X255 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X256 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X257 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X258 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X259 a_29974_13220# a_34102_12620# vss ppolyf_u_1k r_width=1u r_length=20u
X260 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X261 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X262 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X263 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X264 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=2.6079p ps=9.38u w=4.38u l=0.5u
X265 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X266 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X267 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X268 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X269 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X270 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X271 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X272 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X273 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X274 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X275 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X276 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X277 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X278 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X279 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X280 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X281 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X282 ota_0.cm_nmos_0.iout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X283 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X284 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X285 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X286 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X287 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X288 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X289 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X290 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X291 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X292 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X293 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X294 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X295 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X296 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X297 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X298 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X299 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X300 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X301 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X302 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X303 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X304 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X305 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X306 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X307 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X308 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X309 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X310 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X311 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X312 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X313 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X314 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X315 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X316 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X317 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X318 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X319 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X320 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X321 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X322 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X323 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X324 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X325 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X326 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X327 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X328 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X329 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X330 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X331 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X332 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X333 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X334 vss vss vss ppolyf_u_1k r_width=1u r_length=20u
X335 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X336 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X337 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X338 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X339 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X340 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X341 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X342 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X343 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X344 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X345 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X346 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X347 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X348 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X349 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X350 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X351 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X352 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X353 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X354 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X355 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X356 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X357 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X358 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X359 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X360 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X361 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X362 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X363 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X364 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X365 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X366 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X367 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X368 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X369 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X370 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X371 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X372 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X373 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X374 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X375 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X376 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X377 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X378 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X379 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X380 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X381 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X382 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X383 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X384 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X385 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X386 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X387 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X388 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X389 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X390 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X391 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X392 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X393 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X394 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=0 ps=0 w=2.5u l=1u
X395 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X396 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X397 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X398 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X399 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X400 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X401 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X402 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=3.2335p ps=9.38u w=4.38u l=0.5u
X403 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X404 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X405 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X406 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X407 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X408 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X409 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X410 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X411 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X412 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X413 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X414 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X415 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X416 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X417 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X418 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X419 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X420 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X421 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X422 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X423 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X424 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X425 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X426 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X427 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X428 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X429 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X430 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X431 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X432 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X433 vdd a_30505_n7588# ota_0.vout vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X434 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X435 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X436 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X437 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X438 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X439 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X440 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X441 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X442 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X443 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X444 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X445 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X446 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X447 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X448 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X449 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X450 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X451 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X452 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X453 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X454 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X455 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X456 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X457 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X458 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X459 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X460 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X461 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X462 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X463 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X464 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X465 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X466 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X467 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X468 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X469 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X470 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X471 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X472 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X473 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X474 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X475 a_29974_8420# a_34102_10220# vss ppolyf_u_1k r_width=1u r_length=20u
X476 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X477 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X478 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X479 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X480 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X481 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X482 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X483 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X484 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X485 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X486 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X487 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X488 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X489 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X490 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X491 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X492 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X493 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X494 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X495 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X496 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X497 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X498 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X499 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X500 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X501 ota_0.vout a_30505_n7588# vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X502 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X503 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X504 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X505 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X506 iref iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X507 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X508 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X509 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X510 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X511 a_29974_9020# a_34102_9620# vss ppolyf_u_1k r_width=1u r_length=20u
X512 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X513 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X514 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X515 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X516 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X517 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X518 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X519 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X520 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X521 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X522 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X523 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X524 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X525 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X526 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X527 ota_0.cm_nmos_0.iout ref a_34724_n8101# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X528 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X529 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X530 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X531 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X532 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X533 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X534 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X535 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X536 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X537 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X538 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X539 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X540 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X541 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X542 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X543 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X544 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X545 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X546 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X547 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X548 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X549 a_29974_13820# a_34102_12020# vss ppolyf_u_1k r_width=1u r_length=20u
X550 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X551 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X552 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X553 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X554 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X555 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X556 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X557 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X558 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X559 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X560 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X561 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X562 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X563 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X564 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X565 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X566 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X567 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X568 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X569 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X570 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X571 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X572 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X573 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X574 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X575 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X576 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X577 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X578 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X579 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X580 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X581 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X582 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X583 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X584 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X585 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X586 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X587 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X588 vdd a_34724_n8101# a_30505_n7588# vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X589 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X590 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X591 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X592 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X593 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X594 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X595 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X596 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X597 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X598 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X599 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X600 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X601 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X602 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X603 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X604 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X605 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X606 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X607 vss vss vss ppolyf_u_1k r_width=1u r_length=5u
X608 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X609 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X610 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X611 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X612 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X613 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X614 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X615 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X616 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X617 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X618 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X619 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X620 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X621 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X622 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X623 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X624 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X625 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X626 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X627 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X628 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X629 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X630 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X631 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X632 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X633 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X634 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X635 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X636 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X637 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X638 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X639 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X640 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X641 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X642 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X643 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X644 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X645 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X646 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X647 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X648 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X649 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X650 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X651 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X652 ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X653 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X654 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X655 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X656 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X657 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X658 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X659 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X660 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X661 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X662 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X663 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X664 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X665 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X666 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X667 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X668 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X669 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X670 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X671 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X672 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X673 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X674 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X675 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X676 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X677 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X678 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X679 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X680 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X681 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X682 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X683 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X684 vdd vdd vdd vdd pfet_03v3 ad=3.25p pd=11.299999u as=6.366214n ps=0.01721 w=5u l=1u
X685 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X686 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X687 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X688 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X689 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X690 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X691 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X692 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X693 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X694 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X695 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X696 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X697 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X698 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X699 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X700 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X701 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X702 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X703 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X704 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X705 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X706 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X707 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X708 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X709 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X710 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X711 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X712 vss vss vss ppolyf_u_1k r_width=1u r_length=20u
X713 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X714 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X715 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X716 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X717 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X718 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X719 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X720 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X721 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X722 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X723 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X724 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X725 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X726 vss iref ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X727 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X728 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X729 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X730 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X731 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X732 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X733 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X734 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X735 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X736 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X737 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X738 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X739 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X740 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X741 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X742 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X743 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=3.2335p ps=9.38u w=4.38u l=0.5u
X744 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X745 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X746 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X747 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X748 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X749 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X750 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X751 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X752 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X753 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X754 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X755 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X756 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X757 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X758 a_29974_10820# a_34102_10220# vss ppolyf_u_1k r_width=1u r_length=20u
X759 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X760 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X761 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X762 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X763 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X764 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X765 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X766 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X767 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X768 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X769 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X770 vdd vdd vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=0 ps=0 w=5u l=1u
X771 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X772 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X773 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X774 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X775 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X776 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X777 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X778 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X779 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X780 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X781 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X782 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X783 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X784 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X785 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X786 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X787 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X788 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X789 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X790 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X791 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X792 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X793 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X794 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X795 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X796 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X797 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X798 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X799 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X800 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X801 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X802 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X803 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X804 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X805 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X806 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X807 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X808 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X809 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X810 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X811 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X812 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X813 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X814 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X815 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X816 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X817 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X818 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X819 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X820 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X821 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X822 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X823 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X824 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X825 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X826 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X827 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X828 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X829 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X830 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X831 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X832 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X833 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X834 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X835 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X836 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X837 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X838 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X839 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X840 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X841 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X842 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X843 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X844 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X845 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X846 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X847 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X848 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X849 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X850 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X851 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X852 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X853 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X854 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X855 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X856 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X857 ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X858 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X859 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X860 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X861 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X862 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X863 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X864 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X865 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X866 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X867 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X868 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X869 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X870 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X871 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X872 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X873 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X874 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X875 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X876 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X877 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X878 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X879 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X880 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X881 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X882 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X883 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X884 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X885 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X886 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X887 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X888 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X889 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X890 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X891 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X892 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X893 ota_0.vout a_29905_n7588# cap_mim_2f0_m4m5_noshield c_width=22u c_length=22u
X894 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X895 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X896 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X897 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X898 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X899 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X900 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X901 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X902 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X903 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X904 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X905 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X906 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X907 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X908 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X909 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X910 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X911 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X912 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X913 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X914 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X915 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X916 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X917 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X918 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X919 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X920 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X921 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X922 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X923 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X924 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X925 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X926 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X927 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X928 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X929 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X930 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X931 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X932 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X933 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X934 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X935 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X936 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X937 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X938 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X939 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X940 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X941 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X942 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X943 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X944 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X945 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X946 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X947 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X948 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X949 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X950 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X951 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X952 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X953 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X954 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X955 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X956 a_29974_13820# a_34102_14420# vss ppolyf_u_1k r_width=1u r_length=20u
X957 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X958 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X959 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X960 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X961 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X962 ota_0.cm_nmos_0.iout vin_p a_30505_n7588# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X963 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X964 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X965 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X966 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X967 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X968 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X969 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X970 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X971 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X972 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X973 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X974 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X975 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X976 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X977 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X978 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X979 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X980 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X981 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X982 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X983 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X984 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X985 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X986 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X987 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X988 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X989 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X990 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X991 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X992 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X993 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X994 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X995 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X996 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X997 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X998 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X999 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1000 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1001 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1002 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1003 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1004 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1005 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1006 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1007 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1008 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1009 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1010 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1011 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1012 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1013 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1014 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1015 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1016 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1017 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1018 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1019 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1020 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1021 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1022 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1023 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1024 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1025 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1026 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1027 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1028 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1029 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1030 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1031 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1032 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1033 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1034 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1035 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1036 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1037 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1038 vdd vdd vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=0 ps=0 w=25u l=1u
X1039 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1040 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1041 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1042 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1043 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1044 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1045 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1046 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1047 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1048 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1049 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1050 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1051 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1052 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1053 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1054 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1055 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1056 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1057 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1058 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1059 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1060 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1061 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1062 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1063 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1064 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1065 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1066 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1067 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1068 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1069 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1070 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1071 a_29905_n6460# a_30505_n7588# vss ppolyf_u_1k r_width=1u r_length=5u
X1072 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1073 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1074 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1075 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1076 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1077 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1078 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1079 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1080 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1081 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1082 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1083 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1084 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1085 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1086 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1087 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1088 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1089 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1090 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1091 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1092 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1093 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1094 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1095 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1096 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1097 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1098 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1099 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1100 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1101 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1102 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1103 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1104 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1105 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1106 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1107 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1108 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1109 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1110 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1111 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1112 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1113 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1114 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1115 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1116 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1117 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1118 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1119 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1120 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1121 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1122 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1123 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1124 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1125 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1126 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1127 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1128 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1129 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1130 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1131 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1132 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1133 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1134 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1135 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1136 vss iref ota_0.cm_nmos_0.iout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1137 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1138 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1139 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1140 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1141 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1142 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1143 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1144 a_29974_7220# feedback vss ppolyf_u_1k r_width=1u r_length=20u
X1145 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1146 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1147 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1148 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1149 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1150 ota_0.vout a_30505_n7588# vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X1151 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1152 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1153 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1154 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1155 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1156 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1157 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1158 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1159 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1160 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1161 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1162 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1163 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1164 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1165 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1166 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1167 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1168 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1169 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1170 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1171 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1172 a_34724_n8101# a_34724_n8101# vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1173 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1174 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1175 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1176 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1177 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1178 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1179 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1180 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1181 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1182 a_29974_11420# a_34102_9620# vss ppolyf_u_1k r_width=1u r_length=20u
X1183 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1184 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1185 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1186 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1187 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1188 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1189 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1190 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1191 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1192 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1193 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1194 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1195 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1196 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1197 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1198 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1199 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1200 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1201 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1202 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1203 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1204 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1205 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1206 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1207 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1208 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1209 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1210 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1211 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1212 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1213 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1214 vdd vdd vdd vdd pfet_03v3 ad=16.25p pd=51.3u as=0 ps=0 w=25u l=1u
X1215 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1216 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1217 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1218 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1219 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1220 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1221 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1222 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1223 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1224 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1225 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1226 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1227 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1228 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1229 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1230 vss iref ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1231 out ota_0.vout vdd vdd pfet_03v3 ad=2.6079p pd=9.38u as=4.814p ps=13.61u w=4.38u l=0.5u
X1232 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1233 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1234 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1235 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1236 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1237 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1238 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1239 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1240 ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1241 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1242 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1243 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1244 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1245 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1246 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1247 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1248 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1249 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1250 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1251 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1252 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1253 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1254 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1255 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1256 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1257 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1258 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1259 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1260 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1261 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1262 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1263 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1264 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1265 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1266 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1267 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1268 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1269 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1270 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1271 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1272 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1273 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1274 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1275 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1276 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1277 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1278 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1279 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1280 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1281 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1282 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1283 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1284 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1285 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1286 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1287 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1288 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1289 ota_0.cm_nmos_0.iout vss vss vss nfet_03v3 ad=1.3p pd=5.52u as=3.05p ps=11.219999u w=5u l=1u
X1290 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1291 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1292 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1293 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1294 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1295 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1296 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1297 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1298 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1299 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1300 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1301 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1302 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1303 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1304 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1305 vss iref ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1306 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1307 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1308 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1309 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1310 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1311 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1312 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1313 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1314 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1315 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1316 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1317 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1318 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1319 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1320 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1321 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1322 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1323 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1324 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1325 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1326 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1327 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1328 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1329 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1330 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1331 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1332 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1333 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1334 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1335 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1336 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1337 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1338 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1339 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1340 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1341 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1342 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1343 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1344 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1345 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1346 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1347 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1348 vss iref iref vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1349 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1350 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1351 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1352 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1353 a_29974_13220# vss vss ppolyf_u_1k r_width=1u r_length=20u
X1354 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1355 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1356 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1357 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1358 vdd ota_0.vout out vdd pfet_03v3 ad=3.2335p pd=9.38u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1359 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1360 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1361 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1362 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1363 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1364 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1365 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1366 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1367 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1368 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1369 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1370 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1371 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1372 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1373 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1374 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1375 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1376 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1377 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1378 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1379 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1380 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1381 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1382 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1383 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1384 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1385 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1386 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1387 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1388 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1389 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1390 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1391 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1392 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1393 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1394 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1395 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1396 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1397 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1398 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1399 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1400 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1401 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1402 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1403 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1404 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1405 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1406 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1407 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1408 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1409 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1410 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1411 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1412 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1413 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1414 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1415 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1416 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1417 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1418 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1419 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1420 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1421 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1422 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1423 a_29974_7220# a_34102_7820# vss ppolyf_u_1k r_width=1u r_length=20u
X1424 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1425 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1426 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1427 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1428 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1429 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1430 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1431 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1432 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1433 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1434 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1435 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1436 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1437 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1438 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1439 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1440 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1441 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1442 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1443 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1444 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1445 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1446 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1447 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1448 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1449 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1450 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1451 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1452 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1453 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1454 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1455 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1456 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1457 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1458 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1459 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1460 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1461 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1462 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1463 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1464 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1465 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1466 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1467 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1468 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1469 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1470 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1471 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1472 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1473 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1474 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1475 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1476 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1477 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1478 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1479 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1480 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1481 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1482 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1483 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1484 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1485 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1486 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1487 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1488 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1489 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1490 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1491 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1492 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1493 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1494 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1495 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1496 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1497 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1498 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1499 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1500 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1501 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1502 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1503 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1504 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1505 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1506 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1507 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1508 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1509 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1510 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1511 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1512 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1513 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1514 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1515 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1516 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1517 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1518 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1519 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1520 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1521 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1522 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1523 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1524 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1525 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1526 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1527 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1528 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1529 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1530 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1531 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1532 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1533 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1534 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1535 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1536 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1537 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1538 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1539 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1540 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1541 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1542 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1543 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1544 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1545 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1546 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1547 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1548 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1549 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1550 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1551 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1552 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1553 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1554 a_29905_n6460# a_29905_n7588# vss ppolyf_u_1k r_width=1u r_length=5u
X1555 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1556 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1557 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1558 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1559 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1560 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1561 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1562 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1563 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1564 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1565 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1566 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1567 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1568 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1569 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1570 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1571 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1572 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1573 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1574 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1575 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1576 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1577 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1578 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1579 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1580 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1581 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1582 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1583 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1584 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1585 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1586 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1587 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1588 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1589 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1590 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1591 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1592 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1593 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1594 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1595 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1596 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1597 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1598 a_29974_11420# a_34102_12020# vss ppolyf_u_1k r_width=1u r_length=20u
X1599 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1600 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1601 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1602 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1603 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1604 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1605 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1606 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1607 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1608 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1609 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1610 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1611 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1612 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1613 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1614 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1615 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1616 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1617 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1618 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1619 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1620 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1621 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1622 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1623 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1624 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1625 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1626 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1627 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1628 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1629 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1630 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1631 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1632 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1633 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1634 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1635 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1636 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1637 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1638 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1639 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1640 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1641 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1642 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1643 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1644 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1645 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1646 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1647 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1648 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1649 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1650 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1651 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1652 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1653 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1654 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1655 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1656 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1657 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1658 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1659 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1660 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1661 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1662 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1663 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1664 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1665 a_29974_15620# a_34102_14420# vss ppolyf_u_1k r_width=1u r_length=20u
X1666 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1667 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1668 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1669 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1670 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1671 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1672 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1673 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1674 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1675 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1676 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1677 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1678 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1679 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1680 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1681 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1682 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1683 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1684 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1685 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1686 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1687 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1688 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1689 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1690 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1691 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1692 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1693 vss vss ota_0.cm_nmos_0.iout vss nfet_03v3 ad=3.075p pd=11.23u as=1.3p ps=5.52u w=5u l=1u
X1694 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1695 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1696 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1697 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1698 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1699 ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1700 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1701 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1702 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1703 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1704 vss iref ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1705 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1706 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1707 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1708 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1709 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1710 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1711 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1712 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1713 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1714 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1715 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1716 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1717 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1718 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1719 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1720 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1721 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1722 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1723 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1724 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1725 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1726 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1727 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1728 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1729 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1730 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1731 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1732 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1733 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1734 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1735 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1736 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1737 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1738 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1739 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1740 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1741 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1742 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1743 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1744 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1745 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1746 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1747 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1748 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1749 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1750 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1751 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1752 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1753 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1754 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1755 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1756 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1757 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1758 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1759 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1760 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1761 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1762 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1763 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1764 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1765 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1766 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1767 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1768 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1769 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1770 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1771 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1772 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1773 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1774 vss vss vss ppolyf_u_1k r_width=1u r_length=5u
X1775 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1776 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1777 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1778 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1779 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1780 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1781 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1782 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1783 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1784 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1785 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1786 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1787 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1788 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1789 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1790 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1791 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1792 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1793 out ota_0.vout vdd vdd pfet_03v3 ad=2.6079p pd=9.38u as=4.814p ps=13.61u w=4.38u l=0.5u
X1794 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1795 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1796 a_30505_n7588# a_34724_n8101# vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1797 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1798 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1799 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1800 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1801 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=2.6079p ps=9.38u w=4.38u l=0.5u
X1802 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1803 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1804 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1805 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1806 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1807 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1808 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1809 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1810 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1811 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1812 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1813 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1814 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1815 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1816 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1817 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1818 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1819 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1820 vss iref ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1821 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1822 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1823 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1824 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1825 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1826 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1827 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1828 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1829 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1830 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1831 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1832 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1833 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1834 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1835 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1836 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1837 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1838 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1839 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1840 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1841 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1842 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1843 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1844 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1845 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1846 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1847 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1848 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1849 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1850 a_29974_8420# feedback vss ppolyf_u_1k r_width=1u r_length=20u
X1851 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1852 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1853 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1854 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1855 a_30505_n7588# vin_p ota_0.cm_nmos_0.iout vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1856 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1857 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1858 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1859 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1860 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1861 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=0 ps=0 w=2.5u l=1u
X1862 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1863 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1864 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1865 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1866 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1867 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1868 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1869 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1870 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1871 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1872 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1873 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1874 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1875 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1876 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1877 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1878 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1879 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1880 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1881 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1882 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1883 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1884 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1885 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1886 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1887 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1888 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1889 a_29974_10820# a_34102_12620# vss ppolyf_u_1k r_width=1u r_length=20u
X1890 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1891 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1892 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1893 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1894 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1895 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1896 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1897 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1898 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1899 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1900 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1901 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1902 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1903 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1904 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1905 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1906 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1907 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1908 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1909 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1910 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1911 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1912 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1913 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1914 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1915 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1916 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1917 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1918 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1919 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1920 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1921 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1922 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1923 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1924 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1925 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1926 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1927 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1928 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1929 vdd a_30505_n7588# ota_0.vout vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X1930 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1931 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1932 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1933 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1934 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1935 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1936 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1937 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1938 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1939 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1940 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1941 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1942 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1943 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1944 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1945 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1946 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1947 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1948 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1949 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1950 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1951 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1952 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1953 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1954 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1955 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1956 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1957 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1958 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1959 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1960 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1961 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1962 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1963 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1964 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1965 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1966 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1967 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1968 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1969 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1970 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1971 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1972 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1973 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1974 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1975 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1976 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1977 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1978 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1979 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1980 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1981 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1982 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1983 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1984 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1985 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1986 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1987 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1988 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1989 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1990 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1991 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1992 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1993 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1994 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1995 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1996 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1997 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1998 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1999 out ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X2000 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2001 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2002 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2003 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2004 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2005 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2006 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2007 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2008 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2009 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2010 vdd ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2011 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2012 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2013 a_34724_n8101# ref ota_0.cm_nmos_0.iout vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X2014 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2015 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2016 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2017 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2018 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2019 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2020 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2021 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2022 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2023 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2024 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2025 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2026 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2027 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2028 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2029 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2030 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2031 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2032 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2033 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2034 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2035 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2036 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2037 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2038 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2039 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2040 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2041 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2042 out ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2043 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2044 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2045 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2046 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2047 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2048 vdd ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
C0 ota_0.vout iref 1.63363f
C1 vdd a_34724_n8101# 3.29537f
C2 feedback m1_35032_7810# 0.10346f
C3 a_29974_13220# a_29974_15620# 0.120932f
C4 ota_0.vout a_29905_n7588# 2.74789f
C5 ota_0.cm_nmos_0.iout a_34724_n8101# 0.250752f
C6 a_34102_12020# a_34102_14420# 0.14109f
C7 ota_0.vout a_30505_n7588# 2.87172f
C8 a_29974_13220# a_29974_10820# 0.14109f
C9 feedback a_34102_7820# 0.592967f
C10 a_29974_10820# a_29974_8420# 0.14109f
C11 vdd ota_0.cm_nmos_0.iout 1.60493f
C12 a_30505_n7588# a_29905_n7588# 0.332743f
C13 out vdd 2.32064p
C14 vin_p a_30505_n7588# 1.11127f
C15 a_29974_10820# a_29974_11420# 0.864964f
C16 a_29974_8420# a_29974_9020# 0.864964f
C17 vdd iref 0.457403f
C18 a_34724_n8101# ref 1.11601f
C19 vdd ota_0.vout 1.76674p
C20 a_29974_13820# a_29974_13220# 0.864964f
C21 vdd ref 0.449627f
C22 ota_0.cm_nmos_0.iout iref 0.340145f
C23 a_34102_9620# a_34102_10220# 0.802011f
C24 vdd a_29905_n7588# 0.270536f
C25 a_30505_n7588# a_34724_n8101# 0.915286f
C26 vin_p a_34724_n8101# 0.41246f
C27 ota_0.cm_nmos_0.iout ref 2.52489f
C28 vdd a_30505_n7588# 9.19771f
C29 out a_34102_14420# 0.120238f
C30 a_34102_9620# a_34102_7820# 0.14109f
C31 out ota_0.vout 1.31651p
C32 ota_0.cm_nmos_0.iout a_30505_n7588# 0.514834f
C33 vin_p ota_0.cm_nmos_0.iout 1.25837f
C34 a_34102_12020# a_34102_9620# 0.14109f
C35 a_34102_12020# a_34102_12620# 0.802011f
C36 a_29974_8420# a_29974_7220# 0.120932f
C37 vin_p vss 9.57911f
C38 ref vss 4.07884f
C39 iref vss 10.2837f
C40 feedback vss 9.031231f
C41 out vss 0.134212p
C42 vdd vss 4.84609p
C43 m1_35032_6610# vss 0.262201f $ **FLOATING
C44 m1_34632_6610# vss 0.31235f $ **FLOATING
C45 m1_29300_6610# vss 0.26928f $ **FLOATING
C46 m1_28900_6610# vss 0.25079f $ **FLOATING
C47 m1_35032_7810# vss 0.195149f $ **FLOATING
C48 m1_35032_9010# vss 0.205536f $ **FLOATING
C49 m1_35032_9610# vss 0.205536f $ **FLOATING
C50 m1_35032_11410# vss 0.205536f $ **FLOATING
C51 m1_28900_8410# vss 0.205536f $ **FLOATING
C52 m1_28900_10210# vss 0.205536f $ **FLOATING
C53 m1_35032_12010# vss 0.205536f $ **FLOATING
C54 m1_35032_13810# vss 0.205536f $ **FLOATING
C55 m1_28900_10810# vss 0.205536f $ **FLOATING
C56 m1_28900_12610# vss 0.205536f $ **FLOATING
C57 m1_35032_14410# vss 0.269682f $ **FLOATING
C58 m1_35032_15610# vss 0.267473f $ **FLOATING
C59 m1_28900_13210# vss 0.205536f $ **FLOATING
C60 m1_28900_15010# vss 0.205536f $ **FLOATING
C61 m1_35032_16810# vss 0.245969f $ **FLOATING
C62 m1_34632_16810# vss 0.289052f $ **FLOATING
C63 m1_29300_16810# vss 0.26928f $ **FLOATING
C64 m1_28900_16810# vss 0.25079f $ **FLOATING
C65 a_29905_n7588# vss 3.67203f
C66 a_29905_n6460# vss 1.30871f
C67 a_30505_n7588# vss 3.7114f
C68 a_34724_n8101# vss 1.53696f
C69 ota_0.cm_nmos_0.iout vss 5.20193f
C70 ota_0.vout vss 0.13008p
C71 a_29974_7220# vss 1.84618f
C72 a_34102_7820# vss 2.16629f
C73 a_29974_9020# vss 1.55313f
C74 a_29974_8420# vss 1.94188f
C75 a_34102_10220# vss 1.80662f
C76 a_34102_9620# vss 2.46883f
C77 a_29974_11420# vss 1.55691f
C78 a_29974_10820# vss 1.92754f
C79 a_34102_12620# vss 1.81178f
C80 a_34102_12020# vss 2.46883f
C81 a_29974_13820# vss 1.55313f
C82 a_29974_13220# vss 1.94188f
C83 a_34102_14420# vss 2.67952f
C84 a_29974_15620# vss 1.84618f
.ends


* NGSPICE file created from resistor.ext - technology: gf180mcuD

.subckt polyf_res_inst_d09b0e8d a_4000_0# a_n376_0# a_n132_0#
X0 a_n132_0# a_4000_0# a_n376_0# ppolyf_u r_width=1u r_length=20u
.ends

.subckt res_dev polyf_res_inst_d09b0e8d_0/a_n132_0# polyf_res_inst_d09b0e8d_0/a_4000_0#
+ VSUBS
Xpolyf_res_inst_d09b0e8d_0 polyf_res_inst_d09b0e8d_0/a_4000_0# VSUBS polyf_res_inst_d09b0e8d_0/a_n132_0#
+ polyf_res_inst_d09b0e8d
.ends

.subckt resistor B IN1 IN2 OUT1 OUT2
Xres_dev_0[0] B B B res_dev
Xres_dev_0[1] OUT1 m1_3956_590# B res_dev
Xres_dev_0[2] m1_n776_1190# m1_3956_590# B res_dev
Xres_dev_0[3] OUT2 m1_3956_1790# B res_dev
Xres_dev_0[4] m1_n776_1190# m1_3956_2390# B res_dev
Xres_dev_0[5] m1_n776_2990# m1_3956_2390# B res_dev
Xres_dev_0[6] m1_n1176_3590# m1_3956_1790# B res_dev
Xres_dev_0[7] m1_n1176_3590# m1_3956_4190# B res_dev
Xres_dev_0[8] m1_n776_2990# m1_3956_4790# B res_dev
Xres_dev_0[9] m1_n776_5390# m1_3956_4790# B res_dev
Xres_dev_0[10] m1_n1176_5990# m1_3956_4190# B res_dev
Xres_dev_0[11] m1_n1176_5990# m1_3956_6590# B res_dev
Xres_dev_0[12] m1_n776_5390# m1_3956_7190# B res_dev
Xres_dev_0[13] m1_n776_7790# m1_3956_7190# B res_dev
Xres_dev_0[14] IN2 m1_3956_6590# B res_dev
Xres_dev_0[15] m1_n776_7790# m1_3956_8990# B res_dev
Xres_dev_0[16] IN1 m1_3956_8990# B res_dev
Xres_dev_0[17] B B B res_dev
.ends


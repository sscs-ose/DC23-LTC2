** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/test/inv_sample/inv_sample-test.sch

.include /home/designer/.volare/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_statistical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice bjt_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical


.control
write
set appendwrite
.endc


**.subckt inv_sample-test
x1 VDD out in GND inv_sample
vvdd VDD GND 3.3
vin in GND pulse(0 3.3 100p 100p 1n 4n 10n)
**** begin user architecture code


.control
save all

tran 0.01n 100n
*plot in out

set curplotname=transient
write
.endc




.control
save all

dc vin 0 3.3 0.01
*plot out vs in in

set curplotname=transfer_curve
write
.endc




.include inv_sample_pex.spice
* inv_sample_pex vdd vss out in
XDUT VDD GND out_pex in inv_sample_pex


**** end user architecture code
**.ends

* expanding   symbol:  /workspaces/DC23-LTC2-LDO/LDO/xschem/test/inv_sample/inv_sample.sym # of
*+ pins=4
** sym_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/test/inv_sample/inv_sample.sym
** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/test/inv_sample/inv_sample.sch
.subckt inv_sample vdd out in vss
*.iopin vdd
*.iopin out
*.iopin vss
*.iopin in
XM1 out in vdd vdd pfet_03v3 L=0.28u W=1.26u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 out in vss vss nfet_03v3 L=0.28u W=0.42u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end

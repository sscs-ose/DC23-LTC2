* Extracted by KLayout with GF180MCU LVS runset on : 30/12/2023 06:00

.SUBCKT cap_mim_2f IN2 IN1
C$1 IN2 IN1 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
.ENDS cap_mim_2f

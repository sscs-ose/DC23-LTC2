* NGSPICE file created from resistor_pex.ext - technology: gf180mcuD

.subckt resistor_pex B IN1 IN2 OUT1 OUT2
X0 OUT2.t0 a_4000_1800.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X1 a_n132_5400.t0 a_4000_4800.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X2 a_n132_7800.t1 a_4000_9000.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X3 a_n132_1200.t1 a_4000_2400.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X4 a_n132_6000.t1 a_4000_4200.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X5 IN1.t0 a_4000_9000.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X6 a_n132_3000.t0 a_4000_2400.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X7 B.t3 B.t4 B.t0 ppolyf_u r_width=1u r_length=20u
X8 a_n132_6000.t0 a_4000_6600.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X9 OUT1.t0 a_4000_600.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X10 a_n132_3600.t0 a_4000_1800.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X11 a_n132_5400.t1 a_4000_7200.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X12 a_n132_3600.t1 a_4000_4200.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X13 a_n132_7800.t0 a_4000_7200.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X14 a_n132_1200.t0 a_4000_600.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X15 a_n132_3000.t1 a_4000_4800.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X16 IN2.t0 a_4000_6600.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X17 B.t1 B.t2 B.t0 ppolyf_u r_width=1u r_length=20u
R0 OUT2 OUT2.t0 11.9413
R1 a_4000_1800.t0 a_4000_1800.t1 26.5088
R2 B.n1 B.t0 675.453
R3 B.n0 B.t1 12.3094
R4 B B.t3 11.4364
R5 B.n0 B.t2 10.4095
R6 B.n2 B.t4 10.4095
R7 B.n1 B.n0 2.3841
R8 B.n2 B.n1 2.37125
R9 B B.n2 0.8735
R10 a_n132_5400.t0 a_n132_5400.t1 26.5082
R11 a_4000_4800.t0 a_4000_4800.t1 26.3444
R12 a_n132_7800.t0 a_n132_7800.t1 26.2628
R13 a_4000_9000.t0 a_4000_9000.t1 26.3451
R14 a_n132_1200.t0 a_n132_1200.t1 26.2628
R15 a_4000_2400.t0 a_4000_2400.t1 26.3451
R16 a_n132_6000.t0 a_n132_6000.t1 26.3446
R17 a_4000_4200.t0 a_4000_4200.t1 26.5088
R18 IN1 IN1.t0 11.949
R19 a_n132_3000.t0 a_n132_3000.t1 26.5082
R20 a_4000_6600.t0 a_4000_6600.t1 26.508
R21 OUT1 OUT1.t0 11.9438
R22 a_4000_600.t0 a_4000_600.t1 26.3444
R23 a_n132_3600.t0 a_n132_3600.t1 26.3446
R24 a_4000_7200.t0 a_4000_7200.t1 26.3451
R25 IN2 IN2.t0 11.9454
C0 m1_4956_5990# m1_4956_6590# 0.048f
C1 m1_4956_4190# m1_4956_3590# 0.048f
C2 m1_n1176_7790# IN2 0.048f
C3 m1_n1176_8990# IN2 0.048f
C4 m1_n1176_n10# OUT1 0.048f
C5 m1_n1176_7190# m1_n1176_7790# 0.048f
C6 m1_n1176_8990# IN1 0.048f
C7 m1_n1176_1190# OUT1 0.048f
C8 m1_n1176_4790# m1_n1176_5390# 0.048f
C9 m1_n1176_10190# m1_n776_10190# 0.097131f
C10 IN1 m1_n776_10190# 0.027147f
C11 m1_n776_n10# m1_n1176_n10# 0.097131f
C12 m1_n1176_1190# OUT2 0.048f
C13 m1_n1176_2390# m1_n1176_2990# 0.048f
C14 m1_4956_n10# m1_4556_n10# 0.097131f
C15 m1_4956_10190# m1_4556_10190# 0.097131f
C16 IN2 IN1 0.008167f
C17 m1_n1176_10190# IN1 0.048f
C18 OUT1 OUT2 0.008167f
C19 m1_n1176_2390# OUT2 0.048f
C20 m1_n776_n10# OUT1 0.027147f
C21 OUT1 B 1.06247f
C22 OUT2 B 0.874969f
C23 IN2 B 0.874969f
C24 IN1 B 1.06247f
C25 m1_4956_n10# B 0.250822f $ **FLOATING
C26 m1_4556_n10# B 0.269428f $ **FLOATING
C27 m1_n776_n10# B 0.290488f $ **FLOATING
C28 m1_n1176_n10# B 0.250822f $ **FLOATING
C29 m1_4956_1790# B 0.205536f $ **FLOATING
C30 m1_4956_3590# B 0.205536f $ **FLOATING
C31 m1_n1176_1190# B 0.205536f $ **FLOATING
C32 m1_n1176_2390# B 0.205536f $ **FLOATING
C33 m1_4956_4190# B 0.205536f $ **FLOATING
C34 m1_4956_5990# B 0.205536f $ **FLOATING
C35 m1_n1176_2990# B 0.205536f $ **FLOATING
C36 m1_n1176_4790# B 0.205536f $ **FLOATING
C37 m1_4956_6590# B 0.205536f $ **FLOATING
C38 m1_4956_8390# B 0.205536f $ **FLOATING
C39 m1_n1176_5390# B 0.205536f $ **FLOATING
C40 m1_n1176_7190# B 0.205536f $ **FLOATING
C41 m1_n1176_7790# B 0.205536f $ **FLOATING
C42 m1_n1176_8990# B 0.205536f $ **FLOATING
C43 m1_4956_10190# B 0.250822f $ **FLOATING
C44 m1_4556_10190# B 0.269428f $ **FLOATING
C45 m1_n776_10190# B 0.290488f $ **FLOATING
C46 m1_n1176_10190# B 0.250822f $ **FLOATING
.ends


** sch_path: /workspaces/DC23-LTC2-LDO/LDO/xschem/ota-ldo/
**.subckt
**.ends
.end

* NGSPICE file created from sar.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VPW nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends 

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 VDD ZN B A1 A2 VSS A3 VNW VPW
X0 a_468_497# A1 ZN VNW pfet_06v0 ad=0.58035p pd=2.155u as=0.4012p ps=1.85u w=1.095u l=0.5u
X1 a_244_69# A2 ZN VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.4137p ps=1.9u w=0.815u l=0.6u
X2 a_780_497# A2 a_468_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.58035p ps=2.155u w=1.095u l=0.5u
X3 ZN A1 a_244_69# VPW nfet_06v0 ad=0.4137p pd=1.9u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4 VDD A3 a_780_497# VNW pfet_06v0 ad=0.5913p pd=3.27u as=0.2847p ps=1.615u w=1.095u l=0.5u
X5 a_244_69# B VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.4012p pd=1.85u as=0.4972p ps=3.14u w=1.13u l=0.5u
X7 ZN A3 a_244_69# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VNW VPW
X0 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VNW VPW
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VPW nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_68# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X5 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6 VSS a_36_68# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD a_36_68# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VPW nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VPW nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VPW nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VPW nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 Z VSS VDD I VNW VPW
X0 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X1 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X3 a_224_552# I VSS VPW nfet_06v0 ad=0.2662p pd=2.09u as=0.2662p ps=2.09u w=0.605u l=0.6u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X8 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.2002p ps=1.79u w=0.455u l=0.6u
X9 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X10 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VNW VPW
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VPW nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VPW nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_455_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 VDD Q CLK VSS D VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2304_115# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X3 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X5 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X6 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X7 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X10 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X12 Q a_2304_115# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X13 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X14 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X15 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X18 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X19 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X20 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X21 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X22 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X23 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VPW nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 Z VSS VDD I VNW VPW
X0 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3 a_224_552# I VDD VNW pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X4 VDD I a_224_552# VNW pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X7 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X10 VSS a_224_552# Z VPW nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X11 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X12 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X13 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X15 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X16 VDD I a_224_552# VNW pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X17 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X18 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X19 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X20 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X21 a_224_552# I VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X22 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 B C VDD VSS ZN A1 A2 VNW VPW
X0 a_692_68# B a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X3 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4016p ps=1.94u w=0.985u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4016p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.44325p pd=2.87u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS C a_692_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 VDD VSS Z I VNW VPW
X0 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X11 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X12 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X13 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X15 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X16 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X17 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X18 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X19 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X20 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X21 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X22 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X23 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X24 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X25 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X26 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X27 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X28 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X29 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X30 a_224_552# I VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X31 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X32 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X33 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X34 VSS a_224_552# Z VPW nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X35 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X36 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X37 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X38 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X39 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X40 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X41 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X42 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X43 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X44 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X45 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D VDD VSS CLK Q VNW VPW
X0 VSS a_2304_115# Q VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2 Q a_2304_115# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X4 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X8 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 VDD a_2304_115# Q VNW pfet_06v0 ad=0.854p pd=3.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X12 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 Q a_2304_115# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X15 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X16 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X17 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X18 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X19 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X21 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X22 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X23 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X24 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X25 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A3 A4 VDD VSS Z A1 A2 VNW VPW
X0 VSS A4 a_56_604# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1 Z a_56_604# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.218p ps=1.52u w=0.82u l=0.6u
X2 Z a_56_604# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.389p ps=2.02u w=1.22u l=0.5u
X3 VSS A2 a_56_604# VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X4 VDD A4 a_708_604# VNW pfet_06v0 ad=0.389p pd=2.02u as=0.1736p ps=1.18u w=0.56u l=0.5u
X5 a_244_604# A1 a_56_604# VNW pfet_06v0 ad=0.196p pd=1.26u as=0.2464p ps=2u w=0.56u l=0.5u
X6 a_56_604# A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7 a_56_604# A3 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X8 a_708_604# A3 a_484_604# VNW pfet_06v0 ad=0.1736p pd=1.18u as=0.1736p ps=1.18u w=0.56u l=0.5u
X9 a_484_604# A2 a_244_604# VNW pfet_06v0 ad=0.1736p pd=1.18u as=0.196p ps=1.26u w=0.56u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A2 a_448_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 VSS A1 ZN VPW nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2 VSS A3 ZN VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3 a_244_472# A4 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 a_448_472# A3 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6 ZN A4 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7 ZN A1 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VNW VPW
X0 VSS B a_36_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VNW VPW
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.4488p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VPW nfet_06v0 ad=0.151p pd=1.185u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VPW nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 Z a_36_160# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.151p ps=1.185u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D Q VDD VSS CLK VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VDD a_2011_527# a_2304_115# VNW pfet_06v0 ad=0.38575p pd=1.92u as=0.2457p ps=1.465u w=0.945u l=0.5u
X2 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VSS a_2304_115# Q VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.2333p ps=1.555u w=0.815u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X8 Q a_2304_115# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.38575p ps=1.92u w=1.22u l=0.5u
X9 VSS a_2304_115# Q VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X10 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X11 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X12 VDD a_2304_115# Q VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X13 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X14 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X15 Q a_2304_115# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X16 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X17 Q a_2304_115# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X18 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X19 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.2333p pd=1.555u as=43.199997f ps=0.6u w=0.36u l=0.6u
X20 Q a_2304_115# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.2608p ps=1.455u w=0.815u l=0.6u
X21 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X25 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X26 VDD a_2304_115# Q VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X27 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X28 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X29 VSS a_2011_527# a_2304_115# VPW nfet_06v0 ad=0.2608p pd=1.455u as=0.2119p ps=1.335u w=0.815u l=0.6u
X30 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.2619p pd=1.685u as=50.399998f ps=0.64u w=0.36u l=0.5u
X31 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.2457p pd=1.465u as=0.2619p ps=1.685u w=0.945u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VNW VPW
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VNW VPW
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VPW nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VNW VPW
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2 ZN A3 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X11 ZN A2 a_36_68# VPW nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X13 a_36_68# B VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VPW nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VPW nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 Z I VDD VSS VNW VPW
X0 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7 VSS a_224_472# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VNW VPW
X0 ZN A1 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VNW VPW
X0 ZN B1 a_257_69# VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A3 A4 VDD VSS Z A1 A2 VNW VPW
X0 VSS a_244_72# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 Z a_244_72# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.23375p ps=1.52u w=0.82u l=0.6u
X2 a_458_472# A3 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X3 VDD a_244_72# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS A4 a_244_72# VPW nfet_06v0 ad=0.23375p pd=1.52u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 Z a_244_72# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 VSS A2 a_244_72# VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 VDD A4 a_1578_472# VNW pfet_06v0 ad=0.5185p pd=2.07u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 a_244_472# A4 VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X9 a_244_72# A1 a_682_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4087p ps=1.89u w=1.22u l=0.5u
X10 VSS A1 a_244_72# VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_1578_472# A3 a_1364_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X12 VDD a_244_72# Z VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3477p ps=1.79u w=1.22u l=0.5u
X13 VSS A3 a_244_72# VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X14 a_1120_472# A1 a_244_72# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_244_72# A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X16 a_1364_472# A2 a_1120_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X17 Z a_244_72# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X18 a_682_472# A2 a_458_472# VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3782p ps=1.84u w=1.22u l=0.5u
X19 a_244_72# A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 a_244_72# A4 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 Z a_244_72# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5185p ps=2.07u w=1.22u l=0.5u
X22 VSS a_244_72# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X23 a_244_72# A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VNW VPW
X0 VSS A2 a_1133_69# VPW nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3 a_741_69# A2 VSS VPW nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X9 VSS B ZN VPW nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VPW nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VPW nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 VDD VSS Z A1 A2 VNW VPW
X0 VSS a_730_497# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 a_954_497# A1 a_730_497# VNW pfet_06v0 ad=0.5256p pd=2.055u as=0.33945p ps=1.715u w=1.095u l=0.5u
X2 a_286_93# A2 a_78_93# VPW nfet_06v0 ad=57.599995f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3 Z a_730_497# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_730_497# a_78_93# VDD VNW pfet_06v0 ad=0.33945p pd=1.715u as=0.344375p ps=1.895u w=1.095u l=0.5u
X5 Z a_730_497# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6 a_78_93# A2 VDD VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X7 a_730_497# A1 a_730_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VDD A1 a_78_93# VNW pfet_06v0 ad=0.344375p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X9 VDD a_730_497# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X10 VSS A1 a_286_93# VPW nfet_06v0 ad=0.218p pd=1.52u as=57.599995f ps=0.68u w=0.36u l=0.6u
X11 a_730_68# A2 a_730_497# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X12 a_730_68# a_78_93# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X13 VDD A2 a_954_497# VNW pfet_06v0 ad=0.4818p pd=3.07u as=0.5256p ps=2.055u w=1.095u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A4 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X1 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4 a_275_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_673_68# A2 a_469_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X6 a_469_68# A3 a_275_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X7 ZN A1 a_673_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
.ends

.subckt sar_logic VDD VSS clk comp current_state[0] current_state[1] dbot[0] dbot[10] dbot[11]
+ dbot[1] dbot[2] dbot[3] dbot[4] dbot[5] dbot[6] dbot[7] dbot[8] dbot[9] dtop[0]
+ dtop[10] dtop[11] dtop[1] dtop[2] dtop[3] dtop[4] dtop[5] dtop[6] dtop[7] dtop[8]
+ dtop[9] rst
XFILLER_0_18_18 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_131_ _093_ VDD VSS _096_ _076_ _088_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_200_ VDD _020_ _065_ current_bit\[3\] _036_ VSS _064_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_9_16 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_114_ VDD VSS net1 _080_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_95 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_72 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_150 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_84 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 dtop[1] VSS VDD net20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput7 VSS dbot[11] net7 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_131 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_142 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_130_ _093_ VDD VSS _095_ _076_ _088_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_113_ VDD VSS net35 _079_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_107 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput10 VSS dbot[3] net10 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput21 VSS dtop[2] net21 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput8 VSS dbot[1] net8 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_189_ VDD VSS _015_ _094_ _059_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_149 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_112_ VDD VSS current_bit\[1\] _078_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_16_31 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 VSS dtop[3] net22 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput11 dbot[4] VSS VDD net11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput9 VSS dbot[2] net9 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_122 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_188_ VDD VSS _014_ _036_ _059_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_18_150 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_111_ VSS _077_ current_bit\[0\] VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_1_64 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput12 VSS dbot[5] net12 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput23 VSS dtop[4] net23 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_187_ _059_ VDD VSS _013_ _086_ _030_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_110_ VDD VSS net4 _076_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_239_ VDD net10 clknet_2_2_0_clk VSS _019_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput24 VSS dtop[5] net24 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput13 VSS dbot[6] net13 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_186_ VDD VSS _012_ current_bit\[0\] _059_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_68 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_169_ _087_ VDD VSS _047_ current_bit\[3\] _079_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_238_ VDD net9 clknet_2_0_0_clk VSS _018_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_100 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput14 VSS dbot[7] net14 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput25 VSS dtop[6] net25 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_185_ VDD VSS _059_ net3 _076_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_168_ _046_ VDD VSS _007_ net31 _045_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_237_ VDD net8 clknet_2_2_0_clk VSS _017_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_104 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput26 VSS dtop[7] net26 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput15 dbot[8] VSS VDD net15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xclkbuf_2_3_0_clk clknet_2_3_0_clk VSS VDD clknet_1_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_184_ _058_ net30 VDD VSS _011_ _083_ _056_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_236_ VDD net5 clknet_2_0_0_clk VSS _016_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_167_ VDD _046_ net26 net33 _030_ VSS _035_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_21_36 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_135 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_138 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_219_ VDD VSS _029_ _085_ net32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput16 VSS dbot[9] net16 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput27 VSS dtop[8] net27 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_0_clk VDD VSS clknet_0_clk clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_2_2_0_clk clknet_2_2_0_clk VSS VDD clknet_1_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_183_ net29 VDD VSS _058_ net36 _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_235_ _015_ VDD VSS clknet_2_1_0_clk current_bit\[3\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_166_ _030_ _035_ VDD VSS _045_ net1 net33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_149_ VDD _032_ net22 current_bit\[2\] net33 VSS _030_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_218_ net2 _088_ VDD VSS _028_ net3 net4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xoutput17 VSS dtop[0] net17 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput28 dtop[9] VSS VDD net28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_11_150 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout30 net30 VSS VDD net32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_182_ net29 VDD VSS _057_ net36 _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_1_26 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_234_ VDD current_bit\[2\] clknet_2_1_0_clk VSS _014_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_165_ _030_ _035_ VDD VSS _044_ net37 net33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
Xclkbuf_2_1_0_clk clknet_2_1_0_clk VSS VDD clknet_1_0_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_148_ VDD VSS _031_ current_bit\[2\] _030_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_12_118 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_217_ VDD net30 _075_ _027_ _057_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput18 VSS dtop[10] net18 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_20_140 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout31 net31 VSS VDD net32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_181_ VDD VSS _056_ _031_ net29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_164_ _043_ net32 VDD VSS _006_ net1 _042_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_233_ _013_ current_bit\[1\] VDD VSS clknet_2_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_21_119 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_147_ VDD VSS _030_ current_bit\[0\] current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_216_ net7 VDD VSS _075_ _031_ _049_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput19 VSS dtop[11] net19 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_2_0_0_clk clknet_2_0_0_clk VSS VDD clknet_1_0_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_180_ _055_ net30 VDD VSS _010_ _082_ _053_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xfanout32 VSS net32 _102_ VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_232_ _012_ current_bit\[0\] VDD VSS clknet_2_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_163_ VDD _043_ net25 net33 _105_ VSS _035_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_146_ _109_ VDD VSS _002_ net30 _107_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_215_ VDD net32 _074_ _026_ _054_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_72 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_129_ VDD VSS _094_ _088_ _093_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_150 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout33 VSS net33 _096_ VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_18 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_162_ _036_ VDD VSS _042_ net34 _104_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_231_ VDD net19 clknet_2_2_0_clk VSS _011_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_18 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput1 net1 VSS VDD comp VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_145_ _106_ VDD VSS _109_ net37 net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_214_ net6 VDD VSS _074_ _106_ net29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_126 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_128_ current_bit\[1\] net35 current_bit\[3\] VDD VSS _093_ current_bit\[0\] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
Xfanout34 VSS net34 _095_ VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_230_ VDD net18 clknet_2_0_0_clk VSS _010_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_161_ _041_ net31 VDD VSS _005_ net1 _040_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_94 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_31 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput2 VSS net2 rst VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_144_ _106_ VDD VSS _108_ net36 net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_213_ VDD net30 _073_ _025_ _051_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_127_ VDD _090_ _092_ _000_ _091_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_8 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout35 net35 current_bit\[2\] VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_1_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_160_ VDD _041_ net24 net33 _098_ VSS _035_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_11_65 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_143_ VDD _107_ net21 net35 net33 VSS _105_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_212_ net16 VDD VSS _073_ _099_ _049_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_126_ VDD VSS _092_ _076_ net17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout36 VSS net36 _080_ VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_142_ net35 VDD VSS _106_ current_bit\[0\] _078_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_211_ _072_ net32 VDD VSS _024_ net35 _064_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_125_ VDD VSS _091_ net3 net4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_110 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout37 net37 VSS VDD _080_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_125 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_141_ VDD VSS _105_ _077_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_210_ VDD VSS _072_ net15 _047_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_124_ _088_ _089_ net17 VDD VSS _090_ net36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_17_66 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_114 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_31 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_148 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_140_ VDD VSS _104_ current_bit\[0\] _078_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_150 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_123_ VDD VSS _089_ net4 _088_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_1_1_0_clk clknet_1_1_0_clk VSS VDD clknet_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_199_ net11 _037_ VDD VSS _065_ net3 _076_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_45 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_122_ current_bit\[3\] net35 VDD VSS _088_ current_bit\[0\] current_bit\[1\] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_0_138 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout29 net29 VSS VDD _049_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_198_ _088_ VDD VSS _064_ net1 _087_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_121_ current_bit\[1\] VDD VSS _087_ net4 current_bit\[0\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_3_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_128 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_1_0_0_clk clknet_1_0_0_clk VSS VDD clknet_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_37 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_80 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_107 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_197_ VDD net31 _063_ _019_ _033_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_120_ VDD VSS _086_ current_bit\[0\] current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_17_26 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_249_ _029_ VDD VSS clknet_2_0_0_clk net4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_19_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_57 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_80 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_121 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_37 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_196_ net10 VDD VSS _063_ _095_ _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_179_ net29 VDD VSS _055_ net36 _106_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_248_ _028_ VDD VSS clknet_2_0_0_clk net3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_195_ VDD net30 _062_ _018_ _108_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_247_ VDD net7 clknet_2_2_0_clk VSS _027_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_178_ net29 VDD VSS _054_ net36 _106_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_194_ net9 VDD VSS _062_ net34 _106_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_18 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_246_ VDD net6 clknet_2_0_0_clk VSS _026_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_177_ VDD VSS _053_ _106_ net29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_229_ VDD net28 clknet_2_2_0_clk VSS _009_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_149 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_193_ VDD net30 _061_ _017_ _100_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_245_ VDD net16 clknet_2_2_0_clk VSS _025_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_176_ _052_ net30 VDD VSS _009_ _081_ _050_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_159_ _036_ VDD VSS _040_ net34 _097_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_228_ VDD net27 clknet_2_1_0_clk VSS _008_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_96 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_192_ net8 VDD VSS _061_ net34 _099_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_101 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_244_ VDD net15 clknet_2_1_0_clk VSS _024_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_175_ net29 VDD VSS _052_ net36 _099_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_227_ VDD net26 clknet_2_3_0_clk VSS _007_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_158_ VDD _004_ _039_ current_bit\[3\] _036_ VSS _038_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_191_ net32 _060_ VDD VSS _016_ _084_ _089_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_243_ VDD net14 clknet_2_3_0_clk VSS _023_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_174_ net29 VDD VSS _051_ net36 _099_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_226_ VDD net25 clknet_2_1_0_clk VSS _006_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_157_ net23 _037_ VDD VSS _039_ net3 _076_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_209_ _071_ VDD VSS _023_ net31 _044_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ VDD VSS _060_ net1 _089_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_242_ VDD net13 clknet_2_1_0_clk VSS _022_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_173_ VDD VSS _050_ _099_ net29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_225_ VDD net24 clknet_2_3_0_clk VSS _005_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_156_ _088_ VDD VSS _038_ net37 _087_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_54 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_208_ VDD _071_ net14 _096_ _030_ VSS _035_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_139_ _103_ VDD VSS _001_ _101_ net30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_98 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_123 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_241_ VDD net12 clknet_2_3_0_clk VSS _021_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_172_ net4 VDD VSS _049_ _088_ _093_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_155_ _079_ _086_ VDD VSS _037_ net4 current_bit\[3\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_224_ VDD net23 clknet_2_0_0_clk VSS _004_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_207_ _070_ VDD VSS _022_ net32 _069_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_20_45 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_138_ VDD _103_ net20 net35 net33 VSS _098_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_20_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_171_ _048_ net32 VDD VSS _008_ net35 _038_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_240_ VDD net11 clknet_2_0_0_clk VSS _020_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_223_ VDD net22 clknet_2_3_0_clk VSS _003_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_154_ VDD VSS _036_ _079_ _086_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_206_ VDD _070_ net13 net33 _105_ VSS _035_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_137_ VDD VSS _102_ net3 _076_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_170_ VDD VSS _048_ net27 _047_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_153_ VDD VSS _035_ net35 _086_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_222_ VDD net21 clknet_2_1_0_clk VSS _002_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_205_ _036_ _066_ VDD VSS _069_ _094_ _104_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_136_ _099_ VDD VSS _101_ net36 net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_9_66 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_119_ VDD VSS net2 _085_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_107 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_152_ _034_ VDD VSS _003_ net30 _032_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_221_ VDD net20 clknet_2_3_0_clk VSS _001_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_204_ _068_ VDD VSS _021_ net31 _067_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_36 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_37 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_135_ _099_ VDD VSS _100_ net36 net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_118_ VDD VSS net5 _084_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput3 VSS current_state[0] net3 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_3_36 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_26 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_151_ _031_ VDD VSS _034_ net37 net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_220_ VDD net17 clknet_2_0_0_clk VSS _000_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_203_ VDD _068_ net12 net33 _098_ VSS _035_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_134_ net35 VDD VSS _099_ _077_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_9_35 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_117_ VDD VSS net19 _083_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_81 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput4 VSS current_state[1] net4 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_150 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_150_ _031_ VDD VSS _033_ net37 net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_0_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_202_ _036_ _066_ VDD VSS _067_ _094_ _097_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_133_ VDD VSS _098_ current_bit\[0\] _078_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_116_ VDD VSS net18 _082_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput5 VSS dbot[0] net5 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_132_ VDD VSS _097_ _077_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_201_ VDD VSS _066_ net4 net37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_115_ VDD VSS net28 _081_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_16 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 VSS dbot[10] net6 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
.ends


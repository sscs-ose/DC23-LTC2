* NGSPICE file created from sar.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 VDD Q CLK VSS D VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2304_115# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X3 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X5 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X6 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X7 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X10 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X12 Q a_2304_115# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X13 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X14 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X15 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X18 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X19 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X20 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X21 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X22 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X23 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A3 a_36_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 VSS A4 a_244_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5 a_1468_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 a_1866_68# A2 a_1662_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A4 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X10 a_3276_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X11 a_652_68# A4 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 a_36_68# A3 a_652_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X13 VDD A2 ZN VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 VSS A4 a_1060_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X16 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X17 a_2372_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X18 a_36_68# A2 a_2372_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X19 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X20 a_1060_68# A3 a_36_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X21 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X22 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X23 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X24 ZN A1 a_2780_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.1312p ps=1.14u w=0.82u l=0.6u
X25 a_2780_68# A2 a_36_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X26 ZN A4 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X27 VDD A1 ZN VNW pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X28 a_36_68# A2 a_3276_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X29 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X30 a_1662_68# A3 a_1468_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X31 ZN A1 a_1866_68# VPW nfet_06v0 ad=0.4161p pd=1.905u as=0.1517p ps=1.19u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_68# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X5 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6 VSS a_36_68# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD a_36_68# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VPW nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VNW VPW
X0 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VNW VPW
X0 VSS B a_36_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 Z VSS VDD I VNW VPW
X0 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X1 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X3 a_224_552# I VSS VPW nfet_06v0 ad=0.2662p pd=2.09u as=0.2662p ps=2.09u w=0.605u l=0.6u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X8 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.2002p ps=1.79u w=0.455u l=0.6u
X9 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X10 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 B C VDD VSS ZN A1 A2 VNW VPW
X0 a_692_68# B a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X3 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4016p ps=1.94u w=0.985u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4016p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.44325p pd=2.87u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS C a_692_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VPW nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VPW nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VPW nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VPW nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 Z VSS VDD I VNW VPW
X0 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3 a_224_552# I VDD VNW pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X4 VDD I a_224_552# VNW pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X7 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X10 VSS a_224_552# Z VPW nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X11 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X12 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X13 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X15 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X16 VDD I a_224_552# VNW pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X17 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X18 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X19 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X20 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X21 a_224_552# I VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X22 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 VDD VSS Z I VNW VPW
X0 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X11 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X12 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X13 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X15 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X16 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X17 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X18 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X19 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X20 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X21 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X22 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X23 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X24 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X25 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X26 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X27 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X28 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X29 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X30 a_224_552# I VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X31 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X32 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X33 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X34 VSS a_224_552# Z VPW nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X35 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X36 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X37 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X38 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X39 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X40 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X41 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X42 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X43 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X44 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X45 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VNW VPW
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VPW nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D Q VDD VSS CLK VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 VDD a_2011_527# a_2304_115# VNW pfet_06v0 ad=0.38575p pd=1.92u as=0.2457p ps=1.465u w=0.945u l=0.5u
X2 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3 VSS a_2304_115# Q VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.2333p ps=1.555u w=0.815u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X8 Q a_2304_115# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.38575p ps=1.92u w=1.22u l=0.5u
X9 VSS a_2304_115# Q VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X10 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X11 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X12 VDD a_2304_115# Q VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X13 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X14 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X15 Q a_2304_115# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X16 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X17 Q a_2304_115# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X18 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X19 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.2333p pd=1.555u as=43.199997f ps=0.6u w=0.36u l=0.6u
X20 Q a_2304_115# VSS VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.2608p ps=1.455u w=0.815u l=0.6u
X21 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X23 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X24 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X25 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X26 VDD a_2304_115# Q VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X27 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X28 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X29 VSS a_2011_527# a_2304_115# VPW nfet_06v0 ad=0.2608p pd=1.455u as=0.2119p ps=1.335u w=0.815u l=0.6u
X30 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.2619p pd=1.685u as=50.399998f ps=0.64u w=0.36u l=0.5u
X31 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.2457p pd=1.465u as=0.2619p ps=1.685u w=0.945u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VPW nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 Z I VDD VSS VNW VPW
X0 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7 VSS a_224_472# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 a_224_604# A1 a_36_88# VNW pfet_06v0 ad=0.1736p pd=1.18u as=0.2464p ps=2u w=0.56u l=0.5u
X1 a_36_88# A2 VSS VPW nfet_06v0 ad=0.14p pd=1.1u as=0.104p ps=0.92u w=0.4u l=0.6u
X2 Z a_36_88# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.389p ps=2.02u w=1.22u l=0.5u
X3 VSS A1 a_36_88# VPW nfet_06v0 ad=0.104p pd=0.92u as=0.176p ps=1.68u w=0.4u l=0.6u
X4 a_448_604# A2 a_224_604# VNW pfet_06v0 ad=0.224p pd=1.36u as=0.1736p ps=1.18u w=0.56u l=0.5u
X5 VSS A3 a_36_88# VPW nfet_06v0 ad=0.224p pd=1.52u as=0.14p ps=1.1u w=0.4u l=0.6u
X6 VDD A3 a_448_604# VNW pfet_06v0 ad=0.389p pd=2.02u as=0.224p ps=1.36u w=0.56u l=0.5u
X7 Z a_36_88# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.224p ps=1.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VNW VPW
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VPW nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VPW nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VNW VPW
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VPW nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 VDD ZN I VSS VNW VPW
X0 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2 VDD I ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 ZN I VSS VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
X4 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VSS I ZN VPW nfet_06v0 ad=0.1248p pd=1u as=0.1248p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VPW nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VPW nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 VSS ZN I VDD VNW VPW
X0 ZN I VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 ZN I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 VSS I ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 ZN I VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6 VSS I ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD I ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 a_1458_68# A3 a_1254_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 VDD VSS ZN I VNW VPW
X0 ZN I VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 VSS I ZN VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
X2 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.1248p ps=1u w=0.48u l=0.6u
X5 ZN I VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6 VDD I ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X7 VSS I ZN VPW nfet_06v0 ad=0.1248p pd=1u as=0.1248p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VNW VPW
X0 ZN B1 a_257_69# VPW nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 a_257_69# B2 VSS VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VPW nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_728_472# a_56_604# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X1 Z A1 a_728_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2 VSS A1 a_56_604# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3 a_728_472# A2 Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 Z a_56_604# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X5 VSS A2 a_952_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 a_244_604# A2 a_56_604# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X7 a_56_604# A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 a_952_68# A1 Z VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 VDD A1 a_244_604# VNW pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VNW VPW
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2 Z a_36_159# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VPW nfet_06v0 ad=0.23405p pd=1.555u as=58.399994f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VPW nfet_06v0 ad=58.399994f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_455_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A4 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X1 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4 a_275_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_673_68# A2 a_469_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X6 a_469_68# A3 a_275_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X7 ZN A1 a_673_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt sar EOC VDD VSS clk comp current_state dbot[0] dbot[10] dbot[11] dbot[1] dbot[2]
+ dbot[3] dbot[4] dbot[5] dbot[6] dbot[7] dbot[8] dbot[9] dtop[0] dtop[10] dtop[11]
+ dtop[1] dtop[2] dtop[3] dtop[4] dtop[5] dtop[6] dtop[7] dtop[8] dtop[9] rst
X_200_ VDD net24 clknet_2_0_0_clk VSS _021_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_131_ _062_ current_bit\[2\] VDD VSS _031_ _060_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_19_114 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_114_ VDD VSS _079_ current_bit\[2\] _064_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput7 VSS dbot[11] net7 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput20 VSS dtop[1] net20 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_130_ VDD VSS _009_ net3 _030_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_61 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_113_ VDD net30 _078_ _004_ _077_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput8 dbot[1] VSS VDD net8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput10 dbot[3] VSS VDD net10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput21 VSS dtop[2] net21 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_189_ VDD net13 clknet_2_0_0_clk VSS _010_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_138 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_112_ VDD VSS _078_ net5 _071_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput11 VSS dbot[4] net11 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput9 VSS dbot[2] net9 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput22 VSS dtop[3] net22 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_188_ VDD net12 clknet_2_0_0_clk VSS _009_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_111_ VDD VSS _077_ net33 _072_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_97 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_53 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput23 VSS dtop[4] net23 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput12 dbot[5] VSS VDD net12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_187_ VDD net11 clknet_2_1_0_clk VSS _008_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_110_ VDD VSS _076_ current_bit\[2\] net33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput24 VSS dtop[5] net24 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput13 VSS dbot[6] net13 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_18_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_186_ VDD net10 clknet_2_3_0_clk VSS _007_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_44 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_169_ _055_ net29 VDD VSS _023_ net33 _033_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xoutput14 VSS dbot[7] net14 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput25 dtop[6] VSS VDD net25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_185_ VDD net9 clknet_2_2_0_clk VSS _006_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_168_ VDD VSS _055_ net26 _033_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_099_ _067_ VDD VSS _001_ net29 _066_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_19_89 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput26 VSS dtop[7] net26 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput15 VSS dbot[8] net15 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_2_3_0_clk clknet_2_3_0_clk VSS VDD clknet_1_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_10_37 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_184_ VDD net8 clknet_2_2_0_clk VSS _005_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_167_ _054_ net29 VDD VSS _022_ net33 _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_098_ VDD VSS _067_ net32 _061_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput27 VSS dtop[8] net27 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_0_clk VDD VSS clknet_0_clk clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput16 dbot[9] VSS VDD net16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_16_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_2_2_0_clk clknet_2_2_0_clk VSS VDD clknet_1_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_166_ VDD VSS _054_ net25 _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_183_ VDD net5 clknet_2_1_0_clk VSS _004_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_097_ VDD VSS _066_ _060_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_36 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput17 VSS dtop[0] net17 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_149_ _076_ VDD VSS _044_ _060_ _061_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xoutput28 VSS dtop[9] net28 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xfanout30 VSS net30 net31 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_182_ _003_ current_bit\[3\] VDD VSS clknet_2_3_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_165_ _053_ net29 VDD VSS _021_ net33 _029_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_096_ VDD VSS _000_ net32 net3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_2_1_0_clk clknet_2_1_0_clk VSS VDD clknet_1_0_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_12_107 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_148_ _084_ VDD VSS _043_ current_bit\[3\] _063_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_18_112 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput18 VSS dtop[10] net18 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_095_ VDD VSS net23 _065_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_164_ VDD VSS _053_ net24 _029_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout31 VSS net31 net4 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_181_ _002_ current_bit\[2\] VDD VSS clknet_2_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_19_16 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput19 dtop[11] VSS VDD net19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_11_72 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_147_ _042_ net29 VDD VSS _014_ _064_ _040_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_2_0_0_clk clknet_2_0_0_clk VSS VDD clknet_1_0_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout32 net32 current_bit\[0\] VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_180_ _001_ current_bit\[1\] VDD VSS clknet_2_2_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_094_ VDD VSS net33 _064_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_163_ _052_ VDD VSS _020_ net3 _088_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_129_ _029_ VDD VSS _030_ net33 net12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_146_ VDD VSS _042_ net6 _040_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout33 net33 VSS VDD net1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_162_ _065_ VDD VSS _052_ current_bit\[2\] _075_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_093_ VDD _063_ current_bit\[2\] VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_1_18 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput1 VSS net1 comp VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_145_ _076_ VDD VSS _041_ current_bit\[0\] _061_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_0_132 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_128_ _062_ current_bit\[2\] VDD VSS _029_ net32 _061_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_092_ VSS _062_ current_bit\[3\] VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
Xinput2 VSS net2 rst VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_161_ VDD VSS _019_ net31 _051_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_127_ VDD net29 _088_ _008_ _087_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_144_ current_bit\[3\] _063_ VDD VSS _040_ _060_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_5_40 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_75 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_091_ VDD VSS _061_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_160_ _044_ _074_ VDD VSS _051_ net22 _085_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_143_ _039_ net30 VDD VSS _013_ _064_ _037_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_126_ _075_ VDD VSS _088_ current_bit\[2\] _064_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_109_ current_bit\[3\] VDD VSS _075_ net32 current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_090_ VDD VSS net29 net3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_125_ net11 VDD VSS _087_ current_bit\[2\] _075_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_142_ VDD VSS _039_ net16 _037_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_108_ VDD VSS _003_ net30 _074_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_141_ _076_ VDD VSS _038_ _060_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_124_ _086_ net30 VDD VSS _007_ _064_ _085_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_107_ VDD VSS _074_ _062_ _068_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_140_ current_bit\[3\] _063_ VDD VSS _037_ net32 _061_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_106_ VDD VSS _073_ current_bit\[3\] _068_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_123_ VDD VSS _086_ net10 _085_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_199_ VDD net23 clknet_2_1_0_clk VSS _020_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_122_ _084_ VDD VSS _085_ _062_ _063_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xclkbuf_1_1_0_clk clknet_1_1_0_clk VSS VDD clknet_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_105_ VDD VSS _072_ _062_ _068_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout29 net29 VSS VDD net31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_198_ VDD net22 clknet_2_3_0_clk VSS _019_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_114 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_104_ VDD VSS _071_ _062_ _068_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_1_0_0_clk clknet_1_0_0_clk VSS VDD clknet_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_121_ VDD VSS _084_ net32 current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_18_90 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_123 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_120_ _083_ VDD VSS _006_ net29 _082_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_197_ VDD net21 clknet_2_2_0_clk VSS _018_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_103_ VDD VSS _070_ _062_ _063_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_196_ VDD net20 clknet_2_2_0_clk VSS _017_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_179_ VDD current_bit\[0\] clknet_2_1_0_clk VSS _000_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_102_ _069_ VDD VSS _002_ net3 _068_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_195_ VDD net17 clknet_2_1_0_clk VSS _016_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_178_ net2 VDD VSS _028_ net30 _071_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_101_ _063_ VDD VSS _069_ _060_ _061_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_82 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_194_ VDD net7 clknet_2_3_0_clk VSS _015_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_100_ current_bit\[2\] VDD VSS _068_ net32 current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_177_ VDD VSS _027_ net31 _059_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_193_ VDD net6 clknet_2_3_0_clk VSS _014_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_176_ _044_ current_bit\[3\] VDD VSS _059_ net19 _043_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_159_ _050_ VDD VSS _018_ net31 _049_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_192_ VDD net16 clknet_2_3_0_clk VSS _013_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_31 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_97 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_175_ VDD VSS _026_ net31 _058_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_158_ VDD net21 _070_ _050_ _066_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_089_ VDD _060_ net32 VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_191_ VDD net15 clknet_2_1_0_clk VSS _012_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_121 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_157_ VDD VSS _049_ _074_ _041_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_174_ _041_ current_bit\[3\] VDD VSS _058_ net18 _040_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_10 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_190_ VDD net14 clknet_2_0_0_clk VSS _011_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_173_ VDD VSS _025_ net31 _057_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_31 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_156_ _048_ VDD VSS _017_ net29 _047_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_139_ VDD net30 _036_ _012_ _035_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_155_ VDD net20 _070_ _048_ _067_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_172_ _038_ current_bit\[3\] VDD VSS _057_ net28 _037_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_138_ net15 VDD VSS _036_ current_bit\[3\] _068_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_207_ VDD net4 clknet_2_1_0_clk VSS _028_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_171_ _056_ net30 VDD VSS _024_ net1 _073_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_154_ VDD VSS _047_ _074_ _038_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_137_ VDD VSS _035_ net33 _073_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_206_ VDD net19 clknet_2_3_0_clk VSS _027_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_130 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_170_ VDD VSS _056_ net27 _073_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_136_ VDD VSS _011_ net3 _034_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_153_ _046_ net30 VDD VSS _016_ net1 _072_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_205_ VDD net18 clknet_2_2_0_clk VSS _026_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_119_ VDD net9 _070_ _083_ _066_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_152_ VDD VSS _046_ net17 _072_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_36 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_135_ _033_ VDD VSS _034_ net33 net14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_34 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_118_ _062_ _079_ VDD VSS _082_ _060_ current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_204_ VDD net28 clknet_2_3_0_clk VSS _025_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput3 VSS EOC net3 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_203_ VDD net27 clknet_2_1_0_clk VSS _024_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_134_ _062_ current_bit\[2\] VDD VSS _033_ net32 current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_151_ _045_ net30 VDD VSS _015_ _064_ _043_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_16_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_117_ _081_ VDD VSS _005_ net29 _080_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput4 current_state VSS VDD net30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_5_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_150_ VDD VSS _045_ net7 _043_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_16 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_202_ VDD net26 clknet_2_0_0_clk VSS _023_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_133_ VDD VSS _010_ net3 _032_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_70 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_116_ VDD net8 _070_ _081_ _067_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput5 dbot[0] VSS VDD net5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_201_ VDD net25 clknet_2_0_0_clk VSS _022_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_132_ _031_ VDD VSS _032_ net33 net13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_115_ _062_ _079_ VDD VSS _080_ net32 _061_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_6_16 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 VSS dbot[10] net6 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
.ends


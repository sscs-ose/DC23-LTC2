* Extracted by KLayout with GF180MCU LVS runset on : 05/01/2024 21:32

.SUBCKT cs-vth-ref
X$1 \$1 \$6 \$1 \$6 \$1 \$6 \$1 \$6 \$1 \$6 \$6 \$6 \$6 \$6 \$6 \$6 \$6 \$17
+ \$1 pfet$1
X$2 \$1 \$7 \$1 \$7 \$1 \$7 \$1 \$7 \$1 \$6 \$6 \$6 \$6 \$6 \$6 \$6 \$6 \$18
+ \$1 pfet$1
X$3 \$1 \$I858 \$I879 vdd backgate_n
X$4 \$1 \$I847 \$I868 vdd backgate_n
X$5 \$1 m1_source
X$6 \$1 \$I848 \$18 vdd backgate_n
X$7 \$1 \$I848 \$18 vdd backgate_n
X$8 \$1 m1_source
X$9 \$1 \$I848 \$18 vdd backgate_n
X$10 \$1 \$I848 \$18 vdd backgate_n
X$11 \$1 m1_source
X$12 \$1 \$I848 \$18 vdd backgate_n
X$13 \$1 \$I848 \$18 vdd backgate_n
X$14 \$1 m1_source
X$15 \$1 \$I848 \$18 vdd backgate_n
X$16 \$1 \$I848 \$18 vdd backgate_n
X$17 \$1 m1_source
X$18 \$1 \$I848 \$18 vdd backgate_n
X$19 \$1 \$I848 \$18 vdd backgate_n
X$20 \$12 \$12 \$6 \$7 \$7 \$1 \$12 \$14 \$14 \$51 \$15 nfet
X$21 vss vss \$7 \$12 \$12 \$1 vss \$15 \$15 \$52 \$54 nfet
X$22 \$1 m1_source
X$23 \$1 \$I838 \$17 vdd backgate_n
X$24 \$1 \$I838 \$17 vdd backgate_n
X$25 \$1 m1_source
X$26 \$1 \$I838 \$17 vdd backgate_n
X$27 \$1 \$I838 \$17 vdd backgate_n
X$28 \$1 m1_source
X$29 \$1 \$I838 \$17 vdd backgate_n
X$30 \$1 \$I838 \$17 vdd backgate_n
X$31 \$1 m1_source
X$32 \$1 \$I838 \$17 vdd backgate_n
X$33 \$1 \$I838 \$17 vdd backgate_n
X$34 \$1 m1_source
X$35 \$1 \$I838 \$17 vdd backgate_n
X$36 \$1 \$I838 \$17 vdd backgate_n
X$37 vss \$1 vdd pg_mesh
X$38 vss \$1 vdd pg_mesh
X$39 vss \$1 vdd pg_mesh
X$40 vss \$1 vdd pg_mesh
X$41 vss \$1 vdd pg_mesh
X$42 vss \$1 vdd pg_mesh
X$43 vss \$1 vdd pg_mesh
X$44 vss \$1 vdd pg_mesh
X$45 vss \$1 vdd pg_mesh
X$46 vss \$1 vdd pg_mesh
X$47 vss \$1 vdd pg_mesh
X$48 vss \$1 vdd pg_mesh
X$49 vss \$1 vdd pg_mesh
X$50 vss \$1 vdd pg_mesh
X$51 vss \$1 vdd pg_mesh
X$52 vss \$1 vdd pg_mesh
X$53 vss \$1 vdd pg_mesh
X$54 vss \$1 vdd pg_mesh
X$55 vss \$1 vdd pg_mesh
X$56 vss \$1 vdd pg_mesh
X$57 vss \$1 vdd pg_mesh
X$58 vss \$1 vdd pg_mesh
X$59 vss \$1 vdd pg_mesh
X$60 vss \$1 vdd pg_mesh
X$61 vss \$1 vdd pg_mesh
X$62 vss \$1 vdd pg_mesh
X$63 vss \$1 vdd pg_mesh
X$64 vss \$1 vdd pg_mesh
X$65 vss \$1 vdd pg_mesh
X$66 vss \$1 vdd pg_mesh
X$67 vss \$1 vdd pg_mesh
X$68 vss \$1 vdd pg_mesh
X$69 vss \$1 vdd pg_mesh
X$70 vss \$1 vdd pg_mesh
X$71 vss \$1 vdd pg_mesh
X$72 vss \$1 vdd pg_mesh
X$73 vss \$1 vdd pg_mesh
X$74 vss \$1 vdd pg_mesh
X$75 vss \$1 vdd pg_mesh
X$76 vss \$1 vdd pg_mesh
X$77 vss \$1 vdd pg_mesh
X$78 vss \$1 vdd pg_mesh
X$79 vss \$1 vdd pg_mesh
X$80 vss \$1 vdd pg_mesh
X$81 vss \$1 vdd pg_mesh
X$82 vss \$1 vdd pg_mesh
X$83 vss \$1 vdd pg_mesh
X$84 vss \$1 vdd pg_mesh
X$85 vss \$1 vdd pg_mesh
X$86 vss \$1 vdd pg_mesh
X$87 vss \$1 vdd pg_mesh
X$88 vss \$1 vdd pg_mesh
X$89 vss \$1 vdd pg_mesh
X$90 vss \$1 vdd pg_mesh
X$91 vss \$1 vdd pg_mesh
X$92 vss \$1 vdd pg_mesh
X$93 vss \$1 vdd pg_mesh
X$94 vss \$1 vdd pg_mesh
X$95 vss \$1 vdd pg_mesh
X$96 vss \$1 vdd pg_mesh
X$97 vss \$1 vdd pg_mesh
X$98 vss \$1 vdd pg_mesh
X$99 vss \$1 vdd pg_mesh
X$100 vss \$1 vdd pg_mesh
X$101 vss \$1 vdd pg_mesh
X$102 vss \$1 vdd pg_mesh
X$103 vss \$1 vdd pg_mesh
X$104 vss \$1 vdd pg_mesh
X$105 vss \$1 vdd pg_mesh
X$106 vss \$1 vdd pg_mesh
X$107 vss \$1 vdd pg_mesh
X$108 vss \$1 vdd pg_mesh
X$109 vss \$1 vdd pg_mesh
X$110 vss \$1 vdd pg_mesh
X$111 vss \$1 vdd pg_mesh
X$112 vss \$1 vdd pg_mesh
X$113 vss \$1 vdd pg_mesh
X$114 vss \$1 vdd pg_mesh
X$115 vss \$1 vdd pg_mesh
X$116 vss \$1 vdd pg_mesh
X$117 vss \$1 vdd pg_mesh
X$118 vss \$1 vdd pg_mesh
X$119 vss \$1 vdd pg_mesh
X$120 vss \$1 vdd pg_mesh
X$121 vss \$1 vdd pg_mesh
X$122 vss \$1 vdd pg_mesh
X$123 vss \$1 vdd pg_mesh
X$124 vss \$1 vdd pg_mesh
X$125 vss \$1 vdd pg_mesh
X$126 vss \$1 vdd pg_mesh
X$127 vss \$1 vdd pg_mesh
X$128 vss \$1 vdd pg_mesh
X$129 vss \$1 vdd pg_mesh
X$130 vss \$1 vdd pg_mesh
X$131 vss \$1 vdd pg_mesh
X$132 vss \$1 vdd pg_mesh
X$133 vss \$1 vdd pg_mesh
X$134 vss \$1 vdd pg_mesh
X$135 vss \$1 vdd pg_mesh
X$136 vss \$1 vdd pg_mesh
X$137 vss \$1 vdd pg_mesh
X$138 vss \$1 vdd pg_mesh
X$139 vss \$1 vdd pg_mesh
X$140 vss \$1 vdd pg_mesh
X$141 vss \$1 vdd pg_mesh
X$142 vss \$1 vdd pg_mesh
X$143 vss \$1 vdd pg_mesh
X$144 vss \$1 vdd pg_mesh
X$145 vss \$1 vdd pg_mesh
X$146 vss \$1 vdd pg_mesh
X$147 vss \$1 vdd pg_mesh
X$148 vss \$1 vdd pg_mesh
X$149 vss \$1 vdd pg_mesh
X$150 vss \$1 vdd pg_mesh
X$151 vss \$1 vdd pg_mesh
X$152 vss \$1 vdd pg_mesh
X$153 vss \$1 vdd pg_mesh
X$154 vss \$1 vdd pg_mesh
X$155 vss \$1 vdd pg_mesh
X$156 vss \$1 vdd pg_mesh
X$157 vss \$1 vdd pg_mesh
X$158 vss \$1 vdd pg_mesh
X$159 vss \$1 vdd pg_mesh
X$160 vss \$1 vdd pg_mesh
X$161 vss \$1 vdd pg_mesh
X$162 vss \$1 vdd pg_mesh
X$163 vss \$1 vdd pg_mesh
X$164 vss \$1 vdd pg_mesh
X$165 vss \$1 vdd pg_mesh
X$166 vss \$1 vdd pg_mesh
X$167 vss \$1 vdd pg_mesh
X$168 vss \$1 vdd pg_mesh
X$169 vss \$1 vdd pg_mesh
X$170 vss \$1 vdd pg_mesh
X$171 vss \$1 vdd pg_mesh
X$172 vss \$1 vdd pg_mesh
X$173 vss \$1 vdd pg_mesh
X$174 vss \$1 vdd pg_mesh
X$175 vss \$1 vdd pg_mesh
X$176 vss \$1 vdd pg_mesh
X$177 vss \$1 vdd pg_mesh
X$178 vss \$1 vdd pg_mesh
X$179 vss \$1 vdd pg_mesh
X$180 vss \$1 vdd pg_mesh
X$181 vss \$1 vdd pg_mesh
X$182 vss \$1 vdd pg_mesh
X$183 vss \$1 vdd pg_mesh
X$184 vss \$1 vdd pg_mesh
X$185 vss \$1 vdd pg_mesh
X$186 vss \$1 vdd pg_mesh
X$187 vss \$1 vdd pg_mesh
X$188 vss \$1 vdd pg_mesh
X$189 vss \$1 vdd pg_mesh
X$190 vss \$1 vdd pg_mesh
X$191 vss \$1 vdd pg_mesh
X$192 vss \$1 vdd pg_mesh
X$193 vss \$1 vdd pg_mesh
X$194 vss \$1 vdd pg_mesh
X$195 vss \$1 vdd pg_mesh
X$196 vss \$1 vdd pg_mesh
X$197 vss \$1 vdd pg_mesh
X$198 vss \$1 vdd pg_mesh
X$199 vss \$1 vdd pg_mesh
X$200 vss \$1 vdd pg_mesh
X$201 vss \$1 vdd pg_mesh
X$202 vss \$1 vdd pg_mesh
X$203 vss \$1 vdd pg_mesh
X$204 vss \$1 vdd pg_mesh
X$205 vss \$1 vdd pg_mesh
X$206 vss \$1 vdd pg_mesh
X$207 vss \$1 vdd pg_mesh
X$208 vss \$1 vdd pg_mesh
X$209 vss \$1 vdd pg_mesh
X$210 vss \$1 vdd pg_mesh
X$211 vss \$1 vdd pg_mesh
X$212 vss \$1 vdd pg_mesh
X$213 vss \$1 vdd pg_mesh
X$214 vss \$1 vdd pg_mesh
X$215 vss \$1 vdd pg_mesh
X$216 vss \$1 vdd pg_mesh
X$217 \$6 vb m12_sd
X$218 \$6 vb m12_sd
X$219 \$6 vb m12_sd
X$220 \$6 vb m12_sd
X$221 \$6 vb m12_sd
X$222 \$6 vb m12_sd
X$223 \$7 \$57 m12_sd
X$224 \$7 \$57 m12_sd
X$225 \$7 \$57 m12_sd
X$226 \$7 \$57 m12_sd
X$227 \$7 \$57 m12_sd
X$228 \$7 \$57 m12_sd
X$229 vss \$I769 tap_psub
X$230 vss \$I769 tap_psub
X$231 vss \$I769 tap_psub
X$232 vss \$I769 tap_psub
X$233 vss \$I769 tap_psub
X$234 vss \$I769 tap_psub
X$235 vss \$I769 tap_psub
X$236 vss \$I769 tap_psub
X$237 vss \$I769 tap_psub
X$238 vss \$I769 tap_psub
X$239 vss \$I769 tap_psub
X$240 vss \$I769 tap_psub
X$241 vss \$I769 tap_psub
X$242 vss \$I769 tap_psub
X$243 vss \$I769 tap_psub
X$244 vss \$I769 tap_psub
X$245 vss \$I769 tap_psub
X$246 vss \$I769 tap_psub
X$247 vss \$I769 tap_psub
X$248 vss \$I769 tap_psub
X$249 vss \$I769 tap_psub
X$250 vss \$I769 tap_psub
X$251 vss \$I769 tap_psub
X$252 vss \$I769 tap_psub
X$253 vss \$I769 tap_psub
X$254 vss \$I769 tap_psub
X$255 vss \$I769 tap_psub
X$256 vss \$I769 tap_psub
X$257 vss \$I769 tap_psub
X$258 vss \$I769 tap_psub
X$259 vss \$I769 tap_psub
X$260 vss \$I769 tap_psub
X$261 vss \$I769 tap_psub
X$262 vss \$I769 tap_psub
X$263 vss \$I769 tap_psub
X$264 vss \$I769 tap_psub
X$265 vss \$I769 tap_psub
X$266 vss \$I769 tap_psub
X$267 vss \$I769 tap_psub
X$268 vss \$I769 tap_psub
X$269 vss \$I769 tap_psub
X$270 vss \$I769 tap_psub
X$271 vss \$I769 tap_psub
X$272 vss \$I769 tap_psub
X$273 vss \$I769 tap_psub
X$274 vss \$I769 tap_psub
X$275 vss \$I769 tap_psub
X$276 vss \$I769 tap_psub
X$277 vss \$I769 tap_psub
X$278 vss \$I769 tap_psub
X$279 vss \$I769 tap_psub
X$280 vss \$I769 tap_psub
X$281 vss \$I769 tap_psub
X$282 vss \$I769 tap_psub
X$283 vss \$I769 tap_psub
X$284 vss \$I769 tap_psub
X$285 vss \$I769 tap_psub
X$286 vss \$I769 tap_psub
X$287 vss \$I769 tap_psub
X$288 vss \$I769 tap_psub
X$289 vss \$I769 tap_psub
X$290 vss \$I769 tap_psub
X$291 vss \$I769 tap_psub
X$292 vss \$I769 tap_psub
X$293 vss \$I769 tap_psub
X$294 vss \$I769 tap_psub
X$295 vss \$I769 tap_psub
X$296 vss \$I769 tap_psub
X$297 vss \$I769 tap_psub
X$298 vss \$I769 tap_psub
X$299 vss \$I769 tap_psub
X$300 vss \$I769 tap_psub
X$301 vss \$I769 tap_psub
X$302 vss \$I769 tap_psub
X$303 vss \$I769 tap_psub
X$304 vss \$I769 tap_psub
X$305 vss \$I769 tap_psub
X$306 vss \$I769 tap_psub
X$307 vss \$I769 tap_psub
X$308 vss \$I769 tap_psub
X$309 vss \$I769 tap_psub
X$310 vss \$I769 tap_psub
X$311 vss \$I769 tap_psub
X$312 vss \$I769 tap_psub
X$313 vss \$I769 tap_psub
X$314 vss \$I769 tap_psub
X$315 vss \$I769 tap_psub
X$316 vss \$I769 tap_psub
X$317 vss \$I769 tap_psub
X$318 vss \$I769 tap_psub
X$319 vss \$I769 tap_psub
X$320 vss \$I769 tap_psub
X$321 vss \$I769 tap_psub
X$322 vss \$I769 tap_psub
X$323 vss \$I769 tap_psub
X$324 vss \$I769 tap_psub
X$325 vss \$I769 tap_psub
X$326 vss \$I769 tap_psub
X$327 vss \$I769 tap_psub
X$328 vss \$I828 \$I833 backgate_p
X$329 vss \$I828 \$I833 backgate_p
X$330 vss \$I828 \$I833 backgate_p
X$331 vss m1_source
X$332 vss m1_source
X$333 vss \$36 vss \$I24 GND ppolyf_u_resistor$1
X$334 vss \$I24 ptap
X$335 vss \$I23 ptap
X$336 vss \$I22 ptap
X$337 vss \$I21 ptap
X$338 vss \$I20 ptap
X$339 vss \$35 \$12 \$I16 GND ppolyf_u_resistor$1
X$340 vss \$I16 ptap
X$341 vss \$35 \$37 \$I15 GND ppolyf_u_resistor$1
X$342 vss \$I15 ptap
X$343 vss \$36 \$37 \$I14 GND ppolyf_u_resistor$1
X$344 vss \$I14 ptap
X$345 \$12 \$I830 \$16 backgate_p
X$346 \$12 m1_source
X$347 \$12 \$I830 \$16 backgate_p
X$348 \$12 \$I830 \$16 backgate_p
X$349 \$12 m1_source
X$350 \$12 via1
X$351 \$12 via1
.ENDS cs-vth-ref

.SUBCKT m12_sd \$1 \$2
X$1 \$1 via1
X$2 \$1 via1
X$3 \$1 via1
X$4 \$1 via1
X$5 \$1 via1
.ENDS m12_sd

.SUBCKT m1_source \$1
.ENDS m1_source

.SUBCKT backgate_n \$1 \$2 \$3 \$5
X$1 \$1 via1
.ENDS backgate_n

.SUBCKT tap_psub \$1 \$2
.ENDS tap_psub

.SUBCKT pfet$1 \$2 \$3 \$4 \$5 \$6 \$7 \$8 \$9 \$10 \$11 \$12 \$13 \$14 \$15
+ \$16 \$17 \$18 \$19 \$20
M$1 \$3 \$11 \$2 \$20 pfet_03v3 L=0.56U W=5.6U AS=3.64P AD=1.456P PS=12.5U
+ PD=6.12U
M$2 \$4 \$12 \$3 \$20 pfet_03v3 L=0.56U W=5.6U AS=1.456P AD=1.456P PS=6.12U
+ PD=6.12U
M$3 \$5 \$13 \$4 \$20 pfet_03v3 L=0.56U W=5.6U AS=1.456P AD=1.456P PS=6.12U
+ PD=6.12U
M$4 \$6 \$14 \$5 \$20 pfet_03v3 L=0.56U W=5.6U AS=1.456P AD=1.456P PS=6.12U
+ PD=6.12U
M$5 \$7 \$15 \$6 \$20 pfet_03v3 L=0.56U W=5.6U AS=1.456P AD=1.456P PS=6.12U
+ PD=6.12U
M$6 \$8 \$16 \$7 \$20 pfet_03v3 L=0.56U W=5.6U AS=1.456P AD=1.456P PS=6.12U
+ PD=6.12U
M$7 \$9 \$17 \$8 \$20 pfet_03v3 L=0.56U W=5.6U AS=1.456P AD=1.456P PS=6.12U
+ PD=6.12U
M$8 \$10 \$18 \$9 \$20 pfet_03v3 L=0.56U W=5.6U AS=1.456P AD=3.64P PS=6.12U
+ PD=12.5U
.ENDS pfet$1

.SUBCKT ptap \$1 \$2
.ENDS ptap

.SUBCKT backgate_p \$1 \$2 \$5
X$1 \$1 cnt
X$2 \$1 cnt
X$3 \$1 via1
.ENDS backgate_p

.SUBCKT nfet \$2 \$3 \$4 \$5 \$6 \$7 \$8 \$9 \$10 \$11 \$13
M$1 \$4 \$5 \$2 \$8 nfet_03v3_dn L=0.56U W=5.6U AS=3.416P AD=1.456P PS=12.42U
+ PD=6.12U
M$2 \$3 \$6 \$4 \$8 nfet_03v3_dn L=0.56U W=5.6U AS=1.456P AD=3.416P PS=6.12U
+ PD=12.42U
.ENDS nfet

.SUBCKT pg_mesh \$1 \$2 \$3
.ENDS pg_mesh

.SUBCKT ppolyf_u_resistor$1 \$1 \$2 \$3 \$4 GND
R$1 \$2 \$3 GND 9625 ppolyf_u L=22U W=0.8U
.ENDS ppolyf_u_resistor$1

.SUBCKT via1 \$1
.ENDS via1

.SUBCKT cnt \$1
.ENDS cnt

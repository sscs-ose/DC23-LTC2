.subckt DELETE_padring_side_top
+ tail_DVDD tail_VDD tail_DVSS tail_VSS
+ head_DVDD head_VDD head_DVSS head_VSS

X_cor_0  tail_DVDD  tail_DVSS tail_VDD  tail_VSS  gf180mcu_fd_io__cor

X_fill10_3   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_4   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_5   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_6   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_7   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_8   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_9   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_40  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_41  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_30  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_31  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_20  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_42  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_10  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_43  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_32  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_21  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_11  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_33  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_22  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_12  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_34  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_23  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_13  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_35  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_24  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_14  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_36  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_25  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_15  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_37  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_26  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_16  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_38  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_27  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_0   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_17  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_39  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_28  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_1   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_18  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_29  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_2   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10
X_fill10_19  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill10

X_fill5_11   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_22   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_33   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_44   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_55   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_99   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_88   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_77   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_66   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_289  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_278  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_267  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_256  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_245  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_234  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_223  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_212  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_201  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_12   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_23   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_34   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_45   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_56   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_89   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_78   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_67   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_279  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_268  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_257  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_246  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_235  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_224  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_213  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_202  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_13   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_24   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_35   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_46   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_57   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_79   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_68   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_269  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_258  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_247  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_236  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_225  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_214  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_203  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_14   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_25   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_36   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_47   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_69   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_58   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_259  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_248  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_237  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_226  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_215  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_204  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_15   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_26   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_37   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_48   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_59   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_238  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_227  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_216  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_205  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_249  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_16   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_27   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_38   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_49   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_239  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_228  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_217  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_206  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_17   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_28   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_39   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_229  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_218  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_207  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_18   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_29   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_219  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_208  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_0    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_19   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_209  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_1    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_2    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_190  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_3    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_350  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_191  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_180  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_4    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_351  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_340  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_192  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_181  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_170  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_5    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_341  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_330  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_193  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_182  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_171  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_160  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_6    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_331  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_320  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_342  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_150  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_194  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_183  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_172  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_161  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_7    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_343  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_332  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_321  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_310  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_151  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_140  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_195  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_184  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_173  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_162  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_8    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_344  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_333  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_322  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_311  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_300  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_152  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_130  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_141  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_196  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_185  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_174  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_163  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_9    tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_345  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_334  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_323  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_312  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_301  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_153  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_120  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_131  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_142  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_197  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_186  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_175  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_164  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_346  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_335  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_324  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_313  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_302  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_154  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_121  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_132  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_143  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_110  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_198  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_187  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_176  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_165  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_347  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_336  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_325  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_314  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_303  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_144  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_155  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_122  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_133  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_111  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_100  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_199  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_188  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_177  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_166  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_348  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_337  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_326  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_315  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_304  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_145  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_156  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_123  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_134  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_112  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_101  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_189  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_178  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_167  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_349  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_338  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_327  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_316  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_305  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_113  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_102  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_146  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_124  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_135  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_179  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_168  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_157  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_339  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_328  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_317  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_306  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_147  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_125  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_136  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_114  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_103  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_169  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_158  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_329  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_318  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_307  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_148  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_126  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_137  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_115  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_104  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_159  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_319  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_308  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_149  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_127  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_138  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_116  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_105  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_309  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_128  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_139  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_117  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_106  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_118  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_107  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_129  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_290  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_119  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_108  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_90   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_291  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_280  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_109  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_91   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_80   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_292  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_281  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_270  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_92   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_81   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_70   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_293  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_282  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_271  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_260  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_60   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_93   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_82   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_71   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_294  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_283  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_272  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_261  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_250  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_50   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_94   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_83   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_72   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_61   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_295  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_284  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_273  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_262  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_251  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_240  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_40   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_51   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_95   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_84   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_73   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_62   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_296  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_285  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_274  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_263  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_252  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_241  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_230  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_30   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_41   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_52   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_96   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_85   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_74   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_63   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_297  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_286  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_275  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_264  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_253  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_242  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_231  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_220  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_20   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_31   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_42   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_53   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_97   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_86   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_75   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_64   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_298  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_287  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_276  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_265  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_254  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_243  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_232  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_221  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_210  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_10   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_21   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_32   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_43   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_54   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_76   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_65   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_98   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_87   tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_222  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_211  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_200  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_299  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_288  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_277  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_266  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_255  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_244  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5
X_fill5_233  tail_DVDD  tail_DVSS  tail_VDD  tail_VSS  gf180mcu_fd_io__fill5

.ends
magic
tech sky130A
timestamp 1699286806
<< nwell >>
rect -1125 -1175 14375 14325
<< pwell >>
rect -5925 14325 19175 19125
rect -5925 -1175 -1125 14325
rect 14375 -1175 19175 14325
rect -5925 -5975 19175 -1175
<< mvpmos >>
rect 0 13231 50 13669
rect 550 13231 600 13669
rect 1100 13231 1150 13669
rect 1650 13231 1700 13669
rect 2200 13231 2250 13669
rect 2750 13231 2800 13669
rect 3300 13231 3350 13669
rect 3850 13231 3900 13669
rect 4400 13231 4450 13669
rect 4950 13231 5000 13669
rect 5500 13231 5550 13669
rect 6050 13231 6100 13669
rect 6600 13231 6650 13669
rect 7150 13231 7200 13669
rect 7700 13231 7750 13669
rect 8250 13231 8300 13669
rect 8800 13231 8850 13669
rect 9350 13231 9400 13669
rect 9900 13231 9950 13669
rect 10450 13231 10500 13669
rect 11000 13231 11050 13669
rect 11550 13231 11600 13669
rect 12100 13231 12150 13669
rect 12650 13231 12700 13669
rect 13200 13231 13250 13669
rect -469 13150 -31 13200
rect 81 13150 519 13200
rect 631 13150 1069 13200
rect 1181 13150 1619 13200
rect 1731 13150 2169 13200
rect 2281 13150 2719 13200
rect 2831 13150 3269 13200
rect 3381 13150 3819 13200
rect 3931 13150 4369 13200
rect 4481 13150 4919 13200
rect 5031 13150 5469 13200
rect 5581 13150 6019 13200
rect 6131 13150 6569 13200
rect 6681 13150 7119 13200
rect 7231 13150 7669 13200
rect 7781 13150 8219 13200
rect 8331 13150 8769 13200
rect 8881 13150 9319 13200
rect 9431 13150 9869 13200
rect 9981 13150 10419 13200
rect 10531 13150 10969 13200
rect 11081 13150 11519 13200
rect 11631 13150 12069 13200
rect 12181 13150 12619 13200
rect 12731 13150 13169 13200
rect 13281 13150 13719 13200
rect 0 12681 50 13119
rect 550 12681 600 13119
rect 1100 12681 1150 13119
rect 1650 12681 1700 13119
rect 2200 12681 2250 13119
rect 2750 12681 2800 13119
rect 3300 12681 3350 13119
rect 3850 12681 3900 13119
rect 4400 12681 4450 13119
rect 4950 12681 5000 13119
rect 5500 12681 5550 13119
rect 6050 12681 6100 13119
rect 6600 12681 6650 13119
rect 7150 12681 7200 13119
rect 7700 12681 7750 13119
rect 8250 12681 8300 13119
rect 8800 12681 8850 13119
rect 9350 12681 9400 13119
rect 9900 12681 9950 13119
rect 10450 12681 10500 13119
rect 11000 12681 11050 13119
rect 11550 12681 11600 13119
rect 12100 12681 12150 13119
rect 12650 12681 12700 13119
rect 13200 12681 13250 13119
rect -469 12600 -31 12650
rect 81 12600 519 12650
rect 631 12600 1069 12650
rect 1181 12600 1619 12650
rect 1731 12600 2169 12650
rect 2281 12600 2719 12650
rect 2831 12600 3269 12650
rect 3381 12600 3819 12650
rect 3931 12600 4369 12650
rect 4481 12600 4919 12650
rect 5031 12600 5469 12650
rect 5581 12600 6019 12650
rect 6131 12600 6569 12650
rect 6681 12600 7119 12650
rect 7231 12600 7669 12650
rect 7781 12600 8219 12650
rect 8331 12600 8769 12650
rect 8881 12600 9319 12650
rect 9431 12600 9869 12650
rect 9981 12600 10419 12650
rect 10531 12600 10969 12650
rect 11081 12600 11519 12650
rect 11631 12600 12069 12650
rect 12181 12600 12619 12650
rect 12731 12600 13169 12650
rect 13281 12600 13719 12650
rect 0 12131 50 12569
rect 550 12131 600 12569
rect 1100 12131 1150 12569
rect 1650 12131 1700 12569
rect 2200 12131 2250 12569
rect 2750 12131 2800 12569
rect 3300 12131 3350 12569
rect 3850 12131 3900 12569
rect 4400 12131 4450 12569
rect 4950 12131 5000 12569
rect 5500 12131 5550 12569
rect 6050 12131 6100 12569
rect 6600 12131 6650 12569
rect 7150 12131 7200 12569
rect 7700 12131 7750 12569
rect 8250 12131 8300 12569
rect 8800 12131 8850 12569
rect 9350 12131 9400 12569
rect 9900 12131 9950 12569
rect 10450 12131 10500 12569
rect 11000 12131 11050 12569
rect 11550 12131 11600 12569
rect 12100 12131 12150 12569
rect 12650 12131 12700 12569
rect 13200 12131 13250 12569
rect -469 12050 -31 12100
rect 81 12050 519 12100
rect 631 12050 1069 12100
rect 1181 12050 1619 12100
rect 1731 12050 2169 12100
rect 2281 12050 2719 12100
rect 2831 12050 3269 12100
rect 3381 12050 3819 12100
rect 3931 12050 4369 12100
rect 4481 12050 4919 12100
rect 5031 12050 5469 12100
rect 5581 12050 6019 12100
rect 6131 12050 6569 12100
rect 6681 12050 7119 12100
rect 7231 12050 7669 12100
rect 7781 12050 8219 12100
rect 8331 12050 8769 12100
rect 8881 12050 9319 12100
rect 9431 12050 9869 12100
rect 9981 12050 10419 12100
rect 10531 12050 10969 12100
rect 11081 12050 11519 12100
rect 11631 12050 12069 12100
rect 12181 12050 12619 12100
rect 12731 12050 13169 12100
rect 13281 12050 13719 12100
rect 0 11581 50 12019
rect 550 11581 600 12019
rect 1100 11581 1150 12019
rect 1650 11581 1700 12019
rect 2200 11581 2250 12019
rect 2750 11581 2800 12019
rect 3300 11581 3350 12019
rect 3850 11581 3900 12019
rect 4400 11581 4450 12019
rect 4950 11581 5000 12019
rect 5500 11581 5550 12019
rect 6050 11581 6100 12019
rect 6600 11581 6650 12019
rect 7150 11581 7200 12019
rect 7700 11581 7750 12019
rect 8250 11581 8300 12019
rect 8800 11581 8850 12019
rect 9350 11581 9400 12019
rect 9900 11581 9950 12019
rect 10450 11581 10500 12019
rect 11000 11581 11050 12019
rect 11550 11581 11600 12019
rect 12100 11581 12150 12019
rect 12650 11581 12700 12019
rect 13200 11581 13250 12019
rect -469 11500 -31 11550
rect 81 11500 519 11550
rect 631 11500 1069 11550
rect 1181 11500 1619 11550
rect 1731 11500 2169 11550
rect 2281 11500 2719 11550
rect 2831 11500 3269 11550
rect 3381 11500 3819 11550
rect 3931 11500 4369 11550
rect 4481 11500 4919 11550
rect 5031 11500 5469 11550
rect 5581 11500 6019 11550
rect 6131 11500 6569 11550
rect 6681 11500 7119 11550
rect 7231 11500 7669 11550
rect 7781 11500 8219 11550
rect 8331 11500 8769 11550
rect 8881 11500 9319 11550
rect 9431 11500 9869 11550
rect 9981 11500 10419 11550
rect 10531 11500 10969 11550
rect 11081 11500 11519 11550
rect 11631 11500 12069 11550
rect 12181 11500 12619 11550
rect 12731 11500 13169 11550
rect 13281 11500 13719 11550
rect 0 11031 50 11469
rect 550 11031 600 11469
rect 1100 11031 1150 11469
rect 1650 11031 1700 11469
rect 2200 11031 2250 11469
rect 2750 11031 2800 11469
rect 3300 11031 3350 11469
rect 3850 11031 3900 11469
rect 4400 11031 4450 11469
rect 4950 11031 5000 11469
rect 5500 11031 5550 11469
rect 6050 11031 6100 11469
rect 6600 11031 6650 11469
rect 7150 11031 7200 11469
rect 7700 11031 7750 11469
rect 8250 11031 8300 11469
rect 8800 11031 8850 11469
rect 9350 11031 9400 11469
rect 9900 11031 9950 11469
rect 10450 11031 10500 11469
rect 11000 11031 11050 11469
rect 11550 11031 11600 11469
rect 12100 11031 12150 11469
rect 12650 11031 12700 11469
rect 13200 11031 13250 11469
rect -469 10950 -31 11000
rect 81 10950 519 11000
rect 631 10950 1069 11000
rect 1181 10950 1619 11000
rect 1731 10950 2169 11000
rect 2281 10950 2719 11000
rect 2831 10950 3269 11000
rect 3381 10950 3819 11000
rect 3931 10950 4369 11000
rect 4481 10950 4919 11000
rect 5031 10950 5469 11000
rect 5581 10950 6019 11000
rect 6131 10950 6569 11000
rect 6681 10950 7119 11000
rect 7231 10950 7669 11000
rect 7781 10950 8219 11000
rect 8331 10950 8769 11000
rect 8881 10950 9319 11000
rect 9431 10950 9869 11000
rect 9981 10950 10419 11000
rect 10531 10950 10969 11000
rect 11081 10950 11519 11000
rect 11631 10950 12069 11000
rect 12181 10950 12619 11000
rect 12731 10950 13169 11000
rect 13281 10950 13719 11000
rect 0 10481 50 10919
rect 550 10481 600 10919
rect 1100 10481 1150 10919
rect 1650 10481 1700 10919
rect 2200 10481 2250 10919
rect 2750 10481 2800 10919
rect 3300 10481 3350 10919
rect 3850 10481 3900 10919
rect 4400 10481 4450 10919
rect 4950 10481 5000 10919
rect 5500 10481 5550 10919
rect 6050 10481 6100 10919
rect 6600 10481 6650 10919
rect 7150 10481 7200 10919
rect 7700 10481 7750 10919
rect 8250 10481 8300 10919
rect 8800 10481 8850 10919
rect 9350 10481 9400 10919
rect 9900 10481 9950 10919
rect 10450 10481 10500 10919
rect 11000 10481 11050 10919
rect 11550 10481 11600 10919
rect 12100 10481 12150 10919
rect 12650 10481 12700 10919
rect 13200 10481 13250 10919
rect -469 10400 -31 10450
rect 81 10400 519 10450
rect 631 10400 1069 10450
rect 1181 10400 1619 10450
rect 1731 10400 2169 10450
rect 2281 10400 2719 10450
rect 2831 10400 3269 10450
rect 3381 10400 3819 10450
rect 3931 10400 4369 10450
rect 4481 10400 4919 10450
rect 5031 10400 5469 10450
rect 5581 10400 6019 10450
rect 6131 10400 6569 10450
rect 6681 10400 7119 10450
rect 7231 10400 7669 10450
rect 7781 10400 8219 10450
rect 8331 10400 8769 10450
rect 8881 10400 9319 10450
rect 9431 10400 9869 10450
rect 9981 10400 10419 10450
rect 10531 10400 10969 10450
rect 11081 10400 11519 10450
rect 11631 10400 12069 10450
rect 12181 10400 12619 10450
rect 12731 10400 13169 10450
rect 13281 10400 13719 10450
rect 0 9931 50 10369
rect 550 9931 600 10369
rect 1100 9931 1150 10369
rect 1650 9931 1700 10369
rect 2200 9931 2250 10369
rect 2750 9931 2800 10369
rect 3300 9931 3350 10369
rect 3850 9931 3900 10369
rect 4400 9931 4450 10369
rect 4950 9931 5000 10369
rect 5500 9931 5550 10369
rect 6050 9931 6100 10369
rect 6600 9931 6650 10369
rect 7150 9931 7200 10369
rect 7700 9931 7750 10369
rect 8250 9931 8300 10369
rect 8800 9931 8850 10369
rect 9350 9931 9400 10369
rect 9900 9931 9950 10369
rect 10450 9931 10500 10369
rect 11000 9931 11050 10369
rect 11550 9931 11600 10369
rect 12100 9931 12150 10369
rect 12650 9931 12700 10369
rect 13200 9931 13250 10369
rect -469 9850 -31 9900
rect 81 9850 519 9900
rect 631 9850 1069 9900
rect 1181 9850 1619 9900
rect 1731 9850 2169 9900
rect 2281 9850 2719 9900
rect 2831 9850 3269 9900
rect 3381 9850 3819 9900
rect 3931 9850 4369 9900
rect 4481 9850 4919 9900
rect 5031 9850 5469 9900
rect 5581 9850 6019 9900
rect 6131 9850 6569 9900
rect 6681 9850 7119 9900
rect 7231 9850 7669 9900
rect 7781 9850 8219 9900
rect 8331 9850 8769 9900
rect 8881 9850 9319 9900
rect 9431 9850 9869 9900
rect 9981 9850 10419 9900
rect 10531 9850 10969 9900
rect 11081 9850 11519 9900
rect 11631 9850 12069 9900
rect 12181 9850 12619 9900
rect 12731 9850 13169 9900
rect 13281 9850 13719 9900
rect 0 9381 50 9819
rect 550 9381 600 9819
rect 1100 9381 1150 9819
rect 1650 9381 1700 9819
rect 2200 9381 2250 9819
rect 2750 9381 2800 9819
rect 3300 9381 3350 9819
rect 3850 9381 3900 9819
rect 4400 9381 4450 9819
rect 4950 9381 5000 9819
rect 5500 9381 5550 9819
rect 6050 9381 6100 9819
rect 6600 9381 6650 9819
rect 7150 9381 7200 9819
rect 7700 9381 7750 9819
rect 8250 9381 8300 9819
rect 8800 9381 8850 9819
rect 9350 9381 9400 9819
rect 9900 9381 9950 9819
rect 10450 9381 10500 9819
rect 11000 9381 11050 9819
rect 11550 9381 11600 9819
rect 12100 9381 12150 9819
rect 12650 9381 12700 9819
rect 13200 9381 13250 9819
rect -469 9300 -31 9350
rect 81 9300 519 9350
rect 631 9300 1069 9350
rect 1181 9300 1619 9350
rect 1731 9300 2169 9350
rect 2281 9300 2719 9350
rect 2831 9300 3269 9350
rect 3381 9300 3819 9350
rect 3931 9300 4369 9350
rect 4481 9300 4919 9350
rect 5031 9300 5469 9350
rect 5581 9300 6019 9350
rect 6131 9300 6569 9350
rect 6681 9300 7119 9350
rect 7231 9300 7669 9350
rect 7781 9300 8219 9350
rect 8331 9300 8769 9350
rect 8881 9300 9319 9350
rect 9431 9300 9869 9350
rect 9981 9300 10419 9350
rect 10531 9300 10969 9350
rect 11081 9300 11519 9350
rect 11631 9300 12069 9350
rect 12181 9300 12619 9350
rect 12731 9300 13169 9350
rect 13281 9300 13719 9350
rect 0 8831 50 9269
rect 550 8831 600 9269
rect 1100 8831 1150 9269
rect 1650 8831 1700 9269
rect 2200 8831 2250 9269
rect 2750 8831 2800 9269
rect 3300 8831 3350 9269
rect 3850 8831 3900 9269
rect 4400 8831 4450 9269
rect 4950 8831 5000 9269
rect 5500 8831 5550 9269
rect 6050 8831 6100 9269
rect 6600 8831 6650 9269
rect 7150 8831 7200 9269
rect 7700 8831 7750 9269
rect 8250 8831 8300 9269
rect 8800 8831 8850 9269
rect 9350 8831 9400 9269
rect 9900 8831 9950 9269
rect 10450 8831 10500 9269
rect 11000 8831 11050 9269
rect 11550 8831 11600 9269
rect 12100 8831 12150 9269
rect 12650 8831 12700 9269
rect 13200 8831 13250 9269
rect -469 8750 -31 8800
rect 81 8750 519 8800
rect 631 8750 1069 8800
rect 1181 8750 1619 8800
rect 1731 8750 2169 8800
rect 2281 8750 2719 8800
rect 2831 8750 3269 8800
rect 3381 8750 3819 8800
rect 3931 8750 4369 8800
rect 4481 8750 4919 8800
rect 5031 8750 5469 8800
rect 5581 8750 6019 8800
rect 6131 8750 6569 8800
rect 6681 8750 7119 8800
rect 7231 8750 7669 8800
rect 7781 8750 8219 8800
rect 8331 8750 8769 8800
rect 8881 8750 9319 8800
rect 9431 8750 9869 8800
rect 9981 8750 10419 8800
rect 10531 8750 10969 8800
rect 11081 8750 11519 8800
rect 11631 8750 12069 8800
rect 12181 8750 12619 8800
rect 12731 8750 13169 8800
rect 13281 8750 13719 8800
rect 0 8281 50 8719
rect 550 8281 600 8719
rect 1100 8281 1150 8719
rect 1650 8281 1700 8719
rect 2200 8281 2250 8719
rect 2750 8281 2800 8719
rect 3300 8281 3350 8719
rect 3850 8281 3900 8719
rect 4400 8281 4450 8719
rect 4950 8281 5000 8719
rect 5500 8281 5550 8719
rect 6050 8281 6100 8719
rect 6600 8281 6650 8719
rect 7150 8281 7200 8719
rect 7700 8281 7750 8719
rect 8250 8281 8300 8719
rect 8800 8281 8850 8719
rect 9350 8281 9400 8719
rect 9900 8281 9950 8719
rect 10450 8281 10500 8719
rect 11000 8281 11050 8719
rect 11550 8281 11600 8719
rect 12100 8281 12150 8719
rect 12650 8281 12700 8719
rect 13200 8281 13250 8719
rect -469 8200 -31 8250
rect 81 8200 519 8250
rect 631 8200 1069 8250
rect 1181 8200 1619 8250
rect 1731 8200 2169 8250
rect 2281 8200 2719 8250
rect 2831 8200 3269 8250
rect 3381 8200 3819 8250
rect 3931 8200 4369 8250
rect 4481 8200 4919 8250
rect 5031 8200 5469 8250
rect 5581 8200 6019 8250
rect 6131 8200 6569 8250
rect 6681 8200 7119 8250
rect 7231 8200 7669 8250
rect 7781 8200 8219 8250
rect 8331 8200 8769 8250
rect 8881 8200 9319 8250
rect 9431 8200 9869 8250
rect 9981 8200 10419 8250
rect 10531 8200 10969 8250
rect 11081 8200 11519 8250
rect 11631 8200 12069 8250
rect 12181 8200 12619 8250
rect 12731 8200 13169 8250
rect 13281 8200 13719 8250
rect 0 7731 50 8169
rect 550 7731 600 8169
rect 1100 7731 1150 8169
rect 1650 7731 1700 8169
rect 2200 7731 2250 8169
rect 2750 7731 2800 8169
rect 3300 7731 3350 8169
rect 3850 7731 3900 8169
rect 4400 7731 4450 8169
rect 4950 7731 5000 8169
rect 5500 7731 5550 8169
rect 6050 7731 6100 8169
rect 6600 7731 6650 8169
rect 7150 7731 7200 8169
rect 7700 7731 7750 8169
rect 8250 7731 8300 8169
rect 8800 7731 8850 8169
rect 9350 7731 9400 8169
rect 9900 7731 9950 8169
rect 10450 7731 10500 8169
rect 11000 7731 11050 8169
rect 11550 7731 11600 8169
rect 12100 7731 12150 8169
rect 12650 7731 12700 8169
rect 13200 7731 13250 8169
rect -469 7650 -31 7700
rect 81 7650 519 7700
rect 631 7650 1069 7700
rect 1181 7650 1619 7700
rect 1731 7650 2169 7700
rect 2281 7650 2719 7700
rect 2831 7650 3269 7700
rect 3381 7650 3819 7700
rect 3931 7650 4369 7700
rect 4481 7650 4919 7700
rect 5031 7650 5469 7700
rect 5581 7650 6019 7700
rect 6131 7650 6569 7700
rect 6681 7650 7119 7700
rect 7231 7650 7669 7700
rect 7781 7650 8219 7700
rect 8331 7650 8769 7700
rect 8881 7650 9319 7700
rect 9431 7650 9869 7700
rect 9981 7650 10419 7700
rect 10531 7650 10969 7700
rect 11081 7650 11519 7700
rect 11631 7650 12069 7700
rect 12181 7650 12619 7700
rect 12731 7650 13169 7700
rect 13281 7650 13719 7700
rect 0 7181 50 7619
rect 550 7181 600 7619
rect 1100 7181 1150 7619
rect 1650 7181 1700 7619
rect 2200 7181 2250 7619
rect 2750 7181 2800 7619
rect 3300 7181 3350 7619
rect 3850 7181 3900 7619
rect 4400 7181 4450 7619
rect 4950 7181 5000 7619
rect 5500 7181 5550 7619
rect 6050 7181 6100 7619
rect 6600 7181 6650 7619
rect 7150 7181 7200 7619
rect 7700 7181 7750 7619
rect 8250 7181 8300 7619
rect 8800 7181 8850 7619
rect 9350 7181 9400 7619
rect 9900 7181 9950 7619
rect 10450 7181 10500 7619
rect 11000 7181 11050 7619
rect 11550 7181 11600 7619
rect 12100 7181 12150 7619
rect 12650 7181 12700 7619
rect 13200 7181 13250 7619
rect -469 7100 -31 7150
rect 81 7100 519 7150
rect 631 7100 1069 7150
rect 1181 7100 1619 7150
rect 1731 7100 2169 7150
rect 2281 7100 2719 7150
rect 2831 7100 3269 7150
rect 3381 7100 3819 7150
rect 3931 7100 4369 7150
rect 4481 7100 4919 7150
rect 5031 7100 5469 7150
rect 5581 7100 6019 7150
rect 6131 7100 6569 7150
rect 6681 7100 7119 7150
rect 7231 7100 7669 7150
rect 7781 7100 8219 7150
rect 8331 7100 8769 7150
rect 8881 7100 9319 7150
rect 9431 7100 9869 7150
rect 9981 7100 10419 7150
rect 10531 7100 10969 7150
rect 11081 7100 11519 7150
rect 11631 7100 12069 7150
rect 12181 7100 12619 7150
rect 12731 7100 13169 7150
rect 13281 7100 13719 7150
rect 0 6631 50 7069
rect 550 6631 600 7069
rect 1100 6631 1150 7069
rect 1650 6631 1700 7069
rect 2200 6631 2250 7069
rect 2750 6631 2800 7069
rect 3300 6631 3350 7069
rect 3850 6631 3900 7069
rect 4400 6631 4450 7069
rect 4950 6631 5000 7069
rect 5500 6631 5550 7069
rect 6050 6631 6100 7069
rect 6600 6631 6650 7069
rect 7150 6631 7200 7069
rect 7700 6631 7750 7069
rect 8250 6631 8300 7069
rect 8800 6631 8850 7069
rect 9350 6631 9400 7069
rect 9900 6631 9950 7069
rect 10450 6631 10500 7069
rect 11000 6631 11050 7069
rect 11550 6631 11600 7069
rect 12100 6631 12150 7069
rect 12650 6631 12700 7069
rect 13200 6631 13250 7069
rect -469 6550 -31 6600
rect 81 6550 519 6600
rect 631 6550 1069 6600
rect 1181 6550 1619 6600
rect 1731 6550 2169 6600
rect 2281 6550 2719 6600
rect 2831 6550 3269 6600
rect 3381 6550 3819 6600
rect 3931 6550 4369 6600
rect 4481 6550 4919 6600
rect 5031 6550 5469 6600
rect 5581 6550 6019 6600
rect 6131 6550 6569 6600
rect 6681 6550 7119 6600
rect 7231 6550 7669 6600
rect 7781 6550 8219 6600
rect 8331 6550 8769 6600
rect 8881 6550 9319 6600
rect 9431 6550 9869 6600
rect 9981 6550 10419 6600
rect 10531 6550 10969 6600
rect 11081 6550 11519 6600
rect 11631 6550 12069 6600
rect 12181 6550 12619 6600
rect 12731 6550 13169 6600
rect 13281 6550 13719 6600
rect 0 6081 50 6519
rect 550 6081 600 6519
rect 1100 6081 1150 6519
rect 1650 6081 1700 6519
rect 2200 6081 2250 6519
rect 2750 6081 2800 6519
rect 3300 6081 3350 6519
rect 3850 6081 3900 6519
rect 4400 6081 4450 6519
rect 4950 6081 5000 6519
rect 5500 6081 5550 6519
rect 6050 6081 6100 6519
rect 6600 6081 6650 6519
rect 7150 6081 7200 6519
rect 7700 6081 7750 6519
rect 8250 6081 8300 6519
rect 8800 6081 8850 6519
rect 9350 6081 9400 6519
rect 9900 6081 9950 6519
rect 10450 6081 10500 6519
rect 11000 6081 11050 6519
rect 11550 6081 11600 6519
rect 12100 6081 12150 6519
rect 12650 6081 12700 6519
rect 13200 6081 13250 6519
rect -469 6000 -31 6050
rect 81 6000 519 6050
rect 631 6000 1069 6050
rect 1181 6000 1619 6050
rect 1731 6000 2169 6050
rect 2281 6000 2719 6050
rect 2831 6000 3269 6050
rect 3381 6000 3819 6050
rect 3931 6000 4369 6050
rect 4481 6000 4919 6050
rect 5031 6000 5469 6050
rect 5581 6000 6019 6050
rect 6131 6000 6569 6050
rect 6681 6000 7119 6050
rect 7231 6000 7669 6050
rect 7781 6000 8219 6050
rect 8331 6000 8769 6050
rect 8881 6000 9319 6050
rect 9431 6000 9869 6050
rect 9981 6000 10419 6050
rect 10531 6000 10969 6050
rect 11081 6000 11519 6050
rect 11631 6000 12069 6050
rect 12181 6000 12619 6050
rect 12731 6000 13169 6050
rect 13281 6000 13719 6050
rect 0 5531 50 5969
rect 550 5531 600 5969
rect 1100 5531 1150 5969
rect 1650 5531 1700 5969
rect 2200 5531 2250 5969
rect 2750 5531 2800 5969
rect 3300 5531 3350 5969
rect 3850 5531 3900 5969
rect 4400 5531 4450 5969
rect 4950 5531 5000 5969
rect 5500 5531 5550 5969
rect 6050 5531 6100 5969
rect 6600 5531 6650 5969
rect 7150 5531 7200 5969
rect 7700 5531 7750 5969
rect 8250 5531 8300 5969
rect 8800 5531 8850 5969
rect 9350 5531 9400 5969
rect 9900 5531 9950 5969
rect 10450 5531 10500 5969
rect 11000 5531 11050 5969
rect 11550 5531 11600 5969
rect 12100 5531 12150 5969
rect 12650 5531 12700 5969
rect 13200 5531 13250 5969
rect -469 5450 -31 5500
rect 81 5450 519 5500
rect 631 5450 1069 5500
rect 1181 5450 1619 5500
rect 1731 5450 2169 5500
rect 2281 5450 2719 5500
rect 2831 5450 3269 5500
rect 3381 5450 3819 5500
rect 3931 5450 4369 5500
rect 4481 5450 4919 5500
rect 5031 5450 5469 5500
rect 5581 5450 6019 5500
rect 6131 5450 6569 5500
rect 6681 5450 7119 5500
rect 7231 5450 7669 5500
rect 7781 5450 8219 5500
rect 8331 5450 8769 5500
rect 8881 5450 9319 5500
rect 9431 5450 9869 5500
rect 9981 5450 10419 5500
rect 10531 5450 10969 5500
rect 11081 5450 11519 5500
rect 11631 5450 12069 5500
rect 12181 5450 12619 5500
rect 12731 5450 13169 5500
rect 13281 5450 13719 5500
rect 0 4981 50 5419
rect 550 4981 600 5419
rect 1100 4981 1150 5419
rect 1650 4981 1700 5419
rect 2200 4981 2250 5419
rect 2750 4981 2800 5419
rect 3300 4981 3350 5419
rect 3850 4981 3900 5419
rect 4400 4981 4450 5419
rect 4950 4981 5000 5419
rect 5500 4981 5550 5419
rect 6050 4981 6100 5419
rect 6600 4981 6650 5419
rect 7150 4981 7200 5419
rect 7700 4981 7750 5419
rect 8250 4981 8300 5419
rect 8800 4981 8850 5419
rect 9350 4981 9400 5419
rect 9900 4981 9950 5419
rect 10450 4981 10500 5419
rect 11000 4981 11050 5419
rect 11550 4981 11600 5419
rect 12100 4981 12150 5419
rect 12650 4981 12700 5419
rect 13200 4981 13250 5419
rect -469 4900 -31 4950
rect 81 4900 519 4950
rect 631 4900 1069 4950
rect 1181 4900 1619 4950
rect 1731 4900 2169 4950
rect 2281 4900 2719 4950
rect 2831 4900 3269 4950
rect 3381 4900 3819 4950
rect 3931 4900 4369 4950
rect 4481 4900 4919 4950
rect 5031 4900 5469 4950
rect 5581 4900 6019 4950
rect 6131 4900 6569 4950
rect 6681 4900 7119 4950
rect 7231 4900 7669 4950
rect 7781 4900 8219 4950
rect 8331 4900 8769 4950
rect 8881 4900 9319 4950
rect 9431 4900 9869 4950
rect 9981 4900 10419 4950
rect 10531 4900 10969 4950
rect 11081 4900 11519 4950
rect 11631 4900 12069 4950
rect 12181 4900 12619 4950
rect 12731 4900 13169 4950
rect 13281 4900 13719 4950
rect 0 4431 50 4869
rect 550 4431 600 4869
rect 1100 4431 1150 4869
rect 1650 4431 1700 4869
rect 2200 4431 2250 4869
rect 2750 4431 2800 4869
rect 3300 4431 3350 4869
rect 3850 4431 3900 4869
rect 4400 4431 4450 4869
rect 4950 4431 5000 4869
rect 5500 4431 5550 4869
rect 6050 4431 6100 4869
rect 6600 4431 6650 4869
rect 7150 4431 7200 4869
rect 7700 4431 7750 4869
rect 8250 4431 8300 4869
rect 8800 4431 8850 4869
rect 9350 4431 9400 4869
rect 9900 4431 9950 4869
rect 10450 4431 10500 4869
rect 11000 4431 11050 4869
rect 11550 4431 11600 4869
rect 12100 4431 12150 4869
rect 12650 4431 12700 4869
rect 13200 4431 13250 4869
rect -469 4350 -31 4400
rect 81 4350 519 4400
rect 631 4350 1069 4400
rect 1181 4350 1619 4400
rect 1731 4350 2169 4400
rect 2281 4350 2719 4400
rect 2831 4350 3269 4400
rect 3381 4350 3819 4400
rect 3931 4350 4369 4400
rect 4481 4350 4919 4400
rect 5031 4350 5469 4400
rect 5581 4350 6019 4400
rect 6131 4350 6569 4400
rect 6681 4350 7119 4400
rect 7231 4350 7669 4400
rect 7781 4350 8219 4400
rect 8331 4350 8769 4400
rect 8881 4350 9319 4400
rect 9431 4350 9869 4400
rect 9981 4350 10419 4400
rect 10531 4350 10969 4400
rect 11081 4350 11519 4400
rect 11631 4350 12069 4400
rect 12181 4350 12619 4400
rect 12731 4350 13169 4400
rect 13281 4350 13719 4400
rect 0 3881 50 4319
rect 550 3881 600 4319
rect 1100 3881 1150 4319
rect 1650 3881 1700 4319
rect 2200 3881 2250 4319
rect 2750 3881 2800 4319
rect 3300 3881 3350 4319
rect 3850 3881 3900 4319
rect 4400 3881 4450 4319
rect 4950 3881 5000 4319
rect 5500 3881 5550 4319
rect 6050 3881 6100 4319
rect 6600 3881 6650 4319
rect 7150 3881 7200 4319
rect 7700 3881 7750 4319
rect 8250 3881 8300 4319
rect 8800 3881 8850 4319
rect 9350 3881 9400 4319
rect 9900 3881 9950 4319
rect 10450 3881 10500 4319
rect 11000 3881 11050 4319
rect 11550 3881 11600 4319
rect 12100 3881 12150 4319
rect 12650 3881 12700 4319
rect 13200 3881 13250 4319
rect -469 3800 -31 3850
rect 81 3800 519 3850
rect 631 3800 1069 3850
rect 1181 3800 1619 3850
rect 1731 3800 2169 3850
rect 2281 3800 2719 3850
rect 2831 3800 3269 3850
rect 3381 3800 3819 3850
rect 3931 3800 4369 3850
rect 4481 3800 4919 3850
rect 5031 3800 5469 3850
rect 5581 3800 6019 3850
rect 6131 3800 6569 3850
rect 6681 3800 7119 3850
rect 7231 3800 7669 3850
rect 7781 3800 8219 3850
rect 8331 3800 8769 3850
rect 8881 3800 9319 3850
rect 9431 3800 9869 3850
rect 9981 3800 10419 3850
rect 10531 3800 10969 3850
rect 11081 3800 11519 3850
rect 11631 3800 12069 3850
rect 12181 3800 12619 3850
rect 12731 3800 13169 3850
rect 13281 3800 13719 3850
rect 0 3331 50 3769
rect 550 3331 600 3769
rect 1100 3331 1150 3769
rect 1650 3331 1700 3769
rect 2200 3331 2250 3769
rect 2750 3331 2800 3769
rect 3300 3331 3350 3769
rect 3850 3331 3900 3769
rect 4400 3331 4450 3769
rect 4950 3331 5000 3769
rect 5500 3331 5550 3769
rect 6050 3331 6100 3769
rect 6600 3331 6650 3769
rect 7150 3331 7200 3769
rect 7700 3331 7750 3769
rect 8250 3331 8300 3769
rect 8800 3331 8850 3769
rect 9350 3331 9400 3769
rect 9900 3331 9950 3769
rect 10450 3331 10500 3769
rect 11000 3331 11050 3769
rect 11550 3331 11600 3769
rect 12100 3331 12150 3769
rect 12650 3331 12700 3769
rect 13200 3331 13250 3769
rect -469 3250 -31 3300
rect 81 3250 519 3300
rect 631 3250 1069 3300
rect 1181 3250 1619 3300
rect 1731 3250 2169 3300
rect 2281 3250 2719 3300
rect 2831 3250 3269 3300
rect 3381 3250 3819 3300
rect 3931 3250 4369 3300
rect 4481 3250 4919 3300
rect 5031 3250 5469 3300
rect 5581 3250 6019 3300
rect 6131 3250 6569 3300
rect 6681 3250 7119 3300
rect 7231 3250 7669 3300
rect 7781 3250 8219 3300
rect 8331 3250 8769 3300
rect 8881 3250 9319 3300
rect 9431 3250 9869 3300
rect 9981 3250 10419 3300
rect 10531 3250 10969 3300
rect 11081 3250 11519 3300
rect 11631 3250 12069 3300
rect 12181 3250 12619 3300
rect 12731 3250 13169 3300
rect 13281 3250 13719 3300
rect 0 2781 50 3219
rect 550 2781 600 3219
rect 1100 2781 1150 3219
rect 1650 2781 1700 3219
rect 2200 2781 2250 3219
rect 2750 2781 2800 3219
rect 3300 2781 3350 3219
rect 3850 2781 3900 3219
rect 4400 2781 4450 3219
rect 4950 2781 5000 3219
rect 5500 2781 5550 3219
rect 6050 2781 6100 3219
rect 6600 2781 6650 3219
rect 7150 2781 7200 3219
rect 7700 2781 7750 3219
rect 8250 2781 8300 3219
rect 8800 2781 8850 3219
rect 9350 2781 9400 3219
rect 9900 2781 9950 3219
rect 10450 2781 10500 3219
rect 11000 2781 11050 3219
rect 11550 2781 11600 3219
rect 12100 2781 12150 3219
rect 12650 2781 12700 3219
rect 13200 2781 13250 3219
rect -469 2700 -31 2750
rect 81 2700 519 2750
rect 631 2700 1069 2750
rect 1181 2700 1619 2750
rect 1731 2700 2169 2750
rect 2281 2700 2719 2750
rect 2831 2700 3269 2750
rect 3381 2700 3819 2750
rect 3931 2700 4369 2750
rect 4481 2700 4919 2750
rect 5031 2700 5469 2750
rect 5581 2700 6019 2750
rect 6131 2700 6569 2750
rect 6681 2700 7119 2750
rect 7231 2700 7669 2750
rect 7781 2700 8219 2750
rect 8331 2700 8769 2750
rect 8881 2700 9319 2750
rect 9431 2700 9869 2750
rect 9981 2700 10419 2750
rect 10531 2700 10969 2750
rect 11081 2700 11519 2750
rect 11631 2700 12069 2750
rect 12181 2700 12619 2750
rect 12731 2700 13169 2750
rect 13281 2700 13719 2750
rect 0 2231 50 2669
rect 550 2231 600 2669
rect 1100 2231 1150 2669
rect 1650 2231 1700 2669
rect 2200 2231 2250 2669
rect 2750 2231 2800 2669
rect 3300 2231 3350 2669
rect 3850 2231 3900 2669
rect 4400 2231 4450 2669
rect 4950 2231 5000 2669
rect 5500 2231 5550 2669
rect 6050 2231 6100 2669
rect 6600 2231 6650 2669
rect 7150 2231 7200 2669
rect 7700 2231 7750 2669
rect 8250 2231 8300 2669
rect 8800 2231 8850 2669
rect 9350 2231 9400 2669
rect 9900 2231 9950 2669
rect 10450 2231 10500 2669
rect 11000 2231 11050 2669
rect 11550 2231 11600 2669
rect 12100 2231 12150 2669
rect 12650 2231 12700 2669
rect 13200 2231 13250 2669
rect -469 2150 -31 2200
rect 81 2150 519 2200
rect 631 2150 1069 2200
rect 1181 2150 1619 2200
rect 1731 2150 2169 2200
rect 2281 2150 2719 2200
rect 2831 2150 3269 2200
rect 3381 2150 3819 2200
rect 3931 2150 4369 2200
rect 4481 2150 4919 2200
rect 5031 2150 5469 2200
rect 5581 2150 6019 2200
rect 6131 2150 6569 2200
rect 6681 2150 7119 2200
rect 7231 2150 7669 2200
rect 7781 2150 8219 2200
rect 8331 2150 8769 2200
rect 8881 2150 9319 2200
rect 9431 2150 9869 2200
rect 9981 2150 10419 2200
rect 10531 2150 10969 2200
rect 11081 2150 11519 2200
rect 11631 2150 12069 2200
rect 12181 2150 12619 2200
rect 12731 2150 13169 2200
rect 13281 2150 13719 2200
rect 0 1681 50 2119
rect 550 1681 600 2119
rect 1100 1681 1150 2119
rect 1650 1681 1700 2119
rect 2200 1681 2250 2119
rect 2750 1681 2800 2119
rect 3300 1681 3350 2119
rect 3850 1681 3900 2119
rect 4400 1681 4450 2119
rect 4950 1681 5000 2119
rect 5500 1681 5550 2119
rect 6050 1681 6100 2119
rect 6600 1681 6650 2119
rect 7150 1681 7200 2119
rect 7700 1681 7750 2119
rect 8250 1681 8300 2119
rect 8800 1681 8850 2119
rect 9350 1681 9400 2119
rect 9900 1681 9950 2119
rect 10450 1681 10500 2119
rect 11000 1681 11050 2119
rect 11550 1681 11600 2119
rect 12100 1681 12150 2119
rect 12650 1681 12700 2119
rect 13200 1681 13250 2119
rect -469 1600 -31 1650
rect 81 1600 519 1650
rect 631 1600 1069 1650
rect 1181 1600 1619 1650
rect 1731 1600 2169 1650
rect 2281 1600 2719 1650
rect 2831 1600 3269 1650
rect 3381 1600 3819 1650
rect 3931 1600 4369 1650
rect 4481 1600 4919 1650
rect 5031 1600 5469 1650
rect 5581 1600 6019 1650
rect 6131 1600 6569 1650
rect 6681 1600 7119 1650
rect 7231 1600 7669 1650
rect 7781 1600 8219 1650
rect 8331 1600 8769 1650
rect 8881 1600 9319 1650
rect 9431 1600 9869 1650
rect 9981 1600 10419 1650
rect 10531 1600 10969 1650
rect 11081 1600 11519 1650
rect 11631 1600 12069 1650
rect 12181 1600 12619 1650
rect 12731 1600 13169 1650
rect 13281 1600 13719 1650
rect 0 1131 50 1569
rect 550 1131 600 1569
rect 1100 1131 1150 1569
rect 1650 1131 1700 1569
rect 2200 1131 2250 1569
rect 2750 1131 2800 1569
rect 3300 1131 3350 1569
rect 3850 1131 3900 1569
rect 4400 1131 4450 1569
rect 4950 1131 5000 1569
rect 5500 1131 5550 1569
rect 6050 1131 6100 1569
rect 6600 1131 6650 1569
rect 7150 1131 7200 1569
rect 7700 1131 7750 1569
rect 8250 1131 8300 1569
rect 8800 1131 8850 1569
rect 9350 1131 9400 1569
rect 9900 1131 9950 1569
rect 10450 1131 10500 1569
rect 11000 1131 11050 1569
rect 11550 1131 11600 1569
rect 12100 1131 12150 1569
rect 12650 1131 12700 1569
rect 13200 1131 13250 1569
rect -469 1050 -31 1100
rect 81 1050 519 1100
rect 631 1050 1069 1100
rect 1181 1050 1619 1100
rect 1731 1050 2169 1100
rect 2281 1050 2719 1100
rect 2831 1050 3269 1100
rect 3381 1050 3819 1100
rect 3931 1050 4369 1100
rect 4481 1050 4919 1100
rect 5031 1050 5469 1100
rect 5581 1050 6019 1100
rect 6131 1050 6569 1100
rect 6681 1050 7119 1100
rect 7231 1050 7669 1100
rect 7781 1050 8219 1100
rect 8331 1050 8769 1100
rect 8881 1050 9319 1100
rect 9431 1050 9869 1100
rect 9981 1050 10419 1100
rect 10531 1050 10969 1100
rect 11081 1050 11519 1100
rect 11631 1050 12069 1100
rect 12181 1050 12619 1100
rect 12731 1050 13169 1100
rect 13281 1050 13719 1100
rect 0 581 50 1019
rect 550 581 600 1019
rect 1100 581 1150 1019
rect 1650 581 1700 1019
rect 2200 581 2250 1019
rect 2750 581 2800 1019
rect 3300 581 3350 1019
rect 3850 581 3900 1019
rect 4400 581 4450 1019
rect 4950 581 5000 1019
rect 5500 581 5550 1019
rect 6050 581 6100 1019
rect 6600 581 6650 1019
rect 7150 581 7200 1019
rect 7700 581 7750 1019
rect 8250 581 8300 1019
rect 8800 581 8850 1019
rect 9350 581 9400 1019
rect 9900 581 9950 1019
rect 10450 581 10500 1019
rect 11000 581 11050 1019
rect 11550 581 11600 1019
rect 12100 581 12150 1019
rect 12650 581 12700 1019
rect 13200 581 13250 1019
rect -469 500 -31 550
rect 81 500 519 550
rect 631 500 1069 550
rect 1181 500 1619 550
rect 1731 500 2169 550
rect 2281 500 2719 550
rect 2831 500 3269 550
rect 3381 500 3819 550
rect 3931 500 4369 550
rect 4481 500 4919 550
rect 5031 500 5469 550
rect 5581 500 6019 550
rect 6131 500 6569 550
rect 6681 500 7119 550
rect 7231 500 7669 550
rect 7781 500 8219 550
rect 8331 500 8769 550
rect 8881 500 9319 550
rect 9431 500 9869 550
rect 9981 500 10419 550
rect 10531 500 10969 550
rect 11081 500 11519 550
rect 11631 500 12069 550
rect 12181 500 12619 550
rect 12731 500 13169 550
rect 13281 500 13719 550
rect 0 31 50 469
rect 550 31 600 469
rect 1100 31 1150 469
rect 1650 31 1700 469
rect 2200 31 2250 469
rect 2750 31 2800 469
rect 3300 31 3350 469
rect 3850 31 3900 469
rect 4400 31 4450 469
rect 4950 31 5000 469
rect 5500 31 5550 469
rect 6050 31 6100 469
rect 6600 31 6650 469
rect 7150 31 7200 469
rect 7700 31 7750 469
rect 8250 31 8300 469
rect 8800 31 8850 469
rect 9350 31 9400 469
rect 9900 31 9950 469
rect 10450 31 10500 469
rect 11000 31 11050 469
rect 11550 31 11600 469
rect 12100 31 12150 469
rect 12650 31 12700 469
rect 13200 31 13250 469
rect -469 -50 -31 0
rect 81 -50 519 0
rect 631 -50 1069 0
rect 1181 -50 1619 0
rect 1731 -50 2169 0
rect 2281 -50 2719 0
rect 2831 -50 3269 0
rect 3381 -50 3819 0
rect 3931 -50 4369 0
rect 4481 -50 4919 0
rect 5031 -50 5469 0
rect 5581 -50 6019 0
rect 6131 -50 6569 0
rect 6681 -50 7119 0
rect 7231 -50 7669 0
rect 7781 -50 8219 0
rect 8331 -50 8769 0
rect 8881 -50 9319 0
rect 9431 -50 9869 0
rect 9981 -50 10419 0
rect 10531 -50 10969 0
rect 11081 -50 11519 0
rect 11631 -50 12069 0
rect 12181 -50 12619 0
rect 12731 -50 13169 0
rect 13281 -50 13719 0
rect 0 -519 50 -81
rect 550 -519 600 -81
rect 1100 -519 1150 -81
rect 1650 -519 1700 -81
rect 2200 -519 2250 -81
rect 2750 -519 2800 -81
rect 3300 -519 3350 -81
rect 3850 -519 3900 -81
rect 4400 -519 4450 -81
rect 4950 -519 5000 -81
rect 5500 -519 5550 -81
rect 6050 -519 6100 -81
rect 6600 -519 6650 -81
rect 7150 -519 7200 -81
rect 7700 -519 7750 -81
rect 8250 -519 8300 -81
rect 8800 -519 8850 -81
rect 9350 -519 9400 -81
rect 9900 -519 9950 -81
rect 10450 -519 10500 -81
rect 11000 -519 11050 -81
rect 11550 -519 11600 -81
rect 12100 -519 12150 -81
rect 12650 -519 12700 -81
rect 13200 -519 13250 -81
<< mvpdiff >>
rect 79 13669 521 13671
rect 1179 13669 1621 13671
rect 2279 13669 2721 13671
rect 3379 13669 3821 13671
rect 4479 13669 4921 13671
rect 5579 13669 6021 13671
rect 6679 13669 7121 13671
rect 7779 13669 8221 13671
rect 8879 13669 9321 13671
rect 9979 13669 10421 13671
rect 11079 13669 11521 13671
rect 12179 13669 12621 13671
rect 13279 13669 13721 13671
rect -29 13663 0 13669
rect -29 13264 -23 13663
rect -64 13237 -23 13264
rect -6 13237 0 13663
rect -64 13231 0 13237
rect 50 13663 550 13669
rect 50 13237 56 13663
rect 73 13615 527 13663
rect 73 13285 135 13615
rect 465 13285 527 13615
rect 73 13237 527 13285
rect 544 13237 550 13663
rect 50 13231 550 13237
rect 600 13663 629 13669
rect 600 13237 606 13663
rect 623 13264 629 13663
rect 1071 13663 1100 13669
rect 1071 13264 1077 13663
rect 623 13237 664 13264
rect 600 13231 664 13237
rect -64 13229 -31 13231
rect -469 13223 -31 13229
rect -469 13206 -463 13223
rect -37 13206 -31 13223
rect -469 13200 -31 13206
rect 79 13229 521 13231
rect 81 13223 519 13229
rect 81 13206 87 13223
rect 513 13206 519 13223
rect 81 13200 519 13206
rect 631 13229 664 13231
rect 1036 13237 1077 13264
rect 1094 13237 1100 13663
rect 1036 13231 1100 13237
rect 1150 13663 1650 13669
rect 1150 13237 1156 13663
rect 1173 13615 1627 13663
rect 1173 13285 1235 13615
rect 1565 13285 1627 13615
rect 1173 13237 1627 13285
rect 1644 13237 1650 13663
rect 1150 13231 1650 13237
rect 1700 13663 1729 13669
rect 1700 13237 1706 13663
rect 1723 13264 1729 13663
rect 2171 13663 2200 13669
rect 2171 13264 2177 13663
rect 1723 13237 1764 13264
rect 1700 13231 1764 13237
rect 1036 13229 1069 13231
rect 631 13223 1069 13229
rect 631 13206 637 13223
rect 1063 13206 1069 13223
rect 631 13200 1069 13206
rect 1179 13229 1621 13231
rect 1181 13223 1619 13229
rect 1181 13206 1187 13223
rect 1613 13206 1619 13223
rect 1181 13200 1619 13206
rect 1731 13229 1764 13231
rect 2136 13237 2177 13264
rect 2194 13237 2200 13663
rect 2136 13231 2200 13237
rect 2250 13663 2750 13669
rect 2250 13237 2256 13663
rect 2273 13615 2727 13663
rect 2273 13285 2335 13615
rect 2665 13285 2727 13615
rect 2273 13237 2727 13285
rect 2744 13237 2750 13663
rect 2250 13231 2750 13237
rect 2800 13663 2829 13669
rect 2800 13237 2806 13663
rect 2823 13264 2829 13663
rect 3271 13663 3300 13669
rect 3271 13264 3277 13663
rect 2823 13237 2864 13264
rect 2800 13231 2864 13237
rect 2136 13229 2169 13231
rect 1731 13223 2169 13229
rect 1731 13206 1737 13223
rect 2163 13206 2169 13223
rect 1731 13200 2169 13206
rect 2279 13229 2721 13231
rect 2281 13223 2719 13229
rect 2281 13206 2287 13223
rect 2713 13206 2719 13223
rect 2281 13200 2719 13206
rect 2831 13229 2864 13231
rect 3236 13237 3277 13264
rect 3294 13237 3300 13663
rect 3236 13231 3300 13237
rect 3350 13663 3850 13669
rect 3350 13237 3356 13663
rect 3373 13615 3827 13663
rect 3373 13285 3435 13615
rect 3765 13285 3827 13615
rect 3373 13237 3827 13285
rect 3844 13237 3850 13663
rect 3350 13231 3850 13237
rect 3900 13663 3929 13669
rect 3900 13237 3906 13663
rect 3923 13264 3929 13663
rect 4371 13663 4400 13669
rect 4371 13264 4377 13663
rect 3923 13237 3964 13264
rect 3900 13231 3964 13237
rect 3236 13229 3269 13231
rect 2831 13223 3269 13229
rect 2831 13206 2837 13223
rect 3263 13206 3269 13223
rect 2831 13200 3269 13206
rect 3379 13229 3821 13231
rect 3381 13223 3819 13229
rect 3381 13206 3387 13223
rect 3813 13206 3819 13223
rect 3381 13200 3819 13206
rect 3931 13229 3964 13231
rect 4336 13237 4377 13264
rect 4394 13237 4400 13663
rect 4336 13231 4400 13237
rect 4450 13663 4950 13669
rect 4450 13237 4456 13663
rect 4473 13615 4927 13663
rect 4473 13285 4535 13615
rect 4865 13285 4927 13615
rect 4473 13237 4927 13285
rect 4944 13237 4950 13663
rect 4450 13231 4950 13237
rect 5000 13663 5029 13669
rect 5000 13237 5006 13663
rect 5023 13264 5029 13663
rect 5471 13663 5500 13669
rect 5471 13264 5477 13663
rect 5023 13237 5064 13264
rect 5000 13231 5064 13237
rect 4336 13229 4369 13231
rect 3931 13223 4369 13229
rect 3931 13206 3937 13223
rect 4363 13206 4369 13223
rect 3931 13200 4369 13206
rect 4479 13229 4921 13231
rect 4481 13223 4919 13229
rect 4481 13206 4487 13223
rect 4913 13206 4919 13223
rect 4481 13200 4919 13206
rect 5031 13229 5064 13231
rect 5436 13237 5477 13264
rect 5494 13237 5500 13663
rect 5436 13231 5500 13237
rect 5550 13663 6050 13669
rect 5550 13237 5556 13663
rect 5573 13615 6027 13663
rect 5573 13285 5635 13615
rect 5965 13285 6027 13615
rect 5573 13237 6027 13285
rect 6044 13237 6050 13663
rect 5550 13231 6050 13237
rect 6100 13663 6129 13669
rect 6100 13237 6106 13663
rect 6123 13264 6129 13663
rect 6571 13663 6600 13669
rect 6571 13264 6577 13663
rect 6123 13237 6164 13264
rect 6100 13231 6164 13237
rect 5436 13229 5469 13231
rect 5031 13223 5469 13229
rect 5031 13206 5037 13223
rect 5463 13206 5469 13223
rect 5031 13200 5469 13206
rect 5579 13229 6021 13231
rect 5581 13223 6019 13229
rect 5581 13206 5587 13223
rect 6013 13206 6019 13223
rect 5581 13200 6019 13206
rect 6131 13229 6164 13231
rect 6536 13237 6577 13264
rect 6594 13237 6600 13663
rect 6536 13231 6600 13237
rect 6650 13663 7150 13669
rect 6650 13237 6656 13663
rect 6673 13615 7127 13663
rect 6673 13285 6735 13615
rect 7065 13285 7127 13615
rect 6673 13237 7127 13285
rect 7144 13237 7150 13663
rect 6650 13231 7150 13237
rect 7200 13663 7229 13669
rect 7200 13237 7206 13663
rect 7223 13264 7229 13663
rect 7671 13663 7700 13669
rect 7671 13264 7677 13663
rect 7223 13237 7264 13264
rect 7200 13231 7264 13237
rect 6536 13229 6569 13231
rect 6131 13223 6569 13229
rect 6131 13206 6137 13223
rect 6563 13206 6569 13223
rect 6131 13200 6569 13206
rect 6679 13229 7121 13231
rect 6681 13223 7119 13229
rect 6681 13206 6687 13223
rect 7113 13206 7119 13223
rect 6681 13200 7119 13206
rect 7231 13229 7264 13231
rect 7636 13237 7677 13264
rect 7694 13237 7700 13663
rect 7636 13231 7700 13237
rect 7750 13663 8250 13669
rect 7750 13237 7756 13663
rect 7773 13615 8227 13663
rect 7773 13285 7835 13615
rect 8165 13285 8227 13615
rect 7773 13237 8227 13285
rect 8244 13237 8250 13663
rect 7750 13231 8250 13237
rect 8300 13663 8329 13669
rect 8300 13237 8306 13663
rect 8323 13264 8329 13663
rect 8771 13663 8800 13669
rect 8771 13264 8777 13663
rect 8323 13237 8364 13264
rect 8300 13231 8364 13237
rect 7636 13229 7669 13231
rect 7231 13223 7669 13229
rect 7231 13206 7237 13223
rect 7663 13206 7669 13223
rect 7231 13200 7669 13206
rect 7779 13229 8221 13231
rect 7781 13223 8219 13229
rect 7781 13206 7787 13223
rect 8213 13206 8219 13223
rect 7781 13200 8219 13206
rect 8331 13229 8364 13231
rect 8736 13237 8777 13264
rect 8794 13237 8800 13663
rect 8736 13231 8800 13237
rect 8850 13663 9350 13669
rect 8850 13237 8856 13663
rect 8873 13615 9327 13663
rect 8873 13285 8935 13615
rect 9265 13285 9327 13615
rect 8873 13237 9327 13285
rect 9344 13237 9350 13663
rect 8850 13231 9350 13237
rect 9400 13663 9429 13669
rect 9400 13237 9406 13663
rect 9423 13264 9429 13663
rect 9871 13663 9900 13669
rect 9871 13264 9877 13663
rect 9423 13237 9464 13264
rect 9400 13231 9464 13237
rect 8736 13229 8769 13231
rect 8331 13223 8769 13229
rect 8331 13206 8337 13223
rect 8763 13206 8769 13223
rect 8331 13200 8769 13206
rect 8879 13229 9321 13231
rect 8881 13223 9319 13229
rect 8881 13206 8887 13223
rect 9313 13206 9319 13223
rect 8881 13200 9319 13206
rect 9431 13229 9464 13231
rect 9836 13237 9877 13264
rect 9894 13237 9900 13663
rect 9836 13231 9900 13237
rect 9950 13663 10450 13669
rect 9950 13237 9956 13663
rect 9973 13615 10427 13663
rect 9973 13285 10035 13615
rect 10365 13285 10427 13615
rect 9973 13237 10427 13285
rect 10444 13237 10450 13663
rect 9950 13231 10450 13237
rect 10500 13663 10529 13669
rect 10500 13237 10506 13663
rect 10523 13264 10529 13663
rect 10971 13663 11000 13669
rect 10971 13264 10977 13663
rect 10523 13237 10564 13264
rect 10500 13231 10564 13237
rect 9836 13229 9869 13231
rect 9431 13223 9869 13229
rect 9431 13206 9437 13223
rect 9863 13206 9869 13223
rect 9431 13200 9869 13206
rect 9979 13229 10421 13231
rect 9981 13223 10419 13229
rect 9981 13206 9987 13223
rect 10413 13206 10419 13223
rect 9981 13200 10419 13206
rect 10531 13229 10564 13231
rect 10936 13237 10977 13264
rect 10994 13237 11000 13663
rect 10936 13231 11000 13237
rect 11050 13663 11550 13669
rect 11050 13237 11056 13663
rect 11073 13615 11527 13663
rect 11073 13285 11135 13615
rect 11465 13285 11527 13615
rect 11073 13237 11527 13285
rect 11544 13237 11550 13663
rect 11050 13231 11550 13237
rect 11600 13663 11629 13669
rect 11600 13237 11606 13663
rect 11623 13264 11629 13663
rect 12071 13663 12100 13669
rect 12071 13264 12077 13663
rect 11623 13237 11664 13264
rect 11600 13231 11664 13237
rect 10936 13229 10969 13231
rect 10531 13223 10969 13229
rect 10531 13206 10537 13223
rect 10963 13206 10969 13223
rect 10531 13200 10969 13206
rect 11079 13229 11521 13231
rect 11081 13223 11519 13229
rect 11081 13206 11087 13223
rect 11513 13206 11519 13223
rect 11081 13200 11519 13206
rect 11631 13229 11664 13231
rect 12036 13237 12077 13264
rect 12094 13237 12100 13663
rect 12036 13231 12100 13237
rect 12150 13663 12650 13669
rect 12150 13237 12156 13663
rect 12173 13615 12627 13663
rect 12173 13285 12235 13615
rect 12565 13285 12627 13615
rect 12173 13237 12627 13285
rect 12644 13237 12650 13663
rect 12150 13231 12650 13237
rect 12700 13663 12729 13669
rect 12700 13237 12706 13663
rect 12723 13264 12729 13663
rect 13171 13663 13200 13669
rect 13171 13264 13177 13663
rect 12723 13237 12764 13264
rect 12700 13231 12764 13237
rect 12036 13229 12069 13231
rect 11631 13223 12069 13229
rect 11631 13206 11637 13223
rect 12063 13206 12069 13223
rect 11631 13200 12069 13206
rect 12179 13229 12621 13231
rect 12181 13223 12619 13229
rect 12181 13206 12187 13223
rect 12613 13206 12619 13223
rect 12181 13200 12619 13206
rect 12731 13229 12764 13231
rect 13136 13237 13177 13264
rect 13194 13237 13200 13663
rect 13136 13231 13200 13237
rect 13250 13663 13721 13669
rect 13250 13237 13256 13663
rect 13273 13615 13721 13663
rect 13273 13285 13335 13615
rect 13665 13285 13721 13615
rect 13273 13237 13721 13285
rect 13250 13231 13721 13237
rect 13136 13229 13169 13231
rect 12731 13223 13169 13229
rect 12731 13206 12737 13223
rect 13163 13206 13169 13223
rect 12731 13200 13169 13206
rect 13279 13229 13721 13231
rect 13281 13223 13719 13229
rect 13281 13206 13287 13223
rect 13713 13206 13719 13223
rect 13281 13200 13719 13206
rect -469 13144 -31 13150
rect -469 13127 -463 13144
rect -37 13127 -31 13144
rect -469 13121 -31 13127
rect -471 13119 -29 13121
rect 81 13144 519 13150
rect 81 13127 87 13144
rect 513 13127 519 13144
rect 81 13121 519 13127
rect 81 13119 114 13121
rect -471 13113 0 13119
rect -471 13065 -23 13113
rect -471 12735 -415 13065
rect -85 12735 -23 13065
rect -471 12687 -23 12735
rect -6 12687 0 13113
rect -471 12681 0 12687
rect 50 13113 114 13119
rect 50 12687 56 13113
rect 73 13086 114 13113
rect 486 13119 519 13121
rect 631 13144 1069 13150
rect 631 13127 637 13144
rect 1063 13127 1069 13144
rect 631 13121 1069 13127
rect 629 13119 1071 13121
rect 1181 13144 1619 13150
rect 1181 13127 1187 13144
rect 1613 13127 1619 13144
rect 1181 13121 1619 13127
rect 1181 13119 1214 13121
rect 486 13113 550 13119
rect 486 13086 527 13113
rect 73 12714 79 13086
rect 521 12714 527 13086
rect 73 12687 114 12714
rect 50 12681 114 12687
rect -471 12679 -29 12681
rect -469 12673 -31 12679
rect -469 12656 -463 12673
rect -37 12656 -31 12673
rect -469 12650 -31 12656
rect 81 12679 114 12681
rect 486 12687 527 12714
rect 544 12687 550 13113
rect 486 12681 550 12687
rect 600 13113 1100 13119
rect 600 12687 606 13113
rect 623 13065 1077 13113
rect 623 12735 685 13065
rect 1015 12735 1077 13065
rect 623 12687 1077 12735
rect 1094 12687 1100 13113
rect 600 12681 1100 12687
rect 1150 13113 1214 13119
rect 1150 12687 1156 13113
rect 1173 13086 1214 13113
rect 1586 13119 1619 13121
rect 1731 13144 2169 13150
rect 1731 13127 1737 13144
rect 2163 13127 2169 13144
rect 1731 13121 2169 13127
rect 1729 13119 2171 13121
rect 2281 13144 2719 13150
rect 2281 13127 2287 13144
rect 2713 13127 2719 13144
rect 2281 13121 2719 13127
rect 2281 13119 2314 13121
rect 1586 13113 1650 13119
rect 1586 13086 1627 13113
rect 1173 12714 1179 13086
rect 1621 12714 1627 13086
rect 1173 12687 1214 12714
rect 1150 12681 1214 12687
rect 486 12679 519 12681
rect 81 12673 519 12679
rect 81 12656 87 12673
rect 513 12656 519 12673
rect 81 12650 519 12656
rect 629 12679 1071 12681
rect 631 12673 1069 12679
rect 631 12656 637 12673
rect 1063 12656 1069 12673
rect 631 12650 1069 12656
rect 1181 12679 1214 12681
rect 1586 12687 1627 12714
rect 1644 12687 1650 13113
rect 1586 12681 1650 12687
rect 1700 13113 2200 13119
rect 1700 12687 1706 13113
rect 1723 13065 2177 13113
rect 1723 12735 1785 13065
rect 2115 12735 2177 13065
rect 1723 12687 2177 12735
rect 2194 12687 2200 13113
rect 1700 12681 2200 12687
rect 2250 13113 2314 13119
rect 2250 12687 2256 13113
rect 2273 13086 2314 13113
rect 2686 13119 2719 13121
rect 2831 13144 3269 13150
rect 2831 13127 2837 13144
rect 3263 13127 3269 13144
rect 2831 13121 3269 13127
rect 2829 13119 3271 13121
rect 3381 13144 3819 13150
rect 3381 13127 3387 13144
rect 3813 13127 3819 13144
rect 3381 13121 3819 13127
rect 3381 13119 3414 13121
rect 2686 13113 2750 13119
rect 2686 13086 2727 13113
rect 2273 12714 2279 13086
rect 2721 12714 2727 13086
rect 2273 12687 2314 12714
rect 2250 12681 2314 12687
rect 1586 12679 1619 12681
rect 1181 12673 1619 12679
rect 1181 12656 1187 12673
rect 1613 12656 1619 12673
rect 1181 12650 1619 12656
rect 1729 12679 2171 12681
rect 1731 12673 2169 12679
rect 1731 12656 1737 12673
rect 2163 12656 2169 12673
rect 1731 12650 2169 12656
rect 2281 12679 2314 12681
rect 2686 12687 2727 12714
rect 2744 12687 2750 13113
rect 2686 12681 2750 12687
rect 2800 13113 3300 13119
rect 2800 12687 2806 13113
rect 2823 13065 3277 13113
rect 2823 12735 2885 13065
rect 3215 12735 3277 13065
rect 2823 12687 3277 12735
rect 3294 12687 3300 13113
rect 2800 12681 3300 12687
rect 3350 13113 3414 13119
rect 3350 12687 3356 13113
rect 3373 13086 3414 13113
rect 3786 13119 3819 13121
rect 3931 13144 4369 13150
rect 3931 13127 3937 13144
rect 4363 13127 4369 13144
rect 3931 13121 4369 13127
rect 3929 13119 4371 13121
rect 4481 13144 4919 13150
rect 4481 13127 4487 13144
rect 4913 13127 4919 13144
rect 4481 13121 4919 13127
rect 4481 13119 4514 13121
rect 3786 13113 3850 13119
rect 3786 13086 3827 13113
rect 3373 12714 3379 13086
rect 3821 12714 3827 13086
rect 3373 12687 3414 12714
rect 3350 12681 3414 12687
rect 2686 12679 2719 12681
rect 2281 12673 2719 12679
rect 2281 12656 2287 12673
rect 2713 12656 2719 12673
rect 2281 12650 2719 12656
rect 2829 12679 3271 12681
rect 2831 12673 3269 12679
rect 2831 12656 2837 12673
rect 3263 12656 3269 12673
rect 2831 12650 3269 12656
rect 3381 12679 3414 12681
rect 3786 12687 3827 12714
rect 3844 12687 3850 13113
rect 3786 12681 3850 12687
rect 3900 13113 4400 13119
rect 3900 12687 3906 13113
rect 3923 13065 4377 13113
rect 3923 12735 3985 13065
rect 4315 12735 4377 13065
rect 3923 12687 4377 12735
rect 4394 12687 4400 13113
rect 3900 12681 4400 12687
rect 4450 13113 4514 13119
rect 4450 12687 4456 13113
rect 4473 13086 4514 13113
rect 4886 13119 4919 13121
rect 5031 13144 5469 13150
rect 5031 13127 5037 13144
rect 5463 13127 5469 13144
rect 5031 13121 5469 13127
rect 5029 13119 5471 13121
rect 5581 13144 6019 13150
rect 5581 13127 5587 13144
rect 6013 13127 6019 13144
rect 5581 13121 6019 13127
rect 5581 13119 5614 13121
rect 4886 13113 4950 13119
rect 4886 13086 4927 13113
rect 4473 12714 4479 13086
rect 4921 12714 4927 13086
rect 4473 12687 4514 12714
rect 4450 12681 4514 12687
rect 3786 12679 3819 12681
rect 3381 12673 3819 12679
rect 3381 12656 3387 12673
rect 3813 12656 3819 12673
rect 3381 12650 3819 12656
rect 3929 12679 4371 12681
rect 3931 12673 4369 12679
rect 3931 12656 3937 12673
rect 4363 12656 4369 12673
rect 3931 12650 4369 12656
rect 4481 12679 4514 12681
rect 4886 12687 4927 12714
rect 4944 12687 4950 13113
rect 4886 12681 4950 12687
rect 5000 13113 5500 13119
rect 5000 12687 5006 13113
rect 5023 13065 5477 13113
rect 5023 12735 5085 13065
rect 5415 12735 5477 13065
rect 5023 12687 5477 12735
rect 5494 12687 5500 13113
rect 5000 12681 5500 12687
rect 5550 13113 5614 13119
rect 5550 12687 5556 13113
rect 5573 13086 5614 13113
rect 5986 13119 6019 13121
rect 6131 13144 6569 13150
rect 6131 13127 6137 13144
rect 6563 13127 6569 13144
rect 6131 13121 6569 13127
rect 6129 13119 6571 13121
rect 6681 13144 7119 13150
rect 6681 13127 6687 13144
rect 7113 13127 7119 13144
rect 6681 13121 7119 13127
rect 6681 13119 6714 13121
rect 5986 13113 6050 13119
rect 5986 13086 6027 13113
rect 5573 12714 5579 13086
rect 6021 12714 6027 13086
rect 5573 12687 5614 12714
rect 5550 12681 5614 12687
rect 4886 12679 4919 12681
rect 4481 12673 4919 12679
rect 4481 12656 4487 12673
rect 4913 12656 4919 12673
rect 4481 12650 4919 12656
rect 5029 12679 5471 12681
rect 5031 12673 5469 12679
rect 5031 12656 5037 12673
rect 5463 12656 5469 12673
rect 5031 12650 5469 12656
rect 5581 12679 5614 12681
rect 5986 12687 6027 12714
rect 6044 12687 6050 13113
rect 5986 12681 6050 12687
rect 6100 13113 6600 13119
rect 6100 12687 6106 13113
rect 6123 13065 6577 13113
rect 6123 12735 6185 13065
rect 6515 12735 6577 13065
rect 6123 12687 6577 12735
rect 6594 12687 6600 13113
rect 6100 12681 6600 12687
rect 6650 13113 6714 13119
rect 6650 12687 6656 13113
rect 6673 13086 6714 13113
rect 7086 13119 7119 13121
rect 7231 13144 7669 13150
rect 7231 13127 7237 13144
rect 7663 13127 7669 13144
rect 7231 13121 7669 13127
rect 7229 13119 7671 13121
rect 7781 13144 8219 13150
rect 7781 13127 7787 13144
rect 8213 13127 8219 13144
rect 7781 13121 8219 13127
rect 7781 13119 7814 13121
rect 7086 13113 7150 13119
rect 7086 13086 7127 13113
rect 6673 12714 6679 13086
rect 7121 12714 7127 13086
rect 6673 12687 6714 12714
rect 6650 12681 6714 12687
rect 5986 12679 6019 12681
rect 5581 12673 6019 12679
rect 5581 12656 5587 12673
rect 6013 12656 6019 12673
rect 5581 12650 6019 12656
rect 6129 12679 6571 12681
rect 6131 12673 6569 12679
rect 6131 12656 6137 12673
rect 6563 12656 6569 12673
rect 6131 12650 6569 12656
rect 6681 12679 6714 12681
rect 7086 12687 7127 12714
rect 7144 12687 7150 13113
rect 7086 12681 7150 12687
rect 7200 13113 7700 13119
rect 7200 12687 7206 13113
rect 7223 13065 7677 13113
rect 7223 12735 7285 13065
rect 7615 12735 7677 13065
rect 7223 12687 7677 12735
rect 7694 12687 7700 13113
rect 7200 12681 7700 12687
rect 7750 13113 7814 13119
rect 7750 12687 7756 13113
rect 7773 13086 7814 13113
rect 8186 13119 8219 13121
rect 8331 13144 8769 13150
rect 8331 13127 8337 13144
rect 8763 13127 8769 13144
rect 8331 13121 8769 13127
rect 8329 13119 8771 13121
rect 8881 13144 9319 13150
rect 8881 13127 8887 13144
rect 9313 13127 9319 13144
rect 8881 13121 9319 13127
rect 8881 13119 8914 13121
rect 8186 13113 8250 13119
rect 8186 13086 8227 13113
rect 7773 12714 7779 13086
rect 8221 12714 8227 13086
rect 7773 12687 7814 12714
rect 7750 12681 7814 12687
rect 7086 12679 7119 12681
rect 6681 12673 7119 12679
rect 6681 12656 6687 12673
rect 7113 12656 7119 12673
rect 6681 12650 7119 12656
rect 7229 12679 7671 12681
rect 7231 12673 7669 12679
rect 7231 12656 7237 12673
rect 7663 12656 7669 12673
rect 7231 12650 7669 12656
rect 7781 12679 7814 12681
rect 8186 12687 8227 12714
rect 8244 12687 8250 13113
rect 8186 12681 8250 12687
rect 8300 13113 8800 13119
rect 8300 12687 8306 13113
rect 8323 13065 8777 13113
rect 8323 12735 8385 13065
rect 8715 12735 8777 13065
rect 8323 12687 8777 12735
rect 8794 12687 8800 13113
rect 8300 12681 8800 12687
rect 8850 13113 8914 13119
rect 8850 12687 8856 13113
rect 8873 13086 8914 13113
rect 9286 13119 9319 13121
rect 9431 13144 9869 13150
rect 9431 13127 9437 13144
rect 9863 13127 9869 13144
rect 9431 13121 9869 13127
rect 9429 13119 9871 13121
rect 9981 13144 10419 13150
rect 9981 13127 9987 13144
rect 10413 13127 10419 13144
rect 9981 13121 10419 13127
rect 9981 13119 10014 13121
rect 9286 13113 9350 13119
rect 9286 13086 9327 13113
rect 8873 12714 8879 13086
rect 9321 12714 9327 13086
rect 8873 12687 8914 12714
rect 8850 12681 8914 12687
rect 8186 12679 8219 12681
rect 7781 12673 8219 12679
rect 7781 12656 7787 12673
rect 8213 12656 8219 12673
rect 7781 12650 8219 12656
rect 8329 12679 8771 12681
rect 8331 12673 8769 12679
rect 8331 12656 8337 12673
rect 8763 12656 8769 12673
rect 8331 12650 8769 12656
rect 8881 12679 8914 12681
rect 9286 12687 9327 12714
rect 9344 12687 9350 13113
rect 9286 12681 9350 12687
rect 9400 13113 9900 13119
rect 9400 12687 9406 13113
rect 9423 13065 9877 13113
rect 9423 12735 9485 13065
rect 9815 12735 9877 13065
rect 9423 12687 9877 12735
rect 9894 12687 9900 13113
rect 9400 12681 9900 12687
rect 9950 13113 10014 13119
rect 9950 12687 9956 13113
rect 9973 13086 10014 13113
rect 10386 13119 10419 13121
rect 10531 13144 10969 13150
rect 10531 13127 10537 13144
rect 10963 13127 10969 13144
rect 10531 13121 10969 13127
rect 10529 13119 10971 13121
rect 11081 13144 11519 13150
rect 11081 13127 11087 13144
rect 11513 13127 11519 13144
rect 11081 13121 11519 13127
rect 11081 13119 11114 13121
rect 10386 13113 10450 13119
rect 10386 13086 10427 13113
rect 9973 12714 9979 13086
rect 10421 12714 10427 13086
rect 9973 12687 10014 12714
rect 9950 12681 10014 12687
rect 9286 12679 9319 12681
rect 8881 12673 9319 12679
rect 8881 12656 8887 12673
rect 9313 12656 9319 12673
rect 8881 12650 9319 12656
rect 9429 12679 9871 12681
rect 9431 12673 9869 12679
rect 9431 12656 9437 12673
rect 9863 12656 9869 12673
rect 9431 12650 9869 12656
rect 9981 12679 10014 12681
rect 10386 12687 10427 12714
rect 10444 12687 10450 13113
rect 10386 12681 10450 12687
rect 10500 13113 11000 13119
rect 10500 12687 10506 13113
rect 10523 13065 10977 13113
rect 10523 12735 10585 13065
rect 10915 12735 10977 13065
rect 10523 12687 10977 12735
rect 10994 12687 11000 13113
rect 10500 12681 11000 12687
rect 11050 13113 11114 13119
rect 11050 12687 11056 13113
rect 11073 13086 11114 13113
rect 11486 13119 11519 13121
rect 11631 13144 12069 13150
rect 11631 13127 11637 13144
rect 12063 13127 12069 13144
rect 11631 13121 12069 13127
rect 11629 13119 12071 13121
rect 12181 13144 12619 13150
rect 12181 13127 12187 13144
rect 12613 13127 12619 13144
rect 12181 13121 12619 13127
rect 12181 13119 12214 13121
rect 11486 13113 11550 13119
rect 11486 13086 11527 13113
rect 11073 12714 11079 13086
rect 11521 12714 11527 13086
rect 11073 12687 11114 12714
rect 11050 12681 11114 12687
rect 10386 12679 10419 12681
rect 9981 12673 10419 12679
rect 9981 12656 9987 12673
rect 10413 12656 10419 12673
rect 9981 12650 10419 12656
rect 10529 12679 10971 12681
rect 10531 12673 10969 12679
rect 10531 12656 10537 12673
rect 10963 12656 10969 12673
rect 10531 12650 10969 12656
rect 11081 12679 11114 12681
rect 11486 12687 11527 12714
rect 11544 12687 11550 13113
rect 11486 12681 11550 12687
rect 11600 13113 12100 13119
rect 11600 12687 11606 13113
rect 11623 13065 12077 13113
rect 11623 12735 11685 13065
rect 12015 12735 12077 13065
rect 11623 12687 12077 12735
rect 12094 12687 12100 13113
rect 11600 12681 12100 12687
rect 12150 13113 12214 13119
rect 12150 12687 12156 13113
rect 12173 13086 12214 13113
rect 12586 13119 12619 13121
rect 12731 13144 13169 13150
rect 12731 13127 12737 13144
rect 13163 13127 13169 13144
rect 12731 13121 13169 13127
rect 12729 13119 13171 13121
rect 13281 13144 13719 13150
rect 13281 13127 13287 13144
rect 13713 13127 13719 13144
rect 13281 13121 13719 13127
rect 13281 13119 13314 13121
rect 12586 13113 12650 13119
rect 12586 13086 12627 13113
rect 12173 12714 12179 13086
rect 12621 12714 12627 13086
rect 12173 12687 12214 12714
rect 12150 12681 12214 12687
rect 11486 12679 11519 12681
rect 11081 12673 11519 12679
rect 11081 12656 11087 12673
rect 11513 12656 11519 12673
rect 11081 12650 11519 12656
rect 11629 12679 12071 12681
rect 11631 12673 12069 12679
rect 11631 12656 11637 12673
rect 12063 12656 12069 12673
rect 11631 12650 12069 12656
rect 12181 12679 12214 12681
rect 12586 12687 12627 12714
rect 12644 12687 12650 13113
rect 12586 12681 12650 12687
rect 12700 13113 13200 13119
rect 12700 12687 12706 13113
rect 12723 13065 13177 13113
rect 12723 12735 12785 13065
rect 13115 12735 13177 13065
rect 12723 12687 13177 12735
rect 13194 12687 13200 13113
rect 12700 12681 13200 12687
rect 13250 13113 13314 13119
rect 13250 12687 13256 13113
rect 13273 13086 13314 13113
rect 13273 12714 13279 13086
rect 13273 12687 13314 12714
rect 13250 12681 13314 12687
rect 12586 12679 12619 12681
rect 12181 12673 12619 12679
rect 12181 12656 12187 12673
rect 12613 12656 12619 12673
rect 12181 12650 12619 12656
rect 12729 12679 13171 12681
rect 12731 12673 13169 12679
rect 12731 12656 12737 12673
rect 13163 12656 13169 12673
rect 12731 12650 13169 12656
rect 13281 12679 13314 12681
rect 13281 12673 13719 12679
rect 13281 12656 13287 12673
rect 13713 12656 13719 12673
rect 13281 12650 13719 12656
rect -469 12594 -31 12600
rect -469 12577 -463 12594
rect -37 12577 -31 12594
rect -469 12571 -31 12577
rect -64 12569 -31 12571
rect 81 12594 519 12600
rect 81 12577 87 12594
rect 513 12577 519 12594
rect 81 12571 519 12577
rect 79 12569 521 12571
rect 631 12594 1069 12600
rect 631 12577 637 12594
rect 1063 12577 1069 12594
rect 631 12571 1069 12577
rect 631 12569 664 12571
rect -64 12563 0 12569
rect -64 12536 -23 12563
rect -29 12164 -23 12536
rect -64 12137 -23 12164
rect -6 12137 0 12563
rect -64 12131 0 12137
rect 50 12563 550 12569
rect 50 12137 56 12563
rect 73 12515 527 12563
rect 73 12185 135 12515
rect 465 12185 527 12515
rect 73 12137 527 12185
rect 544 12137 550 12563
rect 50 12131 550 12137
rect 600 12563 664 12569
rect 600 12137 606 12563
rect 623 12536 664 12563
rect 1036 12569 1069 12571
rect 1181 12594 1619 12600
rect 1181 12577 1187 12594
rect 1613 12577 1619 12594
rect 1181 12571 1619 12577
rect 1179 12569 1621 12571
rect 1731 12594 2169 12600
rect 1731 12577 1737 12594
rect 2163 12577 2169 12594
rect 1731 12571 2169 12577
rect 1731 12569 1764 12571
rect 1036 12563 1100 12569
rect 1036 12536 1077 12563
rect 623 12164 629 12536
rect 1071 12164 1077 12536
rect 623 12137 664 12164
rect 600 12131 664 12137
rect -64 12129 -31 12131
rect -469 12123 -31 12129
rect -469 12106 -463 12123
rect -37 12106 -31 12123
rect -469 12100 -31 12106
rect 79 12129 521 12131
rect 81 12123 519 12129
rect 81 12106 87 12123
rect 513 12106 519 12123
rect 81 12100 519 12106
rect 631 12129 664 12131
rect 1036 12137 1077 12164
rect 1094 12137 1100 12563
rect 1036 12131 1100 12137
rect 1150 12563 1650 12569
rect 1150 12137 1156 12563
rect 1173 12515 1627 12563
rect 1173 12185 1235 12515
rect 1565 12185 1627 12515
rect 1173 12137 1627 12185
rect 1644 12137 1650 12563
rect 1150 12131 1650 12137
rect 1700 12563 1764 12569
rect 1700 12137 1706 12563
rect 1723 12536 1764 12563
rect 2136 12569 2169 12571
rect 2281 12594 2719 12600
rect 2281 12577 2287 12594
rect 2713 12577 2719 12594
rect 2281 12571 2719 12577
rect 2279 12569 2721 12571
rect 2831 12594 3269 12600
rect 2831 12577 2837 12594
rect 3263 12577 3269 12594
rect 2831 12571 3269 12577
rect 2831 12569 2864 12571
rect 2136 12563 2200 12569
rect 2136 12536 2177 12563
rect 1723 12164 1729 12536
rect 2171 12164 2177 12536
rect 1723 12137 1764 12164
rect 1700 12131 1764 12137
rect 1036 12129 1069 12131
rect 631 12123 1069 12129
rect 631 12106 637 12123
rect 1063 12106 1069 12123
rect 631 12100 1069 12106
rect 1179 12129 1621 12131
rect 1181 12123 1619 12129
rect 1181 12106 1187 12123
rect 1613 12106 1619 12123
rect 1181 12100 1619 12106
rect 1731 12129 1764 12131
rect 2136 12137 2177 12164
rect 2194 12137 2200 12563
rect 2136 12131 2200 12137
rect 2250 12563 2750 12569
rect 2250 12137 2256 12563
rect 2273 12515 2727 12563
rect 2273 12185 2335 12515
rect 2665 12185 2727 12515
rect 2273 12137 2727 12185
rect 2744 12137 2750 12563
rect 2250 12131 2750 12137
rect 2800 12563 2864 12569
rect 2800 12137 2806 12563
rect 2823 12536 2864 12563
rect 3236 12569 3269 12571
rect 3381 12594 3819 12600
rect 3381 12577 3387 12594
rect 3813 12577 3819 12594
rect 3381 12571 3819 12577
rect 3379 12569 3821 12571
rect 3931 12594 4369 12600
rect 3931 12577 3937 12594
rect 4363 12577 4369 12594
rect 3931 12571 4369 12577
rect 3931 12569 3964 12571
rect 3236 12563 3300 12569
rect 3236 12536 3277 12563
rect 2823 12164 2829 12536
rect 3271 12164 3277 12536
rect 2823 12137 2864 12164
rect 2800 12131 2864 12137
rect 2136 12129 2169 12131
rect 1731 12123 2169 12129
rect 1731 12106 1737 12123
rect 2163 12106 2169 12123
rect 1731 12100 2169 12106
rect 2279 12129 2721 12131
rect 2281 12123 2719 12129
rect 2281 12106 2287 12123
rect 2713 12106 2719 12123
rect 2281 12100 2719 12106
rect 2831 12129 2864 12131
rect 3236 12137 3277 12164
rect 3294 12137 3300 12563
rect 3236 12131 3300 12137
rect 3350 12563 3850 12569
rect 3350 12137 3356 12563
rect 3373 12515 3827 12563
rect 3373 12185 3435 12515
rect 3765 12185 3827 12515
rect 3373 12137 3827 12185
rect 3844 12137 3850 12563
rect 3350 12131 3850 12137
rect 3900 12563 3964 12569
rect 3900 12137 3906 12563
rect 3923 12536 3964 12563
rect 4336 12569 4369 12571
rect 4481 12594 4919 12600
rect 4481 12577 4487 12594
rect 4913 12577 4919 12594
rect 4481 12571 4919 12577
rect 4479 12569 4921 12571
rect 5031 12594 5469 12600
rect 5031 12577 5037 12594
rect 5463 12577 5469 12594
rect 5031 12571 5469 12577
rect 5031 12569 5064 12571
rect 4336 12563 4400 12569
rect 4336 12536 4377 12563
rect 3923 12164 3929 12536
rect 4371 12164 4377 12536
rect 3923 12137 3964 12164
rect 3900 12131 3964 12137
rect 3236 12129 3269 12131
rect 2831 12123 3269 12129
rect 2831 12106 2837 12123
rect 3263 12106 3269 12123
rect 2831 12100 3269 12106
rect 3379 12129 3821 12131
rect 3381 12123 3819 12129
rect 3381 12106 3387 12123
rect 3813 12106 3819 12123
rect 3381 12100 3819 12106
rect 3931 12129 3964 12131
rect 4336 12137 4377 12164
rect 4394 12137 4400 12563
rect 4336 12131 4400 12137
rect 4450 12563 4950 12569
rect 4450 12137 4456 12563
rect 4473 12515 4927 12563
rect 4473 12185 4535 12515
rect 4865 12185 4927 12515
rect 4473 12137 4927 12185
rect 4944 12137 4950 12563
rect 4450 12131 4950 12137
rect 5000 12563 5064 12569
rect 5000 12137 5006 12563
rect 5023 12536 5064 12563
rect 5436 12569 5469 12571
rect 5581 12594 6019 12600
rect 5581 12577 5587 12594
rect 6013 12577 6019 12594
rect 5581 12571 6019 12577
rect 5579 12569 6021 12571
rect 6131 12594 6569 12600
rect 6131 12577 6137 12594
rect 6563 12577 6569 12594
rect 6131 12571 6569 12577
rect 6131 12569 6164 12571
rect 5436 12563 5500 12569
rect 5436 12536 5477 12563
rect 5023 12164 5029 12536
rect 5471 12164 5477 12536
rect 5023 12137 5064 12164
rect 5000 12131 5064 12137
rect 4336 12129 4369 12131
rect 3931 12123 4369 12129
rect 3931 12106 3937 12123
rect 4363 12106 4369 12123
rect 3931 12100 4369 12106
rect 4479 12129 4921 12131
rect 4481 12123 4919 12129
rect 4481 12106 4487 12123
rect 4913 12106 4919 12123
rect 4481 12100 4919 12106
rect 5031 12129 5064 12131
rect 5436 12137 5477 12164
rect 5494 12137 5500 12563
rect 5436 12131 5500 12137
rect 5550 12563 6050 12569
rect 5550 12137 5556 12563
rect 5573 12515 6027 12563
rect 5573 12185 5635 12515
rect 5965 12185 6027 12515
rect 5573 12137 6027 12185
rect 6044 12137 6050 12563
rect 5550 12131 6050 12137
rect 6100 12563 6164 12569
rect 6100 12137 6106 12563
rect 6123 12536 6164 12563
rect 6536 12569 6569 12571
rect 6681 12594 7119 12600
rect 6681 12577 6687 12594
rect 7113 12577 7119 12594
rect 6681 12571 7119 12577
rect 6679 12569 7121 12571
rect 7231 12594 7669 12600
rect 7231 12577 7237 12594
rect 7663 12577 7669 12594
rect 7231 12571 7669 12577
rect 7231 12569 7264 12571
rect 6536 12563 6600 12569
rect 6536 12536 6577 12563
rect 6123 12164 6129 12536
rect 6571 12164 6577 12536
rect 6123 12137 6164 12164
rect 6100 12131 6164 12137
rect 5436 12129 5469 12131
rect 5031 12123 5469 12129
rect 5031 12106 5037 12123
rect 5463 12106 5469 12123
rect 5031 12100 5469 12106
rect 5579 12129 6021 12131
rect 5581 12123 6019 12129
rect 5581 12106 5587 12123
rect 6013 12106 6019 12123
rect 5581 12100 6019 12106
rect 6131 12129 6164 12131
rect 6536 12137 6577 12164
rect 6594 12137 6600 12563
rect 6536 12131 6600 12137
rect 6650 12563 7150 12569
rect 6650 12137 6656 12563
rect 6673 12515 7127 12563
rect 6673 12185 6735 12515
rect 7065 12185 7127 12515
rect 6673 12137 7127 12185
rect 7144 12137 7150 12563
rect 6650 12131 7150 12137
rect 7200 12563 7264 12569
rect 7200 12137 7206 12563
rect 7223 12536 7264 12563
rect 7636 12569 7669 12571
rect 7781 12594 8219 12600
rect 7781 12577 7787 12594
rect 8213 12577 8219 12594
rect 7781 12571 8219 12577
rect 7779 12569 8221 12571
rect 8331 12594 8769 12600
rect 8331 12577 8337 12594
rect 8763 12577 8769 12594
rect 8331 12571 8769 12577
rect 8331 12569 8364 12571
rect 7636 12563 7700 12569
rect 7636 12536 7677 12563
rect 7223 12164 7229 12536
rect 7671 12164 7677 12536
rect 7223 12137 7264 12164
rect 7200 12131 7264 12137
rect 6536 12129 6569 12131
rect 6131 12123 6569 12129
rect 6131 12106 6137 12123
rect 6563 12106 6569 12123
rect 6131 12100 6569 12106
rect 6679 12129 7121 12131
rect 6681 12123 7119 12129
rect 6681 12106 6687 12123
rect 7113 12106 7119 12123
rect 6681 12100 7119 12106
rect 7231 12129 7264 12131
rect 7636 12137 7677 12164
rect 7694 12137 7700 12563
rect 7636 12131 7700 12137
rect 7750 12563 8250 12569
rect 7750 12137 7756 12563
rect 7773 12515 8227 12563
rect 7773 12185 7835 12515
rect 8165 12185 8227 12515
rect 7773 12137 8227 12185
rect 8244 12137 8250 12563
rect 7750 12131 8250 12137
rect 8300 12563 8364 12569
rect 8300 12137 8306 12563
rect 8323 12536 8364 12563
rect 8736 12569 8769 12571
rect 8881 12594 9319 12600
rect 8881 12577 8887 12594
rect 9313 12577 9319 12594
rect 8881 12571 9319 12577
rect 8879 12569 9321 12571
rect 9431 12594 9869 12600
rect 9431 12577 9437 12594
rect 9863 12577 9869 12594
rect 9431 12571 9869 12577
rect 9431 12569 9464 12571
rect 8736 12563 8800 12569
rect 8736 12536 8777 12563
rect 8323 12164 8329 12536
rect 8771 12164 8777 12536
rect 8323 12137 8364 12164
rect 8300 12131 8364 12137
rect 7636 12129 7669 12131
rect 7231 12123 7669 12129
rect 7231 12106 7237 12123
rect 7663 12106 7669 12123
rect 7231 12100 7669 12106
rect 7779 12129 8221 12131
rect 7781 12123 8219 12129
rect 7781 12106 7787 12123
rect 8213 12106 8219 12123
rect 7781 12100 8219 12106
rect 8331 12129 8364 12131
rect 8736 12137 8777 12164
rect 8794 12137 8800 12563
rect 8736 12131 8800 12137
rect 8850 12563 9350 12569
rect 8850 12137 8856 12563
rect 8873 12515 9327 12563
rect 8873 12185 8935 12515
rect 9265 12185 9327 12515
rect 8873 12137 9327 12185
rect 9344 12137 9350 12563
rect 8850 12131 9350 12137
rect 9400 12563 9464 12569
rect 9400 12137 9406 12563
rect 9423 12536 9464 12563
rect 9836 12569 9869 12571
rect 9981 12594 10419 12600
rect 9981 12577 9987 12594
rect 10413 12577 10419 12594
rect 9981 12571 10419 12577
rect 9979 12569 10421 12571
rect 10531 12594 10969 12600
rect 10531 12577 10537 12594
rect 10963 12577 10969 12594
rect 10531 12571 10969 12577
rect 10531 12569 10564 12571
rect 9836 12563 9900 12569
rect 9836 12536 9877 12563
rect 9423 12164 9429 12536
rect 9871 12164 9877 12536
rect 9423 12137 9464 12164
rect 9400 12131 9464 12137
rect 8736 12129 8769 12131
rect 8331 12123 8769 12129
rect 8331 12106 8337 12123
rect 8763 12106 8769 12123
rect 8331 12100 8769 12106
rect 8879 12129 9321 12131
rect 8881 12123 9319 12129
rect 8881 12106 8887 12123
rect 9313 12106 9319 12123
rect 8881 12100 9319 12106
rect 9431 12129 9464 12131
rect 9836 12137 9877 12164
rect 9894 12137 9900 12563
rect 9836 12131 9900 12137
rect 9950 12563 10450 12569
rect 9950 12137 9956 12563
rect 9973 12515 10427 12563
rect 9973 12185 10035 12515
rect 10365 12185 10427 12515
rect 9973 12137 10427 12185
rect 10444 12137 10450 12563
rect 9950 12131 10450 12137
rect 10500 12563 10564 12569
rect 10500 12137 10506 12563
rect 10523 12536 10564 12563
rect 10936 12569 10969 12571
rect 11081 12594 11519 12600
rect 11081 12577 11087 12594
rect 11513 12577 11519 12594
rect 11081 12571 11519 12577
rect 11079 12569 11521 12571
rect 11631 12594 12069 12600
rect 11631 12577 11637 12594
rect 12063 12577 12069 12594
rect 11631 12571 12069 12577
rect 11631 12569 11664 12571
rect 10936 12563 11000 12569
rect 10936 12536 10977 12563
rect 10523 12164 10529 12536
rect 10971 12164 10977 12536
rect 10523 12137 10564 12164
rect 10500 12131 10564 12137
rect 9836 12129 9869 12131
rect 9431 12123 9869 12129
rect 9431 12106 9437 12123
rect 9863 12106 9869 12123
rect 9431 12100 9869 12106
rect 9979 12129 10421 12131
rect 9981 12123 10419 12129
rect 9981 12106 9987 12123
rect 10413 12106 10419 12123
rect 9981 12100 10419 12106
rect 10531 12129 10564 12131
rect 10936 12137 10977 12164
rect 10994 12137 11000 12563
rect 10936 12131 11000 12137
rect 11050 12563 11550 12569
rect 11050 12137 11056 12563
rect 11073 12515 11527 12563
rect 11073 12185 11135 12515
rect 11465 12185 11527 12515
rect 11073 12137 11527 12185
rect 11544 12137 11550 12563
rect 11050 12131 11550 12137
rect 11600 12563 11664 12569
rect 11600 12137 11606 12563
rect 11623 12536 11664 12563
rect 12036 12569 12069 12571
rect 12181 12594 12619 12600
rect 12181 12577 12187 12594
rect 12613 12577 12619 12594
rect 12181 12571 12619 12577
rect 12179 12569 12621 12571
rect 12731 12594 13169 12600
rect 12731 12577 12737 12594
rect 13163 12577 13169 12594
rect 12731 12571 13169 12577
rect 12731 12569 12764 12571
rect 12036 12563 12100 12569
rect 12036 12536 12077 12563
rect 11623 12164 11629 12536
rect 12071 12164 12077 12536
rect 11623 12137 11664 12164
rect 11600 12131 11664 12137
rect 10936 12129 10969 12131
rect 10531 12123 10969 12129
rect 10531 12106 10537 12123
rect 10963 12106 10969 12123
rect 10531 12100 10969 12106
rect 11079 12129 11521 12131
rect 11081 12123 11519 12129
rect 11081 12106 11087 12123
rect 11513 12106 11519 12123
rect 11081 12100 11519 12106
rect 11631 12129 11664 12131
rect 12036 12137 12077 12164
rect 12094 12137 12100 12563
rect 12036 12131 12100 12137
rect 12150 12563 12650 12569
rect 12150 12137 12156 12563
rect 12173 12515 12627 12563
rect 12173 12185 12235 12515
rect 12565 12185 12627 12515
rect 12173 12137 12627 12185
rect 12644 12137 12650 12563
rect 12150 12131 12650 12137
rect 12700 12563 12764 12569
rect 12700 12137 12706 12563
rect 12723 12536 12764 12563
rect 13136 12569 13169 12571
rect 13281 12594 13719 12600
rect 13281 12577 13287 12594
rect 13713 12577 13719 12594
rect 13281 12571 13719 12577
rect 13279 12569 13721 12571
rect 13136 12563 13200 12569
rect 13136 12536 13177 12563
rect 12723 12164 12729 12536
rect 13171 12164 13177 12536
rect 12723 12137 12764 12164
rect 12700 12131 12764 12137
rect 12036 12129 12069 12131
rect 11631 12123 12069 12129
rect 11631 12106 11637 12123
rect 12063 12106 12069 12123
rect 11631 12100 12069 12106
rect 12179 12129 12621 12131
rect 12181 12123 12619 12129
rect 12181 12106 12187 12123
rect 12613 12106 12619 12123
rect 12181 12100 12619 12106
rect 12731 12129 12764 12131
rect 13136 12137 13177 12164
rect 13194 12137 13200 12563
rect 13136 12131 13200 12137
rect 13250 12563 13721 12569
rect 13250 12137 13256 12563
rect 13273 12515 13721 12563
rect 13273 12185 13335 12515
rect 13665 12185 13721 12515
rect 13273 12137 13721 12185
rect 13250 12131 13721 12137
rect 13136 12129 13169 12131
rect 12731 12123 13169 12129
rect 12731 12106 12737 12123
rect 13163 12106 13169 12123
rect 12731 12100 13169 12106
rect 13279 12129 13721 12131
rect 13281 12123 13719 12129
rect 13281 12106 13287 12123
rect 13713 12106 13719 12123
rect 13281 12100 13719 12106
rect -469 12044 -31 12050
rect -469 12027 -463 12044
rect -37 12027 -31 12044
rect -469 12021 -31 12027
rect -471 12019 -29 12021
rect 81 12044 519 12050
rect 81 12027 87 12044
rect 513 12027 519 12044
rect 81 12021 519 12027
rect 81 12019 114 12021
rect -471 12013 0 12019
rect -471 11965 -23 12013
rect -471 11635 -415 11965
rect -85 11635 -23 11965
rect -471 11587 -23 11635
rect -6 11587 0 12013
rect -471 11581 0 11587
rect 50 12013 114 12019
rect 50 11587 56 12013
rect 73 11986 114 12013
rect 486 12019 519 12021
rect 631 12044 1069 12050
rect 631 12027 637 12044
rect 1063 12027 1069 12044
rect 631 12021 1069 12027
rect 629 12019 1071 12021
rect 1181 12044 1619 12050
rect 1181 12027 1187 12044
rect 1613 12027 1619 12044
rect 1181 12021 1619 12027
rect 1181 12019 1214 12021
rect 486 12013 550 12019
rect 486 11986 527 12013
rect 73 11614 79 11986
rect 521 11614 527 11986
rect 73 11587 114 11614
rect 50 11581 114 11587
rect -471 11579 -29 11581
rect -469 11573 -31 11579
rect -469 11556 -463 11573
rect -37 11556 -31 11573
rect -469 11550 -31 11556
rect 81 11579 114 11581
rect 486 11587 527 11614
rect 544 11587 550 12013
rect 486 11581 550 11587
rect 600 12013 1100 12019
rect 600 11587 606 12013
rect 623 11965 1077 12013
rect 623 11635 685 11965
rect 1015 11635 1077 11965
rect 623 11587 1077 11635
rect 1094 11587 1100 12013
rect 600 11581 1100 11587
rect 1150 12013 1214 12019
rect 1150 11587 1156 12013
rect 1173 11986 1214 12013
rect 1586 12019 1619 12021
rect 1731 12044 2169 12050
rect 1731 12027 1737 12044
rect 2163 12027 2169 12044
rect 1731 12021 2169 12027
rect 1729 12019 2171 12021
rect 2281 12044 2719 12050
rect 2281 12027 2287 12044
rect 2713 12027 2719 12044
rect 2281 12021 2719 12027
rect 2281 12019 2314 12021
rect 1586 12013 1650 12019
rect 1586 11986 1627 12013
rect 1173 11614 1179 11986
rect 1621 11614 1627 11986
rect 1173 11587 1214 11614
rect 1150 11581 1214 11587
rect 486 11579 519 11581
rect 81 11573 519 11579
rect 81 11556 87 11573
rect 513 11556 519 11573
rect 81 11550 519 11556
rect 629 11579 1071 11581
rect 631 11573 1069 11579
rect 631 11556 637 11573
rect 1063 11556 1069 11573
rect 631 11550 1069 11556
rect 1181 11579 1214 11581
rect 1586 11587 1627 11614
rect 1644 11587 1650 12013
rect 1586 11581 1650 11587
rect 1700 12013 2200 12019
rect 1700 11587 1706 12013
rect 1723 11965 2177 12013
rect 1723 11635 1785 11965
rect 2115 11635 2177 11965
rect 1723 11587 2177 11635
rect 2194 11587 2200 12013
rect 1700 11581 2200 11587
rect 2250 12013 2314 12019
rect 2250 11587 2256 12013
rect 2273 11986 2314 12013
rect 2686 12019 2719 12021
rect 2831 12044 3269 12050
rect 2831 12027 2837 12044
rect 3263 12027 3269 12044
rect 2831 12021 3269 12027
rect 2829 12019 3271 12021
rect 3381 12044 3819 12050
rect 3381 12027 3387 12044
rect 3813 12027 3819 12044
rect 3381 12021 3819 12027
rect 3381 12019 3414 12021
rect 2686 12013 2750 12019
rect 2686 11986 2727 12013
rect 2273 11614 2279 11986
rect 2721 11614 2727 11986
rect 2273 11587 2314 11614
rect 2250 11581 2314 11587
rect 1586 11579 1619 11581
rect 1181 11573 1619 11579
rect 1181 11556 1187 11573
rect 1613 11556 1619 11573
rect 1181 11550 1619 11556
rect 1729 11579 2171 11581
rect 1731 11573 2169 11579
rect 1731 11556 1737 11573
rect 2163 11556 2169 11573
rect 1731 11550 2169 11556
rect 2281 11579 2314 11581
rect 2686 11587 2727 11614
rect 2744 11587 2750 12013
rect 2686 11581 2750 11587
rect 2800 12013 3300 12019
rect 2800 11587 2806 12013
rect 2823 11965 3277 12013
rect 2823 11635 2885 11965
rect 3215 11635 3277 11965
rect 2823 11587 3277 11635
rect 3294 11587 3300 12013
rect 2800 11581 3300 11587
rect 3350 12013 3414 12019
rect 3350 11587 3356 12013
rect 3373 11986 3414 12013
rect 3786 12019 3819 12021
rect 3931 12044 4369 12050
rect 3931 12027 3937 12044
rect 4363 12027 4369 12044
rect 3931 12021 4369 12027
rect 3929 12019 4371 12021
rect 4481 12044 4919 12050
rect 4481 12027 4487 12044
rect 4913 12027 4919 12044
rect 4481 12021 4919 12027
rect 4481 12019 4514 12021
rect 3786 12013 3850 12019
rect 3786 11986 3827 12013
rect 3373 11614 3379 11986
rect 3821 11614 3827 11986
rect 3373 11587 3414 11614
rect 3350 11581 3414 11587
rect 2686 11579 2719 11581
rect 2281 11573 2719 11579
rect 2281 11556 2287 11573
rect 2713 11556 2719 11573
rect 2281 11550 2719 11556
rect 2829 11579 3271 11581
rect 2831 11573 3269 11579
rect 2831 11556 2837 11573
rect 3263 11556 3269 11573
rect 2831 11550 3269 11556
rect 3381 11579 3414 11581
rect 3786 11587 3827 11614
rect 3844 11587 3850 12013
rect 3786 11581 3850 11587
rect 3900 12013 4400 12019
rect 3900 11587 3906 12013
rect 3923 11965 4377 12013
rect 3923 11635 3985 11965
rect 4315 11635 4377 11965
rect 3923 11587 4377 11635
rect 4394 11587 4400 12013
rect 3900 11581 4400 11587
rect 4450 12013 4514 12019
rect 4450 11587 4456 12013
rect 4473 11986 4514 12013
rect 4886 12019 4919 12021
rect 5031 12044 5469 12050
rect 5031 12027 5037 12044
rect 5463 12027 5469 12044
rect 5031 12021 5469 12027
rect 5029 12019 5471 12021
rect 5581 12044 6019 12050
rect 5581 12027 5587 12044
rect 6013 12027 6019 12044
rect 5581 12021 6019 12027
rect 5581 12019 5614 12021
rect 4886 12013 4950 12019
rect 4886 11986 4927 12013
rect 4473 11614 4479 11986
rect 4921 11614 4927 11986
rect 4473 11587 4514 11614
rect 4450 11581 4514 11587
rect 3786 11579 3819 11581
rect 3381 11573 3819 11579
rect 3381 11556 3387 11573
rect 3813 11556 3819 11573
rect 3381 11550 3819 11556
rect 3929 11579 4371 11581
rect 3931 11573 4369 11579
rect 3931 11556 3937 11573
rect 4363 11556 4369 11573
rect 3931 11550 4369 11556
rect 4481 11579 4514 11581
rect 4886 11587 4927 11614
rect 4944 11587 4950 12013
rect 4886 11581 4950 11587
rect 5000 12013 5500 12019
rect 5000 11587 5006 12013
rect 5023 11965 5477 12013
rect 5023 11635 5085 11965
rect 5415 11635 5477 11965
rect 5023 11587 5477 11635
rect 5494 11587 5500 12013
rect 5000 11581 5500 11587
rect 5550 12013 5614 12019
rect 5550 11587 5556 12013
rect 5573 11986 5614 12013
rect 5986 12019 6019 12021
rect 6131 12044 6569 12050
rect 6131 12027 6137 12044
rect 6563 12027 6569 12044
rect 6131 12021 6569 12027
rect 6129 12019 6571 12021
rect 6681 12044 7119 12050
rect 6681 12027 6687 12044
rect 7113 12027 7119 12044
rect 6681 12021 7119 12027
rect 6681 12019 6714 12021
rect 5986 12013 6050 12019
rect 5986 11986 6027 12013
rect 5573 11614 5579 11986
rect 6021 11614 6027 11986
rect 5573 11587 5614 11614
rect 5550 11581 5614 11587
rect 4886 11579 4919 11581
rect 4481 11573 4919 11579
rect 4481 11556 4487 11573
rect 4913 11556 4919 11573
rect 4481 11550 4919 11556
rect 5029 11579 5471 11581
rect 5031 11573 5469 11579
rect 5031 11556 5037 11573
rect 5463 11556 5469 11573
rect 5031 11550 5469 11556
rect 5581 11579 5614 11581
rect 5986 11587 6027 11614
rect 6044 11587 6050 12013
rect 5986 11581 6050 11587
rect 6100 12013 6600 12019
rect 6100 11587 6106 12013
rect 6123 11965 6577 12013
rect 6123 11635 6185 11965
rect 6515 11635 6577 11965
rect 6123 11587 6577 11635
rect 6594 11587 6600 12013
rect 6100 11581 6600 11587
rect 6650 12013 6714 12019
rect 6650 11587 6656 12013
rect 6673 11986 6714 12013
rect 7086 12019 7119 12021
rect 7231 12044 7669 12050
rect 7231 12027 7237 12044
rect 7663 12027 7669 12044
rect 7231 12021 7669 12027
rect 7229 12019 7671 12021
rect 7781 12044 8219 12050
rect 7781 12027 7787 12044
rect 8213 12027 8219 12044
rect 7781 12021 8219 12027
rect 7781 12019 7814 12021
rect 7086 12013 7150 12019
rect 7086 11986 7127 12013
rect 6673 11614 6679 11986
rect 7121 11614 7127 11986
rect 6673 11587 6714 11614
rect 6650 11581 6714 11587
rect 5986 11579 6019 11581
rect 5581 11573 6019 11579
rect 5581 11556 5587 11573
rect 6013 11556 6019 11573
rect 5581 11550 6019 11556
rect 6129 11579 6571 11581
rect 6131 11573 6569 11579
rect 6131 11556 6137 11573
rect 6563 11556 6569 11573
rect 6131 11550 6569 11556
rect 6681 11579 6714 11581
rect 7086 11587 7127 11614
rect 7144 11587 7150 12013
rect 7086 11581 7150 11587
rect 7200 12013 7700 12019
rect 7200 11587 7206 12013
rect 7223 11965 7677 12013
rect 7223 11635 7285 11965
rect 7615 11635 7677 11965
rect 7223 11587 7677 11635
rect 7694 11587 7700 12013
rect 7200 11581 7700 11587
rect 7750 12013 7814 12019
rect 7750 11587 7756 12013
rect 7773 11986 7814 12013
rect 8186 12019 8219 12021
rect 8331 12044 8769 12050
rect 8331 12027 8337 12044
rect 8763 12027 8769 12044
rect 8331 12021 8769 12027
rect 8329 12019 8771 12021
rect 8881 12044 9319 12050
rect 8881 12027 8887 12044
rect 9313 12027 9319 12044
rect 8881 12021 9319 12027
rect 8881 12019 8914 12021
rect 8186 12013 8250 12019
rect 8186 11986 8227 12013
rect 7773 11614 7779 11986
rect 8221 11614 8227 11986
rect 7773 11587 7814 11614
rect 7750 11581 7814 11587
rect 7086 11579 7119 11581
rect 6681 11573 7119 11579
rect 6681 11556 6687 11573
rect 7113 11556 7119 11573
rect 6681 11550 7119 11556
rect 7229 11579 7671 11581
rect 7231 11573 7669 11579
rect 7231 11556 7237 11573
rect 7663 11556 7669 11573
rect 7231 11550 7669 11556
rect 7781 11579 7814 11581
rect 8186 11587 8227 11614
rect 8244 11587 8250 12013
rect 8186 11581 8250 11587
rect 8300 12013 8800 12019
rect 8300 11587 8306 12013
rect 8323 11965 8777 12013
rect 8323 11635 8385 11965
rect 8715 11635 8777 11965
rect 8323 11587 8777 11635
rect 8794 11587 8800 12013
rect 8300 11581 8800 11587
rect 8850 12013 8914 12019
rect 8850 11587 8856 12013
rect 8873 11986 8914 12013
rect 9286 12019 9319 12021
rect 9431 12044 9869 12050
rect 9431 12027 9437 12044
rect 9863 12027 9869 12044
rect 9431 12021 9869 12027
rect 9429 12019 9871 12021
rect 9981 12044 10419 12050
rect 9981 12027 9987 12044
rect 10413 12027 10419 12044
rect 9981 12021 10419 12027
rect 9981 12019 10014 12021
rect 9286 12013 9350 12019
rect 9286 11986 9327 12013
rect 8873 11614 8879 11986
rect 9321 11614 9327 11986
rect 8873 11587 8914 11614
rect 8850 11581 8914 11587
rect 8186 11579 8219 11581
rect 7781 11573 8219 11579
rect 7781 11556 7787 11573
rect 8213 11556 8219 11573
rect 7781 11550 8219 11556
rect 8329 11579 8771 11581
rect 8331 11573 8769 11579
rect 8331 11556 8337 11573
rect 8763 11556 8769 11573
rect 8331 11550 8769 11556
rect 8881 11579 8914 11581
rect 9286 11587 9327 11614
rect 9344 11587 9350 12013
rect 9286 11581 9350 11587
rect 9400 12013 9900 12019
rect 9400 11587 9406 12013
rect 9423 11965 9877 12013
rect 9423 11635 9485 11965
rect 9815 11635 9877 11965
rect 9423 11587 9877 11635
rect 9894 11587 9900 12013
rect 9400 11581 9900 11587
rect 9950 12013 10014 12019
rect 9950 11587 9956 12013
rect 9973 11986 10014 12013
rect 10386 12019 10419 12021
rect 10531 12044 10969 12050
rect 10531 12027 10537 12044
rect 10963 12027 10969 12044
rect 10531 12021 10969 12027
rect 10529 12019 10971 12021
rect 11081 12044 11519 12050
rect 11081 12027 11087 12044
rect 11513 12027 11519 12044
rect 11081 12021 11519 12027
rect 11081 12019 11114 12021
rect 10386 12013 10450 12019
rect 10386 11986 10427 12013
rect 9973 11614 9979 11986
rect 10421 11614 10427 11986
rect 9973 11587 10014 11614
rect 9950 11581 10014 11587
rect 9286 11579 9319 11581
rect 8881 11573 9319 11579
rect 8881 11556 8887 11573
rect 9313 11556 9319 11573
rect 8881 11550 9319 11556
rect 9429 11579 9871 11581
rect 9431 11573 9869 11579
rect 9431 11556 9437 11573
rect 9863 11556 9869 11573
rect 9431 11550 9869 11556
rect 9981 11579 10014 11581
rect 10386 11587 10427 11614
rect 10444 11587 10450 12013
rect 10386 11581 10450 11587
rect 10500 12013 11000 12019
rect 10500 11587 10506 12013
rect 10523 11965 10977 12013
rect 10523 11635 10585 11965
rect 10915 11635 10977 11965
rect 10523 11587 10977 11635
rect 10994 11587 11000 12013
rect 10500 11581 11000 11587
rect 11050 12013 11114 12019
rect 11050 11587 11056 12013
rect 11073 11986 11114 12013
rect 11486 12019 11519 12021
rect 11631 12044 12069 12050
rect 11631 12027 11637 12044
rect 12063 12027 12069 12044
rect 11631 12021 12069 12027
rect 11629 12019 12071 12021
rect 12181 12044 12619 12050
rect 12181 12027 12187 12044
rect 12613 12027 12619 12044
rect 12181 12021 12619 12027
rect 12181 12019 12214 12021
rect 11486 12013 11550 12019
rect 11486 11986 11527 12013
rect 11073 11614 11079 11986
rect 11521 11614 11527 11986
rect 11073 11587 11114 11614
rect 11050 11581 11114 11587
rect 10386 11579 10419 11581
rect 9981 11573 10419 11579
rect 9981 11556 9987 11573
rect 10413 11556 10419 11573
rect 9981 11550 10419 11556
rect 10529 11579 10971 11581
rect 10531 11573 10969 11579
rect 10531 11556 10537 11573
rect 10963 11556 10969 11573
rect 10531 11550 10969 11556
rect 11081 11579 11114 11581
rect 11486 11587 11527 11614
rect 11544 11587 11550 12013
rect 11486 11581 11550 11587
rect 11600 12013 12100 12019
rect 11600 11587 11606 12013
rect 11623 11965 12077 12013
rect 11623 11635 11685 11965
rect 12015 11635 12077 11965
rect 11623 11587 12077 11635
rect 12094 11587 12100 12013
rect 11600 11581 12100 11587
rect 12150 12013 12214 12019
rect 12150 11587 12156 12013
rect 12173 11986 12214 12013
rect 12586 12019 12619 12021
rect 12731 12044 13169 12050
rect 12731 12027 12737 12044
rect 13163 12027 13169 12044
rect 12731 12021 13169 12027
rect 12729 12019 13171 12021
rect 13281 12044 13719 12050
rect 13281 12027 13287 12044
rect 13713 12027 13719 12044
rect 13281 12021 13719 12027
rect 13281 12019 13314 12021
rect 12586 12013 12650 12019
rect 12586 11986 12627 12013
rect 12173 11614 12179 11986
rect 12621 11614 12627 11986
rect 12173 11587 12214 11614
rect 12150 11581 12214 11587
rect 11486 11579 11519 11581
rect 11081 11573 11519 11579
rect 11081 11556 11087 11573
rect 11513 11556 11519 11573
rect 11081 11550 11519 11556
rect 11629 11579 12071 11581
rect 11631 11573 12069 11579
rect 11631 11556 11637 11573
rect 12063 11556 12069 11573
rect 11631 11550 12069 11556
rect 12181 11579 12214 11581
rect 12586 11587 12627 11614
rect 12644 11587 12650 12013
rect 12586 11581 12650 11587
rect 12700 12013 13200 12019
rect 12700 11587 12706 12013
rect 12723 11965 13177 12013
rect 12723 11635 12785 11965
rect 13115 11635 13177 11965
rect 12723 11587 13177 11635
rect 13194 11587 13200 12013
rect 12700 11581 13200 11587
rect 13250 12013 13314 12019
rect 13250 11587 13256 12013
rect 13273 11986 13314 12013
rect 13273 11614 13279 11986
rect 13273 11587 13314 11614
rect 13250 11581 13314 11587
rect 12586 11579 12619 11581
rect 12181 11573 12619 11579
rect 12181 11556 12187 11573
rect 12613 11556 12619 11573
rect 12181 11550 12619 11556
rect 12729 11579 13171 11581
rect 12731 11573 13169 11579
rect 12731 11556 12737 11573
rect 13163 11556 13169 11573
rect 12731 11550 13169 11556
rect 13281 11579 13314 11581
rect 13281 11573 13719 11579
rect 13281 11556 13287 11573
rect 13713 11556 13719 11573
rect 13281 11550 13719 11556
rect -469 11494 -31 11500
rect -469 11477 -463 11494
rect -37 11477 -31 11494
rect -469 11471 -31 11477
rect -64 11469 -31 11471
rect 81 11494 519 11500
rect 81 11477 87 11494
rect 513 11477 519 11494
rect 81 11471 519 11477
rect 79 11469 521 11471
rect 631 11494 1069 11500
rect 631 11477 637 11494
rect 1063 11477 1069 11494
rect 631 11471 1069 11477
rect 631 11469 664 11471
rect -64 11463 0 11469
rect -64 11436 -23 11463
rect -29 11064 -23 11436
rect -64 11037 -23 11064
rect -6 11037 0 11463
rect -64 11031 0 11037
rect 50 11463 550 11469
rect 50 11037 56 11463
rect 73 11415 527 11463
rect 73 11085 135 11415
rect 465 11085 527 11415
rect 73 11037 527 11085
rect 544 11037 550 11463
rect 50 11031 550 11037
rect 600 11463 664 11469
rect 600 11037 606 11463
rect 623 11436 664 11463
rect 1036 11469 1069 11471
rect 1181 11494 1619 11500
rect 1181 11477 1187 11494
rect 1613 11477 1619 11494
rect 1181 11471 1619 11477
rect 1179 11469 1621 11471
rect 1731 11494 2169 11500
rect 1731 11477 1737 11494
rect 2163 11477 2169 11494
rect 1731 11471 2169 11477
rect 1731 11469 1764 11471
rect 1036 11463 1100 11469
rect 1036 11436 1077 11463
rect 623 11064 629 11436
rect 1071 11064 1077 11436
rect 623 11037 664 11064
rect 600 11031 664 11037
rect -64 11029 -31 11031
rect -469 11023 -31 11029
rect -469 11006 -463 11023
rect -37 11006 -31 11023
rect -469 11000 -31 11006
rect 79 11029 521 11031
rect 81 11023 519 11029
rect 81 11006 87 11023
rect 513 11006 519 11023
rect 81 11000 519 11006
rect 631 11029 664 11031
rect 1036 11037 1077 11064
rect 1094 11037 1100 11463
rect 1036 11031 1100 11037
rect 1150 11463 1650 11469
rect 1150 11037 1156 11463
rect 1173 11415 1627 11463
rect 1173 11085 1235 11415
rect 1565 11085 1627 11415
rect 1173 11037 1627 11085
rect 1644 11037 1650 11463
rect 1150 11031 1650 11037
rect 1700 11463 1764 11469
rect 1700 11037 1706 11463
rect 1723 11436 1764 11463
rect 2136 11469 2169 11471
rect 2281 11494 2719 11500
rect 2281 11477 2287 11494
rect 2713 11477 2719 11494
rect 2281 11471 2719 11477
rect 2279 11469 2721 11471
rect 2831 11494 3269 11500
rect 2831 11477 2837 11494
rect 3263 11477 3269 11494
rect 2831 11471 3269 11477
rect 2831 11469 2864 11471
rect 2136 11463 2200 11469
rect 2136 11436 2177 11463
rect 1723 11064 1729 11436
rect 2171 11064 2177 11436
rect 1723 11037 1764 11064
rect 1700 11031 1764 11037
rect 1036 11029 1069 11031
rect 631 11023 1069 11029
rect 631 11006 637 11023
rect 1063 11006 1069 11023
rect 631 11000 1069 11006
rect 1179 11029 1621 11031
rect 1181 11023 1619 11029
rect 1181 11006 1187 11023
rect 1613 11006 1619 11023
rect 1181 11000 1619 11006
rect 1731 11029 1764 11031
rect 2136 11037 2177 11064
rect 2194 11037 2200 11463
rect 2136 11031 2200 11037
rect 2250 11463 2750 11469
rect 2250 11037 2256 11463
rect 2273 11415 2727 11463
rect 2273 11085 2335 11415
rect 2665 11085 2727 11415
rect 2273 11037 2727 11085
rect 2744 11037 2750 11463
rect 2250 11031 2750 11037
rect 2800 11463 2864 11469
rect 2800 11037 2806 11463
rect 2823 11436 2864 11463
rect 3236 11469 3269 11471
rect 3381 11494 3819 11500
rect 3381 11477 3387 11494
rect 3813 11477 3819 11494
rect 3381 11471 3819 11477
rect 3379 11469 3821 11471
rect 3931 11494 4369 11500
rect 3931 11477 3937 11494
rect 4363 11477 4369 11494
rect 3931 11471 4369 11477
rect 3931 11469 3964 11471
rect 3236 11463 3300 11469
rect 3236 11436 3277 11463
rect 2823 11064 2829 11436
rect 3271 11064 3277 11436
rect 2823 11037 2864 11064
rect 2800 11031 2864 11037
rect 2136 11029 2169 11031
rect 1731 11023 2169 11029
rect 1731 11006 1737 11023
rect 2163 11006 2169 11023
rect 1731 11000 2169 11006
rect 2279 11029 2721 11031
rect 2281 11023 2719 11029
rect 2281 11006 2287 11023
rect 2713 11006 2719 11023
rect 2281 11000 2719 11006
rect 2831 11029 2864 11031
rect 3236 11037 3277 11064
rect 3294 11037 3300 11463
rect 3236 11031 3300 11037
rect 3350 11463 3850 11469
rect 3350 11037 3356 11463
rect 3373 11415 3827 11463
rect 3373 11085 3435 11415
rect 3765 11085 3827 11415
rect 3373 11037 3827 11085
rect 3844 11037 3850 11463
rect 3350 11031 3850 11037
rect 3900 11463 3964 11469
rect 3900 11037 3906 11463
rect 3923 11436 3964 11463
rect 4336 11469 4369 11471
rect 4481 11494 4919 11500
rect 4481 11477 4487 11494
rect 4913 11477 4919 11494
rect 4481 11471 4919 11477
rect 4479 11469 4921 11471
rect 5031 11494 5469 11500
rect 5031 11477 5037 11494
rect 5463 11477 5469 11494
rect 5031 11471 5469 11477
rect 5031 11469 5064 11471
rect 4336 11463 4400 11469
rect 4336 11436 4377 11463
rect 3923 11064 3929 11436
rect 4371 11064 4377 11436
rect 3923 11037 3964 11064
rect 3900 11031 3964 11037
rect 3236 11029 3269 11031
rect 2831 11023 3269 11029
rect 2831 11006 2837 11023
rect 3263 11006 3269 11023
rect 2831 11000 3269 11006
rect 3379 11029 3821 11031
rect 3381 11023 3819 11029
rect 3381 11006 3387 11023
rect 3813 11006 3819 11023
rect 3381 11000 3819 11006
rect 3931 11029 3964 11031
rect 4336 11037 4377 11064
rect 4394 11037 4400 11463
rect 4336 11031 4400 11037
rect 4450 11463 4950 11469
rect 4450 11037 4456 11463
rect 4473 11415 4927 11463
rect 4473 11085 4535 11415
rect 4865 11085 4927 11415
rect 4473 11037 4927 11085
rect 4944 11037 4950 11463
rect 4450 11031 4950 11037
rect 5000 11463 5064 11469
rect 5000 11037 5006 11463
rect 5023 11436 5064 11463
rect 5436 11469 5469 11471
rect 5581 11494 6019 11500
rect 5581 11477 5587 11494
rect 6013 11477 6019 11494
rect 5581 11471 6019 11477
rect 5579 11469 6021 11471
rect 6131 11494 6569 11500
rect 6131 11477 6137 11494
rect 6563 11477 6569 11494
rect 6131 11471 6569 11477
rect 6131 11469 6164 11471
rect 5436 11463 5500 11469
rect 5436 11436 5477 11463
rect 5023 11064 5029 11436
rect 5471 11064 5477 11436
rect 5023 11037 5064 11064
rect 5000 11031 5064 11037
rect 4336 11029 4369 11031
rect 3931 11023 4369 11029
rect 3931 11006 3937 11023
rect 4363 11006 4369 11023
rect 3931 11000 4369 11006
rect 4479 11029 4921 11031
rect 4481 11023 4919 11029
rect 4481 11006 4487 11023
rect 4913 11006 4919 11023
rect 4481 11000 4919 11006
rect 5031 11029 5064 11031
rect 5436 11037 5477 11064
rect 5494 11037 5500 11463
rect 5436 11031 5500 11037
rect 5550 11463 6050 11469
rect 5550 11037 5556 11463
rect 5573 11415 6027 11463
rect 5573 11085 5635 11415
rect 5965 11085 6027 11415
rect 5573 11037 6027 11085
rect 6044 11037 6050 11463
rect 5550 11031 6050 11037
rect 6100 11463 6164 11469
rect 6100 11037 6106 11463
rect 6123 11436 6164 11463
rect 6536 11469 6569 11471
rect 6681 11494 7119 11500
rect 6681 11477 6687 11494
rect 7113 11477 7119 11494
rect 6681 11471 7119 11477
rect 6679 11469 7121 11471
rect 7231 11494 7669 11500
rect 7231 11477 7237 11494
rect 7663 11477 7669 11494
rect 7231 11471 7669 11477
rect 7231 11469 7264 11471
rect 6536 11463 6600 11469
rect 6536 11436 6577 11463
rect 6123 11064 6129 11436
rect 6571 11064 6577 11436
rect 6123 11037 6164 11064
rect 6100 11031 6164 11037
rect 5436 11029 5469 11031
rect 5031 11023 5469 11029
rect 5031 11006 5037 11023
rect 5463 11006 5469 11023
rect 5031 11000 5469 11006
rect 5579 11029 6021 11031
rect 5581 11023 6019 11029
rect 5581 11006 5587 11023
rect 6013 11006 6019 11023
rect 5581 11000 6019 11006
rect 6131 11029 6164 11031
rect 6536 11037 6577 11064
rect 6594 11037 6600 11463
rect 6536 11031 6600 11037
rect 6650 11463 7150 11469
rect 6650 11037 6656 11463
rect 6673 11415 7127 11463
rect 6673 11085 6735 11415
rect 7065 11085 7127 11415
rect 6673 11037 7127 11085
rect 7144 11037 7150 11463
rect 6650 11031 7150 11037
rect 7200 11463 7264 11469
rect 7200 11037 7206 11463
rect 7223 11436 7264 11463
rect 7636 11469 7669 11471
rect 7781 11494 8219 11500
rect 7781 11477 7787 11494
rect 8213 11477 8219 11494
rect 7781 11471 8219 11477
rect 7779 11469 8221 11471
rect 8331 11494 8769 11500
rect 8331 11477 8337 11494
rect 8763 11477 8769 11494
rect 8331 11471 8769 11477
rect 8331 11469 8364 11471
rect 7636 11463 7700 11469
rect 7636 11436 7677 11463
rect 7223 11064 7229 11436
rect 7671 11064 7677 11436
rect 7223 11037 7264 11064
rect 7200 11031 7264 11037
rect 6536 11029 6569 11031
rect 6131 11023 6569 11029
rect 6131 11006 6137 11023
rect 6563 11006 6569 11023
rect 6131 11000 6569 11006
rect 6679 11029 7121 11031
rect 6681 11023 7119 11029
rect 6681 11006 6687 11023
rect 7113 11006 7119 11023
rect 6681 11000 7119 11006
rect 7231 11029 7264 11031
rect 7636 11037 7677 11064
rect 7694 11037 7700 11463
rect 7636 11031 7700 11037
rect 7750 11463 8250 11469
rect 7750 11037 7756 11463
rect 7773 11415 8227 11463
rect 7773 11085 7835 11415
rect 8165 11085 8227 11415
rect 7773 11037 8227 11085
rect 8244 11037 8250 11463
rect 7750 11031 8250 11037
rect 8300 11463 8364 11469
rect 8300 11037 8306 11463
rect 8323 11436 8364 11463
rect 8736 11469 8769 11471
rect 8881 11494 9319 11500
rect 8881 11477 8887 11494
rect 9313 11477 9319 11494
rect 8881 11471 9319 11477
rect 8879 11469 9321 11471
rect 9431 11494 9869 11500
rect 9431 11477 9437 11494
rect 9863 11477 9869 11494
rect 9431 11471 9869 11477
rect 9431 11469 9464 11471
rect 8736 11463 8800 11469
rect 8736 11436 8777 11463
rect 8323 11064 8329 11436
rect 8771 11064 8777 11436
rect 8323 11037 8364 11064
rect 8300 11031 8364 11037
rect 7636 11029 7669 11031
rect 7231 11023 7669 11029
rect 7231 11006 7237 11023
rect 7663 11006 7669 11023
rect 7231 11000 7669 11006
rect 7779 11029 8221 11031
rect 7781 11023 8219 11029
rect 7781 11006 7787 11023
rect 8213 11006 8219 11023
rect 7781 11000 8219 11006
rect 8331 11029 8364 11031
rect 8736 11037 8777 11064
rect 8794 11037 8800 11463
rect 8736 11031 8800 11037
rect 8850 11463 9350 11469
rect 8850 11037 8856 11463
rect 8873 11415 9327 11463
rect 8873 11085 8935 11415
rect 9265 11085 9327 11415
rect 8873 11037 9327 11085
rect 9344 11037 9350 11463
rect 8850 11031 9350 11037
rect 9400 11463 9464 11469
rect 9400 11037 9406 11463
rect 9423 11436 9464 11463
rect 9836 11469 9869 11471
rect 9981 11494 10419 11500
rect 9981 11477 9987 11494
rect 10413 11477 10419 11494
rect 9981 11471 10419 11477
rect 9979 11469 10421 11471
rect 10531 11494 10969 11500
rect 10531 11477 10537 11494
rect 10963 11477 10969 11494
rect 10531 11471 10969 11477
rect 10531 11469 10564 11471
rect 9836 11463 9900 11469
rect 9836 11436 9877 11463
rect 9423 11064 9429 11436
rect 9871 11064 9877 11436
rect 9423 11037 9464 11064
rect 9400 11031 9464 11037
rect 8736 11029 8769 11031
rect 8331 11023 8769 11029
rect 8331 11006 8337 11023
rect 8763 11006 8769 11023
rect 8331 11000 8769 11006
rect 8879 11029 9321 11031
rect 8881 11023 9319 11029
rect 8881 11006 8887 11023
rect 9313 11006 9319 11023
rect 8881 11000 9319 11006
rect 9431 11029 9464 11031
rect 9836 11037 9877 11064
rect 9894 11037 9900 11463
rect 9836 11031 9900 11037
rect 9950 11463 10450 11469
rect 9950 11037 9956 11463
rect 9973 11415 10427 11463
rect 9973 11085 10035 11415
rect 10365 11085 10427 11415
rect 9973 11037 10427 11085
rect 10444 11037 10450 11463
rect 9950 11031 10450 11037
rect 10500 11463 10564 11469
rect 10500 11037 10506 11463
rect 10523 11436 10564 11463
rect 10936 11469 10969 11471
rect 11081 11494 11519 11500
rect 11081 11477 11087 11494
rect 11513 11477 11519 11494
rect 11081 11471 11519 11477
rect 11079 11469 11521 11471
rect 11631 11494 12069 11500
rect 11631 11477 11637 11494
rect 12063 11477 12069 11494
rect 11631 11471 12069 11477
rect 11631 11469 11664 11471
rect 10936 11463 11000 11469
rect 10936 11436 10977 11463
rect 10523 11064 10529 11436
rect 10971 11064 10977 11436
rect 10523 11037 10564 11064
rect 10500 11031 10564 11037
rect 9836 11029 9869 11031
rect 9431 11023 9869 11029
rect 9431 11006 9437 11023
rect 9863 11006 9869 11023
rect 9431 11000 9869 11006
rect 9979 11029 10421 11031
rect 9981 11023 10419 11029
rect 9981 11006 9987 11023
rect 10413 11006 10419 11023
rect 9981 11000 10419 11006
rect 10531 11029 10564 11031
rect 10936 11037 10977 11064
rect 10994 11037 11000 11463
rect 10936 11031 11000 11037
rect 11050 11463 11550 11469
rect 11050 11037 11056 11463
rect 11073 11415 11527 11463
rect 11073 11085 11135 11415
rect 11465 11085 11527 11415
rect 11073 11037 11527 11085
rect 11544 11037 11550 11463
rect 11050 11031 11550 11037
rect 11600 11463 11664 11469
rect 11600 11037 11606 11463
rect 11623 11436 11664 11463
rect 12036 11469 12069 11471
rect 12181 11494 12619 11500
rect 12181 11477 12187 11494
rect 12613 11477 12619 11494
rect 12181 11471 12619 11477
rect 12179 11469 12621 11471
rect 12731 11494 13169 11500
rect 12731 11477 12737 11494
rect 13163 11477 13169 11494
rect 12731 11471 13169 11477
rect 12731 11469 12764 11471
rect 12036 11463 12100 11469
rect 12036 11436 12077 11463
rect 11623 11064 11629 11436
rect 12071 11064 12077 11436
rect 11623 11037 11664 11064
rect 11600 11031 11664 11037
rect 10936 11029 10969 11031
rect 10531 11023 10969 11029
rect 10531 11006 10537 11023
rect 10963 11006 10969 11023
rect 10531 11000 10969 11006
rect 11079 11029 11521 11031
rect 11081 11023 11519 11029
rect 11081 11006 11087 11023
rect 11513 11006 11519 11023
rect 11081 11000 11519 11006
rect 11631 11029 11664 11031
rect 12036 11037 12077 11064
rect 12094 11037 12100 11463
rect 12036 11031 12100 11037
rect 12150 11463 12650 11469
rect 12150 11037 12156 11463
rect 12173 11415 12627 11463
rect 12173 11085 12235 11415
rect 12565 11085 12627 11415
rect 12173 11037 12627 11085
rect 12644 11037 12650 11463
rect 12150 11031 12650 11037
rect 12700 11463 12764 11469
rect 12700 11037 12706 11463
rect 12723 11436 12764 11463
rect 13136 11469 13169 11471
rect 13281 11494 13719 11500
rect 13281 11477 13287 11494
rect 13713 11477 13719 11494
rect 13281 11471 13719 11477
rect 13279 11469 13721 11471
rect 13136 11463 13200 11469
rect 13136 11436 13177 11463
rect 12723 11064 12729 11436
rect 13171 11064 13177 11436
rect 12723 11037 12764 11064
rect 12700 11031 12764 11037
rect 12036 11029 12069 11031
rect 11631 11023 12069 11029
rect 11631 11006 11637 11023
rect 12063 11006 12069 11023
rect 11631 11000 12069 11006
rect 12179 11029 12621 11031
rect 12181 11023 12619 11029
rect 12181 11006 12187 11023
rect 12613 11006 12619 11023
rect 12181 11000 12619 11006
rect 12731 11029 12764 11031
rect 13136 11037 13177 11064
rect 13194 11037 13200 11463
rect 13136 11031 13200 11037
rect 13250 11463 13721 11469
rect 13250 11037 13256 11463
rect 13273 11415 13721 11463
rect 13273 11085 13335 11415
rect 13665 11085 13721 11415
rect 13273 11037 13721 11085
rect 13250 11031 13721 11037
rect 13136 11029 13169 11031
rect 12731 11023 13169 11029
rect 12731 11006 12737 11023
rect 13163 11006 13169 11023
rect 12731 11000 13169 11006
rect 13279 11029 13721 11031
rect 13281 11023 13719 11029
rect 13281 11006 13287 11023
rect 13713 11006 13719 11023
rect 13281 11000 13719 11006
rect -469 10944 -31 10950
rect -469 10927 -463 10944
rect -37 10927 -31 10944
rect -469 10921 -31 10927
rect -471 10919 -29 10921
rect 81 10944 519 10950
rect 81 10927 87 10944
rect 513 10927 519 10944
rect 81 10921 519 10927
rect 81 10919 114 10921
rect -471 10913 0 10919
rect -471 10865 -23 10913
rect -471 10535 -415 10865
rect -85 10535 -23 10865
rect -471 10487 -23 10535
rect -6 10487 0 10913
rect -471 10481 0 10487
rect 50 10913 114 10919
rect 50 10487 56 10913
rect 73 10886 114 10913
rect 486 10919 519 10921
rect 631 10944 1069 10950
rect 631 10927 637 10944
rect 1063 10927 1069 10944
rect 631 10921 1069 10927
rect 629 10919 1071 10921
rect 1181 10944 1619 10950
rect 1181 10927 1187 10944
rect 1613 10927 1619 10944
rect 1181 10921 1619 10927
rect 1181 10919 1214 10921
rect 486 10913 550 10919
rect 486 10886 527 10913
rect 73 10514 79 10886
rect 521 10514 527 10886
rect 73 10487 114 10514
rect 50 10481 114 10487
rect -471 10479 -29 10481
rect -469 10473 -31 10479
rect -469 10456 -463 10473
rect -37 10456 -31 10473
rect -469 10450 -31 10456
rect 81 10479 114 10481
rect 486 10487 527 10514
rect 544 10487 550 10913
rect 486 10481 550 10487
rect 600 10913 1100 10919
rect 600 10487 606 10913
rect 623 10865 1077 10913
rect 623 10535 685 10865
rect 1015 10535 1077 10865
rect 623 10487 1077 10535
rect 1094 10487 1100 10913
rect 600 10481 1100 10487
rect 1150 10913 1214 10919
rect 1150 10487 1156 10913
rect 1173 10886 1214 10913
rect 1586 10919 1619 10921
rect 1731 10944 2169 10950
rect 1731 10927 1737 10944
rect 2163 10927 2169 10944
rect 1731 10921 2169 10927
rect 1729 10919 2171 10921
rect 2281 10944 2719 10950
rect 2281 10927 2287 10944
rect 2713 10927 2719 10944
rect 2281 10921 2719 10927
rect 2281 10919 2314 10921
rect 1586 10913 1650 10919
rect 1586 10886 1627 10913
rect 1173 10514 1179 10886
rect 1621 10514 1627 10886
rect 1173 10487 1214 10514
rect 1150 10481 1214 10487
rect 486 10479 519 10481
rect 81 10473 519 10479
rect 81 10456 87 10473
rect 513 10456 519 10473
rect 81 10450 519 10456
rect 629 10479 1071 10481
rect 631 10473 1069 10479
rect 631 10456 637 10473
rect 1063 10456 1069 10473
rect 631 10450 1069 10456
rect 1181 10479 1214 10481
rect 1586 10487 1627 10514
rect 1644 10487 1650 10913
rect 1586 10481 1650 10487
rect 1700 10913 2200 10919
rect 1700 10487 1706 10913
rect 1723 10865 2177 10913
rect 1723 10535 1785 10865
rect 2115 10535 2177 10865
rect 1723 10487 2177 10535
rect 2194 10487 2200 10913
rect 1700 10481 2200 10487
rect 2250 10913 2314 10919
rect 2250 10487 2256 10913
rect 2273 10886 2314 10913
rect 2686 10919 2719 10921
rect 2831 10944 3269 10950
rect 2831 10927 2837 10944
rect 3263 10927 3269 10944
rect 2831 10921 3269 10927
rect 2829 10919 3271 10921
rect 3381 10944 3819 10950
rect 3381 10927 3387 10944
rect 3813 10927 3819 10944
rect 3381 10921 3819 10927
rect 3381 10919 3414 10921
rect 2686 10913 2750 10919
rect 2686 10886 2727 10913
rect 2273 10514 2279 10886
rect 2721 10514 2727 10886
rect 2273 10487 2314 10514
rect 2250 10481 2314 10487
rect 1586 10479 1619 10481
rect 1181 10473 1619 10479
rect 1181 10456 1187 10473
rect 1613 10456 1619 10473
rect 1181 10450 1619 10456
rect 1729 10479 2171 10481
rect 1731 10473 2169 10479
rect 1731 10456 1737 10473
rect 2163 10456 2169 10473
rect 1731 10450 2169 10456
rect 2281 10479 2314 10481
rect 2686 10487 2727 10514
rect 2744 10487 2750 10913
rect 2686 10481 2750 10487
rect 2800 10913 3300 10919
rect 2800 10487 2806 10913
rect 2823 10865 3277 10913
rect 2823 10535 2885 10865
rect 3215 10535 3277 10865
rect 2823 10487 3277 10535
rect 3294 10487 3300 10913
rect 2800 10481 3300 10487
rect 3350 10913 3414 10919
rect 3350 10487 3356 10913
rect 3373 10886 3414 10913
rect 3786 10919 3819 10921
rect 3931 10944 4369 10950
rect 3931 10927 3937 10944
rect 4363 10927 4369 10944
rect 3931 10921 4369 10927
rect 3929 10919 4371 10921
rect 4481 10944 4919 10950
rect 4481 10927 4487 10944
rect 4913 10927 4919 10944
rect 4481 10921 4919 10927
rect 4481 10919 4514 10921
rect 3786 10913 3850 10919
rect 3786 10886 3827 10913
rect 3373 10514 3379 10886
rect 3821 10514 3827 10886
rect 3373 10487 3414 10514
rect 3350 10481 3414 10487
rect 2686 10479 2719 10481
rect 2281 10473 2719 10479
rect 2281 10456 2287 10473
rect 2713 10456 2719 10473
rect 2281 10450 2719 10456
rect 2829 10479 3271 10481
rect 2831 10473 3269 10479
rect 2831 10456 2837 10473
rect 3263 10456 3269 10473
rect 2831 10450 3269 10456
rect 3381 10479 3414 10481
rect 3786 10487 3827 10514
rect 3844 10487 3850 10913
rect 3786 10481 3850 10487
rect 3900 10913 4400 10919
rect 3900 10487 3906 10913
rect 3923 10865 4377 10913
rect 3923 10535 3985 10865
rect 4315 10535 4377 10865
rect 3923 10487 4377 10535
rect 4394 10487 4400 10913
rect 3900 10481 4400 10487
rect 4450 10913 4514 10919
rect 4450 10487 4456 10913
rect 4473 10886 4514 10913
rect 4886 10919 4919 10921
rect 5031 10944 5469 10950
rect 5031 10927 5037 10944
rect 5463 10927 5469 10944
rect 5031 10921 5469 10927
rect 5029 10919 5471 10921
rect 5581 10944 6019 10950
rect 5581 10927 5587 10944
rect 6013 10927 6019 10944
rect 5581 10921 6019 10927
rect 5581 10919 5614 10921
rect 4886 10913 4950 10919
rect 4886 10886 4927 10913
rect 4473 10514 4479 10886
rect 4921 10514 4927 10886
rect 4473 10487 4514 10514
rect 4450 10481 4514 10487
rect 3786 10479 3819 10481
rect 3381 10473 3819 10479
rect 3381 10456 3387 10473
rect 3813 10456 3819 10473
rect 3381 10450 3819 10456
rect 3929 10479 4371 10481
rect 3931 10473 4369 10479
rect 3931 10456 3937 10473
rect 4363 10456 4369 10473
rect 3931 10450 4369 10456
rect 4481 10479 4514 10481
rect 4886 10487 4927 10514
rect 4944 10487 4950 10913
rect 4886 10481 4950 10487
rect 5000 10913 5500 10919
rect 5000 10487 5006 10913
rect 5023 10865 5477 10913
rect 5023 10535 5085 10865
rect 5415 10535 5477 10865
rect 5023 10487 5477 10535
rect 5494 10487 5500 10913
rect 5000 10481 5500 10487
rect 5550 10913 5614 10919
rect 5550 10487 5556 10913
rect 5573 10886 5614 10913
rect 5986 10919 6019 10921
rect 6131 10944 6569 10950
rect 6131 10927 6137 10944
rect 6563 10927 6569 10944
rect 6131 10921 6569 10927
rect 6129 10919 6571 10921
rect 6681 10944 7119 10950
rect 6681 10927 6687 10944
rect 7113 10927 7119 10944
rect 6681 10921 7119 10927
rect 6681 10919 6714 10921
rect 5986 10913 6050 10919
rect 5986 10886 6027 10913
rect 5573 10514 5579 10886
rect 6021 10514 6027 10886
rect 5573 10487 5614 10514
rect 5550 10481 5614 10487
rect 4886 10479 4919 10481
rect 4481 10473 4919 10479
rect 4481 10456 4487 10473
rect 4913 10456 4919 10473
rect 4481 10450 4919 10456
rect 5029 10479 5471 10481
rect 5031 10473 5469 10479
rect 5031 10456 5037 10473
rect 5463 10456 5469 10473
rect 5031 10450 5469 10456
rect 5581 10479 5614 10481
rect 5986 10487 6027 10514
rect 6044 10487 6050 10913
rect 5986 10481 6050 10487
rect 6100 10913 6600 10919
rect 6100 10487 6106 10913
rect 6123 10865 6577 10913
rect 6123 10535 6185 10865
rect 6515 10535 6577 10865
rect 6123 10487 6577 10535
rect 6594 10487 6600 10913
rect 6100 10481 6600 10487
rect 6650 10913 6714 10919
rect 6650 10487 6656 10913
rect 6673 10886 6714 10913
rect 7086 10919 7119 10921
rect 7231 10944 7669 10950
rect 7231 10927 7237 10944
rect 7663 10927 7669 10944
rect 7231 10921 7669 10927
rect 7229 10919 7671 10921
rect 7781 10944 8219 10950
rect 7781 10927 7787 10944
rect 8213 10927 8219 10944
rect 7781 10921 8219 10927
rect 7781 10919 7814 10921
rect 7086 10913 7150 10919
rect 7086 10886 7127 10913
rect 6673 10514 6679 10886
rect 7121 10514 7127 10886
rect 6673 10487 6714 10514
rect 6650 10481 6714 10487
rect 5986 10479 6019 10481
rect 5581 10473 6019 10479
rect 5581 10456 5587 10473
rect 6013 10456 6019 10473
rect 5581 10450 6019 10456
rect 6129 10479 6571 10481
rect 6131 10473 6569 10479
rect 6131 10456 6137 10473
rect 6563 10456 6569 10473
rect 6131 10450 6569 10456
rect 6681 10479 6714 10481
rect 7086 10487 7127 10514
rect 7144 10487 7150 10913
rect 7086 10481 7150 10487
rect 7200 10913 7700 10919
rect 7200 10487 7206 10913
rect 7223 10865 7677 10913
rect 7223 10535 7285 10865
rect 7615 10535 7677 10865
rect 7223 10487 7677 10535
rect 7694 10487 7700 10913
rect 7200 10481 7700 10487
rect 7750 10913 7814 10919
rect 7750 10487 7756 10913
rect 7773 10886 7814 10913
rect 8186 10919 8219 10921
rect 8331 10944 8769 10950
rect 8331 10927 8337 10944
rect 8763 10927 8769 10944
rect 8331 10921 8769 10927
rect 8329 10919 8771 10921
rect 8881 10944 9319 10950
rect 8881 10927 8887 10944
rect 9313 10927 9319 10944
rect 8881 10921 9319 10927
rect 8881 10919 8914 10921
rect 8186 10913 8250 10919
rect 8186 10886 8227 10913
rect 7773 10514 7779 10886
rect 8221 10514 8227 10886
rect 7773 10487 7814 10514
rect 7750 10481 7814 10487
rect 7086 10479 7119 10481
rect 6681 10473 7119 10479
rect 6681 10456 6687 10473
rect 7113 10456 7119 10473
rect 6681 10450 7119 10456
rect 7229 10479 7671 10481
rect 7231 10473 7669 10479
rect 7231 10456 7237 10473
rect 7663 10456 7669 10473
rect 7231 10450 7669 10456
rect 7781 10479 7814 10481
rect 8186 10487 8227 10514
rect 8244 10487 8250 10913
rect 8186 10481 8250 10487
rect 8300 10913 8800 10919
rect 8300 10487 8306 10913
rect 8323 10865 8777 10913
rect 8323 10535 8385 10865
rect 8715 10535 8777 10865
rect 8323 10487 8777 10535
rect 8794 10487 8800 10913
rect 8300 10481 8800 10487
rect 8850 10913 8914 10919
rect 8850 10487 8856 10913
rect 8873 10886 8914 10913
rect 9286 10919 9319 10921
rect 9431 10944 9869 10950
rect 9431 10927 9437 10944
rect 9863 10927 9869 10944
rect 9431 10921 9869 10927
rect 9429 10919 9871 10921
rect 9981 10944 10419 10950
rect 9981 10927 9987 10944
rect 10413 10927 10419 10944
rect 9981 10921 10419 10927
rect 9981 10919 10014 10921
rect 9286 10913 9350 10919
rect 9286 10886 9327 10913
rect 8873 10514 8879 10886
rect 9321 10514 9327 10886
rect 8873 10487 8914 10514
rect 8850 10481 8914 10487
rect 8186 10479 8219 10481
rect 7781 10473 8219 10479
rect 7781 10456 7787 10473
rect 8213 10456 8219 10473
rect 7781 10450 8219 10456
rect 8329 10479 8771 10481
rect 8331 10473 8769 10479
rect 8331 10456 8337 10473
rect 8763 10456 8769 10473
rect 8331 10450 8769 10456
rect 8881 10479 8914 10481
rect 9286 10487 9327 10514
rect 9344 10487 9350 10913
rect 9286 10481 9350 10487
rect 9400 10913 9900 10919
rect 9400 10487 9406 10913
rect 9423 10865 9877 10913
rect 9423 10535 9485 10865
rect 9815 10535 9877 10865
rect 9423 10487 9877 10535
rect 9894 10487 9900 10913
rect 9400 10481 9900 10487
rect 9950 10913 10014 10919
rect 9950 10487 9956 10913
rect 9973 10886 10014 10913
rect 10386 10919 10419 10921
rect 10531 10944 10969 10950
rect 10531 10927 10537 10944
rect 10963 10927 10969 10944
rect 10531 10921 10969 10927
rect 10529 10919 10971 10921
rect 11081 10944 11519 10950
rect 11081 10927 11087 10944
rect 11513 10927 11519 10944
rect 11081 10921 11519 10927
rect 11081 10919 11114 10921
rect 10386 10913 10450 10919
rect 10386 10886 10427 10913
rect 9973 10514 9979 10886
rect 10421 10514 10427 10886
rect 9973 10487 10014 10514
rect 9950 10481 10014 10487
rect 9286 10479 9319 10481
rect 8881 10473 9319 10479
rect 8881 10456 8887 10473
rect 9313 10456 9319 10473
rect 8881 10450 9319 10456
rect 9429 10479 9871 10481
rect 9431 10473 9869 10479
rect 9431 10456 9437 10473
rect 9863 10456 9869 10473
rect 9431 10450 9869 10456
rect 9981 10479 10014 10481
rect 10386 10487 10427 10514
rect 10444 10487 10450 10913
rect 10386 10481 10450 10487
rect 10500 10913 11000 10919
rect 10500 10487 10506 10913
rect 10523 10865 10977 10913
rect 10523 10535 10585 10865
rect 10915 10535 10977 10865
rect 10523 10487 10977 10535
rect 10994 10487 11000 10913
rect 10500 10481 11000 10487
rect 11050 10913 11114 10919
rect 11050 10487 11056 10913
rect 11073 10886 11114 10913
rect 11486 10919 11519 10921
rect 11631 10944 12069 10950
rect 11631 10927 11637 10944
rect 12063 10927 12069 10944
rect 11631 10921 12069 10927
rect 11629 10919 12071 10921
rect 12181 10944 12619 10950
rect 12181 10927 12187 10944
rect 12613 10927 12619 10944
rect 12181 10921 12619 10927
rect 12181 10919 12214 10921
rect 11486 10913 11550 10919
rect 11486 10886 11527 10913
rect 11073 10514 11079 10886
rect 11521 10514 11527 10886
rect 11073 10487 11114 10514
rect 11050 10481 11114 10487
rect 10386 10479 10419 10481
rect 9981 10473 10419 10479
rect 9981 10456 9987 10473
rect 10413 10456 10419 10473
rect 9981 10450 10419 10456
rect 10529 10479 10971 10481
rect 10531 10473 10969 10479
rect 10531 10456 10537 10473
rect 10963 10456 10969 10473
rect 10531 10450 10969 10456
rect 11081 10479 11114 10481
rect 11486 10487 11527 10514
rect 11544 10487 11550 10913
rect 11486 10481 11550 10487
rect 11600 10913 12100 10919
rect 11600 10487 11606 10913
rect 11623 10865 12077 10913
rect 11623 10535 11685 10865
rect 12015 10535 12077 10865
rect 11623 10487 12077 10535
rect 12094 10487 12100 10913
rect 11600 10481 12100 10487
rect 12150 10913 12214 10919
rect 12150 10487 12156 10913
rect 12173 10886 12214 10913
rect 12586 10919 12619 10921
rect 12731 10944 13169 10950
rect 12731 10927 12737 10944
rect 13163 10927 13169 10944
rect 12731 10921 13169 10927
rect 12729 10919 13171 10921
rect 13281 10944 13719 10950
rect 13281 10927 13287 10944
rect 13713 10927 13719 10944
rect 13281 10921 13719 10927
rect 13281 10919 13314 10921
rect 12586 10913 12650 10919
rect 12586 10886 12627 10913
rect 12173 10514 12179 10886
rect 12621 10514 12627 10886
rect 12173 10487 12214 10514
rect 12150 10481 12214 10487
rect 11486 10479 11519 10481
rect 11081 10473 11519 10479
rect 11081 10456 11087 10473
rect 11513 10456 11519 10473
rect 11081 10450 11519 10456
rect 11629 10479 12071 10481
rect 11631 10473 12069 10479
rect 11631 10456 11637 10473
rect 12063 10456 12069 10473
rect 11631 10450 12069 10456
rect 12181 10479 12214 10481
rect 12586 10487 12627 10514
rect 12644 10487 12650 10913
rect 12586 10481 12650 10487
rect 12700 10913 13200 10919
rect 12700 10487 12706 10913
rect 12723 10865 13177 10913
rect 12723 10535 12785 10865
rect 13115 10535 13177 10865
rect 12723 10487 13177 10535
rect 13194 10487 13200 10913
rect 12700 10481 13200 10487
rect 13250 10913 13314 10919
rect 13250 10487 13256 10913
rect 13273 10886 13314 10913
rect 13273 10514 13279 10886
rect 13273 10487 13314 10514
rect 13250 10481 13314 10487
rect 12586 10479 12619 10481
rect 12181 10473 12619 10479
rect 12181 10456 12187 10473
rect 12613 10456 12619 10473
rect 12181 10450 12619 10456
rect 12729 10479 13171 10481
rect 12731 10473 13169 10479
rect 12731 10456 12737 10473
rect 13163 10456 13169 10473
rect 12731 10450 13169 10456
rect 13281 10479 13314 10481
rect 13281 10473 13719 10479
rect 13281 10456 13287 10473
rect 13713 10456 13719 10473
rect 13281 10450 13719 10456
rect -469 10394 -31 10400
rect -469 10377 -463 10394
rect -37 10377 -31 10394
rect -469 10371 -31 10377
rect -64 10369 -31 10371
rect 81 10394 519 10400
rect 81 10377 87 10394
rect 513 10377 519 10394
rect 81 10371 519 10377
rect 79 10369 521 10371
rect 631 10394 1069 10400
rect 631 10377 637 10394
rect 1063 10377 1069 10394
rect 631 10371 1069 10377
rect 631 10369 664 10371
rect -64 10363 0 10369
rect -64 10336 -23 10363
rect -29 9964 -23 10336
rect -64 9937 -23 9964
rect -6 9937 0 10363
rect -64 9931 0 9937
rect 50 10363 550 10369
rect 50 9937 56 10363
rect 73 10315 527 10363
rect 73 9985 135 10315
rect 465 9985 527 10315
rect 73 9937 527 9985
rect 544 9937 550 10363
rect 50 9931 550 9937
rect 600 10363 664 10369
rect 600 9937 606 10363
rect 623 10336 664 10363
rect 1036 10369 1069 10371
rect 1181 10394 1619 10400
rect 1181 10377 1187 10394
rect 1613 10377 1619 10394
rect 1181 10371 1619 10377
rect 1179 10369 1621 10371
rect 1731 10394 2169 10400
rect 1731 10377 1737 10394
rect 2163 10377 2169 10394
rect 1731 10371 2169 10377
rect 1731 10369 1764 10371
rect 1036 10363 1100 10369
rect 1036 10336 1077 10363
rect 623 9964 629 10336
rect 1071 9964 1077 10336
rect 623 9937 664 9964
rect 600 9931 664 9937
rect -64 9929 -31 9931
rect -469 9923 -31 9929
rect -469 9906 -463 9923
rect -37 9906 -31 9923
rect -469 9900 -31 9906
rect 79 9929 521 9931
rect 81 9923 519 9929
rect 81 9906 87 9923
rect 513 9906 519 9923
rect 81 9900 519 9906
rect 631 9929 664 9931
rect 1036 9937 1077 9964
rect 1094 9937 1100 10363
rect 1036 9931 1100 9937
rect 1150 10363 1650 10369
rect 1150 9937 1156 10363
rect 1173 10315 1627 10363
rect 1173 9985 1235 10315
rect 1565 9985 1627 10315
rect 1173 9937 1627 9985
rect 1644 9937 1650 10363
rect 1150 9931 1650 9937
rect 1700 10363 1764 10369
rect 1700 9937 1706 10363
rect 1723 10336 1764 10363
rect 2136 10369 2169 10371
rect 2281 10394 2719 10400
rect 2281 10377 2287 10394
rect 2713 10377 2719 10394
rect 2281 10371 2719 10377
rect 2279 10369 2721 10371
rect 2831 10394 3269 10400
rect 2831 10377 2837 10394
rect 3263 10377 3269 10394
rect 2831 10371 3269 10377
rect 2831 10369 2864 10371
rect 2136 10363 2200 10369
rect 2136 10336 2177 10363
rect 1723 9964 1729 10336
rect 2171 9964 2177 10336
rect 1723 9937 1764 9964
rect 1700 9931 1764 9937
rect 1036 9929 1069 9931
rect 631 9923 1069 9929
rect 631 9906 637 9923
rect 1063 9906 1069 9923
rect 631 9900 1069 9906
rect 1179 9929 1621 9931
rect 1181 9923 1619 9929
rect 1181 9906 1187 9923
rect 1613 9906 1619 9923
rect 1181 9900 1619 9906
rect 1731 9929 1764 9931
rect 2136 9937 2177 9964
rect 2194 9937 2200 10363
rect 2136 9931 2200 9937
rect 2250 10363 2750 10369
rect 2250 9937 2256 10363
rect 2273 10315 2727 10363
rect 2273 9985 2335 10315
rect 2665 9985 2727 10315
rect 2273 9937 2727 9985
rect 2744 9937 2750 10363
rect 2250 9931 2750 9937
rect 2800 10363 2864 10369
rect 2800 9937 2806 10363
rect 2823 10336 2864 10363
rect 3236 10369 3269 10371
rect 3381 10394 3819 10400
rect 3381 10377 3387 10394
rect 3813 10377 3819 10394
rect 3381 10371 3819 10377
rect 3379 10369 3821 10371
rect 3931 10394 4369 10400
rect 3931 10377 3937 10394
rect 4363 10377 4369 10394
rect 3931 10371 4369 10377
rect 3931 10369 3964 10371
rect 3236 10363 3300 10369
rect 3236 10336 3277 10363
rect 2823 9964 2829 10336
rect 3271 9964 3277 10336
rect 2823 9937 2864 9964
rect 2800 9931 2864 9937
rect 2136 9929 2169 9931
rect 1731 9923 2169 9929
rect 1731 9906 1737 9923
rect 2163 9906 2169 9923
rect 1731 9900 2169 9906
rect 2279 9929 2721 9931
rect 2281 9923 2719 9929
rect 2281 9906 2287 9923
rect 2713 9906 2719 9923
rect 2281 9900 2719 9906
rect 2831 9929 2864 9931
rect 3236 9937 3277 9964
rect 3294 9937 3300 10363
rect 3236 9931 3300 9937
rect 3350 10363 3850 10369
rect 3350 9937 3356 10363
rect 3373 10315 3827 10363
rect 3373 9985 3435 10315
rect 3765 9985 3827 10315
rect 3373 9937 3827 9985
rect 3844 9937 3850 10363
rect 3350 9931 3850 9937
rect 3900 10363 3964 10369
rect 3900 9937 3906 10363
rect 3923 10336 3964 10363
rect 4336 10369 4369 10371
rect 4481 10394 4919 10400
rect 4481 10377 4487 10394
rect 4913 10377 4919 10394
rect 4481 10371 4919 10377
rect 4479 10369 4921 10371
rect 5031 10394 5469 10400
rect 5031 10377 5037 10394
rect 5463 10377 5469 10394
rect 5031 10371 5469 10377
rect 5031 10369 5064 10371
rect 4336 10363 4400 10369
rect 4336 10336 4377 10363
rect 3923 9964 3929 10336
rect 4371 9964 4377 10336
rect 3923 9937 3964 9964
rect 3900 9931 3964 9937
rect 3236 9929 3269 9931
rect 2831 9923 3269 9929
rect 2831 9906 2837 9923
rect 3263 9906 3269 9923
rect 2831 9900 3269 9906
rect 3379 9929 3821 9931
rect 3381 9923 3819 9929
rect 3381 9906 3387 9923
rect 3813 9906 3819 9923
rect 3381 9900 3819 9906
rect 3931 9929 3964 9931
rect 4336 9937 4377 9964
rect 4394 9937 4400 10363
rect 4336 9931 4400 9937
rect 4450 10363 4950 10369
rect 4450 9937 4456 10363
rect 4473 10315 4927 10363
rect 4473 9985 4535 10315
rect 4865 9985 4927 10315
rect 4473 9937 4927 9985
rect 4944 9937 4950 10363
rect 4450 9931 4950 9937
rect 5000 10363 5064 10369
rect 5000 9937 5006 10363
rect 5023 10336 5064 10363
rect 5436 10369 5469 10371
rect 5581 10394 6019 10400
rect 5581 10377 5587 10394
rect 6013 10377 6019 10394
rect 5581 10371 6019 10377
rect 5579 10369 6021 10371
rect 6131 10394 6569 10400
rect 6131 10377 6137 10394
rect 6563 10377 6569 10394
rect 6131 10371 6569 10377
rect 6131 10369 6164 10371
rect 5436 10363 5500 10369
rect 5436 10336 5477 10363
rect 5023 9964 5029 10336
rect 5471 9964 5477 10336
rect 5023 9937 5064 9964
rect 5000 9931 5064 9937
rect 4336 9929 4369 9931
rect 3931 9923 4369 9929
rect 3931 9906 3937 9923
rect 4363 9906 4369 9923
rect 3931 9900 4369 9906
rect 4479 9929 4921 9931
rect 4481 9923 4919 9929
rect 4481 9906 4487 9923
rect 4913 9906 4919 9923
rect 4481 9900 4919 9906
rect 5031 9929 5064 9931
rect 5436 9937 5477 9964
rect 5494 9937 5500 10363
rect 5436 9931 5500 9937
rect 5550 10363 6050 10369
rect 5550 9937 5556 10363
rect 5573 10315 6027 10363
rect 5573 9985 5635 10315
rect 5965 9985 6027 10315
rect 5573 9937 6027 9985
rect 6044 9937 6050 10363
rect 5550 9931 6050 9937
rect 6100 10363 6164 10369
rect 6100 9937 6106 10363
rect 6123 10336 6164 10363
rect 6536 10369 6569 10371
rect 6681 10394 7119 10400
rect 6681 10377 6687 10394
rect 7113 10377 7119 10394
rect 6681 10371 7119 10377
rect 6679 10369 7121 10371
rect 7231 10394 7669 10400
rect 7231 10377 7237 10394
rect 7663 10377 7669 10394
rect 7231 10371 7669 10377
rect 7231 10369 7264 10371
rect 6536 10363 6600 10369
rect 6536 10336 6577 10363
rect 6123 9964 6129 10336
rect 6571 9964 6577 10336
rect 6123 9937 6164 9964
rect 6100 9931 6164 9937
rect 5436 9929 5469 9931
rect 5031 9923 5469 9929
rect 5031 9906 5037 9923
rect 5463 9906 5469 9923
rect 5031 9900 5469 9906
rect 5579 9929 6021 9931
rect 5581 9923 6019 9929
rect 5581 9906 5587 9923
rect 6013 9906 6019 9923
rect 5581 9900 6019 9906
rect 6131 9929 6164 9931
rect 6536 9937 6577 9964
rect 6594 9937 6600 10363
rect 6536 9931 6600 9937
rect 6650 10363 7150 10369
rect 6650 9937 6656 10363
rect 6673 10315 7127 10363
rect 6673 9985 6735 10315
rect 7065 9985 7127 10315
rect 6673 9937 7127 9985
rect 7144 9937 7150 10363
rect 6650 9931 7150 9937
rect 7200 10363 7264 10369
rect 7200 9937 7206 10363
rect 7223 10336 7264 10363
rect 7636 10369 7669 10371
rect 7781 10394 8219 10400
rect 7781 10377 7787 10394
rect 8213 10377 8219 10394
rect 7781 10371 8219 10377
rect 7779 10369 8221 10371
rect 8331 10394 8769 10400
rect 8331 10377 8337 10394
rect 8763 10377 8769 10394
rect 8331 10371 8769 10377
rect 8331 10369 8364 10371
rect 7636 10363 7700 10369
rect 7636 10336 7677 10363
rect 7223 9964 7229 10336
rect 7671 9964 7677 10336
rect 7223 9937 7264 9964
rect 7200 9931 7264 9937
rect 6536 9929 6569 9931
rect 6131 9923 6569 9929
rect 6131 9906 6137 9923
rect 6563 9906 6569 9923
rect 6131 9900 6569 9906
rect 6679 9929 7121 9931
rect 6681 9923 7119 9929
rect 6681 9906 6687 9923
rect 7113 9906 7119 9923
rect 6681 9900 7119 9906
rect 7231 9929 7264 9931
rect 7636 9937 7677 9964
rect 7694 9937 7700 10363
rect 7636 9931 7700 9937
rect 7750 10363 8250 10369
rect 7750 9937 7756 10363
rect 7773 10315 8227 10363
rect 7773 9985 7835 10315
rect 8165 9985 8227 10315
rect 7773 9937 8227 9985
rect 8244 9937 8250 10363
rect 7750 9931 8250 9937
rect 8300 10363 8364 10369
rect 8300 9937 8306 10363
rect 8323 10336 8364 10363
rect 8736 10369 8769 10371
rect 8881 10394 9319 10400
rect 8881 10377 8887 10394
rect 9313 10377 9319 10394
rect 8881 10371 9319 10377
rect 8879 10369 9321 10371
rect 9431 10394 9869 10400
rect 9431 10377 9437 10394
rect 9863 10377 9869 10394
rect 9431 10371 9869 10377
rect 9431 10369 9464 10371
rect 8736 10363 8800 10369
rect 8736 10336 8777 10363
rect 8323 9964 8329 10336
rect 8771 9964 8777 10336
rect 8323 9937 8364 9964
rect 8300 9931 8364 9937
rect 7636 9929 7669 9931
rect 7231 9923 7669 9929
rect 7231 9906 7237 9923
rect 7663 9906 7669 9923
rect 7231 9900 7669 9906
rect 7779 9929 8221 9931
rect 7781 9923 8219 9929
rect 7781 9906 7787 9923
rect 8213 9906 8219 9923
rect 7781 9900 8219 9906
rect 8331 9929 8364 9931
rect 8736 9937 8777 9964
rect 8794 9937 8800 10363
rect 8736 9931 8800 9937
rect 8850 10363 9350 10369
rect 8850 9937 8856 10363
rect 8873 10315 9327 10363
rect 8873 9985 8935 10315
rect 9265 9985 9327 10315
rect 8873 9937 9327 9985
rect 9344 9937 9350 10363
rect 8850 9931 9350 9937
rect 9400 10363 9464 10369
rect 9400 9937 9406 10363
rect 9423 10336 9464 10363
rect 9836 10369 9869 10371
rect 9981 10394 10419 10400
rect 9981 10377 9987 10394
rect 10413 10377 10419 10394
rect 9981 10371 10419 10377
rect 9979 10369 10421 10371
rect 10531 10394 10969 10400
rect 10531 10377 10537 10394
rect 10963 10377 10969 10394
rect 10531 10371 10969 10377
rect 10531 10369 10564 10371
rect 9836 10363 9900 10369
rect 9836 10336 9877 10363
rect 9423 9964 9429 10336
rect 9871 9964 9877 10336
rect 9423 9937 9464 9964
rect 9400 9931 9464 9937
rect 8736 9929 8769 9931
rect 8331 9923 8769 9929
rect 8331 9906 8337 9923
rect 8763 9906 8769 9923
rect 8331 9900 8769 9906
rect 8879 9929 9321 9931
rect 8881 9923 9319 9929
rect 8881 9906 8887 9923
rect 9313 9906 9319 9923
rect 8881 9900 9319 9906
rect 9431 9929 9464 9931
rect 9836 9937 9877 9964
rect 9894 9937 9900 10363
rect 9836 9931 9900 9937
rect 9950 10363 10450 10369
rect 9950 9937 9956 10363
rect 9973 10315 10427 10363
rect 9973 9985 10035 10315
rect 10365 9985 10427 10315
rect 9973 9937 10427 9985
rect 10444 9937 10450 10363
rect 9950 9931 10450 9937
rect 10500 10363 10564 10369
rect 10500 9937 10506 10363
rect 10523 10336 10564 10363
rect 10936 10369 10969 10371
rect 11081 10394 11519 10400
rect 11081 10377 11087 10394
rect 11513 10377 11519 10394
rect 11081 10371 11519 10377
rect 11079 10369 11521 10371
rect 11631 10394 12069 10400
rect 11631 10377 11637 10394
rect 12063 10377 12069 10394
rect 11631 10371 12069 10377
rect 11631 10369 11664 10371
rect 10936 10363 11000 10369
rect 10936 10336 10977 10363
rect 10523 9964 10529 10336
rect 10971 9964 10977 10336
rect 10523 9937 10564 9964
rect 10500 9931 10564 9937
rect 9836 9929 9869 9931
rect 9431 9923 9869 9929
rect 9431 9906 9437 9923
rect 9863 9906 9869 9923
rect 9431 9900 9869 9906
rect 9979 9929 10421 9931
rect 9981 9923 10419 9929
rect 9981 9906 9987 9923
rect 10413 9906 10419 9923
rect 9981 9900 10419 9906
rect 10531 9929 10564 9931
rect 10936 9937 10977 9964
rect 10994 9937 11000 10363
rect 10936 9931 11000 9937
rect 11050 10363 11550 10369
rect 11050 9937 11056 10363
rect 11073 10315 11527 10363
rect 11073 9985 11135 10315
rect 11465 9985 11527 10315
rect 11073 9937 11527 9985
rect 11544 9937 11550 10363
rect 11050 9931 11550 9937
rect 11600 10363 11664 10369
rect 11600 9937 11606 10363
rect 11623 10336 11664 10363
rect 12036 10369 12069 10371
rect 12181 10394 12619 10400
rect 12181 10377 12187 10394
rect 12613 10377 12619 10394
rect 12181 10371 12619 10377
rect 12179 10369 12621 10371
rect 12731 10394 13169 10400
rect 12731 10377 12737 10394
rect 13163 10377 13169 10394
rect 12731 10371 13169 10377
rect 12731 10369 12764 10371
rect 12036 10363 12100 10369
rect 12036 10336 12077 10363
rect 11623 9964 11629 10336
rect 12071 9964 12077 10336
rect 11623 9937 11664 9964
rect 11600 9931 11664 9937
rect 10936 9929 10969 9931
rect 10531 9923 10969 9929
rect 10531 9906 10537 9923
rect 10963 9906 10969 9923
rect 10531 9900 10969 9906
rect 11079 9929 11521 9931
rect 11081 9923 11519 9929
rect 11081 9906 11087 9923
rect 11513 9906 11519 9923
rect 11081 9900 11519 9906
rect 11631 9929 11664 9931
rect 12036 9937 12077 9964
rect 12094 9937 12100 10363
rect 12036 9931 12100 9937
rect 12150 10363 12650 10369
rect 12150 9937 12156 10363
rect 12173 10315 12627 10363
rect 12173 9985 12235 10315
rect 12565 9985 12627 10315
rect 12173 9937 12627 9985
rect 12644 9937 12650 10363
rect 12150 9931 12650 9937
rect 12700 10363 12764 10369
rect 12700 9937 12706 10363
rect 12723 10336 12764 10363
rect 13136 10369 13169 10371
rect 13281 10394 13719 10400
rect 13281 10377 13287 10394
rect 13713 10377 13719 10394
rect 13281 10371 13719 10377
rect 13279 10369 13721 10371
rect 13136 10363 13200 10369
rect 13136 10336 13177 10363
rect 12723 9964 12729 10336
rect 13171 9964 13177 10336
rect 12723 9937 12764 9964
rect 12700 9931 12764 9937
rect 12036 9929 12069 9931
rect 11631 9923 12069 9929
rect 11631 9906 11637 9923
rect 12063 9906 12069 9923
rect 11631 9900 12069 9906
rect 12179 9929 12621 9931
rect 12181 9923 12619 9929
rect 12181 9906 12187 9923
rect 12613 9906 12619 9923
rect 12181 9900 12619 9906
rect 12731 9929 12764 9931
rect 13136 9937 13177 9964
rect 13194 9937 13200 10363
rect 13136 9931 13200 9937
rect 13250 10363 13721 10369
rect 13250 9937 13256 10363
rect 13273 10315 13721 10363
rect 13273 9985 13335 10315
rect 13665 9985 13721 10315
rect 13273 9937 13721 9985
rect 13250 9931 13721 9937
rect 13136 9929 13169 9931
rect 12731 9923 13169 9929
rect 12731 9906 12737 9923
rect 13163 9906 13169 9923
rect 12731 9900 13169 9906
rect 13279 9929 13721 9931
rect 13281 9923 13719 9929
rect 13281 9906 13287 9923
rect 13713 9906 13719 9923
rect 13281 9900 13719 9906
rect -469 9844 -31 9850
rect -469 9827 -463 9844
rect -37 9827 -31 9844
rect -469 9821 -31 9827
rect -471 9819 -29 9821
rect 81 9844 519 9850
rect 81 9827 87 9844
rect 513 9827 519 9844
rect 81 9821 519 9827
rect 81 9819 114 9821
rect -471 9813 0 9819
rect -471 9765 -23 9813
rect -471 9435 -415 9765
rect -85 9435 -23 9765
rect -471 9387 -23 9435
rect -6 9387 0 9813
rect -471 9381 0 9387
rect 50 9813 114 9819
rect 50 9387 56 9813
rect 73 9786 114 9813
rect 486 9819 519 9821
rect 631 9844 1069 9850
rect 631 9827 637 9844
rect 1063 9827 1069 9844
rect 631 9821 1069 9827
rect 629 9819 1071 9821
rect 1181 9844 1619 9850
rect 1181 9827 1187 9844
rect 1613 9827 1619 9844
rect 1181 9821 1619 9827
rect 1181 9819 1214 9821
rect 486 9813 550 9819
rect 486 9786 527 9813
rect 73 9414 79 9786
rect 521 9414 527 9786
rect 73 9387 114 9414
rect 50 9381 114 9387
rect -471 9379 -29 9381
rect -469 9373 -31 9379
rect -469 9356 -463 9373
rect -37 9356 -31 9373
rect -469 9350 -31 9356
rect 81 9379 114 9381
rect 486 9387 527 9414
rect 544 9387 550 9813
rect 486 9381 550 9387
rect 600 9813 1100 9819
rect 600 9387 606 9813
rect 623 9765 1077 9813
rect 623 9435 685 9765
rect 1015 9435 1077 9765
rect 623 9387 1077 9435
rect 1094 9387 1100 9813
rect 600 9381 1100 9387
rect 1150 9813 1214 9819
rect 1150 9387 1156 9813
rect 1173 9786 1214 9813
rect 1586 9819 1619 9821
rect 1731 9844 2169 9850
rect 1731 9827 1737 9844
rect 2163 9827 2169 9844
rect 1731 9821 2169 9827
rect 1729 9819 2171 9821
rect 2281 9844 2719 9850
rect 2281 9827 2287 9844
rect 2713 9827 2719 9844
rect 2281 9821 2719 9827
rect 2281 9819 2314 9821
rect 1586 9813 1650 9819
rect 1586 9786 1627 9813
rect 1173 9414 1179 9786
rect 1621 9414 1627 9786
rect 1173 9387 1214 9414
rect 1150 9381 1214 9387
rect 486 9379 519 9381
rect 81 9373 519 9379
rect 81 9356 87 9373
rect 513 9356 519 9373
rect 81 9350 519 9356
rect 629 9379 1071 9381
rect 631 9373 1069 9379
rect 631 9356 637 9373
rect 1063 9356 1069 9373
rect 631 9350 1069 9356
rect 1181 9379 1214 9381
rect 1586 9387 1627 9414
rect 1644 9387 1650 9813
rect 1586 9381 1650 9387
rect 1700 9813 2200 9819
rect 1700 9387 1706 9813
rect 1723 9765 2177 9813
rect 1723 9435 1785 9765
rect 2115 9435 2177 9765
rect 1723 9387 2177 9435
rect 2194 9387 2200 9813
rect 1700 9381 2200 9387
rect 2250 9813 2314 9819
rect 2250 9387 2256 9813
rect 2273 9786 2314 9813
rect 2686 9819 2719 9821
rect 2831 9844 3269 9850
rect 2831 9827 2837 9844
rect 3263 9827 3269 9844
rect 2831 9821 3269 9827
rect 2829 9819 3271 9821
rect 3381 9844 3819 9850
rect 3381 9827 3387 9844
rect 3813 9827 3819 9844
rect 3381 9821 3819 9827
rect 3381 9819 3414 9821
rect 2686 9813 2750 9819
rect 2686 9786 2727 9813
rect 2273 9414 2279 9786
rect 2721 9414 2727 9786
rect 2273 9387 2314 9414
rect 2250 9381 2314 9387
rect 1586 9379 1619 9381
rect 1181 9373 1619 9379
rect 1181 9356 1187 9373
rect 1613 9356 1619 9373
rect 1181 9350 1619 9356
rect 1729 9379 2171 9381
rect 1731 9373 2169 9379
rect 1731 9356 1737 9373
rect 2163 9356 2169 9373
rect 1731 9350 2169 9356
rect 2281 9379 2314 9381
rect 2686 9387 2727 9414
rect 2744 9387 2750 9813
rect 2686 9381 2750 9387
rect 2800 9813 3300 9819
rect 2800 9387 2806 9813
rect 2823 9765 3277 9813
rect 2823 9435 2885 9765
rect 3215 9435 3277 9765
rect 2823 9387 3277 9435
rect 3294 9387 3300 9813
rect 2800 9381 3300 9387
rect 3350 9813 3414 9819
rect 3350 9387 3356 9813
rect 3373 9786 3414 9813
rect 3786 9819 3819 9821
rect 3931 9844 4369 9850
rect 3931 9827 3937 9844
rect 4363 9827 4369 9844
rect 3931 9821 4369 9827
rect 3929 9819 4371 9821
rect 4481 9844 4919 9850
rect 4481 9827 4487 9844
rect 4913 9827 4919 9844
rect 4481 9821 4919 9827
rect 4481 9819 4514 9821
rect 3786 9813 3850 9819
rect 3786 9786 3827 9813
rect 3373 9414 3379 9786
rect 3821 9414 3827 9786
rect 3373 9387 3414 9414
rect 3350 9381 3414 9387
rect 2686 9379 2719 9381
rect 2281 9373 2719 9379
rect 2281 9356 2287 9373
rect 2713 9356 2719 9373
rect 2281 9350 2719 9356
rect 2829 9379 3271 9381
rect 2831 9373 3269 9379
rect 2831 9356 2837 9373
rect 3263 9356 3269 9373
rect 2831 9350 3269 9356
rect 3381 9379 3414 9381
rect 3786 9387 3827 9414
rect 3844 9387 3850 9813
rect 3786 9381 3850 9387
rect 3900 9813 4400 9819
rect 3900 9387 3906 9813
rect 3923 9765 4377 9813
rect 3923 9435 3985 9765
rect 4315 9435 4377 9765
rect 3923 9387 4377 9435
rect 4394 9387 4400 9813
rect 3900 9381 4400 9387
rect 4450 9813 4514 9819
rect 4450 9387 4456 9813
rect 4473 9786 4514 9813
rect 4886 9819 4919 9821
rect 5031 9844 5469 9850
rect 5031 9827 5037 9844
rect 5463 9827 5469 9844
rect 5031 9821 5469 9827
rect 5029 9819 5471 9821
rect 5581 9844 6019 9850
rect 5581 9827 5587 9844
rect 6013 9827 6019 9844
rect 5581 9821 6019 9827
rect 5581 9819 5614 9821
rect 4886 9813 4950 9819
rect 4886 9786 4927 9813
rect 4473 9414 4479 9786
rect 4921 9414 4927 9786
rect 4473 9387 4514 9414
rect 4450 9381 4514 9387
rect 3786 9379 3819 9381
rect 3381 9373 3819 9379
rect 3381 9356 3387 9373
rect 3813 9356 3819 9373
rect 3381 9350 3819 9356
rect 3929 9379 4371 9381
rect 3931 9373 4369 9379
rect 3931 9356 3937 9373
rect 4363 9356 4369 9373
rect 3931 9350 4369 9356
rect 4481 9379 4514 9381
rect 4886 9387 4927 9414
rect 4944 9387 4950 9813
rect 4886 9381 4950 9387
rect 5000 9813 5500 9819
rect 5000 9387 5006 9813
rect 5023 9765 5477 9813
rect 5023 9435 5085 9765
rect 5415 9435 5477 9765
rect 5023 9387 5477 9435
rect 5494 9387 5500 9813
rect 5000 9381 5500 9387
rect 5550 9813 5614 9819
rect 5550 9387 5556 9813
rect 5573 9786 5614 9813
rect 5986 9819 6019 9821
rect 6131 9844 6569 9850
rect 6131 9827 6137 9844
rect 6563 9827 6569 9844
rect 6131 9821 6569 9827
rect 6129 9819 6571 9821
rect 6681 9844 7119 9850
rect 6681 9827 6687 9844
rect 7113 9827 7119 9844
rect 6681 9821 7119 9827
rect 6681 9819 6714 9821
rect 5986 9813 6050 9819
rect 5986 9786 6027 9813
rect 5573 9414 5579 9786
rect 6021 9414 6027 9786
rect 5573 9387 5614 9414
rect 5550 9381 5614 9387
rect 4886 9379 4919 9381
rect 4481 9373 4919 9379
rect 4481 9356 4487 9373
rect 4913 9356 4919 9373
rect 4481 9350 4919 9356
rect 5029 9379 5471 9381
rect 5031 9373 5469 9379
rect 5031 9356 5037 9373
rect 5463 9356 5469 9373
rect 5031 9350 5469 9356
rect 5581 9379 5614 9381
rect 5986 9387 6027 9414
rect 6044 9387 6050 9813
rect 5986 9381 6050 9387
rect 6100 9813 6600 9819
rect 6100 9387 6106 9813
rect 6123 9765 6577 9813
rect 6123 9435 6185 9765
rect 6515 9435 6577 9765
rect 6123 9387 6577 9435
rect 6594 9387 6600 9813
rect 6100 9381 6600 9387
rect 6650 9813 6714 9819
rect 6650 9387 6656 9813
rect 6673 9786 6714 9813
rect 7086 9819 7119 9821
rect 7231 9844 7669 9850
rect 7231 9827 7237 9844
rect 7663 9827 7669 9844
rect 7231 9821 7669 9827
rect 7229 9819 7671 9821
rect 7781 9844 8219 9850
rect 7781 9827 7787 9844
rect 8213 9827 8219 9844
rect 7781 9821 8219 9827
rect 7781 9819 7814 9821
rect 7086 9813 7150 9819
rect 7086 9786 7127 9813
rect 6673 9414 6679 9786
rect 7121 9414 7127 9786
rect 6673 9387 6714 9414
rect 6650 9381 6714 9387
rect 5986 9379 6019 9381
rect 5581 9373 6019 9379
rect 5581 9356 5587 9373
rect 6013 9356 6019 9373
rect 5581 9350 6019 9356
rect 6129 9379 6571 9381
rect 6131 9373 6569 9379
rect 6131 9356 6137 9373
rect 6563 9356 6569 9373
rect 6131 9350 6569 9356
rect 6681 9379 6714 9381
rect 7086 9387 7127 9414
rect 7144 9387 7150 9813
rect 7086 9381 7150 9387
rect 7200 9813 7700 9819
rect 7200 9387 7206 9813
rect 7223 9765 7677 9813
rect 7223 9435 7285 9765
rect 7615 9435 7677 9765
rect 7223 9387 7677 9435
rect 7694 9387 7700 9813
rect 7200 9381 7700 9387
rect 7750 9813 7814 9819
rect 7750 9387 7756 9813
rect 7773 9786 7814 9813
rect 8186 9819 8219 9821
rect 8331 9844 8769 9850
rect 8331 9827 8337 9844
rect 8763 9827 8769 9844
rect 8331 9821 8769 9827
rect 8329 9819 8771 9821
rect 8881 9844 9319 9850
rect 8881 9827 8887 9844
rect 9313 9827 9319 9844
rect 8881 9821 9319 9827
rect 8881 9819 8914 9821
rect 8186 9813 8250 9819
rect 8186 9786 8227 9813
rect 7773 9414 7779 9786
rect 8221 9414 8227 9786
rect 7773 9387 7814 9414
rect 7750 9381 7814 9387
rect 7086 9379 7119 9381
rect 6681 9373 7119 9379
rect 6681 9356 6687 9373
rect 7113 9356 7119 9373
rect 6681 9350 7119 9356
rect 7229 9379 7671 9381
rect 7231 9373 7669 9379
rect 7231 9356 7237 9373
rect 7663 9356 7669 9373
rect 7231 9350 7669 9356
rect 7781 9379 7814 9381
rect 8186 9387 8227 9414
rect 8244 9387 8250 9813
rect 8186 9381 8250 9387
rect 8300 9813 8800 9819
rect 8300 9387 8306 9813
rect 8323 9765 8777 9813
rect 8323 9435 8385 9765
rect 8715 9435 8777 9765
rect 8323 9387 8777 9435
rect 8794 9387 8800 9813
rect 8300 9381 8800 9387
rect 8850 9813 8914 9819
rect 8850 9387 8856 9813
rect 8873 9786 8914 9813
rect 9286 9819 9319 9821
rect 9431 9844 9869 9850
rect 9431 9827 9437 9844
rect 9863 9827 9869 9844
rect 9431 9821 9869 9827
rect 9429 9819 9871 9821
rect 9981 9844 10419 9850
rect 9981 9827 9987 9844
rect 10413 9827 10419 9844
rect 9981 9821 10419 9827
rect 9981 9819 10014 9821
rect 9286 9813 9350 9819
rect 9286 9786 9327 9813
rect 8873 9414 8879 9786
rect 9321 9414 9327 9786
rect 8873 9387 8914 9414
rect 8850 9381 8914 9387
rect 8186 9379 8219 9381
rect 7781 9373 8219 9379
rect 7781 9356 7787 9373
rect 8213 9356 8219 9373
rect 7781 9350 8219 9356
rect 8329 9379 8771 9381
rect 8331 9373 8769 9379
rect 8331 9356 8337 9373
rect 8763 9356 8769 9373
rect 8331 9350 8769 9356
rect 8881 9379 8914 9381
rect 9286 9387 9327 9414
rect 9344 9387 9350 9813
rect 9286 9381 9350 9387
rect 9400 9813 9900 9819
rect 9400 9387 9406 9813
rect 9423 9765 9877 9813
rect 9423 9435 9485 9765
rect 9815 9435 9877 9765
rect 9423 9387 9877 9435
rect 9894 9387 9900 9813
rect 9400 9381 9900 9387
rect 9950 9813 10014 9819
rect 9950 9387 9956 9813
rect 9973 9786 10014 9813
rect 10386 9819 10419 9821
rect 10531 9844 10969 9850
rect 10531 9827 10537 9844
rect 10963 9827 10969 9844
rect 10531 9821 10969 9827
rect 10529 9819 10971 9821
rect 11081 9844 11519 9850
rect 11081 9827 11087 9844
rect 11513 9827 11519 9844
rect 11081 9821 11519 9827
rect 11081 9819 11114 9821
rect 10386 9813 10450 9819
rect 10386 9786 10427 9813
rect 9973 9414 9979 9786
rect 10421 9414 10427 9786
rect 9973 9387 10014 9414
rect 9950 9381 10014 9387
rect 9286 9379 9319 9381
rect 8881 9373 9319 9379
rect 8881 9356 8887 9373
rect 9313 9356 9319 9373
rect 8881 9350 9319 9356
rect 9429 9379 9871 9381
rect 9431 9373 9869 9379
rect 9431 9356 9437 9373
rect 9863 9356 9869 9373
rect 9431 9350 9869 9356
rect 9981 9379 10014 9381
rect 10386 9387 10427 9414
rect 10444 9387 10450 9813
rect 10386 9381 10450 9387
rect 10500 9813 11000 9819
rect 10500 9387 10506 9813
rect 10523 9765 10977 9813
rect 10523 9435 10585 9765
rect 10915 9435 10977 9765
rect 10523 9387 10977 9435
rect 10994 9387 11000 9813
rect 10500 9381 11000 9387
rect 11050 9813 11114 9819
rect 11050 9387 11056 9813
rect 11073 9786 11114 9813
rect 11486 9819 11519 9821
rect 11631 9844 12069 9850
rect 11631 9827 11637 9844
rect 12063 9827 12069 9844
rect 11631 9821 12069 9827
rect 11629 9819 12071 9821
rect 12181 9844 12619 9850
rect 12181 9827 12187 9844
rect 12613 9827 12619 9844
rect 12181 9821 12619 9827
rect 12181 9819 12214 9821
rect 11486 9813 11550 9819
rect 11486 9786 11527 9813
rect 11073 9414 11079 9786
rect 11521 9414 11527 9786
rect 11073 9387 11114 9414
rect 11050 9381 11114 9387
rect 10386 9379 10419 9381
rect 9981 9373 10419 9379
rect 9981 9356 9987 9373
rect 10413 9356 10419 9373
rect 9981 9350 10419 9356
rect 10529 9379 10971 9381
rect 10531 9373 10969 9379
rect 10531 9356 10537 9373
rect 10963 9356 10969 9373
rect 10531 9350 10969 9356
rect 11081 9379 11114 9381
rect 11486 9387 11527 9414
rect 11544 9387 11550 9813
rect 11486 9381 11550 9387
rect 11600 9813 12100 9819
rect 11600 9387 11606 9813
rect 11623 9765 12077 9813
rect 11623 9435 11685 9765
rect 12015 9435 12077 9765
rect 11623 9387 12077 9435
rect 12094 9387 12100 9813
rect 11600 9381 12100 9387
rect 12150 9813 12214 9819
rect 12150 9387 12156 9813
rect 12173 9786 12214 9813
rect 12586 9819 12619 9821
rect 12731 9844 13169 9850
rect 12731 9827 12737 9844
rect 13163 9827 13169 9844
rect 12731 9821 13169 9827
rect 12729 9819 13171 9821
rect 13281 9844 13719 9850
rect 13281 9827 13287 9844
rect 13713 9827 13719 9844
rect 13281 9821 13719 9827
rect 13281 9819 13314 9821
rect 12586 9813 12650 9819
rect 12586 9786 12627 9813
rect 12173 9414 12179 9786
rect 12621 9414 12627 9786
rect 12173 9387 12214 9414
rect 12150 9381 12214 9387
rect 11486 9379 11519 9381
rect 11081 9373 11519 9379
rect 11081 9356 11087 9373
rect 11513 9356 11519 9373
rect 11081 9350 11519 9356
rect 11629 9379 12071 9381
rect 11631 9373 12069 9379
rect 11631 9356 11637 9373
rect 12063 9356 12069 9373
rect 11631 9350 12069 9356
rect 12181 9379 12214 9381
rect 12586 9387 12627 9414
rect 12644 9387 12650 9813
rect 12586 9381 12650 9387
rect 12700 9813 13200 9819
rect 12700 9387 12706 9813
rect 12723 9765 13177 9813
rect 12723 9435 12785 9765
rect 13115 9435 13177 9765
rect 12723 9387 13177 9435
rect 13194 9387 13200 9813
rect 12700 9381 13200 9387
rect 13250 9813 13314 9819
rect 13250 9387 13256 9813
rect 13273 9786 13314 9813
rect 13273 9414 13279 9786
rect 13273 9387 13314 9414
rect 13250 9381 13314 9387
rect 12586 9379 12619 9381
rect 12181 9373 12619 9379
rect 12181 9356 12187 9373
rect 12613 9356 12619 9373
rect 12181 9350 12619 9356
rect 12729 9379 13171 9381
rect 12731 9373 13169 9379
rect 12731 9356 12737 9373
rect 13163 9356 13169 9373
rect 12731 9350 13169 9356
rect 13281 9379 13314 9381
rect 13281 9373 13719 9379
rect 13281 9356 13287 9373
rect 13713 9356 13719 9373
rect 13281 9350 13719 9356
rect -469 9294 -31 9300
rect -469 9277 -463 9294
rect -37 9277 -31 9294
rect -469 9271 -31 9277
rect -64 9269 -31 9271
rect 81 9294 519 9300
rect 81 9277 87 9294
rect 513 9277 519 9294
rect 81 9271 519 9277
rect 79 9269 521 9271
rect 631 9294 1069 9300
rect 631 9277 637 9294
rect 1063 9277 1069 9294
rect 631 9271 1069 9277
rect 631 9269 664 9271
rect -64 9263 0 9269
rect -64 9236 -23 9263
rect -29 8864 -23 9236
rect -64 8837 -23 8864
rect -6 8837 0 9263
rect -64 8831 0 8837
rect 50 9263 550 9269
rect 50 8837 56 9263
rect 73 9215 527 9263
rect 73 8885 135 9215
rect 465 8885 527 9215
rect 73 8837 527 8885
rect 544 8837 550 9263
rect 50 8831 550 8837
rect 600 9263 664 9269
rect 600 8837 606 9263
rect 623 9236 664 9263
rect 1036 9269 1069 9271
rect 1181 9294 1619 9300
rect 1181 9277 1187 9294
rect 1613 9277 1619 9294
rect 1181 9271 1619 9277
rect 1179 9269 1621 9271
rect 1731 9294 2169 9300
rect 1731 9277 1737 9294
rect 2163 9277 2169 9294
rect 1731 9271 2169 9277
rect 1731 9269 1764 9271
rect 1036 9263 1100 9269
rect 1036 9236 1077 9263
rect 623 8864 629 9236
rect 1071 8864 1077 9236
rect 623 8837 664 8864
rect 600 8831 664 8837
rect -64 8829 -31 8831
rect -469 8823 -31 8829
rect -469 8806 -463 8823
rect -37 8806 -31 8823
rect -469 8800 -31 8806
rect 79 8829 521 8831
rect 81 8823 519 8829
rect 81 8806 87 8823
rect 513 8806 519 8823
rect 81 8800 519 8806
rect 631 8829 664 8831
rect 1036 8837 1077 8864
rect 1094 8837 1100 9263
rect 1036 8831 1100 8837
rect 1150 9263 1650 9269
rect 1150 8837 1156 9263
rect 1173 9215 1627 9263
rect 1173 8885 1235 9215
rect 1565 8885 1627 9215
rect 1173 8837 1627 8885
rect 1644 8837 1650 9263
rect 1150 8831 1650 8837
rect 1700 9263 1764 9269
rect 1700 8837 1706 9263
rect 1723 9236 1764 9263
rect 2136 9269 2169 9271
rect 2281 9294 2719 9300
rect 2281 9277 2287 9294
rect 2713 9277 2719 9294
rect 2281 9271 2719 9277
rect 2279 9269 2721 9271
rect 2831 9294 3269 9300
rect 2831 9277 2837 9294
rect 3263 9277 3269 9294
rect 2831 9271 3269 9277
rect 2831 9269 2864 9271
rect 2136 9263 2200 9269
rect 2136 9236 2177 9263
rect 1723 8864 1729 9236
rect 2171 8864 2177 9236
rect 1723 8837 1764 8864
rect 1700 8831 1764 8837
rect 1036 8829 1069 8831
rect 631 8823 1069 8829
rect 631 8806 637 8823
rect 1063 8806 1069 8823
rect 631 8800 1069 8806
rect 1179 8829 1621 8831
rect 1181 8823 1619 8829
rect 1181 8806 1187 8823
rect 1613 8806 1619 8823
rect 1181 8800 1619 8806
rect 1731 8829 1764 8831
rect 2136 8837 2177 8864
rect 2194 8837 2200 9263
rect 2136 8831 2200 8837
rect 2250 9263 2750 9269
rect 2250 8837 2256 9263
rect 2273 9215 2727 9263
rect 2273 8885 2335 9215
rect 2665 8885 2727 9215
rect 2273 8837 2727 8885
rect 2744 8837 2750 9263
rect 2250 8831 2750 8837
rect 2800 9263 2864 9269
rect 2800 8837 2806 9263
rect 2823 9236 2864 9263
rect 3236 9269 3269 9271
rect 3381 9294 3819 9300
rect 3381 9277 3387 9294
rect 3813 9277 3819 9294
rect 3381 9271 3819 9277
rect 3379 9269 3821 9271
rect 3931 9294 4369 9300
rect 3931 9277 3937 9294
rect 4363 9277 4369 9294
rect 3931 9271 4369 9277
rect 3931 9269 3964 9271
rect 3236 9263 3300 9269
rect 3236 9236 3277 9263
rect 2823 8864 2829 9236
rect 3271 8864 3277 9236
rect 2823 8837 2864 8864
rect 2800 8831 2864 8837
rect 2136 8829 2169 8831
rect 1731 8823 2169 8829
rect 1731 8806 1737 8823
rect 2163 8806 2169 8823
rect 1731 8800 2169 8806
rect 2279 8829 2721 8831
rect 2281 8823 2719 8829
rect 2281 8806 2287 8823
rect 2713 8806 2719 8823
rect 2281 8800 2719 8806
rect 2831 8829 2864 8831
rect 3236 8837 3277 8864
rect 3294 8837 3300 9263
rect 3236 8831 3300 8837
rect 3350 9263 3850 9269
rect 3350 8837 3356 9263
rect 3373 9215 3827 9263
rect 3373 8885 3435 9215
rect 3765 8885 3827 9215
rect 3373 8837 3827 8885
rect 3844 8837 3850 9263
rect 3350 8831 3850 8837
rect 3900 9263 3964 9269
rect 3900 8837 3906 9263
rect 3923 9236 3964 9263
rect 4336 9269 4369 9271
rect 4481 9294 4919 9300
rect 4481 9277 4487 9294
rect 4913 9277 4919 9294
rect 4481 9271 4919 9277
rect 4479 9269 4921 9271
rect 5031 9294 5469 9300
rect 5031 9277 5037 9294
rect 5463 9277 5469 9294
rect 5031 9271 5469 9277
rect 5031 9269 5064 9271
rect 4336 9263 4400 9269
rect 4336 9236 4377 9263
rect 3923 8864 3929 9236
rect 4371 8864 4377 9236
rect 3923 8837 3964 8864
rect 3900 8831 3964 8837
rect 3236 8829 3269 8831
rect 2831 8823 3269 8829
rect 2831 8806 2837 8823
rect 3263 8806 3269 8823
rect 2831 8800 3269 8806
rect 3379 8829 3821 8831
rect 3381 8823 3819 8829
rect 3381 8806 3387 8823
rect 3813 8806 3819 8823
rect 3381 8800 3819 8806
rect 3931 8829 3964 8831
rect 4336 8837 4377 8864
rect 4394 8837 4400 9263
rect 4336 8831 4400 8837
rect 4450 9263 4950 9269
rect 4450 8837 4456 9263
rect 4473 9215 4927 9263
rect 4473 8885 4535 9215
rect 4865 8885 4927 9215
rect 4473 8837 4927 8885
rect 4944 8837 4950 9263
rect 4450 8831 4950 8837
rect 5000 9263 5064 9269
rect 5000 8837 5006 9263
rect 5023 9236 5064 9263
rect 5436 9269 5469 9271
rect 5581 9294 6019 9300
rect 5581 9277 5587 9294
rect 6013 9277 6019 9294
rect 5581 9271 6019 9277
rect 5579 9269 6021 9271
rect 6131 9294 6569 9300
rect 6131 9277 6137 9294
rect 6563 9277 6569 9294
rect 6131 9271 6569 9277
rect 6131 9269 6164 9271
rect 5436 9263 5500 9269
rect 5436 9236 5477 9263
rect 5023 8864 5029 9236
rect 5471 8864 5477 9236
rect 5023 8837 5064 8864
rect 5000 8831 5064 8837
rect 4336 8829 4369 8831
rect 3931 8823 4369 8829
rect 3931 8806 3937 8823
rect 4363 8806 4369 8823
rect 3931 8800 4369 8806
rect 4479 8829 4921 8831
rect 4481 8823 4919 8829
rect 4481 8806 4487 8823
rect 4913 8806 4919 8823
rect 4481 8800 4919 8806
rect 5031 8829 5064 8831
rect 5436 8837 5477 8864
rect 5494 8837 5500 9263
rect 5436 8831 5500 8837
rect 5550 9263 6050 9269
rect 5550 8837 5556 9263
rect 5573 9215 6027 9263
rect 5573 8885 5635 9215
rect 5965 8885 6027 9215
rect 5573 8837 6027 8885
rect 6044 8837 6050 9263
rect 5550 8831 6050 8837
rect 6100 9263 6164 9269
rect 6100 8837 6106 9263
rect 6123 9236 6164 9263
rect 6536 9269 6569 9271
rect 6681 9294 7119 9300
rect 6681 9277 6687 9294
rect 7113 9277 7119 9294
rect 6681 9271 7119 9277
rect 6679 9269 7121 9271
rect 7231 9294 7669 9300
rect 7231 9277 7237 9294
rect 7663 9277 7669 9294
rect 7231 9271 7669 9277
rect 7231 9269 7264 9271
rect 6536 9263 6600 9269
rect 6536 9236 6577 9263
rect 6123 8864 6129 9236
rect 6571 8864 6577 9236
rect 6123 8837 6164 8864
rect 6100 8831 6164 8837
rect 5436 8829 5469 8831
rect 5031 8823 5469 8829
rect 5031 8806 5037 8823
rect 5463 8806 5469 8823
rect 5031 8800 5469 8806
rect 5579 8829 6021 8831
rect 5581 8823 6019 8829
rect 5581 8806 5587 8823
rect 6013 8806 6019 8823
rect 5581 8800 6019 8806
rect 6131 8829 6164 8831
rect 6536 8837 6577 8864
rect 6594 8837 6600 9263
rect 6536 8831 6600 8837
rect 6650 9263 7150 9269
rect 6650 8837 6656 9263
rect 6673 9215 7127 9263
rect 6673 8885 6735 9215
rect 7065 8885 7127 9215
rect 6673 8837 7127 8885
rect 7144 8837 7150 9263
rect 6650 8831 7150 8837
rect 7200 9263 7264 9269
rect 7200 8837 7206 9263
rect 7223 9236 7264 9263
rect 7636 9269 7669 9271
rect 7781 9294 8219 9300
rect 7781 9277 7787 9294
rect 8213 9277 8219 9294
rect 7781 9271 8219 9277
rect 7779 9269 8221 9271
rect 8331 9294 8769 9300
rect 8331 9277 8337 9294
rect 8763 9277 8769 9294
rect 8331 9271 8769 9277
rect 8331 9269 8364 9271
rect 7636 9263 7700 9269
rect 7636 9236 7677 9263
rect 7223 8864 7229 9236
rect 7671 8864 7677 9236
rect 7223 8837 7264 8864
rect 7200 8831 7264 8837
rect 6536 8829 6569 8831
rect 6131 8823 6569 8829
rect 6131 8806 6137 8823
rect 6563 8806 6569 8823
rect 6131 8800 6569 8806
rect 6679 8829 7121 8831
rect 6681 8823 7119 8829
rect 6681 8806 6687 8823
rect 7113 8806 7119 8823
rect 6681 8800 7119 8806
rect 7231 8829 7264 8831
rect 7636 8837 7677 8864
rect 7694 8837 7700 9263
rect 7636 8831 7700 8837
rect 7750 9263 8250 9269
rect 7750 8837 7756 9263
rect 7773 9215 8227 9263
rect 7773 8885 7835 9215
rect 8165 8885 8227 9215
rect 7773 8837 8227 8885
rect 8244 8837 8250 9263
rect 7750 8831 8250 8837
rect 8300 9263 8364 9269
rect 8300 8837 8306 9263
rect 8323 9236 8364 9263
rect 8736 9269 8769 9271
rect 8881 9294 9319 9300
rect 8881 9277 8887 9294
rect 9313 9277 9319 9294
rect 8881 9271 9319 9277
rect 8879 9269 9321 9271
rect 9431 9294 9869 9300
rect 9431 9277 9437 9294
rect 9863 9277 9869 9294
rect 9431 9271 9869 9277
rect 9431 9269 9464 9271
rect 8736 9263 8800 9269
rect 8736 9236 8777 9263
rect 8323 8864 8329 9236
rect 8771 8864 8777 9236
rect 8323 8837 8364 8864
rect 8300 8831 8364 8837
rect 7636 8829 7669 8831
rect 7231 8823 7669 8829
rect 7231 8806 7237 8823
rect 7663 8806 7669 8823
rect 7231 8800 7669 8806
rect 7779 8829 8221 8831
rect 7781 8823 8219 8829
rect 7781 8806 7787 8823
rect 8213 8806 8219 8823
rect 7781 8800 8219 8806
rect 8331 8829 8364 8831
rect 8736 8837 8777 8864
rect 8794 8837 8800 9263
rect 8736 8831 8800 8837
rect 8850 9263 9350 9269
rect 8850 8837 8856 9263
rect 8873 9215 9327 9263
rect 8873 8885 8935 9215
rect 9265 8885 9327 9215
rect 8873 8837 9327 8885
rect 9344 8837 9350 9263
rect 8850 8831 9350 8837
rect 9400 9263 9464 9269
rect 9400 8837 9406 9263
rect 9423 9236 9464 9263
rect 9836 9269 9869 9271
rect 9981 9294 10419 9300
rect 9981 9277 9987 9294
rect 10413 9277 10419 9294
rect 9981 9271 10419 9277
rect 9979 9269 10421 9271
rect 10531 9294 10969 9300
rect 10531 9277 10537 9294
rect 10963 9277 10969 9294
rect 10531 9271 10969 9277
rect 10531 9269 10564 9271
rect 9836 9263 9900 9269
rect 9836 9236 9877 9263
rect 9423 8864 9429 9236
rect 9871 8864 9877 9236
rect 9423 8837 9464 8864
rect 9400 8831 9464 8837
rect 8736 8829 8769 8831
rect 8331 8823 8769 8829
rect 8331 8806 8337 8823
rect 8763 8806 8769 8823
rect 8331 8800 8769 8806
rect 8879 8829 9321 8831
rect 8881 8823 9319 8829
rect 8881 8806 8887 8823
rect 9313 8806 9319 8823
rect 8881 8800 9319 8806
rect 9431 8829 9464 8831
rect 9836 8837 9877 8864
rect 9894 8837 9900 9263
rect 9836 8831 9900 8837
rect 9950 9263 10450 9269
rect 9950 8837 9956 9263
rect 9973 9215 10427 9263
rect 9973 8885 10035 9215
rect 10365 8885 10427 9215
rect 9973 8837 10427 8885
rect 10444 8837 10450 9263
rect 9950 8831 10450 8837
rect 10500 9263 10564 9269
rect 10500 8837 10506 9263
rect 10523 9236 10564 9263
rect 10936 9269 10969 9271
rect 11081 9294 11519 9300
rect 11081 9277 11087 9294
rect 11513 9277 11519 9294
rect 11081 9271 11519 9277
rect 11079 9269 11521 9271
rect 11631 9294 12069 9300
rect 11631 9277 11637 9294
rect 12063 9277 12069 9294
rect 11631 9271 12069 9277
rect 11631 9269 11664 9271
rect 10936 9263 11000 9269
rect 10936 9236 10977 9263
rect 10523 8864 10529 9236
rect 10971 8864 10977 9236
rect 10523 8837 10564 8864
rect 10500 8831 10564 8837
rect 9836 8829 9869 8831
rect 9431 8823 9869 8829
rect 9431 8806 9437 8823
rect 9863 8806 9869 8823
rect 9431 8800 9869 8806
rect 9979 8829 10421 8831
rect 9981 8823 10419 8829
rect 9981 8806 9987 8823
rect 10413 8806 10419 8823
rect 9981 8800 10419 8806
rect 10531 8829 10564 8831
rect 10936 8837 10977 8864
rect 10994 8837 11000 9263
rect 10936 8831 11000 8837
rect 11050 9263 11550 9269
rect 11050 8837 11056 9263
rect 11073 9215 11527 9263
rect 11073 8885 11135 9215
rect 11465 8885 11527 9215
rect 11073 8837 11527 8885
rect 11544 8837 11550 9263
rect 11050 8831 11550 8837
rect 11600 9263 11664 9269
rect 11600 8837 11606 9263
rect 11623 9236 11664 9263
rect 12036 9269 12069 9271
rect 12181 9294 12619 9300
rect 12181 9277 12187 9294
rect 12613 9277 12619 9294
rect 12181 9271 12619 9277
rect 12179 9269 12621 9271
rect 12731 9294 13169 9300
rect 12731 9277 12737 9294
rect 13163 9277 13169 9294
rect 12731 9271 13169 9277
rect 12731 9269 12764 9271
rect 12036 9263 12100 9269
rect 12036 9236 12077 9263
rect 11623 8864 11629 9236
rect 12071 8864 12077 9236
rect 11623 8837 11664 8864
rect 11600 8831 11664 8837
rect 10936 8829 10969 8831
rect 10531 8823 10969 8829
rect 10531 8806 10537 8823
rect 10963 8806 10969 8823
rect 10531 8800 10969 8806
rect 11079 8829 11521 8831
rect 11081 8823 11519 8829
rect 11081 8806 11087 8823
rect 11513 8806 11519 8823
rect 11081 8800 11519 8806
rect 11631 8829 11664 8831
rect 12036 8837 12077 8864
rect 12094 8837 12100 9263
rect 12036 8831 12100 8837
rect 12150 9263 12650 9269
rect 12150 8837 12156 9263
rect 12173 9215 12627 9263
rect 12173 8885 12235 9215
rect 12565 8885 12627 9215
rect 12173 8837 12627 8885
rect 12644 8837 12650 9263
rect 12150 8831 12650 8837
rect 12700 9263 12764 9269
rect 12700 8837 12706 9263
rect 12723 9236 12764 9263
rect 13136 9269 13169 9271
rect 13281 9294 13719 9300
rect 13281 9277 13287 9294
rect 13713 9277 13719 9294
rect 13281 9271 13719 9277
rect 13279 9269 13721 9271
rect 13136 9263 13200 9269
rect 13136 9236 13177 9263
rect 12723 8864 12729 9236
rect 13171 8864 13177 9236
rect 12723 8837 12764 8864
rect 12700 8831 12764 8837
rect 12036 8829 12069 8831
rect 11631 8823 12069 8829
rect 11631 8806 11637 8823
rect 12063 8806 12069 8823
rect 11631 8800 12069 8806
rect 12179 8829 12621 8831
rect 12181 8823 12619 8829
rect 12181 8806 12187 8823
rect 12613 8806 12619 8823
rect 12181 8800 12619 8806
rect 12731 8829 12764 8831
rect 13136 8837 13177 8864
rect 13194 8837 13200 9263
rect 13136 8831 13200 8837
rect 13250 9263 13721 9269
rect 13250 8837 13256 9263
rect 13273 9215 13721 9263
rect 13273 8885 13335 9215
rect 13665 8885 13721 9215
rect 13273 8837 13721 8885
rect 13250 8831 13721 8837
rect 13136 8829 13169 8831
rect 12731 8823 13169 8829
rect 12731 8806 12737 8823
rect 13163 8806 13169 8823
rect 12731 8800 13169 8806
rect 13279 8829 13721 8831
rect 13281 8823 13719 8829
rect 13281 8806 13287 8823
rect 13713 8806 13719 8823
rect 13281 8800 13719 8806
rect -469 8744 -31 8750
rect -469 8727 -463 8744
rect -37 8727 -31 8744
rect -469 8721 -31 8727
rect -471 8719 -29 8721
rect 81 8744 519 8750
rect 81 8727 87 8744
rect 513 8727 519 8744
rect 81 8721 519 8727
rect 81 8719 114 8721
rect -471 8713 0 8719
rect -471 8665 -23 8713
rect -471 8335 -415 8665
rect -85 8335 -23 8665
rect -471 8287 -23 8335
rect -6 8287 0 8713
rect -471 8281 0 8287
rect 50 8713 114 8719
rect 50 8287 56 8713
rect 73 8686 114 8713
rect 486 8719 519 8721
rect 631 8744 1069 8750
rect 631 8727 637 8744
rect 1063 8727 1069 8744
rect 631 8721 1069 8727
rect 629 8719 1071 8721
rect 1181 8744 1619 8750
rect 1181 8727 1187 8744
rect 1613 8727 1619 8744
rect 1181 8721 1619 8727
rect 1181 8719 1214 8721
rect 486 8713 550 8719
rect 486 8686 527 8713
rect 73 8314 79 8686
rect 521 8314 527 8686
rect 73 8287 114 8314
rect 50 8281 114 8287
rect -471 8279 -29 8281
rect -469 8273 -31 8279
rect -469 8256 -463 8273
rect -37 8256 -31 8273
rect -469 8250 -31 8256
rect 81 8279 114 8281
rect 486 8287 527 8314
rect 544 8287 550 8713
rect 486 8281 550 8287
rect 600 8713 1100 8719
rect 600 8287 606 8713
rect 623 8665 1077 8713
rect 623 8335 685 8665
rect 1015 8335 1077 8665
rect 623 8287 1077 8335
rect 1094 8287 1100 8713
rect 600 8281 1100 8287
rect 1150 8713 1214 8719
rect 1150 8287 1156 8713
rect 1173 8686 1214 8713
rect 1586 8719 1619 8721
rect 1731 8744 2169 8750
rect 1731 8727 1737 8744
rect 2163 8727 2169 8744
rect 1731 8721 2169 8727
rect 1729 8719 2171 8721
rect 2281 8744 2719 8750
rect 2281 8727 2287 8744
rect 2713 8727 2719 8744
rect 2281 8721 2719 8727
rect 2281 8719 2314 8721
rect 1586 8713 1650 8719
rect 1586 8686 1627 8713
rect 1173 8314 1179 8686
rect 1621 8314 1627 8686
rect 1173 8287 1214 8314
rect 1150 8281 1214 8287
rect 486 8279 519 8281
rect 81 8273 519 8279
rect 81 8256 87 8273
rect 513 8256 519 8273
rect 81 8250 519 8256
rect 629 8279 1071 8281
rect 631 8273 1069 8279
rect 631 8256 637 8273
rect 1063 8256 1069 8273
rect 631 8250 1069 8256
rect 1181 8279 1214 8281
rect 1586 8287 1627 8314
rect 1644 8287 1650 8713
rect 1586 8281 1650 8287
rect 1700 8713 2200 8719
rect 1700 8287 1706 8713
rect 1723 8665 2177 8713
rect 1723 8335 1785 8665
rect 2115 8335 2177 8665
rect 1723 8287 2177 8335
rect 2194 8287 2200 8713
rect 1700 8281 2200 8287
rect 2250 8713 2314 8719
rect 2250 8287 2256 8713
rect 2273 8686 2314 8713
rect 2686 8719 2719 8721
rect 2831 8744 3269 8750
rect 2831 8727 2837 8744
rect 3263 8727 3269 8744
rect 2831 8721 3269 8727
rect 2829 8719 3271 8721
rect 3381 8744 3819 8750
rect 3381 8727 3387 8744
rect 3813 8727 3819 8744
rect 3381 8721 3819 8727
rect 3381 8719 3414 8721
rect 2686 8713 2750 8719
rect 2686 8686 2727 8713
rect 2273 8314 2279 8686
rect 2721 8314 2727 8686
rect 2273 8287 2314 8314
rect 2250 8281 2314 8287
rect 1586 8279 1619 8281
rect 1181 8273 1619 8279
rect 1181 8256 1187 8273
rect 1613 8256 1619 8273
rect 1181 8250 1619 8256
rect 1729 8279 2171 8281
rect 1731 8273 2169 8279
rect 1731 8256 1737 8273
rect 2163 8256 2169 8273
rect 1731 8250 2169 8256
rect 2281 8279 2314 8281
rect 2686 8287 2727 8314
rect 2744 8287 2750 8713
rect 2686 8281 2750 8287
rect 2800 8713 3300 8719
rect 2800 8287 2806 8713
rect 2823 8665 3277 8713
rect 2823 8335 2885 8665
rect 3215 8335 3277 8665
rect 2823 8287 3277 8335
rect 3294 8287 3300 8713
rect 2800 8281 3300 8287
rect 3350 8713 3414 8719
rect 3350 8287 3356 8713
rect 3373 8686 3414 8713
rect 3786 8719 3819 8721
rect 3931 8744 4369 8750
rect 3931 8727 3937 8744
rect 4363 8727 4369 8744
rect 3931 8721 4369 8727
rect 3929 8719 4371 8721
rect 4481 8744 4919 8750
rect 4481 8727 4487 8744
rect 4913 8727 4919 8744
rect 4481 8721 4919 8727
rect 4481 8719 4514 8721
rect 3786 8713 3850 8719
rect 3786 8686 3827 8713
rect 3373 8314 3379 8686
rect 3821 8314 3827 8686
rect 3373 8287 3414 8314
rect 3350 8281 3414 8287
rect 2686 8279 2719 8281
rect 2281 8273 2719 8279
rect 2281 8256 2287 8273
rect 2713 8256 2719 8273
rect 2281 8250 2719 8256
rect 2829 8279 3271 8281
rect 2831 8273 3269 8279
rect 2831 8256 2837 8273
rect 3263 8256 3269 8273
rect 2831 8250 3269 8256
rect 3381 8279 3414 8281
rect 3786 8287 3827 8314
rect 3844 8287 3850 8713
rect 3786 8281 3850 8287
rect 3900 8713 4400 8719
rect 3900 8287 3906 8713
rect 3923 8665 4377 8713
rect 3923 8335 3985 8665
rect 4315 8335 4377 8665
rect 3923 8287 4377 8335
rect 4394 8287 4400 8713
rect 3900 8281 4400 8287
rect 4450 8713 4514 8719
rect 4450 8287 4456 8713
rect 4473 8686 4514 8713
rect 4886 8719 4919 8721
rect 5031 8744 5469 8750
rect 5031 8727 5037 8744
rect 5463 8727 5469 8744
rect 5031 8721 5469 8727
rect 5029 8719 5471 8721
rect 5581 8744 6019 8750
rect 5581 8727 5587 8744
rect 6013 8727 6019 8744
rect 5581 8721 6019 8727
rect 5581 8719 5614 8721
rect 4886 8713 4950 8719
rect 4886 8686 4927 8713
rect 4473 8314 4479 8686
rect 4921 8314 4927 8686
rect 4473 8287 4514 8314
rect 4450 8281 4514 8287
rect 3786 8279 3819 8281
rect 3381 8273 3819 8279
rect 3381 8256 3387 8273
rect 3813 8256 3819 8273
rect 3381 8250 3819 8256
rect 3929 8279 4371 8281
rect 3931 8273 4369 8279
rect 3931 8256 3937 8273
rect 4363 8256 4369 8273
rect 3931 8250 4369 8256
rect 4481 8279 4514 8281
rect 4886 8287 4927 8314
rect 4944 8287 4950 8713
rect 4886 8281 4950 8287
rect 5000 8713 5500 8719
rect 5000 8287 5006 8713
rect 5023 8665 5477 8713
rect 5023 8335 5085 8665
rect 5415 8335 5477 8665
rect 5023 8287 5477 8335
rect 5494 8287 5500 8713
rect 5000 8281 5500 8287
rect 5550 8713 5614 8719
rect 5550 8287 5556 8713
rect 5573 8686 5614 8713
rect 5986 8719 6019 8721
rect 6131 8744 6569 8750
rect 6131 8727 6137 8744
rect 6563 8727 6569 8744
rect 6131 8721 6569 8727
rect 6129 8719 6571 8721
rect 6681 8744 7119 8750
rect 6681 8727 6687 8744
rect 7113 8727 7119 8744
rect 6681 8721 7119 8727
rect 6681 8719 6714 8721
rect 5986 8713 6050 8719
rect 5986 8686 6027 8713
rect 5573 8314 5579 8686
rect 6021 8314 6027 8686
rect 5573 8287 5614 8314
rect 5550 8281 5614 8287
rect 4886 8279 4919 8281
rect 4481 8273 4919 8279
rect 4481 8256 4487 8273
rect 4913 8256 4919 8273
rect 4481 8250 4919 8256
rect 5029 8279 5471 8281
rect 5031 8273 5469 8279
rect 5031 8256 5037 8273
rect 5463 8256 5469 8273
rect 5031 8250 5469 8256
rect 5581 8279 5614 8281
rect 5986 8287 6027 8314
rect 6044 8287 6050 8713
rect 5986 8281 6050 8287
rect 6100 8713 6600 8719
rect 6100 8287 6106 8713
rect 6123 8665 6577 8713
rect 6123 8335 6185 8665
rect 6515 8335 6577 8665
rect 6123 8287 6577 8335
rect 6594 8287 6600 8713
rect 6100 8281 6600 8287
rect 6650 8713 6714 8719
rect 6650 8287 6656 8713
rect 6673 8686 6714 8713
rect 7086 8719 7119 8721
rect 7231 8744 7669 8750
rect 7231 8727 7237 8744
rect 7663 8727 7669 8744
rect 7231 8721 7669 8727
rect 7229 8719 7671 8721
rect 7781 8744 8219 8750
rect 7781 8727 7787 8744
rect 8213 8727 8219 8744
rect 7781 8721 8219 8727
rect 7781 8719 7814 8721
rect 7086 8713 7150 8719
rect 7086 8686 7127 8713
rect 6673 8314 6679 8686
rect 7121 8314 7127 8686
rect 6673 8287 6714 8314
rect 6650 8281 6714 8287
rect 5986 8279 6019 8281
rect 5581 8273 6019 8279
rect 5581 8256 5587 8273
rect 6013 8256 6019 8273
rect 5581 8250 6019 8256
rect 6129 8279 6571 8281
rect 6131 8273 6569 8279
rect 6131 8256 6137 8273
rect 6563 8256 6569 8273
rect 6131 8250 6569 8256
rect 6681 8279 6714 8281
rect 7086 8287 7127 8314
rect 7144 8287 7150 8713
rect 7086 8281 7150 8287
rect 7200 8713 7700 8719
rect 7200 8287 7206 8713
rect 7223 8665 7677 8713
rect 7223 8335 7285 8665
rect 7615 8335 7677 8665
rect 7223 8287 7677 8335
rect 7694 8287 7700 8713
rect 7200 8281 7700 8287
rect 7750 8713 7814 8719
rect 7750 8287 7756 8713
rect 7773 8686 7814 8713
rect 8186 8719 8219 8721
rect 8331 8744 8769 8750
rect 8331 8727 8337 8744
rect 8763 8727 8769 8744
rect 8331 8721 8769 8727
rect 8329 8719 8771 8721
rect 8881 8744 9319 8750
rect 8881 8727 8887 8744
rect 9313 8727 9319 8744
rect 8881 8721 9319 8727
rect 8881 8719 8914 8721
rect 8186 8713 8250 8719
rect 8186 8686 8227 8713
rect 7773 8314 7779 8686
rect 8221 8314 8227 8686
rect 7773 8287 7814 8314
rect 7750 8281 7814 8287
rect 7086 8279 7119 8281
rect 6681 8273 7119 8279
rect 6681 8256 6687 8273
rect 7113 8256 7119 8273
rect 6681 8250 7119 8256
rect 7229 8279 7671 8281
rect 7231 8273 7669 8279
rect 7231 8256 7237 8273
rect 7663 8256 7669 8273
rect 7231 8250 7669 8256
rect 7781 8279 7814 8281
rect 8186 8287 8227 8314
rect 8244 8287 8250 8713
rect 8186 8281 8250 8287
rect 8300 8713 8800 8719
rect 8300 8287 8306 8713
rect 8323 8665 8777 8713
rect 8323 8335 8385 8665
rect 8715 8335 8777 8665
rect 8323 8287 8777 8335
rect 8794 8287 8800 8713
rect 8300 8281 8800 8287
rect 8850 8713 8914 8719
rect 8850 8287 8856 8713
rect 8873 8686 8914 8713
rect 9286 8719 9319 8721
rect 9431 8744 9869 8750
rect 9431 8727 9437 8744
rect 9863 8727 9869 8744
rect 9431 8721 9869 8727
rect 9429 8719 9871 8721
rect 9981 8744 10419 8750
rect 9981 8727 9987 8744
rect 10413 8727 10419 8744
rect 9981 8721 10419 8727
rect 9981 8719 10014 8721
rect 9286 8713 9350 8719
rect 9286 8686 9327 8713
rect 8873 8314 8879 8686
rect 9321 8314 9327 8686
rect 8873 8287 8914 8314
rect 8850 8281 8914 8287
rect 8186 8279 8219 8281
rect 7781 8273 8219 8279
rect 7781 8256 7787 8273
rect 8213 8256 8219 8273
rect 7781 8250 8219 8256
rect 8329 8279 8771 8281
rect 8331 8273 8769 8279
rect 8331 8256 8337 8273
rect 8763 8256 8769 8273
rect 8331 8250 8769 8256
rect 8881 8279 8914 8281
rect 9286 8287 9327 8314
rect 9344 8287 9350 8713
rect 9286 8281 9350 8287
rect 9400 8713 9900 8719
rect 9400 8287 9406 8713
rect 9423 8665 9877 8713
rect 9423 8335 9485 8665
rect 9815 8335 9877 8665
rect 9423 8287 9877 8335
rect 9894 8287 9900 8713
rect 9400 8281 9900 8287
rect 9950 8713 10014 8719
rect 9950 8287 9956 8713
rect 9973 8686 10014 8713
rect 10386 8719 10419 8721
rect 10531 8744 10969 8750
rect 10531 8727 10537 8744
rect 10963 8727 10969 8744
rect 10531 8721 10969 8727
rect 10529 8719 10971 8721
rect 11081 8744 11519 8750
rect 11081 8727 11087 8744
rect 11513 8727 11519 8744
rect 11081 8721 11519 8727
rect 11081 8719 11114 8721
rect 10386 8713 10450 8719
rect 10386 8686 10427 8713
rect 9973 8314 9979 8686
rect 10421 8314 10427 8686
rect 9973 8287 10014 8314
rect 9950 8281 10014 8287
rect 9286 8279 9319 8281
rect 8881 8273 9319 8279
rect 8881 8256 8887 8273
rect 9313 8256 9319 8273
rect 8881 8250 9319 8256
rect 9429 8279 9871 8281
rect 9431 8273 9869 8279
rect 9431 8256 9437 8273
rect 9863 8256 9869 8273
rect 9431 8250 9869 8256
rect 9981 8279 10014 8281
rect 10386 8287 10427 8314
rect 10444 8287 10450 8713
rect 10386 8281 10450 8287
rect 10500 8713 11000 8719
rect 10500 8287 10506 8713
rect 10523 8665 10977 8713
rect 10523 8335 10585 8665
rect 10915 8335 10977 8665
rect 10523 8287 10977 8335
rect 10994 8287 11000 8713
rect 10500 8281 11000 8287
rect 11050 8713 11114 8719
rect 11050 8287 11056 8713
rect 11073 8686 11114 8713
rect 11486 8719 11519 8721
rect 11631 8744 12069 8750
rect 11631 8727 11637 8744
rect 12063 8727 12069 8744
rect 11631 8721 12069 8727
rect 11629 8719 12071 8721
rect 12181 8744 12619 8750
rect 12181 8727 12187 8744
rect 12613 8727 12619 8744
rect 12181 8721 12619 8727
rect 12181 8719 12214 8721
rect 11486 8713 11550 8719
rect 11486 8686 11527 8713
rect 11073 8314 11079 8686
rect 11521 8314 11527 8686
rect 11073 8287 11114 8314
rect 11050 8281 11114 8287
rect 10386 8279 10419 8281
rect 9981 8273 10419 8279
rect 9981 8256 9987 8273
rect 10413 8256 10419 8273
rect 9981 8250 10419 8256
rect 10529 8279 10971 8281
rect 10531 8273 10969 8279
rect 10531 8256 10537 8273
rect 10963 8256 10969 8273
rect 10531 8250 10969 8256
rect 11081 8279 11114 8281
rect 11486 8287 11527 8314
rect 11544 8287 11550 8713
rect 11486 8281 11550 8287
rect 11600 8713 12100 8719
rect 11600 8287 11606 8713
rect 11623 8665 12077 8713
rect 11623 8335 11685 8665
rect 12015 8335 12077 8665
rect 11623 8287 12077 8335
rect 12094 8287 12100 8713
rect 11600 8281 12100 8287
rect 12150 8713 12214 8719
rect 12150 8287 12156 8713
rect 12173 8686 12214 8713
rect 12586 8719 12619 8721
rect 12731 8744 13169 8750
rect 12731 8727 12737 8744
rect 13163 8727 13169 8744
rect 12731 8721 13169 8727
rect 12729 8719 13171 8721
rect 13281 8744 13719 8750
rect 13281 8727 13287 8744
rect 13713 8727 13719 8744
rect 13281 8721 13719 8727
rect 13281 8719 13314 8721
rect 12586 8713 12650 8719
rect 12586 8686 12627 8713
rect 12173 8314 12179 8686
rect 12621 8314 12627 8686
rect 12173 8287 12214 8314
rect 12150 8281 12214 8287
rect 11486 8279 11519 8281
rect 11081 8273 11519 8279
rect 11081 8256 11087 8273
rect 11513 8256 11519 8273
rect 11081 8250 11519 8256
rect 11629 8279 12071 8281
rect 11631 8273 12069 8279
rect 11631 8256 11637 8273
rect 12063 8256 12069 8273
rect 11631 8250 12069 8256
rect 12181 8279 12214 8281
rect 12586 8287 12627 8314
rect 12644 8287 12650 8713
rect 12586 8281 12650 8287
rect 12700 8713 13200 8719
rect 12700 8287 12706 8713
rect 12723 8665 13177 8713
rect 12723 8335 12785 8665
rect 13115 8335 13177 8665
rect 12723 8287 13177 8335
rect 13194 8287 13200 8713
rect 12700 8281 13200 8287
rect 13250 8713 13314 8719
rect 13250 8287 13256 8713
rect 13273 8686 13314 8713
rect 13273 8314 13279 8686
rect 13273 8287 13314 8314
rect 13250 8281 13314 8287
rect 12586 8279 12619 8281
rect 12181 8273 12619 8279
rect 12181 8256 12187 8273
rect 12613 8256 12619 8273
rect 12181 8250 12619 8256
rect 12729 8279 13171 8281
rect 12731 8273 13169 8279
rect 12731 8256 12737 8273
rect 13163 8256 13169 8273
rect 12731 8250 13169 8256
rect 13281 8279 13314 8281
rect 13281 8273 13719 8279
rect 13281 8256 13287 8273
rect 13713 8256 13719 8273
rect 13281 8250 13719 8256
rect -469 8194 -31 8200
rect -469 8177 -463 8194
rect -37 8177 -31 8194
rect -469 8171 -31 8177
rect -64 8169 -31 8171
rect 81 8194 519 8200
rect 81 8177 87 8194
rect 513 8177 519 8194
rect 81 8171 519 8177
rect 79 8169 521 8171
rect 631 8194 1069 8200
rect 631 8177 637 8194
rect 1063 8177 1069 8194
rect 631 8171 1069 8177
rect 631 8169 664 8171
rect -64 8163 0 8169
rect -64 8136 -23 8163
rect -29 7764 -23 8136
rect -64 7737 -23 7764
rect -6 7737 0 8163
rect -64 7731 0 7737
rect 50 8163 550 8169
rect 50 7737 56 8163
rect 73 8115 527 8163
rect 73 7785 135 8115
rect 465 7785 527 8115
rect 73 7737 527 7785
rect 544 7737 550 8163
rect 50 7731 550 7737
rect 600 8163 664 8169
rect 600 7737 606 8163
rect 623 8136 664 8163
rect 1036 8169 1069 8171
rect 1181 8194 1619 8200
rect 1181 8177 1187 8194
rect 1613 8177 1619 8194
rect 1181 8171 1619 8177
rect 1179 8169 1621 8171
rect 1731 8194 2169 8200
rect 1731 8177 1737 8194
rect 2163 8177 2169 8194
rect 1731 8171 2169 8177
rect 1731 8169 1764 8171
rect 1036 8163 1100 8169
rect 1036 8136 1077 8163
rect 623 7764 629 8136
rect 1071 7764 1077 8136
rect 623 7737 664 7764
rect 600 7731 664 7737
rect -64 7729 -31 7731
rect -469 7723 -31 7729
rect -469 7706 -463 7723
rect -37 7706 -31 7723
rect -469 7700 -31 7706
rect 79 7729 521 7731
rect 81 7723 519 7729
rect 81 7706 87 7723
rect 513 7706 519 7723
rect 81 7700 519 7706
rect 631 7729 664 7731
rect 1036 7737 1077 7764
rect 1094 7737 1100 8163
rect 1036 7731 1100 7737
rect 1150 8163 1650 8169
rect 1150 7737 1156 8163
rect 1173 8115 1627 8163
rect 1173 7785 1235 8115
rect 1565 7785 1627 8115
rect 1173 7737 1627 7785
rect 1644 7737 1650 8163
rect 1150 7731 1650 7737
rect 1700 8163 1764 8169
rect 1700 7737 1706 8163
rect 1723 8136 1764 8163
rect 2136 8169 2169 8171
rect 2281 8194 2719 8200
rect 2281 8177 2287 8194
rect 2713 8177 2719 8194
rect 2281 8171 2719 8177
rect 2279 8169 2721 8171
rect 2831 8194 3269 8200
rect 2831 8177 2837 8194
rect 3263 8177 3269 8194
rect 2831 8171 3269 8177
rect 2831 8169 2864 8171
rect 2136 8163 2200 8169
rect 2136 8136 2177 8163
rect 1723 7764 1729 8136
rect 2171 7764 2177 8136
rect 1723 7737 1764 7764
rect 1700 7731 1764 7737
rect 1036 7729 1069 7731
rect 631 7723 1069 7729
rect 631 7706 637 7723
rect 1063 7706 1069 7723
rect 631 7700 1069 7706
rect 1179 7729 1621 7731
rect 1181 7723 1619 7729
rect 1181 7706 1187 7723
rect 1613 7706 1619 7723
rect 1181 7700 1619 7706
rect 1731 7729 1764 7731
rect 2136 7737 2177 7764
rect 2194 7737 2200 8163
rect 2136 7731 2200 7737
rect 2250 8163 2750 8169
rect 2250 7737 2256 8163
rect 2273 8115 2727 8163
rect 2273 7785 2335 8115
rect 2665 7785 2727 8115
rect 2273 7737 2727 7785
rect 2744 7737 2750 8163
rect 2250 7731 2750 7737
rect 2800 8163 2864 8169
rect 2800 7737 2806 8163
rect 2823 8136 2864 8163
rect 3236 8169 3269 8171
rect 3381 8194 3819 8200
rect 3381 8177 3387 8194
rect 3813 8177 3819 8194
rect 3381 8171 3819 8177
rect 3379 8169 3821 8171
rect 3931 8194 4369 8200
rect 3931 8177 3937 8194
rect 4363 8177 4369 8194
rect 3931 8171 4369 8177
rect 3931 8169 3964 8171
rect 3236 8163 3300 8169
rect 3236 8136 3277 8163
rect 2823 7764 2829 8136
rect 3271 7764 3277 8136
rect 2823 7737 2864 7764
rect 2800 7731 2864 7737
rect 2136 7729 2169 7731
rect 1731 7723 2169 7729
rect 1731 7706 1737 7723
rect 2163 7706 2169 7723
rect 1731 7700 2169 7706
rect 2279 7729 2721 7731
rect 2281 7723 2719 7729
rect 2281 7706 2287 7723
rect 2713 7706 2719 7723
rect 2281 7700 2719 7706
rect 2831 7729 2864 7731
rect 3236 7737 3277 7764
rect 3294 7737 3300 8163
rect 3236 7731 3300 7737
rect 3350 8163 3850 8169
rect 3350 7737 3356 8163
rect 3373 8115 3827 8163
rect 3373 7785 3435 8115
rect 3765 7785 3827 8115
rect 3373 7737 3827 7785
rect 3844 7737 3850 8163
rect 3350 7731 3850 7737
rect 3900 8163 3964 8169
rect 3900 7737 3906 8163
rect 3923 8136 3964 8163
rect 4336 8169 4369 8171
rect 4481 8194 4919 8200
rect 4481 8177 4487 8194
rect 4913 8177 4919 8194
rect 4481 8171 4919 8177
rect 4479 8169 4921 8171
rect 5031 8194 5469 8200
rect 5031 8177 5037 8194
rect 5463 8177 5469 8194
rect 5031 8171 5469 8177
rect 5031 8169 5064 8171
rect 4336 8163 4400 8169
rect 4336 8136 4377 8163
rect 3923 7764 3929 8136
rect 4371 7764 4377 8136
rect 3923 7737 3964 7764
rect 3900 7731 3964 7737
rect 3236 7729 3269 7731
rect 2831 7723 3269 7729
rect 2831 7706 2837 7723
rect 3263 7706 3269 7723
rect 2831 7700 3269 7706
rect 3379 7729 3821 7731
rect 3381 7723 3819 7729
rect 3381 7706 3387 7723
rect 3813 7706 3819 7723
rect 3381 7700 3819 7706
rect 3931 7729 3964 7731
rect 4336 7737 4377 7764
rect 4394 7737 4400 8163
rect 4336 7731 4400 7737
rect 4450 8163 4950 8169
rect 4450 7737 4456 8163
rect 4473 8115 4927 8163
rect 4473 7785 4535 8115
rect 4865 7785 4927 8115
rect 4473 7737 4927 7785
rect 4944 7737 4950 8163
rect 4450 7731 4950 7737
rect 5000 8163 5064 8169
rect 5000 7737 5006 8163
rect 5023 8136 5064 8163
rect 5436 8169 5469 8171
rect 5581 8194 6019 8200
rect 5581 8177 5587 8194
rect 6013 8177 6019 8194
rect 5581 8171 6019 8177
rect 5579 8169 6021 8171
rect 6131 8194 6569 8200
rect 6131 8177 6137 8194
rect 6563 8177 6569 8194
rect 6131 8171 6569 8177
rect 6131 8169 6164 8171
rect 5436 8163 5500 8169
rect 5436 8136 5477 8163
rect 5023 7764 5029 8136
rect 5471 7764 5477 8136
rect 5023 7737 5064 7764
rect 5000 7731 5064 7737
rect 4336 7729 4369 7731
rect 3931 7723 4369 7729
rect 3931 7706 3937 7723
rect 4363 7706 4369 7723
rect 3931 7700 4369 7706
rect 4479 7729 4921 7731
rect 4481 7723 4919 7729
rect 4481 7706 4487 7723
rect 4913 7706 4919 7723
rect 4481 7700 4919 7706
rect 5031 7729 5064 7731
rect 5436 7737 5477 7764
rect 5494 7737 5500 8163
rect 5436 7731 5500 7737
rect 5550 8163 6050 8169
rect 5550 7737 5556 8163
rect 5573 8115 6027 8163
rect 5573 7785 5635 8115
rect 5965 7785 6027 8115
rect 5573 7737 6027 7785
rect 6044 7737 6050 8163
rect 5550 7731 6050 7737
rect 6100 8163 6164 8169
rect 6100 7737 6106 8163
rect 6123 8136 6164 8163
rect 6536 8169 6569 8171
rect 6681 8194 7119 8200
rect 6681 8177 6687 8194
rect 7113 8177 7119 8194
rect 6681 8171 7119 8177
rect 6679 8169 7121 8171
rect 7231 8194 7669 8200
rect 7231 8177 7237 8194
rect 7663 8177 7669 8194
rect 7231 8171 7669 8177
rect 7231 8169 7264 8171
rect 6536 8163 6600 8169
rect 6536 8136 6577 8163
rect 6123 7764 6129 8136
rect 6571 7764 6577 8136
rect 6123 7737 6164 7764
rect 6100 7731 6164 7737
rect 5436 7729 5469 7731
rect 5031 7723 5469 7729
rect 5031 7706 5037 7723
rect 5463 7706 5469 7723
rect 5031 7700 5469 7706
rect 5579 7729 6021 7731
rect 5581 7723 6019 7729
rect 5581 7706 5587 7723
rect 6013 7706 6019 7723
rect 5581 7700 6019 7706
rect 6131 7729 6164 7731
rect 6536 7737 6577 7764
rect 6594 7737 6600 8163
rect 6536 7731 6600 7737
rect 6650 8163 7150 8169
rect 6650 7737 6656 8163
rect 6673 8115 7127 8163
rect 6673 7785 6735 8115
rect 7065 7785 7127 8115
rect 6673 7737 7127 7785
rect 7144 7737 7150 8163
rect 6650 7731 7150 7737
rect 7200 8163 7264 8169
rect 7200 7737 7206 8163
rect 7223 8136 7264 8163
rect 7636 8169 7669 8171
rect 7781 8194 8219 8200
rect 7781 8177 7787 8194
rect 8213 8177 8219 8194
rect 7781 8171 8219 8177
rect 7779 8169 8221 8171
rect 8331 8194 8769 8200
rect 8331 8177 8337 8194
rect 8763 8177 8769 8194
rect 8331 8171 8769 8177
rect 8331 8169 8364 8171
rect 7636 8163 7700 8169
rect 7636 8136 7677 8163
rect 7223 7764 7229 8136
rect 7671 7764 7677 8136
rect 7223 7737 7264 7764
rect 7200 7731 7264 7737
rect 6536 7729 6569 7731
rect 6131 7723 6569 7729
rect 6131 7706 6137 7723
rect 6563 7706 6569 7723
rect 6131 7700 6569 7706
rect 6679 7729 7121 7731
rect 6681 7723 7119 7729
rect 6681 7706 6687 7723
rect 7113 7706 7119 7723
rect 6681 7700 7119 7706
rect 7231 7729 7264 7731
rect 7636 7737 7677 7764
rect 7694 7737 7700 8163
rect 7636 7731 7700 7737
rect 7750 8163 8250 8169
rect 7750 7737 7756 8163
rect 7773 8115 8227 8163
rect 7773 7785 7835 8115
rect 8165 7785 8227 8115
rect 7773 7737 8227 7785
rect 8244 7737 8250 8163
rect 7750 7731 8250 7737
rect 8300 8163 8364 8169
rect 8300 7737 8306 8163
rect 8323 8136 8364 8163
rect 8736 8169 8769 8171
rect 8881 8194 9319 8200
rect 8881 8177 8887 8194
rect 9313 8177 9319 8194
rect 8881 8171 9319 8177
rect 8879 8169 9321 8171
rect 9431 8194 9869 8200
rect 9431 8177 9437 8194
rect 9863 8177 9869 8194
rect 9431 8171 9869 8177
rect 9431 8169 9464 8171
rect 8736 8163 8800 8169
rect 8736 8136 8777 8163
rect 8323 7764 8329 8136
rect 8771 7764 8777 8136
rect 8323 7737 8364 7764
rect 8300 7731 8364 7737
rect 7636 7729 7669 7731
rect 7231 7723 7669 7729
rect 7231 7706 7237 7723
rect 7663 7706 7669 7723
rect 7231 7700 7669 7706
rect 7779 7729 8221 7731
rect 7781 7723 8219 7729
rect 7781 7706 7787 7723
rect 8213 7706 8219 7723
rect 7781 7700 8219 7706
rect 8331 7729 8364 7731
rect 8736 7737 8777 7764
rect 8794 7737 8800 8163
rect 8736 7731 8800 7737
rect 8850 8163 9350 8169
rect 8850 7737 8856 8163
rect 8873 8115 9327 8163
rect 8873 7785 8935 8115
rect 9265 7785 9327 8115
rect 8873 7737 9327 7785
rect 9344 7737 9350 8163
rect 8850 7731 9350 7737
rect 9400 8163 9464 8169
rect 9400 7737 9406 8163
rect 9423 8136 9464 8163
rect 9836 8169 9869 8171
rect 9981 8194 10419 8200
rect 9981 8177 9987 8194
rect 10413 8177 10419 8194
rect 9981 8171 10419 8177
rect 9979 8169 10421 8171
rect 10531 8194 10969 8200
rect 10531 8177 10537 8194
rect 10963 8177 10969 8194
rect 10531 8171 10969 8177
rect 10531 8169 10564 8171
rect 9836 8163 9900 8169
rect 9836 8136 9877 8163
rect 9423 7764 9429 8136
rect 9871 7764 9877 8136
rect 9423 7737 9464 7764
rect 9400 7731 9464 7737
rect 8736 7729 8769 7731
rect 8331 7723 8769 7729
rect 8331 7706 8337 7723
rect 8763 7706 8769 7723
rect 8331 7700 8769 7706
rect 8879 7729 9321 7731
rect 8881 7723 9319 7729
rect 8881 7706 8887 7723
rect 9313 7706 9319 7723
rect 8881 7700 9319 7706
rect 9431 7729 9464 7731
rect 9836 7737 9877 7764
rect 9894 7737 9900 8163
rect 9836 7731 9900 7737
rect 9950 8163 10450 8169
rect 9950 7737 9956 8163
rect 9973 8115 10427 8163
rect 9973 7785 10035 8115
rect 10365 7785 10427 8115
rect 9973 7737 10427 7785
rect 10444 7737 10450 8163
rect 9950 7731 10450 7737
rect 10500 8163 10564 8169
rect 10500 7737 10506 8163
rect 10523 8136 10564 8163
rect 10936 8169 10969 8171
rect 11081 8194 11519 8200
rect 11081 8177 11087 8194
rect 11513 8177 11519 8194
rect 11081 8171 11519 8177
rect 11079 8169 11521 8171
rect 11631 8194 12069 8200
rect 11631 8177 11637 8194
rect 12063 8177 12069 8194
rect 11631 8171 12069 8177
rect 11631 8169 11664 8171
rect 10936 8163 11000 8169
rect 10936 8136 10977 8163
rect 10523 7764 10529 8136
rect 10971 7764 10977 8136
rect 10523 7737 10564 7764
rect 10500 7731 10564 7737
rect 9836 7729 9869 7731
rect 9431 7723 9869 7729
rect 9431 7706 9437 7723
rect 9863 7706 9869 7723
rect 9431 7700 9869 7706
rect 9979 7729 10421 7731
rect 9981 7723 10419 7729
rect 9981 7706 9987 7723
rect 10413 7706 10419 7723
rect 9981 7700 10419 7706
rect 10531 7729 10564 7731
rect 10936 7737 10977 7764
rect 10994 7737 11000 8163
rect 10936 7731 11000 7737
rect 11050 8163 11550 8169
rect 11050 7737 11056 8163
rect 11073 8115 11527 8163
rect 11073 7785 11135 8115
rect 11465 7785 11527 8115
rect 11073 7737 11527 7785
rect 11544 7737 11550 8163
rect 11050 7731 11550 7737
rect 11600 8163 11664 8169
rect 11600 7737 11606 8163
rect 11623 8136 11664 8163
rect 12036 8169 12069 8171
rect 12181 8194 12619 8200
rect 12181 8177 12187 8194
rect 12613 8177 12619 8194
rect 12181 8171 12619 8177
rect 12179 8169 12621 8171
rect 12731 8194 13169 8200
rect 12731 8177 12737 8194
rect 13163 8177 13169 8194
rect 12731 8171 13169 8177
rect 12731 8169 12764 8171
rect 12036 8163 12100 8169
rect 12036 8136 12077 8163
rect 11623 7764 11629 8136
rect 12071 7764 12077 8136
rect 11623 7737 11664 7764
rect 11600 7731 11664 7737
rect 10936 7729 10969 7731
rect 10531 7723 10969 7729
rect 10531 7706 10537 7723
rect 10963 7706 10969 7723
rect 10531 7700 10969 7706
rect 11079 7729 11521 7731
rect 11081 7723 11519 7729
rect 11081 7706 11087 7723
rect 11513 7706 11519 7723
rect 11081 7700 11519 7706
rect 11631 7729 11664 7731
rect 12036 7737 12077 7764
rect 12094 7737 12100 8163
rect 12036 7731 12100 7737
rect 12150 8163 12650 8169
rect 12150 7737 12156 8163
rect 12173 8115 12627 8163
rect 12173 7785 12235 8115
rect 12565 7785 12627 8115
rect 12173 7737 12627 7785
rect 12644 7737 12650 8163
rect 12150 7731 12650 7737
rect 12700 8163 12764 8169
rect 12700 7737 12706 8163
rect 12723 8136 12764 8163
rect 13136 8169 13169 8171
rect 13281 8194 13719 8200
rect 13281 8177 13287 8194
rect 13713 8177 13719 8194
rect 13281 8171 13719 8177
rect 13279 8169 13721 8171
rect 13136 8163 13200 8169
rect 13136 8136 13177 8163
rect 12723 7764 12729 8136
rect 13171 7764 13177 8136
rect 12723 7737 12764 7764
rect 12700 7731 12764 7737
rect 12036 7729 12069 7731
rect 11631 7723 12069 7729
rect 11631 7706 11637 7723
rect 12063 7706 12069 7723
rect 11631 7700 12069 7706
rect 12179 7729 12621 7731
rect 12181 7723 12619 7729
rect 12181 7706 12187 7723
rect 12613 7706 12619 7723
rect 12181 7700 12619 7706
rect 12731 7729 12764 7731
rect 13136 7737 13177 7764
rect 13194 7737 13200 8163
rect 13136 7731 13200 7737
rect 13250 8163 13721 8169
rect 13250 7737 13256 8163
rect 13273 8115 13721 8163
rect 13273 7785 13335 8115
rect 13665 7785 13721 8115
rect 13273 7737 13721 7785
rect 13250 7731 13721 7737
rect 13136 7729 13169 7731
rect 12731 7723 13169 7729
rect 12731 7706 12737 7723
rect 13163 7706 13169 7723
rect 12731 7700 13169 7706
rect 13279 7729 13721 7731
rect 13281 7723 13719 7729
rect 13281 7706 13287 7723
rect 13713 7706 13719 7723
rect 13281 7700 13719 7706
rect -469 7644 -31 7650
rect -469 7627 -463 7644
rect -37 7627 -31 7644
rect -469 7621 -31 7627
rect -471 7619 -29 7621
rect 81 7644 519 7650
rect 81 7627 87 7644
rect 513 7627 519 7644
rect 81 7621 519 7627
rect 81 7619 114 7621
rect -471 7613 0 7619
rect -471 7565 -23 7613
rect -471 7235 -415 7565
rect -85 7235 -23 7565
rect -471 7187 -23 7235
rect -6 7187 0 7613
rect -471 7181 0 7187
rect 50 7613 114 7619
rect 50 7187 56 7613
rect 73 7586 114 7613
rect 486 7619 519 7621
rect 631 7644 1069 7650
rect 631 7627 637 7644
rect 1063 7627 1069 7644
rect 631 7621 1069 7627
rect 629 7619 1071 7621
rect 1181 7644 1619 7650
rect 1181 7627 1187 7644
rect 1613 7627 1619 7644
rect 1181 7621 1619 7627
rect 1181 7619 1214 7621
rect 486 7613 550 7619
rect 486 7586 527 7613
rect 73 7214 79 7586
rect 521 7214 527 7586
rect 73 7187 114 7214
rect 50 7181 114 7187
rect -471 7179 -29 7181
rect -469 7173 -31 7179
rect -469 7156 -463 7173
rect -37 7156 -31 7173
rect -469 7150 -31 7156
rect 81 7179 114 7181
rect 486 7187 527 7214
rect 544 7187 550 7613
rect 486 7181 550 7187
rect 600 7613 1100 7619
rect 600 7187 606 7613
rect 623 7565 1077 7613
rect 623 7235 685 7565
rect 1015 7235 1077 7565
rect 623 7187 1077 7235
rect 1094 7187 1100 7613
rect 600 7181 1100 7187
rect 1150 7613 1214 7619
rect 1150 7187 1156 7613
rect 1173 7586 1214 7613
rect 1586 7619 1619 7621
rect 1731 7644 2169 7650
rect 1731 7627 1737 7644
rect 2163 7627 2169 7644
rect 1731 7621 2169 7627
rect 1729 7619 2171 7621
rect 2281 7644 2719 7650
rect 2281 7627 2287 7644
rect 2713 7627 2719 7644
rect 2281 7621 2719 7627
rect 2281 7619 2314 7621
rect 1586 7613 1650 7619
rect 1586 7586 1627 7613
rect 1173 7214 1179 7586
rect 1621 7214 1627 7586
rect 1173 7187 1214 7214
rect 1150 7181 1214 7187
rect 486 7179 519 7181
rect 81 7173 519 7179
rect 81 7156 87 7173
rect 513 7156 519 7173
rect 81 7150 519 7156
rect 629 7179 1071 7181
rect 631 7173 1069 7179
rect 631 7156 637 7173
rect 1063 7156 1069 7173
rect 631 7150 1069 7156
rect 1181 7179 1214 7181
rect 1586 7187 1627 7214
rect 1644 7187 1650 7613
rect 1586 7181 1650 7187
rect 1700 7613 2200 7619
rect 1700 7187 1706 7613
rect 1723 7565 2177 7613
rect 1723 7235 1785 7565
rect 2115 7235 2177 7565
rect 1723 7187 2177 7235
rect 2194 7187 2200 7613
rect 1700 7181 2200 7187
rect 2250 7613 2314 7619
rect 2250 7187 2256 7613
rect 2273 7586 2314 7613
rect 2686 7619 2719 7621
rect 2831 7644 3269 7650
rect 2831 7627 2837 7644
rect 3263 7627 3269 7644
rect 2831 7621 3269 7627
rect 2829 7619 3271 7621
rect 3381 7644 3819 7650
rect 3381 7627 3387 7644
rect 3813 7627 3819 7644
rect 3381 7621 3819 7627
rect 3381 7619 3414 7621
rect 2686 7613 2750 7619
rect 2686 7586 2727 7613
rect 2273 7214 2279 7586
rect 2721 7214 2727 7586
rect 2273 7187 2314 7214
rect 2250 7181 2314 7187
rect 1586 7179 1619 7181
rect 1181 7173 1619 7179
rect 1181 7156 1187 7173
rect 1613 7156 1619 7173
rect 1181 7150 1619 7156
rect 1729 7179 2171 7181
rect 1731 7173 2169 7179
rect 1731 7156 1737 7173
rect 2163 7156 2169 7173
rect 1731 7150 2169 7156
rect 2281 7179 2314 7181
rect 2686 7187 2727 7214
rect 2744 7187 2750 7613
rect 2686 7181 2750 7187
rect 2800 7613 3300 7619
rect 2800 7187 2806 7613
rect 2823 7565 3277 7613
rect 2823 7235 2885 7565
rect 3215 7235 3277 7565
rect 2823 7187 3277 7235
rect 3294 7187 3300 7613
rect 2800 7181 3300 7187
rect 3350 7613 3414 7619
rect 3350 7187 3356 7613
rect 3373 7586 3414 7613
rect 3786 7619 3819 7621
rect 3931 7644 4369 7650
rect 3931 7627 3937 7644
rect 4363 7627 4369 7644
rect 3931 7621 4369 7627
rect 3929 7619 4371 7621
rect 4481 7644 4919 7650
rect 4481 7627 4487 7644
rect 4913 7627 4919 7644
rect 4481 7621 4919 7627
rect 4481 7619 4514 7621
rect 3786 7613 3850 7619
rect 3786 7586 3827 7613
rect 3373 7214 3379 7586
rect 3821 7214 3827 7586
rect 3373 7187 3414 7214
rect 3350 7181 3414 7187
rect 2686 7179 2719 7181
rect 2281 7173 2719 7179
rect 2281 7156 2287 7173
rect 2713 7156 2719 7173
rect 2281 7150 2719 7156
rect 2829 7179 3271 7181
rect 2831 7173 3269 7179
rect 2831 7156 2837 7173
rect 3263 7156 3269 7173
rect 2831 7150 3269 7156
rect 3381 7179 3414 7181
rect 3786 7187 3827 7214
rect 3844 7187 3850 7613
rect 3786 7181 3850 7187
rect 3900 7613 4400 7619
rect 3900 7187 3906 7613
rect 3923 7565 4377 7613
rect 3923 7235 3985 7565
rect 4315 7235 4377 7565
rect 3923 7187 4377 7235
rect 4394 7187 4400 7613
rect 3900 7181 4400 7187
rect 4450 7613 4514 7619
rect 4450 7187 4456 7613
rect 4473 7586 4514 7613
rect 4886 7619 4919 7621
rect 5031 7644 5469 7650
rect 5031 7627 5037 7644
rect 5463 7627 5469 7644
rect 5031 7621 5469 7627
rect 5029 7619 5471 7621
rect 5581 7644 6019 7650
rect 5581 7627 5587 7644
rect 6013 7627 6019 7644
rect 5581 7621 6019 7627
rect 5581 7619 5614 7621
rect 4886 7613 4950 7619
rect 4886 7586 4927 7613
rect 4473 7214 4479 7586
rect 4921 7214 4927 7586
rect 4473 7187 4514 7214
rect 4450 7181 4514 7187
rect 3786 7179 3819 7181
rect 3381 7173 3819 7179
rect 3381 7156 3387 7173
rect 3813 7156 3819 7173
rect 3381 7150 3819 7156
rect 3929 7179 4371 7181
rect 3931 7173 4369 7179
rect 3931 7156 3937 7173
rect 4363 7156 4369 7173
rect 3931 7150 4369 7156
rect 4481 7179 4514 7181
rect 4886 7187 4927 7214
rect 4944 7187 4950 7613
rect 4886 7181 4950 7187
rect 5000 7613 5500 7619
rect 5000 7187 5006 7613
rect 5023 7565 5477 7613
rect 5023 7235 5085 7565
rect 5415 7235 5477 7565
rect 5023 7187 5477 7235
rect 5494 7187 5500 7613
rect 5000 7181 5500 7187
rect 5550 7613 5614 7619
rect 5550 7187 5556 7613
rect 5573 7586 5614 7613
rect 5986 7619 6019 7621
rect 6131 7644 6569 7650
rect 6131 7627 6137 7644
rect 6563 7627 6569 7644
rect 6131 7621 6569 7627
rect 6129 7619 6571 7621
rect 6681 7644 7119 7650
rect 6681 7627 6687 7644
rect 7113 7627 7119 7644
rect 6681 7621 7119 7627
rect 6681 7619 6714 7621
rect 5986 7613 6050 7619
rect 5986 7586 6027 7613
rect 5573 7214 5579 7586
rect 6021 7214 6027 7586
rect 5573 7187 5614 7214
rect 5550 7181 5614 7187
rect 4886 7179 4919 7181
rect 4481 7173 4919 7179
rect 4481 7156 4487 7173
rect 4913 7156 4919 7173
rect 4481 7150 4919 7156
rect 5029 7179 5471 7181
rect 5031 7173 5469 7179
rect 5031 7156 5037 7173
rect 5463 7156 5469 7173
rect 5031 7150 5469 7156
rect 5581 7179 5614 7181
rect 5986 7187 6027 7214
rect 6044 7187 6050 7613
rect 5986 7181 6050 7187
rect 6100 7613 6600 7619
rect 6100 7187 6106 7613
rect 6123 7565 6577 7613
rect 6123 7235 6185 7565
rect 6515 7235 6577 7565
rect 6123 7187 6577 7235
rect 6594 7187 6600 7613
rect 6100 7181 6600 7187
rect 6650 7613 6714 7619
rect 6650 7187 6656 7613
rect 6673 7586 6714 7613
rect 7086 7619 7119 7621
rect 7231 7644 7669 7650
rect 7231 7627 7237 7644
rect 7663 7627 7669 7644
rect 7231 7621 7669 7627
rect 7229 7619 7671 7621
rect 7781 7644 8219 7650
rect 7781 7627 7787 7644
rect 8213 7627 8219 7644
rect 7781 7621 8219 7627
rect 7781 7619 7814 7621
rect 7086 7613 7150 7619
rect 7086 7586 7127 7613
rect 6673 7214 6679 7586
rect 7121 7214 7127 7586
rect 6673 7187 6714 7214
rect 6650 7181 6714 7187
rect 5986 7179 6019 7181
rect 5581 7173 6019 7179
rect 5581 7156 5587 7173
rect 6013 7156 6019 7173
rect 5581 7150 6019 7156
rect 6129 7179 6571 7181
rect 6131 7173 6569 7179
rect 6131 7156 6137 7173
rect 6563 7156 6569 7173
rect 6131 7150 6569 7156
rect 6681 7179 6714 7181
rect 7086 7187 7127 7214
rect 7144 7187 7150 7613
rect 7086 7181 7150 7187
rect 7200 7613 7700 7619
rect 7200 7187 7206 7613
rect 7223 7565 7677 7613
rect 7223 7235 7285 7565
rect 7615 7235 7677 7565
rect 7223 7187 7677 7235
rect 7694 7187 7700 7613
rect 7200 7181 7700 7187
rect 7750 7613 7814 7619
rect 7750 7187 7756 7613
rect 7773 7586 7814 7613
rect 8186 7619 8219 7621
rect 8331 7644 8769 7650
rect 8331 7627 8337 7644
rect 8763 7627 8769 7644
rect 8331 7621 8769 7627
rect 8329 7619 8771 7621
rect 8881 7644 9319 7650
rect 8881 7627 8887 7644
rect 9313 7627 9319 7644
rect 8881 7621 9319 7627
rect 8881 7619 8914 7621
rect 8186 7613 8250 7619
rect 8186 7586 8227 7613
rect 7773 7214 7779 7586
rect 8221 7214 8227 7586
rect 7773 7187 7814 7214
rect 7750 7181 7814 7187
rect 7086 7179 7119 7181
rect 6681 7173 7119 7179
rect 6681 7156 6687 7173
rect 7113 7156 7119 7173
rect 6681 7150 7119 7156
rect 7229 7179 7671 7181
rect 7231 7173 7669 7179
rect 7231 7156 7237 7173
rect 7663 7156 7669 7173
rect 7231 7150 7669 7156
rect 7781 7179 7814 7181
rect 8186 7187 8227 7214
rect 8244 7187 8250 7613
rect 8186 7181 8250 7187
rect 8300 7613 8800 7619
rect 8300 7187 8306 7613
rect 8323 7565 8777 7613
rect 8323 7235 8385 7565
rect 8715 7235 8777 7565
rect 8323 7187 8777 7235
rect 8794 7187 8800 7613
rect 8300 7181 8800 7187
rect 8850 7613 8914 7619
rect 8850 7187 8856 7613
rect 8873 7586 8914 7613
rect 9286 7619 9319 7621
rect 9431 7644 9869 7650
rect 9431 7627 9437 7644
rect 9863 7627 9869 7644
rect 9431 7621 9869 7627
rect 9429 7619 9871 7621
rect 9981 7644 10419 7650
rect 9981 7627 9987 7644
rect 10413 7627 10419 7644
rect 9981 7621 10419 7627
rect 9981 7619 10014 7621
rect 9286 7613 9350 7619
rect 9286 7586 9327 7613
rect 8873 7214 8879 7586
rect 9321 7214 9327 7586
rect 8873 7187 8914 7214
rect 8850 7181 8914 7187
rect 8186 7179 8219 7181
rect 7781 7173 8219 7179
rect 7781 7156 7787 7173
rect 8213 7156 8219 7173
rect 7781 7150 8219 7156
rect 8329 7179 8771 7181
rect 8331 7173 8769 7179
rect 8331 7156 8337 7173
rect 8763 7156 8769 7173
rect 8331 7150 8769 7156
rect 8881 7179 8914 7181
rect 9286 7187 9327 7214
rect 9344 7187 9350 7613
rect 9286 7181 9350 7187
rect 9400 7613 9900 7619
rect 9400 7187 9406 7613
rect 9423 7565 9877 7613
rect 9423 7235 9485 7565
rect 9815 7235 9877 7565
rect 9423 7187 9877 7235
rect 9894 7187 9900 7613
rect 9400 7181 9900 7187
rect 9950 7613 10014 7619
rect 9950 7187 9956 7613
rect 9973 7586 10014 7613
rect 10386 7619 10419 7621
rect 10531 7644 10969 7650
rect 10531 7627 10537 7644
rect 10963 7627 10969 7644
rect 10531 7621 10969 7627
rect 10529 7619 10971 7621
rect 11081 7644 11519 7650
rect 11081 7627 11087 7644
rect 11513 7627 11519 7644
rect 11081 7621 11519 7627
rect 11081 7619 11114 7621
rect 10386 7613 10450 7619
rect 10386 7586 10427 7613
rect 9973 7214 9979 7586
rect 10421 7214 10427 7586
rect 9973 7187 10014 7214
rect 9950 7181 10014 7187
rect 9286 7179 9319 7181
rect 8881 7173 9319 7179
rect 8881 7156 8887 7173
rect 9313 7156 9319 7173
rect 8881 7150 9319 7156
rect 9429 7179 9871 7181
rect 9431 7173 9869 7179
rect 9431 7156 9437 7173
rect 9863 7156 9869 7173
rect 9431 7150 9869 7156
rect 9981 7179 10014 7181
rect 10386 7187 10427 7214
rect 10444 7187 10450 7613
rect 10386 7181 10450 7187
rect 10500 7613 11000 7619
rect 10500 7187 10506 7613
rect 10523 7565 10977 7613
rect 10523 7235 10585 7565
rect 10915 7235 10977 7565
rect 10523 7187 10977 7235
rect 10994 7187 11000 7613
rect 10500 7181 11000 7187
rect 11050 7613 11114 7619
rect 11050 7187 11056 7613
rect 11073 7586 11114 7613
rect 11486 7619 11519 7621
rect 11631 7644 12069 7650
rect 11631 7627 11637 7644
rect 12063 7627 12069 7644
rect 11631 7621 12069 7627
rect 11629 7619 12071 7621
rect 12181 7644 12619 7650
rect 12181 7627 12187 7644
rect 12613 7627 12619 7644
rect 12181 7621 12619 7627
rect 12181 7619 12214 7621
rect 11486 7613 11550 7619
rect 11486 7586 11527 7613
rect 11073 7214 11079 7586
rect 11521 7214 11527 7586
rect 11073 7187 11114 7214
rect 11050 7181 11114 7187
rect 10386 7179 10419 7181
rect 9981 7173 10419 7179
rect 9981 7156 9987 7173
rect 10413 7156 10419 7173
rect 9981 7150 10419 7156
rect 10529 7179 10971 7181
rect 10531 7173 10969 7179
rect 10531 7156 10537 7173
rect 10963 7156 10969 7173
rect 10531 7150 10969 7156
rect 11081 7179 11114 7181
rect 11486 7187 11527 7214
rect 11544 7187 11550 7613
rect 11486 7181 11550 7187
rect 11600 7613 12100 7619
rect 11600 7187 11606 7613
rect 11623 7565 12077 7613
rect 11623 7235 11685 7565
rect 12015 7235 12077 7565
rect 11623 7187 12077 7235
rect 12094 7187 12100 7613
rect 11600 7181 12100 7187
rect 12150 7613 12214 7619
rect 12150 7187 12156 7613
rect 12173 7586 12214 7613
rect 12586 7619 12619 7621
rect 12731 7644 13169 7650
rect 12731 7627 12737 7644
rect 13163 7627 13169 7644
rect 12731 7621 13169 7627
rect 12729 7619 13171 7621
rect 13281 7644 13719 7650
rect 13281 7627 13287 7644
rect 13713 7627 13719 7644
rect 13281 7621 13719 7627
rect 13281 7619 13314 7621
rect 12586 7613 12650 7619
rect 12586 7586 12627 7613
rect 12173 7214 12179 7586
rect 12621 7214 12627 7586
rect 12173 7187 12214 7214
rect 12150 7181 12214 7187
rect 11486 7179 11519 7181
rect 11081 7173 11519 7179
rect 11081 7156 11087 7173
rect 11513 7156 11519 7173
rect 11081 7150 11519 7156
rect 11629 7179 12071 7181
rect 11631 7173 12069 7179
rect 11631 7156 11637 7173
rect 12063 7156 12069 7173
rect 11631 7150 12069 7156
rect 12181 7179 12214 7181
rect 12586 7187 12627 7214
rect 12644 7187 12650 7613
rect 12586 7181 12650 7187
rect 12700 7613 13200 7619
rect 12700 7187 12706 7613
rect 12723 7565 13177 7613
rect 12723 7235 12785 7565
rect 13115 7235 13177 7565
rect 12723 7187 13177 7235
rect 13194 7187 13200 7613
rect 12700 7181 13200 7187
rect 13250 7613 13314 7619
rect 13250 7187 13256 7613
rect 13273 7586 13314 7613
rect 13273 7214 13279 7586
rect 13273 7187 13314 7214
rect 13250 7181 13314 7187
rect 12586 7179 12619 7181
rect 12181 7173 12619 7179
rect 12181 7156 12187 7173
rect 12613 7156 12619 7173
rect 12181 7150 12619 7156
rect 12729 7179 13171 7181
rect 12731 7173 13169 7179
rect 12731 7156 12737 7173
rect 13163 7156 13169 7173
rect 12731 7150 13169 7156
rect 13281 7179 13314 7181
rect 13281 7173 13719 7179
rect 13281 7156 13287 7173
rect 13713 7156 13719 7173
rect 13281 7150 13719 7156
rect -469 7094 -31 7100
rect -469 7077 -463 7094
rect -37 7077 -31 7094
rect -469 7071 -31 7077
rect -64 7069 -31 7071
rect 81 7094 519 7100
rect 81 7077 87 7094
rect 513 7077 519 7094
rect 81 7071 519 7077
rect 79 7069 521 7071
rect 631 7094 1069 7100
rect 631 7077 637 7094
rect 1063 7077 1069 7094
rect 631 7071 1069 7077
rect 631 7069 664 7071
rect -64 7063 0 7069
rect -64 7036 -23 7063
rect -29 6664 -23 7036
rect -64 6637 -23 6664
rect -6 6637 0 7063
rect -64 6631 0 6637
rect 50 7063 550 7069
rect 50 6637 56 7063
rect 73 7015 527 7063
rect 73 6685 135 7015
rect 465 6685 527 7015
rect 73 6637 527 6685
rect 544 6637 550 7063
rect 50 6631 550 6637
rect 600 7063 664 7069
rect 600 6637 606 7063
rect 623 7036 664 7063
rect 1036 7069 1069 7071
rect 1181 7094 1619 7100
rect 1181 7077 1187 7094
rect 1613 7077 1619 7094
rect 1181 7071 1619 7077
rect 1179 7069 1621 7071
rect 1731 7094 2169 7100
rect 1731 7077 1737 7094
rect 2163 7077 2169 7094
rect 1731 7071 2169 7077
rect 1731 7069 1764 7071
rect 1036 7063 1100 7069
rect 1036 7036 1077 7063
rect 623 6664 629 7036
rect 1071 6664 1077 7036
rect 623 6637 664 6664
rect 600 6631 664 6637
rect -64 6629 -31 6631
rect -469 6623 -31 6629
rect -469 6606 -463 6623
rect -37 6606 -31 6623
rect -469 6600 -31 6606
rect 79 6629 521 6631
rect 81 6623 519 6629
rect 81 6606 87 6623
rect 513 6606 519 6623
rect 81 6600 519 6606
rect 631 6629 664 6631
rect 1036 6637 1077 6664
rect 1094 6637 1100 7063
rect 1036 6631 1100 6637
rect 1150 7063 1650 7069
rect 1150 6637 1156 7063
rect 1173 7015 1627 7063
rect 1173 6685 1235 7015
rect 1565 6685 1627 7015
rect 1173 6637 1627 6685
rect 1644 6637 1650 7063
rect 1150 6631 1650 6637
rect 1700 7063 1764 7069
rect 1700 6637 1706 7063
rect 1723 7036 1764 7063
rect 2136 7069 2169 7071
rect 2281 7094 2719 7100
rect 2281 7077 2287 7094
rect 2713 7077 2719 7094
rect 2281 7071 2719 7077
rect 2279 7069 2721 7071
rect 2831 7094 3269 7100
rect 2831 7077 2837 7094
rect 3263 7077 3269 7094
rect 2831 7071 3269 7077
rect 2831 7069 2864 7071
rect 2136 7063 2200 7069
rect 2136 7036 2177 7063
rect 1723 6664 1729 7036
rect 2171 6664 2177 7036
rect 1723 6637 1764 6664
rect 1700 6631 1764 6637
rect 1036 6629 1069 6631
rect 631 6623 1069 6629
rect 631 6606 637 6623
rect 1063 6606 1069 6623
rect 631 6600 1069 6606
rect 1179 6629 1621 6631
rect 1181 6623 1619 6629
rect 1181 6606 1187 6623
rect 1613 6606 1619 6623
rect 1181 6600 1619 6606
rect 1731 6629 1764 6631
rect 2136 6637 2177 6664
rect 2194 6637 2200 7063
rect 2136 6631 2200 6637
rect 2250 7063 2750 7069
rect 2250 6637 2256 7063
rect 2273 7015 2727 7063
rect 2273 6685 2335 7015
rect 2665 6685 2727 7015
rect 2273 6637 2727 6685
rect 2744 6637 2750 7063
rect 2250 6631 2750 6637
rect 2800 7063 2864 7069
rect 2800 6637 2806 7063
rect 2823 7036 2864 7063
rect 3236 7069 3269 7071
rect 3381 7094 3819 7100
rect 3381 7077 3387 7094
rect 3813 7077 3819 7094
rect 3381 7071 3819 7077
rect 3379 7069 3821 7071
rect 3931 7094 4369 7100
rect 3931 7077 3937 7094
rect 4363 7077 4369 7094
rect 3931 7071 4369 7077
rect 3931 7069 3964 7071
rect 3236 7063 3300 7069
rect 3236 7036 3277 7063
rect 2823 6664 2829 7036
rect 3271 6664 3277 7036
rect 2823 6637 2864 6664
rect 2800 6631 2864 6637
rect 2136 6629 2169 6631
rect 1731 6623 2169 6629
rect 1731 6606 1737 6623
rect 2163 6606 2169 6623
rect 1731 6600 2169 6606
rect 2279 6629 2721 6631
rect 2281 6623 2719 6629
rect 2281 6606 2287 6623
rect 2713 6606 2719 6623
rect 2281 6600 2719 6606
rect 2831 6629 2864 6631
rect 3236 6637 3277 6664
rect 3294 6637 3300 7063
rect 3236 6631 3300 6637
rect 3350 7063 3850 7069
rect 3350 6637 3356 7063
rect 3373 7015 3827 7063
rect 3373 6685 3435 7015
rect 3765 6685 3827 7015
rect 3373 6637 3827 6685
rect 3844 6637 3850 7063
rect 3350 6631 3850 6637
rect 3900 7063 3964 7069
rect 3900 6637 3906 7063
rect 3923 7036 3964 7063
rect 4336 7069 4369 7071
rect 4481 7094 4919 7100
rect 4481 7077 4487 7094
rect 4913 7077 4919 7094
rect 4481 7071 4919 7077
rect 4479 7069 4921 7071
rect 5031 7094 5469 7100
rect 5031 7077 5037 7094
rect 5463 7077 5469 7094
rect 5031 7071 5469 7077
rect 5031 7069 5064 7071
rect 4336 7063 4400 7069
rect 4336 7036 4377 7063
rect 3923 6664 3929 7036
rect 4371 6664 4377 7036
rect 3923 6637 3964 6664
rect 3900 6631 3964 6637
rect 3236 6629 3269 6631
rect 2831 6623 3269 6629
rect 2831 6606 2837 6623
rect 3263 6606 3269 6623
rect 2831 6600 3269 6606
rect 3379 6629 3821 6631
rect 3381 6623 3819 6629
rect 3381 6606 3387 6623
rect 3813 6606 3819 6623
rect 3381 6600 3819 6606
rect 3931 6629 3964 6631
rect 4336 6637 4377 6664
rect 4394 6637 4400 7063
rect 4336 6631 4400 6637
rect 4450 7063 4950 7069
rect 4450 6637 4456 7063
rect 4473 7015 4927 7063
rect 4473 6685 4535 7015
rect 4865 6685 4927 7015
rect 4473 6637 4927 6685
rect 4944 6637 4950 7063
rect 4450 6631 4950 6637
rect 5000 7063 5064 7069
rect 5000 6637 5006 7063
rect 5023 7036 5064 7063
rect 5436 7069 5469 7071
rect 5581 7094 6019 7100
rect 5581 7077 5587 7094
rect 6013 7077 6019 7094
rect 5581 7071 6019 7077
rect 5579 7069 6021 7071
rect 6131 7094 6569 7100
rect 6131 7077 6137 7094
rect 6563 7077 6569 7094
rect 6131 7071 6569 7077
rect 6131 7069 6164 7071
rect 5436 7063 5500 7069
rect 5436 7036 5477 7063
rect 5023 6664 5029 7036
rect 5471 6664 5477 7036
rect 5023 6637 5064 6664
rect 5000 6631 5064 6637
rect 4336 6629 4369 6631
rect 3931 6623 4369 6629
rect 3931 6606 3937 6623
rect 4363 6606 4369 6623
rect 3931 6600 4369 6606
rect 4479 6629 4921 6631
rect 4481 6623 4919 6629
rect 4481 6606 4487 6623
rect 4913 6606 4919 6623
rect 4481 6600 4919 6606
rect 5031 6629 5064 6631
rect 5436 6637 5477 6664
rect 5494 6637 5500 7063
rect 5436 6631 5500 6637
rect 5550 7063 6050 7069
rect 5550 6637 5556 7063
rect 5573 7015 6027 7063
rect 5573 6685 5635 7015
rect 5965 6685 6027 7015
rect 5573 6637 6027 6685
rect 6044 6637 6050 7063
rect 5550 6631 6050 6637
rect 6100 7063 6164 7069
rect 6100 6637 6106 7063
rect 6123 7036 6164 7063
rect 6536 7069 6569 7071
rect 6681 7094 7119 7100
rect 6681 7077 6687 7094
rect 7113 7077 7119 7094
rect 6681 7071 7119 7077
rect 6679 7069 7121 7071
rect 7231 7094 7669 7100
rect 7231 7077 7237 7094
rect 7663 7077 7669 7094
rect 7231 7071 7669 7077
rect 7231 7069 7264 7071
rect 6536 7063 6600 7069
rect 6536 7036 6577 7063
rect 6123 6664 6129 7036
rect 6571 6664 6577 7036
rect 6123 6637 6164 6664
rect 6100 6631 6164 6637
rect 5436 6629 5469 6631
rect 5031 6623 5469 6629
rect 5031 6606 5037 6623
rect 5463 6606 5469 6623
rect 5031 6600 5469 6606
rect 5579 6629 6021 6631
rect 5581 6623 6019 6629
rect 5581 6606 5587 6623
rect 6013 6606 6019 6623
rect 5581 6600 6019 6606
rect 6131 6629 6164 6631
rect 6536 6637 6577 6664
rect 6594 6637 6600 7063
rect 6536 6631 6600 6637
rect 6650 7063 7150 7069
rect 6650 6637 6656 7063
rect 6673 7015 7127 7063
rect 6673 6685 6735 7015
rect 7065 6685 7127 7015
rect 6673 6637 7127 6685
rect 7144 6637 7150 7063
rect 6650 6631 7150 6637
rect 7200 7063 7264 7069
rect 7200 6637 7206 7063
rect 7223 7036 7264 7063
rect 7636 7069 7669 7071
rect 7781 7094 8219 7100
rect 7781 7077 7787 7094
rect 8213 7077 8219 7094
rect 7781 7071 8219 7077
rect 7779 7069 8221 7071
rect 8331 7094 8769 7100
rect 8331 7077 8337 7094
rect 8763 7077 8769 7094
rect 8331 7071 8769 7077
rect 8331 7069 8364 7071
rect 7636 7063 7700 7069
rect 7636 7036 7677 7063
rect 7223 6664 7229 7036
rect 7671 6664 7677 7036
rect 7223 6637 7264 6664
rect 7200 6631 7264 6637
rect 6536 6629 6569 6631
rect 6131 6623 6569 6629
rect 6131 6606 6137 6623
rect 6563 6606 6569 6623
rect 6131 6600 6569 6606
rect 6679 6629 7121 6631
rect 6681 6623 7119 6629
rect 6681 6606 6687 6623
rect 7113 6606 7119 6623
rect 6681 6600 7119 6606
rect 7231 6629 7264 6631
rect 7636 6637 7677 6664
rect 7694 6637 7700 7063
rect 7636 6631 7700 6637
rect 7750 7063 8250 7069
rect 7750 6637 7756 7063
rect 7773 7015 8227 7063
rect 7773 6685 7835 7015
rect 8165 6685 8227 7015
rect 7773 6637 8227 6685
rect 8244 6637 8250 7063
rect 7750 6631 8250 6637
rect 8300 7063 8364 7069
rect 8300 6637 8306 7063
rect 8323 7036 8364 7063
rect 8736 7069 8769 7071
rect 8881 7094 9319 7100
rect 8881 7077 8887 7094
rect 9313 7077 9319 7094
rect 8881 7071 9319 7077
rect 8879 7069 9321 7071
rect 9431 7094 9869 7100
rect 9431 7077 9437 7094
rect 9863 7077 9869 7094
rect 9431 7071 9869 7077
rect 9431 7069 9464 7071
rect 8736 7063 8800 7069
rect 8736 7036 8777 7063
rect 8323 6664 8329 7036
rect 8771 6664 8777 7036
rect 8323 6637 8364 6664
rect 8300 6631 8364 6637
rect 7636 6629 7669 6631
rect 7231 6623 7669 6629
rect 7231 6606 7237 6623
rect 7663 6606 7669 6623
rect 7231 6600 7669 6606
rect 7779 6629 8221 6631
rect 7781 6623 8219 6629
rect 7781 6606 7787 6623
rect 8213 6606 8219 6623
rect 7781 6600 8219 6606
rect 8331 6629 8364 6631
rect 8736 6637 8777 6664
rect 8794 6637 8800 7063
rect 8736 6631 8800 6637
rect 8850 7063 9350 7069
rect 8850 6637 8856 7063
rect 8873 7015 9327 7063
rect 8873 6685 8935 7015
rect 9265 6685 9327 7015
rect 8873 6637 9327 6685
rect 9344 6637 9350 7063
rect 8850 6631 9350 6637
rect 9400 7063 9464 7069
rect 9400 6637 9406 7063
rect 9423 7036 9464 7063
rect 9836 7069 9869 7071
rect 9981 7094 10419 7100
rect 9981 7077 9987 7094
rect 10413 7077 10419 7094
rect 9981 7071 10419 7077
rect 9979 7069 10421 7071
rect 10531 7094 10969 7100
rect 10531 7077 10537 7094
rect 10963 7077 10969 7094
rect 10531 7071 10969 7077
rect 10531 7069 10564 7071
rect 9836 7063 9900 7069
rect 9836 7036 9877 7063
rect 9423 6664 9429 7036
rect 9871 6664 9877 7036
rect 9423 6637 9464 6664
rect 9400 6631 9464 6637
rect 8736 6629 8769 6631
rect 8331 6623 8769 6629
rect 8331 6606 8337 6623
rect 8763 6606 8769 6623
rect 8331 6600 8769 6606
rect 8879 6629 9321 6631
rect 8881 6623 9319 6629
rect 8881 6606 8887 6623
rect 9313 6606 9319 6623
rect 8881 6600 9319 6606
rect 9431 6629 9464 6631
rect 9836 6637 9877 6664
rect 9894 6637 9900 7063
rect 9836 6631 9900 6637
rect 9950 7063 10450 7069
rect 9950 6637 9956 7063
rect 9973 7015 10427 7063
rect 9973 6685 10035 7015
rect 10365 6685 10427 7015
rect 9973 6637 10427 6685
rect 10444 6637 10450 7063
rect 9950 6631 10450 6637
rect 10500 7063 10564 7069
rect 10500 6637 10506 7063
rect 10523 7036 10564 7063
rect 10936 7069 10969 7071
rect 11081 7094 11519 7100
rect 11081 7077 11087 7094
rect 11513 7077 11519 7094
rect 11081 7071 11519 7077
rect 11079 7069 11521 7071
rect 11631 7094 12069 7100
rect 11631 7077 11637 7094
rect 12063 7077 12069 7094
rect 11631 7071 12069 7077
rect 11631 7069 11664 7071
rect 10936 7063 11000 7069
rect 10936 7036 10977 7063
rect 10523 6664 10529 7036
rect 10971 6664 10977 7036
rect 10523 6637 10564 6664
rect 10500 6631 10564 6637
rect 9836 6629 9869 6631
rect 9431 6623 9869 6629
rect 9431 6606 9437 6623
rect 9863 6606 9869 6623
rect 9431 6600 9869 6606
rect 9979 6629 10421 6631
rect 9981 6623 10419 6629
rect 9981 6606 9987 6623
rect 10413 6606 10419 6623
rect 9981 6600 10419 6606
rect 10531 6629 10564 6631
rect 10936 6637 10977 6664
rect 10994 6637 11000 7063
rect 10936 6631 11000 6637
rect 11050 7063 11550 7069
rect 11050 6637 11056 7063
rect 11073 7015 11527 7063
rect 11073 6685 11135 7015
rect 11465 6685 11527 7015
rect 11073 6637 11527 6685
rect 11544 6637 11550 7063
rect 11050 6631 11550 6637
rect 11600 7063 11664 7069
rect 11600 6637 11606 7063
rect 11623 7036 11664 7063
rect 12036 7069 12069 7071
rect 12181 7094 12619 7100
rect 12181 7077 12187 7094
rect 12613 7077 12619 7094
rect 12181 7071 12619 7077
rect 12179 7069 12621 7071
rect 12731 7094 13169 7100
rect 12731 7077 12737 7094
rect 13163 7077 13169 7094
rect 12731 7071 13169 7077
rect 12731 7069 12764 7071
rect 12036 7063 12100 7069
rect 12036 7036 12077 7063
rect 11623 6664 11629 7036
rect 12071 6664 12077 7036
rect 11623 6637 11664 6664
rect 11600 6631 11664 6637
rect 10936 6629 10969 6631
rect 10531 6623 10969 6629
rect 10531 6606 10537 6623
rect 10963 6606 10969 6623
rect 10531 6600 10969 6606
rect 11079 6629 11521 6631
rect 11081 6623 11519 6629
rect 11081 6606 11087 6623
rect 11513 6606 11519 6623
rect 11081 6600 11519 6606
rect 11631 6629 11664 6631
rect 12036 6637 12077 6664
rect 12094 6637 12100 7063
rect 12036 6631 12100 6637
rect 12150 7063 12650 7069
rect 12150 6637 12156 7063
rect 12173 7015 12627 7063
rect 12173 6685 12235 7015
rect 12565 6685 12627 7015
rect 12173 6637 12627 6685
rect 12644 6637 12650 7063
rect 12150 6631 12650 6637
rect 12700 7063 12764 7069
rect 12700 6637 12706 7063
rect 12723 7036 12764 7063
rect 13136 7069 13169 7071
rect 13281 7094 13719 7100
rect 13281 7077 13287 7094
rect 13713 7077 13719 7094
rect 13281 7071 13719 7077
rect 13279 7069 13721 7071
rect 13136 7063 13200 7069
rect 13136 7036 13177 7063
rect 12723 6664 12729 7036
rect 13171 6664 13177 7036
rect 12723 6637 12764 6664
rect 12700 6631 12764 6637
rect 12036 6629 12069 6631
rect 11631 6623 12069 6629
rect 11631 6606 11637 6623
rect 12063 6606 12069 6623
rect 11631 6600 12069 6606
rect 12179 6629 12621 6631
rect 12181 6623 12619 6629
rect 12181 6606 12187 6623
rect 12613 6606 12619 6623
rect 12181 6600 12619 6606
rect 12731 6629 12764 6631
rect 13136 6637 13177 6664
rect 13194 6637 13200 7063
rect 13136 6631 13200 6637
rect 13250 7063 13721 7069
rect 13250 6637 13256 7063
rect 13273 7015 13721 7063
rect 13273 6685 13335 7015
rect 13665 6685 13721 7015
rect 13273 6637 13721 6685
rect 13250 6631 13721 6637
rect 13136 6629 13169 6631
rect 12731 6623 13169 6629
rect 12731 6606 12737 6623
rect 13163 6606 13169 6623
rect 12731 6600 13169 6606
rect 13279 6629 13721 6631
rect 13281 6623 13719 6629
rect 13281 6606 13287 6623
rect 13713 6606 13719 6623
rect 13281 6600 13719 6606
rect -469 6544 -31 6550
rect -469 6527 -463 6544
rect -37 6527 -31 6544
rect -469 6521 -31 6527
rect -471 6519 -29 6521
rect 81 6544 519 6550
rect 81 6527 87 6544
rect 513 6527 519 6544
rect 81 6521 519 6527
rect 81 6519 114 6521
rect -471 6513 0 6519
rect -471 6465 -23 6513
rect -471 6135 -415 6465
rect -85 6135 -23 6465
rect -471 6087 -23 6135
rect -6 6087 0 6513
rect -471 6081 0 6087
rect 50 6513 114 6519
rect 50 6087 56 6513
rect 73 6486 114 6513
rect 486 6519 519 6521
rect 631 6544 1069 6550
rect 631 6527 637 6544
rect 1063 6527 1069 6544
rect 631 6521 1069 6527
rect 629 6519 1071 6521
rect 1181 6544 1619 6550
rect 1181 6527 1187 6544
rect 1613 6527 1619 6544
rect 1181 6521 1619 6527
rect 1181 6519 1214 6521
rect 486 6513 550 6519
rect 486 6486 527 6513
rect 73 6114 79 6486
rect 521 6114 527 6486
rect 73 6087 114 6114
rect 50 6081 114 6087
rect -471 6079 -29 6081
rect -469 6073 -31 6079
rect -469 6056 -463 6073
rect -37 6056 -31 6073
rect -469 6050 -31 6056
rect 81 6079 114 6081
rect 486 6087 527 6114
rect 544 6087 550 6513
rect 486 6081 550 6087
rect 600 6513 1100 6519
rect 600 6087 606 6513
rect 623 6465 1077 6513
rect 623 6135 685 6465
rect 1015 6135 1077 6465
rect 623 6087 1077 6135
rect 1094 6087 1100 6513
rect 600 6081 1100 6087
rect 1150 6513 1214 6519
rect 1150 6087 1156 6513
rect 1173 6486 1214 6513
rect 1586 6519 1619 6521
rect 1731 6544 2169 6550
rect 1731 6527 1737 6544
rect 2163 6527 2169 6544
rect 1731 6521 2169 6527
rect 1729 6519 2171 6521
rect 2281 6544 2719 6550
rect 2281 6527 2287 6544
rect 2713 6527 2719 6544
rect 2281 6521 2719 6527
rect 2281 6519 2314 6521
rect 1586 6513 1650 6519
rect 1586 6486 1627 6513
rect 1173 6114 1179 6486
rect 1621 6114 1627 6486
rect 1173 6087 1214 6114
rect 1150 6081 1214 6087
rect 486 6079 519 6081
rect 81 6073 519 6079
rect 81 6056 87 6073
rect 513 6056 519 6073
rect 81 6050 519 6056
rect 629 6079 1071 6081
rect 631 6073 1069 6079
rect 631 6056 637 6073
rect 1063 6056 1069 6073
rect 631 6050 1069 6056
rect 1181 6079 1214 6081
rect 1586 6087 1627 6114
rect 1644 6087 1650 6513
rect 1586 6081 1650 6087
rect 1700 6513 2200 6519
rect 1700 6087 1706 6513
rect 1723 6465 2177 6513
rect 1723 6135 1785 6465
rect 2115 6135 2177 6465
rect 1723 6087 2177 6135
rect 2194 6087 2200 6513
rect 1700 6081 2200 6087
rect 2250 6513 2314 6519
rect 2250 6087 2256 6513
rect 2273 6486 2314 6513
rect 2686 6519 2719 6521
rect 2831 6544 3269 6550
rect 2831 6527 2837 6544
rect 3263 6527 3269 6544
rect 2831 6521 3269 6527
rect 2829 6519 3271 6521
rect 3381 6544 3819 6550
rect 3381 6527 3387 6544
rect 3813 6527 3819 6544
rect 3381 6521 3819 6527
rect 3381 6519 3414 6521
rect 2686 6513 2750 6519
rect 2686 6486 2727 6513
rect 2273 6114 2279 6486
rect 2721 6114 2727 6486
rect 2273 6087 2314 6114
rect 2250 6081 2314 6087
rect 1586 6079 1619 6081
rect 1181 6073 1619 6079
rect 1181 6056 1187 6073
rect 1613 6056 1619 6073
rect 1181 6050 1619 6056
rect 1729 6079 2171 6081
rect 1731 6073 2169 6079
rect 1731 6056 1737 6073
rect 2163 6056 2169 6073
rect 1731 6050 2169 6056
rect 2281 6079 2314 6081
rect 2686 6087 2727 6114
rect 2744 6087 2750 6513
rect 2686 6081 2750 6087
rect 2800 6513 3300 6519
rect 2800 6087 2806 6513
rect 2823 6465 3277 6513
rect 2823 6135 2885 6465
rect 3215 6135 3277 6465
rect 2823 6087 3277 6135
rect 3294 6087 3300 6513
rect 2800 6081 3300 6087
rect 3350 6513 3414 6519
rect 3350 6087 3356 6513
rect 3373 6486 3414 6513
rect 3786 6519 3819 6521
rect 3931 6544 4369 6550
rect 3931 6527 3937 6544
rect 4363 6527 4369 6544
rect 3931 6521 4369 6527
rect 3929 6519 4371 6521
rect 4481 6544 4919 6550
rect 4481 6527 4487 6544
rect 4913 6527 4919 6544
rect 4481 6521 4919 6527
rect 4481 6519 4514 6521
rect 3786 6513 3850 6519
rect 3786 6486 3827 6513
rect 3373 6114 3379 6486
rect 3821 6114 3827 6486
rect 3373 6087 3414 6114
rect 3350 6081 3414 6087
rect 2686 6079 2719 6081
rect 2281 6073 2719 6079
rect 2281 6056 2287 6073
rect 2713 6056 2719 6073
rect 2281 6050 2719 6056
rect 2829 6079 3271 6081
rect 2831 6073 3269 6079
rect 2831 6056 2837 6073
rect 3263 6056 3269 6073
rect 2831 6050 3269 6056
rect 3381 6079 3414 6081
rect 3786 6087 3827 6114
rect 3844 6087 3850 6513
rect 3786 6081 3850 6087
rect 3900 6513 4400 6519
rect 3900 6087 3906 6513
rect 3923 6465 4377 6513
rect 3923 6135 3985 6465
rect 4315 6135 4377 6465
rect 3923 6087 4377 6135
rect 4394 6087 4400 6513
rect 3900 6081 4400 6087
rect 4450 6513 4514 6519
rect 4450 6087 4456 6513
rect 4473 6486 4514 6513
rect 4886 6519 4919 6521
rect 5031 6544 5469 6550
rect 5031 6527 5037 6544
rect 5463 6527 5469 6544
rect 5031 6521 5469 6527
rect 5029 6519 5471 6521
rect 5581 6544 6019 6550
rect 5581 6527 5587 6544
rect 6013 6527 6019 6544
rect 5581 6521 6019 6527
rect 5581 6519 5614 6521
rect 4886 6513 4950 6519
rect 4886 6486 4927 6513
rect 4473 6114 4479 6486
rect 4921 6114 4927 6486
rect 4473 6087 4514 6114
rect 4450 6081 4514 6087
rect 3786 6079 3819 6081
rect 3381 6073 3819 6079
rect 3381 6056 3387 6073
rect 3813 6056 3819 6073
rect 3381 6050 3819 6056
rect 3929 6079 4371 6081
rect 3931 6073 4369 6079
rect 3931 6056 3937 6073
rect 4363 6056 4369 6073
rect 3931 6050 4369 6056
rect 4481 6079 4514 6081
rect 4886 6087 4927 6114
rect 4944 6087 4950 6513
rect 4886 6081 4950 6087
rect 5000 6513 5500 6519
rect 5000 6087 5006 6513
rect 5023 6465 5477 6513
rect 5023 6135 5085 6465
rect 5415 6135 5477 6465
rect 5023 6087 5477 6135
rect 5494 6087 5500 6513
rect 5000 6081 5500 6087
rect 5550 6513 5614 6519
rect 5550 6087 5556 6513
rect 5573 6486 5614 6513
rect 5986 6519 6019 6521
rect 6131 6544 6569 6550
rect 6131 6527 6137 6544
rect 6563 6527 6569 6544
rect 6131 6521 6569 6527
rect 6129 6519 6571 6521
rect 6681 6544 7119 6550
rect 6681 6527 6687 6544
rect 7113 6527 7119 6544
rect 6681 6521 7119 6527
rect 6681 6519 6714 6521
rect 5986 6513 6050 6519
rect 5986 6486 6027 6513
rect 5573 6114 5579 6486
rect 6021 6114 6027 6486
rect 5573 6087 5614 6114
rect 5550 6081 5614 6087
rect 4886 6079 4919 6081
rect 4481 6073 4919 6079
rect 4481 6056 4487 6073
rect 4913 6056 4919 6073
rect 4481 6050 4919 6056
rect 5029 6079 5471 6081
rect 5031 6073 5469 6079
rect 5031 6056 5037 6073
rect 5463 6056 5469 6073
rect 5031 6050 5469 6056
rect 5581 6079 5614 6081
rect 5986 6087 6027 6114
rect 6044 6087 6050 6513
rect 5986 6081 6050 6087
rect 6100 6513 6600 6519
rect 6100 6087 6106 6513
rect 6123 6465 6577 6513
rect 6123 6135 6185 6465
rect 6515 6135 6577 6465
rect 6123 6087 6577 6135
rect 6594 6087 6600 6513
rect 6100 6081 6600 6087
rect 6650 6513 6714 6519
rect 6650 6087 6656 6513
rect 6673 6486 6714 6513
rect 7086 6519 7119 6521
rect 7231 6544 7669 6550
rect 7231 6527 7237 6544
rect 7663 6527 7669 6544
rect 7231 6521 7669 6527
rect 7229 6519 7671 6521
rect 7781 6544 8219 6550
rect 7781 6527 7787 6544
rect 8213 6527 8219 6544
rect 7781 6521 8219 6527
rect 7781 6519 7814 6521
rect 7086 6513 7150 6519
rect 7086 6486 7127 6513
rect 6673 6114 6679 6486
rect 7121 6114 7127 6486
rect 6673 6087 6714 6114
rect 6650 6081 6714 6087
rect 5986 6079 6019 6081
rect 5581 6073 6019 6079
rect 5581 6056 5587 6073
rect 6013 6056 6019 6073
rect 5581 6050 6019 6056
rect 6129 6079 6571 6081
rect 6131 6073 6569 6079
rect 6131 6056 6137 6073
rect 6563 6056 6569 6073
rect 6131 6050 6569 6056
rect 6681 6079 6714 6081
rect 7086 6087 7127 6114
rect 7144 6087 7150 6513
rect 7086 6081 7150 6087
rect 7200 6513 7700 6519
rect 7200 6087 7206 6513
rect 7223 6465 7677 6513
rect 7223 6135 7285 6465
rect 7615 6135 7677 6465
rect 7223 6087 7677 6135
rect 7694 6087 7700 6513
rect 7200 6081 7700 6087
rect 7750 6513 7814 6519
rect 7750 6087 7756 6513
rect 7773 6486 7814 6513
rect 8186 6519 8219 6521
rect 8331 6544 8769 6550
rect 8331 6527 8337 6544
rect 8763 6527 8769 6544
rect 8331 6521 8769 6527
rect 8329 6519 8771 6521
rect 8881 6544 9319 6550
rect 8881 6527 8887 6544
rect 9313 6527 9319 6544
rect 8881 6521 9319 6527
rect 8881 6519 8914 6521
rect 8186 6513 8250 6519
rect 8186 6486 8227 6513
rect 7773 6114 7779 6486
rect 8221 6114 8227 6486
rect 7773 6087 7814 6114
rect 7750 6081 7814 6087
rect 7086 6079 7119 6081
rect 6681 6073 7119 6079
rect 6681 6056 6687 6073
rect 7113 6056 7119 6073
rect 6681 6050 7119 6056
rect 7229 6079 7671 6081
rect 7231 6073 7669 6079
rect 7231 6056 7237 6073
rect 7663 6056 7669 6073
rect 7231 6050 7669 6056
rect 7781 6079 7814 6081
rect 8186 6087 8227 6114
rect 8244 6087 8250 6513
rect 8186 6081 8250 6087
rect 8300 6513 8800 6519
rect 8300 6087 8306 6513
rect 8323 6465 8777 6513
rect 8323 6135 8385 6465
rect 8715 6135 8777 6465
rect 8323 6087 8777 6135
rect 8794 6087 8800 6513
rect 8300 6081 8800 6087
rect 8850 6513 8914 6519
rect 8850 6087 8856 6513
rect 8873 6486 8914 6513
rect 9286 6519 9319 6521
rect 9431 6544 9869 6550
rect 9431 6527 9437 6544
rect 9863 6527 9869 6544
rect 9431 6521 9869 6527
rect 9429 6519 9871 6521
rect 9981 6544 10419 6550
rect 9981 6527 9987 6544
rect 10413 6527 10419 6544
rect 9981 6521 10419 6527
rect 9981 6519 10014 6521
rect 9286 6513 9350 6519
rect 9286 6486 9327 6513
rect 8873 6114 8879 6486
rect 9321 6114 9327 6486
rect 8873 6087 8914 6114
rect 8850 6081 8914 6087
rect 8186 6079 8219 6081
rect 7781 6073 8219 6079
rect 7781 6056 7787 6073
rect 8213 6056 8219 6073
rect 7781 6050 8219 6056
rect 8329 6079 8771 6081
rect 8331 6073 8769 6079
rect 8331 6056 8337 6073
rect 8763 6056 8769 6073
rect 8331 6050 8769 6056
rect 8881 6079 8914 6081
rect 9286 6087 9327 6114
rect 9344 6087 9350 6513
rect 9286 6081 9350 6087
rect 9400 6513 9900 6519
rect 9400 6087 9406 6513
rect 9423 6465 9877 6513
rect 9423 6135 9485 6465
rect 9815 6135 9877 6465
rect 9423 6087 9877 6135
rect 9894 6087 9900 6513
rect 9400 6081 9900 6087
rect 9950 6513 10014 6519
rect 9950 6087 9956 6513
rect 9973 6486 10014 6513
rect 10386 6519 10419 6521
rect 10531 6544 10969 6550
rect 10531 6527 10537 6544
rect 10963 6527 10969 6544
rect 10531 6521 10969 6527
rect 10529 6519 10971 6521
rect 11081 6544 11519 6550
rect 11081 6527 11087 6544
rect 11513 6527 11519 6544
rect 11081 6521 11519 6527
rect 11081 6519 11114 6521
rect 10386 6513 10450 6519
rect 10386 6486 10427 6513
rect 9973 6114 9979 6486
rect 10421 6114 10427 6486
rect 9973 6087 10014 6114
rect 9950 6081 10014 6087
rect 9286 6079 9319 6081
rect 8881 6073 9319 6079
rect 8881 6056 8887 6073
rect 9313 6056 9319 6073
rect 8881 6050 9319 6056
rect 9429 6079 9871 6081
rect 9431 6073 9869 6079
rect 9431 6056 9437 6073
rect 9863 6056 9869 6073
rect 9431 6050 9869 6056
rect 9981 6079 10014 6081
rect 10386 6087 10427 6114
rect 10444 6087 10450 6513
rect 10386 6081 10450 6087
rect 10500 6513 11000 6519
rect 10500 6087 10506 6513
rect 10523 6465 10977 6513
rect 10523 6135 10585 6465
rect 10915 6135 10977 6465
rect 10523 6087 10977 6135
rect 10994 6087 11000 6513
rect 10500 6081 11000 6087
rect 11050 6513 11114 6519
rect 11050 6087 11056 6513
rect 11073 6486 11114 6513
rect 11486 6519 11519 6521
rect 11631 6544 12069 6550
rect 11631 6527 11637 6544
rect 12063 6527 12069 6544
rect 11631 6521 12069 6527
rect 11629 6519 12071 6521
rect 12181 6544 12619 6550
rect 12181 6527 12187 6544
rect 12613 6527 12619 6544
rect 12181 6521 12619 6527
rect 12181 6519 12214 6521
rect 11486 6513 11550 6519
rect 11486 6486 11527 6513
rect 11073 6114 11079 6486
rect 11521 6114 11527 6486
rect 11073 6087 11114 6114
rect 11050 6081 11114 6087
rect 10386 6079 10419 6081
rect 9981 6073 10419 6079
rect 9981 6056 9987 6073
rect 10413 6056 10419 6073
rect 9981 6050 10419 6056
rect 10529 6079 10971 6081
rect 10531 6073 10969 6079
rect 10531 6056 10537 6073
rect 10963 6056 10969 6073
rect 10531 6050 10969 6056
rect 11081 6079 11114 6081
rect 11486 6087 11527 6114
rect 11544 6087 11550 6513
rect 11486 6081 11550 6087
rect 11600 6513 12100 6519
rect 11600 6087 11606 6513
rect 11623 6465 12077 6513
rect 11623 6135 11685 6465
rect 12015 6135 12077 6465
rect 11623 6087 12077 6135
rect 12094 6087 12100 6513
rect 11600 6081 12100 6087
rect 12150 6513 12214 6519
rect 12150 6087 12156 6513
rect 12173 6486 12214 6513
rect 12586 6519 12619 6521
rect 12731 6544 13169 6550
rect 12731 6527 12737 6544
rect 13163 6527 13169 6544
rect 12731 6521 13169 6527
rect 12729 6519 13171 6521
rect 13281 6544 13719 6550
rect 13281 6527 13287 6544
rect 13713 6527 13719 6544
rect 13281 6521 13719 6527
rect 13281 6519 13314 6521
rect 12586 6513 12650 6519
rect 12586 6486 12627 6513
rect 12173 6114 12179 6486
rect 12621 6114 12627 6486
rect 12173 6087 12214 6114
rect 12150 6081 12214 6087
rect 11486 6079 11519 6081
rect 11081 6073 11519 6079
rect 11081 6056 11087 6073
rect 11513 6056 11519 6073
rect 11081 6050 11519 6056
rect 11629 6079 12071 6081
rect 11631 6073 12069 6079
rect 11631 6056 11637 6073
rect 12063 6056 12069 6073
rect 11631 6050 12069 6056
rect 12181 6079 12214 6081
rect 12586 6087 12627 6114
rect 12644 6087 12650 6513
rect 12586 6081 12650 6087
rect 12700 6513 13200 6519
rect 12700 6087 12706 6513
rect 12723 6465 13177 6513
rect 12723 6135 12785 6465
rect 13115 6135 13177 6465
rect 12723 6087 13177 6135
rect 13194 6087 13200 6513
rect 12700 6081 13200 6087
rect 13250 6513 13314 6519
rect 13250 6087 13256 6513
rect 13273 6486 13314 6513
rect 13273 6114 13279 6486
rect 13273 6087 13314 6114
rect 13250 6081 13314 6087
rect 12586 6079 12619 6081
rect 12181 6073 12619 6079
rect 12181 6056 12187 6073
rect 12613 6056 12619 6073
rect 12181 6050 12619 6056
rect 12729 6079 13171 6081
rect 12731 6073 13169 6079
rect 12731 6056 12737 6073
rect 13163 6056 13169 6073
rect 12731 6050 13169 6056
rect 13281 6079 13314 6081
rect 13281 6073 13719 6079
rect 13281 6056 13287 6073
rect 13713 6056 13719 6073
rect 13281 6050 13719 6056
rect -469 5994 -31 6000
rect -469 5977 -463 5994
rect -37 5977 -31 5994
rect -469 5971 -31 5977
rect -64 5969 -31 5971
rect 81 5994 519 6000
rect 81 5977 87 5994
rect 513 5977 519 5994
rect 81 5971 519 5977
rect 79 5969 521 5971
rect 631 5994 1069 6000
rect 631 5977 637 5994
rect 1063 5977 1069 5994
rect 631 5971 1069 5977
rect 631 5969 664 5971
rect -64 5963 0 5969
rect -64 5936 -23 5963
rect -29 5564 -23 5936
rect -64 5537 -23 5564
rect -6 5537 0 5963
rect -64 5531 0 5537
rect 50 5963 550 5969
rect 50 5537 56 5963
rect 73 5915 527 5963
rect 73 5585 135 5915
rect 465 5585 527 5915
rect 73 5537 527 5585
rect 544 5537 550 5963
rect 50 5531 550 5537
rect 600 5963 664 5969
rect 600 5537 606 5963
rect 623 5936 664 5963
rect 1036 5969 1069 5971
rect 1181 5994 1619 6000
rect 1181 5977 1187 5994
rect 1613 5977 1619 5994
rect 1181 5971 1619 5977
rect 1179 5969 1621 5971
rect 1731 5994 2169 6000
rect 1731 5977 1737 5994
rect 2163 5977 2169 5994
rect 1731 5971 2169 5977
rect 1731 5969 1764 5971
rect 1036 5963 1100 5969
rect 1036 5936 1077 5963
rect 623 5564 629 5936
rect 1071 5564 1077 5936
rect 623 5537 664 5564
rect 600 5531 664 5537
rect -64 5529 -31 5531
rect -469 5523 -31 5529
rect -469 5506 -463 5523
rect -37 5506 -31 5523
rect -469 5500 -31 5506
rect 79 5529 521 5531
rect 81 5523 519 5529
rect 81 5506 87 5523
rect 513 5506 519 5523
rect 81 5500 519 5506
rect 631 5529 664 5531
rect 1036 5537 1077 5564
rect 1094 5537 1100 5963
rect 1036 5531 1100 5537
rect 1150 5963 1650 5969
rect 1150 5537 1156 5963
rect 1173 5915 1627 5963
rect 1173 5585 1235 5915
rect 1565 5585 1627 5915
rect 1173 5537 1627 5585
rect 1644 5537 1650 5963
rect 1150 5531 1650 5537
rect 1700 5963 1764 5969
rect 1700 5537 1706 5963
rect 1723 5936 1764 5963
rect 2136 5969 2169 5971
rect 2281 5994 2719 6000
rect 2281 5977 2287 5994
rect 2713 5977 2719 5994
rect 2281 5971 2719 5977
rect 2279 5969 2721 5971
rect 2831 5994 3269 6000
rect 2831 5977 2837 5994
rect 3263 5977 3269 5994
rect 2831 5971 3269 5977
rect 2831 5969 2864 5971
rect 2136 5963 2200 5969
rect 2136 5936 2177 5963
rect 1723 5564 1729 5936
rect 2171 5564 2177 5936
rect 1723 5537 1764 5564
rect 1700 5531 1764 5537
rect 1036 5529 1069 5531
rect 631 5523 1069 5529
rect 631 5506 637 5523
rect 1063 5506 1069 5523
rect 631 5500 1069 5506
rect 1179 5529 1621 5531
rect 1181 5523 1619 5529
rect 1181 5506 1187 5523
rect 1613 5506 1619 5523
rect 1181 5500 1619 5506
rect 1731 5529 1764 5531
rect 2136 5537 2177 5564
rect 2194 5537 2200 5963
rect 2136 5531 2200 5537
rect 2250 5963 2750 5969
rect 2250 5537 2256 5963
rect 2273 5915 2727 5963
rect 2273 5585 2335 5915
rect 2665 5585 2727 5915
rect 2273 5537 2727 5585
rect 2744 5537 2750 5963
rect 2250 5531 2750 5537
rect 2800 5963 2864 5969
rect 2800 5537 2806 5963
rect 2823 5936 2864 5963
rect 3236 5969 3269 5971
rect 3381 5994 3819 6000
rect 3381 5977 3387 5994
rect 3813 5977 3819 5994
rect 3381 5971 3819 5977
rect 3379 5969 3821 5971
rect 3931 5994 4369 6000
rect 3931 5977 3937 5994
rect 4363 5977 4369 5994
rect 3931 5971 4369 5977
rect 3931 5969 3964 5971
rect 3236 5963 3300 5969
rect 3236 5936 3277 5963
rect 2823 5564 2829 5936
rect 3271 5564 3277 5936
rect 2823 5537 2864 5564
rect 2800 5531 2864 5537
rect 2136 5529 2169 5531
rect 1731 5523 2169 5529
rect 1731 5506 1737 5523
rect 2163 5506 2169 5523
rect 1731 5500 2169 5506
rect 2279 5529 2721 5531
rect 2281 5523 2719 5529
rect 2281 5506 2287 5523
rect 2713 5506 2719 5523
rect 2281 5500 2719 5506
rect 2831 5529 2864 5531
rect 3236 5537 3277 5564
rect 3294 5537 3300 5963
rect 3236 5531 3300 5537
rect 3350 5963 3850 5969
rect 3350 5537 3356 5963
rect 3373 5915 3827 5963
rect 3373 5585 3435 5915
rect 3765 5585 3827 5915
rect 3373 5537 3827 5585
rect 3844 5537 3850 5963
rect 3350 5531 3850 5537
rect 3900 5963 3964 5969
rect 3900 5537 3906 5963
rect 3923 5936 3964 5963
rect 4336 5969 4369 5971
rect 4481 5994 4919 6000
rect 4481 5977 4487 5994
rect 4913 5977 4919 5994
rect 4481 5971 4919 5977
rect 4479 5969 4921 5971
rect 5031 5994 5469 6000
rect 5031 5977 5037 5994
rect 5463 5977 5469 5994
rect 5031 5971 5469 5977
rect 5031 5969 5064 5971
rect 4336 5963 4400 5969
rect 4336 5936 4377 5963
rect 3923 5564 3929 5936
rect 4371 5564 4377 5936
rect 3923 5537 3964 5564
rect 3900 5531 3964 5537
rect 3236 5529 3269 5531
rect 2831 5523 3269 5529
rect 2831 5506 2837 5523
rect 3263 5506 3269 5523
rect 2831 5500 3269 5506
rect 3379 5529 3821 5531
rect 3381 5523 3819 5529
rect 3381 5506 3387 5523
rect 3813 5506 3819 5523
rect 3381 5500 3819 5506
rect 3931 5529 3964 5531
rect 4336 5537 4377 5564
rect 4394 5537 4400 5963
rect 4336 5531 4400 5537
rect 4450 5963 4950 5969
rect 4450 5537 4456 5963
rect 4473 5915 4927 5963
rect 4473 5585 4535 5915
rect 4865 5585 4927 5915
rect 4473 5537 4927 5585
rect 4944 5537 4950 5963
rect 4450 5531 4950 5537
rect 5000 5963 5064 5969
rect 5000 5537 5006 5963
rect 5023 5936 5064 5963
rect 5436 5969 5469 5971
rect 5581 5994 6019 6000
rect 5581 5977 5587 5994
rect 6013 5977 6019 5994
rect 5581 5971 6019 5977
rect 5579 5969 6021 5971
rect 6131 5994 6569 6000
rect 6131 5977 6137 5994
rect 6563 5977 6569 5994
rect 6131 5971 6569 5977
rect 6131 5969 6164 5971
rect 5436 5963 5500 5969
rect 5436 5936 5477 5963
rect 5023 5564 5029 5936
rect 5471 5564 5477 5936
rect 5023 5537 5064 5564
rect 5000 5531 5064 5537
rect 4336 5529 4369 5531
rect 3931 5523 4369 5529
rect 3931 5506 3937 5523
rect 4363 5506 4369 5523
rect 3931 5500 4369 5506
rect 4479 5529 4921 5531
rect 4481 5523 4919 5529
rect 4481 5506 4487 5523
rect 4913 5506 4919 5523
rect 4481 5500 4919 5506
rect 5031 5529 5064 5531
rect 5436 5537 5477 5564
rect 5494 5537 5500 5963
rect 5436 5531 5500 5537
rect 5550 5963 6050 5969
rect 5550 5537 5556 5963
rect 5573 5915 6027 5963
rect 5573 5585 5635 5915
rect 5965 5585 6027 5915
rect 5573 5537 6027 5585
rect 6044 5537 6050 5963
rect 5550 5531 6050 5537
rect 6100 5963 6164 5969
rect 6100 5537 6106 5963
rect 6123 5936 6164 5963
rect 6536 5969 6569 5971
rect 6681 5994 7119 6000
rect 6681 5977 6687 5994
rect 7113 5977 7119 5994
rect 6681 5971 7119 5977
rect 6679 5969 7121 5971
rect 7231 5994 7669 6000
rect 7231 5977 7237 5994
rect 7663 5977 7669 5994
rect 7231 5971 7669 5977
rect 7231 5969 7264 5971
rect 6536 5963 6600 5969
rect 6536 5936 6577 5963
rect 6123 5564 6129 5936
rect 6571 5564 6577 5936
rect 6123 5537 6164 5564
rect 6100 5531 6164 5537
rect 5436 5529 5469 5531
rect 5031 5523 5469 5529
rect 5031 5506 5037 5523
rect 5463 5506 5469 5523
rect 5031 5500 5469 5506
rect 5579 5529 6021 5531
rect 5581 5523 6019 5529
rect 5581 5506 5587 5523
rect 6013 5506 6019 5523
rect 5581 5500 6019 5506
rect 6131 5529 6164 5531
rect 6536 5537 6577 5564
rect 6594 5537 6600 5963
rect 6536 5531 6600 5537
rect 6650 5963 7150 5969
rect 6650 5537 6656 5963
rect 6673 5915 7127 5963
rect 6673 5585 6735 5915
rect 7065 5585 7127 5915
rect 6673 5537 7127 5585
rect 7144 5537 7150 5963
rect 6650 5531 7150 5537
rect 7200 5963 7264 5969
rect 7200 5537 7206 5963
rect 7223 5936 7264 5963
rect 7636 5969 7669 5971
rect 7781 5994 8219 6000
rect 7781 5977 7787 5994
rect 8213 5977 8219 5994
rect 7781 5971 8219 5977
rect 7779 5969 8221 5971
rect 8331 5994 8769 6000
rect 8331 5977 8337 5994
rect 8763 5977 8769 5994
rect 8331 5971 8769 5977
rect 8331 5969 8364 5971
rect 7636 5963 7700 5969
rect 7636 5936 7677 5963
rect 7223 5564 7229 5936
rect 7671 5564 7677 5936
rect 7223 5537 7264 5564
rect 7200 5531 7264 5537
rect 6536 5529 6569 5531
rect 6131 5523 6569 5529
rect 6131 5506 6137 5523
rect 6563 5506 6569 5523
rect 6131 5500 6569 5506
rect 6679 5529 7121 5531
rect 6681 5523 7119 5529
rect 6681 5506 6687 5523
rect 7113 5506 7119 5523
rect 6681 5500 7119 5506
rect 7231 5529 7264 5531
rect 7636 5537 7677 5564
rect 7694 5537 7700 5963
rect 7636 5531 7700 5537
rect 7750 5963 8250 5969
rect 7750 5537 7756 5963
rect 7773 5915 8227 5963
rect 7773 5585 7835 5915
rect 8165 5585 8227 5915
rect 7773 5537 8227 5585
rect 8244 5537 8250 5963
rect 7750 5531 8250 5537
rect 8300 5963 8364 5969
rect 8300 5537 8306 5963
rect 8323 5936 8364 5963
rect 8736 5969 8769 5971
rect 8881 5994 9319 6000
rect 8881 5977 8887 5994
rect 9313 5977 9319 5994
rect 8881 5971 9319 5977
rect 8879 5969 9321 5971
rect 9431 5994 9869 6000
rect 9431 5977 9437 5994
rect 9863 5977 9869 5994
rect 9431 5971 9869 5977
rect 9431 5969 9464 5971
rect 8736 5963 8800 5969
rect 8736 5936 8777 5963
rect 8323 5564 8329 5936
rect 8771 5564 8777 5936
rect 8323 5537 8364 5564
rect 8300 5531 8364 5537
rect 7636 5529 7669 5531
rect 7231 5523 7669 5529
rect 7231 5506 7237 5523
rect 7663 5506 7669 5523
rect 7231 5500 7669 5506
rect 7779 5529 8221 5531
rect 7781 5523 8219 5529
rect 7781 5506 7787 5523
rect 8213 5506 8219 5523
rect 7781 5500 8219 5506
rect 8331 5529 8364 5531
rect 8736 5537 8777 5564
rect 8794 5537 8800 5963
rect 8736 5531 8800 5537
rect 8850 5963 9350 5969
rect 8850 5537 8856 5963
rect 8873 5915 9327 5963
rect 8873 5585 8935 5915
rect 9265 5585 9327 5915
rect 8873 5537 9327 5585
rect 9344 5537 9350 5963
rect 8850 5531 9350 5537
rect 9400 5963 9464 5969
rect 9400 5537 9406 5963
rect 9423 5936 9464 5963
rect 9836 5969 9869 5971
rect 9981 5994 10419 6000
rect 9981 5977 9987 5994
rect 10413 5977 10419 5994
rect 9981 5971 10419 5977
rect 9979 5969 10421 5971
rect 10531 5994 10969 6000
rect 10531 5977 10537 5994
rect 10963 5977 10969 5994
rect 10531 5971 10969 5977
rect 10531 5969 10564 5971
rect 9836 5963 9900 5969
rect 9836 5936 9877 5963
rect 9423 5564 9429 5936
rect 9871 5564 9877 5936
rect 9423 5537 9464 5564
rect 9400 5531 9464 5537
rect 8736 5529 8769 5531
rect 8331 5523 8769 5529
rect 8331 5506 8337 5523
rect 8763 5506 8769 5523
rect 8331 5500 8769 5506
rect 8879 5529 9321 5531
rect 8881 5523 9319 5529
rect 8881 5506 8887 5523
rect 9313 5506 9319 5523
rect 8881 5500 9319 5506
rect 9431 5529 9464 5531
rect 9836 5537 9877 5564
rect 9894 5537 9900 5963
rect 9836 5531 9900 5537
rect 9950 5963 10450 5969
rect 9950 5537 9956 5963
rect 9973 5915 10427 5963
rect 9973 5585 10035 5915
rect 10365 5585 10427 5915
rect 9973 5537 10427 5585
rect 10444 5537 10450 5963
rect 9950 5531 10450 5537
rect 10500 5963 10564 5969
rect 10500 5537 10506 5963
rect 10523 5936 10564 5963
rect 10936 5969 10969 5971
rect 11081 5994 11519 6000
rect 11081 5977 11087 5994
rect 11513 5977 11519 5994
rect 11081 5971 11519 5977
rect 11079 5969 11521 5971
rect 11631 5994 12069 6000
rect 11631 5977 11637 5994
rect 12063 5977 12069 5994
rect 11631 5971 12069 5977
rect 11631 5969 11664 5971
rect 10936 5963 11000 5969
rect 10936 5936 10977 5963
rect 10523 5564 10529 5936
rect 10971 5564 10977 5936
rect 10523 5537 10564 5564
rect 10500 5531 10564 5537
rect 9836 5529 9869 5531
rect 9431 5523 9869 5529
rect 9431 5506 9437 5523
rect 9863 5506 9869 5523
rect 9431 5500 9869 5506
rect 9979 5529 10421 5531
rect 9981 5523 10419 5529
rect 9981 5506 9987 5523
rect 10413 5506 10419 5523
rect 9981 5500 10419 5506
rect 10531 5529 10564 5531
rect 10936 5537 10977 5564
rect 10994 5537 11000 5963
rect 10936 5531 11000 5537
rect 11050 5963 11550 5969
rect 11050 5537 11056 5963
rect 11073 5915 11527 5963
rect 11073 5585 11135 5915
rect 11465 5585 11527 5915
rect 11073 5537 11527 5585
rect 11544 5537 11550 5963
rect 11050 5531 11550 5537
rect 11600 5963 11664 5969
rect 11600 5537 11606 5963
rect 11623 5936 11664 5963
rect 12036 5969 12069 5971
rect 12181 5994 12619 6000
rect 12181 5977 12187 5994
rect 12613 5977 12619 5994
rect 12181 5971 12619 5977
rect 12179 5969 12621 5971
rect 12731 5994 13169 6000
rect 12731 5977 12737 5994
rect 13163 5977 13169 5994
rect 12731 5971 13169 5977
rect 12731 5969 12764 5971
rect 12036 5963 12100 5969
rect 12036 5936 12077 5963
rect 11623 5564 11629 5936
rect 12071 5564 12077 5936
rect 11623 5537 11664 5564
rect 11600 5531 11664 5537
rect 10936 5529 10969 5531
rect 10531 5523 10969 5529
rect 10531 5506 10537 5523
rect 10963 5506 10969 5523
rect 10531 5500 10969 5506
rect 11079 5529 11521 5531
rect 11081 5523 11519 5529
rect 11081 5506 11087 5523
rect 11513 5506 11519 5523
rect 11081 5500 11519 5506
rect 11631 5529 11664 5531
rect 12036 5537 12077 5564
rect 12094 5537 12100 5963
rect 12036 5531 12100 5537
rect 12150 5963 12650 5969
rect 12150 5537 12156 5963
rect 12173 5915 12627 5963
rect 12173 5585 12235 5915
rect 12565 5585 12627 5915
rect 12173 5537 12627 5585
rect 12644 5537 12650 5963
rect 12150 5531 12650 5537
rect 12700 5963 12764 5969
rect 12700 5537 12706 5963
rect 12723 5936 12764 5963
rect 13136 5969 13169 5971
rect 13281 5994 13719 6000
rect 13281 5977 13287 5994
rect 13713 5977 13719 5994
rect 13281 5971 13719 5977
rect 13279 5969 13721 5971
rect 13136 5963 13200 5969
rect 13136 5936 13177 5963
rect 12723 5564 12729 5936
rect 13171 5564 13177 5936
rect 12723 5537 12764 5564
rect 12700 5531 12764 5537
rect 12036 5529 12069 5531
rect 11631 5523 12069 5529
rect 11631 5506 11637 5523
rect 12063 5506 12069 5523
rect 11631 5500 12069 5506
rect 12179 5529 12621 5531
rect 12181 5523 12619 5529
rect 12181 5506 12187 5523
rect 12613 5506 12619 5523
rect 12181 5500 12619 5506
rect 12731 5529 12764 5531
rect 13136 5537 13177 5564
rect 13194 5537 13200 5963
rect 13136 5531 13200 5537
rect 13250 5963 13721 5969
rect 13250 5537 13256 5963
rect 13273 5915 13721 5963
rect 13273 5585 13335 5915
rect 13665 5585 13721 5915
rect 13273 5537 13721 5585
rect 13250 5531 13721 5537
rect 13136 5529 13169 5531
rect 12731 5523 13169 5529
rect 12731 5506 12737 5523
rect 13163 5506 13169 5523
rect 12731 5500 13169 5506
rect 13279 5529 13721 5531
rect 13281 5523 13719 5529
rect 13281 5506 13287 5523
rect 13713 5506 13719 5523
rect 13281 5500 13719 5506
rect -469 5444 -31 5450
rect -469 5427 -463 5444
rect -37 5427 -31 5444
rect -469 5421 -31 5427
rect -471 5419 -29 5421
rect 81 5444 519 5450
rect 81 5427 87 5444
rect 513 5427 519 5444
rect 81 5421 519 5427
rect 81 5419 114 5421
rect -471 5413 0 5419
rect -471 5365 -23 5413
rect -471 5035 -415 5365
rect -85 5035 -23 5365
rect -471 4987 -23 5035
rect -6 4987 0 5413
rect -471 4981 0 4987
rect 50 5413 114 5419
rect 50 4987 56 5413
rect 73 5386 114 5413
rect 486 5419 519 5421
rect 631 5444 1069 5450
rect 631 5427 637 5444
rect 1063 5427 1069 5444
rect 631 5421 1069 5427
rect 629 5419 1071 5421
rect 1181 5444 1619 5450
rect 1181 5427 1187 5444
rect 1613 5427 1619 5444
rect 1181 5421 1619 5427
rect 1181 5419 1214 5421
rect 486 5413 550 5419
rect 486 5386 527 5413
rect 73 5014 79 5386
rect 521 5014 527 5386
rect 73 4987 114 5014
rect 50 4981 114 4987
rect -471 4979 -29 4981
rect -469 4973 -31 4979
rect -469 4956 -463 4973
rect -37 4956 -31 4973
rect -469 4950 -31 4956
rect 81 4979 114 4981
rect 486 4987 527 5014
rect 544 4987 550 5413
rect 486 4981 550 4987
rect 600 5413 1100 5419
rect 600 4987 606 5413
rect 623 5365 1077 5413
rect 623 5035 685 5365
rect 1015 5035 1077 5365
rect 623 4987 1077 5035
rect 1094 4987 1100 5413
rect 600 4981 1100 4987
rect 1150 5413 1214 5419
rect 1150 4987 1156 5413
rect 1173 5386 1214 5413
rect 1586 5419 1619 5421
rect 1731 5444 2169 5450
rect 1731 5427 1737 5444
rect 2163 5427 2169 5444
rect 1731 5421 2169 5427
rect 1729 5419 2171 5421
rect 2281 5444 2719 5450
rect 2281 5427 2287 5444
rect 2713 5427 2719 5444
rect 2281 5421 2719 5427
rect 2281 5419 2314 5421
rect 1586 5413 1650 5419
rect 1586 5386 1627 5413
rect 1173 5014 1179 5386
rect 1621 5014 1627 5386
rect 1173 4987 1214 5014
rect 1150 4981 1214 4987
rect 486 4979 519 4981
rect 81 4973 519 4979
rect 81 4956 87 4973
rect 513 4956 519 4973
rect 81 4950 519 4956
rect 629 4979 1071 4981
rect 631 4973 1069 4979
rect 631 4956 637 4973
rect 1063 4956 1069 4973
rect 631 4950 1069 4956
rect 1181 4979 1214 4981
rect 1586 4987 1627 5014
rect 1644 4987 1650 5413
rect 1586 4981 1650 4987
rect 1700 5413 2200 5419
rect 1700 4987 1706 5413
rect 1723 5365 2177 5413
rect 1723 5035 1785 5365
rect 2115 5035 2177 5365
rect 1723 4987 2177 5035
rect 2194 4987 2200 5413
rect 1700 4981 2200 4987
rect 2250 5413 2314 5419
rect 2250 4987 2256 5413
rect 2273 5386 2314 5413
rect 2686 5419 2719 5421
rect 2831 5444 3269 5450
rect 2831 5427 2837 5444
rect 3263 5427 3269 5444
rect 2831 5421 3269 5427
rect 2829 5419 3271 5421
rect 3381 5444 3819 5450
rect 3381 5427 3387 5444
rect 3813 5427 3819 5444
rect 3381 5421 3819 5427
rect 3381 5419 3414 5421
rect 2686 5413 2750 5419
rect 2686 5386 2727 5413
rect 2273 5014 2279 5386
rect 2721 5014 2727 5386
rect 2273 4987 2314 5014
rect 2250 4981 2314 4987
rect 1586 4979 1619 4981
rect 1181 4973 1619 4979
rect 1181 4956 1187 4973
rect 1613 4956 1619 4973
rect 1181 4950 1619 4956
rect 1729 4979 2171 4981
rect 1731 4973 2169 4979
rect 1731 4956 1737 4973
rect 2163 4956 2169 4973
rect 1731 4950 2169 4956
rect 2281 4979 2314 4981
rect 2686 4987 2727 5014
rect 2744 4987 2750 5413
rect 2686 4981 2750 4987
rect 2800 5413 3300 5419
rect 2800 4987 2806 5413
rect 2823 5365 3277 5413
rect 2823 5035 2885 5365
rect 3215 5035 3277 5365
rect 2823 4987 3277 5035
rect 3294 4987 3300 5413
rect 2800 4981 3300 4987
rect 3350 5413 3414 5419
rect 3350 4987 3356 5413
rect 3373 5386 3414 5413
rect 3786 5419 3819 5421
rect 3931 5444 4369 5450
rect 3931 5427 3937 5444
rect 4363 5427 4369 5444
rect 3931 5421 4369 5427
rect 3929 5419 4371 5421
rect 4481 5444 4919 5450
rect 4481 5427 4487 5444
rect 4913 5427 4919 5444
rect 4481 5421 4919 5427
rect 4481 5419 4514 5421
rect 3786 5413 3850 5419
rect 3786 5386 3827 5413
rect 3373 5014 3379 5386
rect 3821 5014 3827 5386
rect 3373 4987 3414 5014
rect 3350 4981 3414 4987
rect 2686 4979 2719 4981
rect 2281 4973 2719 4979
rect 2281 4956 2287 4973
rect 2713 4956 2719 4973
rect 2281 4950 2719 4956
rect 2829 4979 3271 4981
rect 2831 4973 3269 4979
rect 2831 4956 2837 4973
rect 3263 4956 3269 4973
rect 2831 4950 3269 4956
rect 3381 4979 3414 4981
rect 3786 4987 3827 5014
rect 3844 4987 3850 5413
rect 3786 4981 3850 4987
rect 3900 5413 4400 5419
rect 3900 4987 3906 5413
rect 3923 5365 4377 5413
rect 3923 5035 3985 5365
rect 4315 5035 4377 5365
rect 3923 4987 4377 5035
rect 4394 4987 4400 5413
rect 3900 4981 4400 4987
rect 4450 5413 4514 5419
rect 4450 4987 4456 5413
rect 4473 5386 4514 5413
rect 4886 5419 4919 5421
rect 5031 5444 5469 5450
rect 5031 5427 5037 5444
rect 5463 5427 5469 5444
rect 5031 5421 5469 5427
rect 5029 5419 5471 5421
rect 5581 5444 6019 5450
rect 5581 5427 5587 5444
rect 6013 5427 6019 5444
rect 5581 5421 6019 5427
rect 5581 5419 5614 5421
rect 4886 5413 4950 5419
rect 4886 5386 4927 5413
rect 4473 5014 4479 5386
rect 4921 5014 4927 5386
rect 4473 4987 4514 5014
rect 4450 4981 4514 4987
rect 3786 4979 3819 4981
rect 3381 4973 3819 4979
rect 3381 4956 3387 4973
rect 3813 4956 3819 4973
rect 3381 4950 3819 4956
rect 3929 4979 4371 4981
rect 3931 4973 4369 4979
rect 3931 4956 3937 4973
rect 4363 4956 4369 4973
rect 3931 4950 4369 4956
rect 4481 4979 4514 4981
rect 4886 4987 4927 5014
rect 4944 4987 4950 5413
rect 4886 4981 4950 4987
rect 5000 5413 5500 5419
rect 5000 4987 5006 5413
rect 5023 5365 5477 5413
rect 5023 5035 5085 5365
rect 5415 5035 5477 5365
rect 5023 4987 5477 5035
rect 5494 4987 5500 5413
rect 5000 4981 5500 4987
rect 5550 5413 5614 5419
rect 5550 4987 5556 5413
rect 5573 5386 5614 5413
rect 5986 5419 6019 5421
rect 6131 5444 6569 5450
rect 6131 5427 6137 5444
rect 6563 5427 6569 5444
rect 6131 5421 6569 5427
rect 6129 5419 6571 5421
rect 6681 5444 7119 5450
rect 6681 5427 6687 5444
rect 7113 5427 7119 5444
rect 6681 5421 7119 5427
rect 6681 5419 6714 5421
rect 5986 5413 6050 5419
rect 5986 5386 6027 5413
rect 5573 5014 5579 5386
rect 6021 5014 6027 5386
rect 5573 4987 5614 5014
rect 5550 4981 5614 4987
rect 4886 4979 4919 4981
rect 4481 4973 4919 4979
rect 4481 4956 4487 4973
rect 4913 4956 4919 4973
rect 4481 4950 4919 4956
rect 5029 4979 5471 4981
rect 5031 4973 5469 4979
rect 5031 4956 5037 4973
rect 5463 4956 5469 4973
rect 5031 4950 5469 4956
rect 5581 4979 5614 4981
rect 5986 4987 6027 5014
rect 6044 4987 6050 5413
rect 5986 4981 6050 4987
rect 6100 5413 6600 5419
rect 6100 4987 6106 5413
rect 6123 5365 6577 5413
rect 6123 5035 6185 5365
rect 6515 5035 6577 5365
rect 6123 4987 6577 5035
rect 6594 4987 6600 5413
rect 6100 4981 6600 4987
rect 6650 5413 6714 5419
rect 6650 4987 6656 5413
rect 6673 5386 6714 5413
rect 7086 5419 7119 5421
rect 7231 5444 7669 5450
rect 7231 5427 7237 5444
rect 7663 5427 7669 5444
rect 7231 5421 7669 5427
rect 7229 5419 7671 5421
rect 7781 5444 8219 5450
rect 7781 5427 7787 5444
rect 8213 5427 8219 5444
rect 7781 5421 8219 5427
rect 7781 5419 7814 5421
rect 7086 5413 7150 5419
rect 7086 5386 7127 5413
rect 6673 5014 6679 5386
rect 7121 5014 7127 5386
rect 6673 4987 6714 5014
rect 6650 4981 6714 4987
rect 5986 4979 6019 4981
rect 5581 4973 6019 4979
rect 5581 4956 5587 4973
rect 6013 4956 6019 4973
rect 5581 4950 6019 4956
rect 6129 4979 6571 4981
rect 6131 4973 6569 4979
rect 6131 4956 6137 4973
rect 6563 4956 6569 4973
rect 6131 4950 6569 4956
rect 6681 4979 6714 4981
rect 7086 4987 7127 5014
rect 7144 4987 7150 5413
rect 7086 4981 7150 4987
rect 7200 5413 7700 5419
rect 7200 4987 7206 5413
rect 7223 5365 7677 5413
rect 7223 5035 7285 5365
rect 7615 5035 7677 5365
rect 7223 4987 7677 5035
rect 7694 4987 7700 5413
rect 7200 4981 7700 4987
rect 7750 5413 7814 5419
rect 7750 4987 7756 5413
rect 7773 5386 7814 5413
rect 8186 5419 8219 5421
rect 8331 5444 8769 5450
rect 8331 5427 8337 5444
rect 8763 5427 8769 5444
rect 8331 5421 8769 5427
rect 8329 5419 8771 5421
rect 8881 5444 9319 5450
rect 8881 5427 8887 5444
rect 9313 5427 9319 5444
rect 8881 5421 9319 5427
rect 8881 5419 8914 5421
rect 8186 5413 8250 5419
rect 8186 5386 8227 5413
rect 7773 5014 7779 5386
rect 8221 5014 8227 5386
rect 7773 4987 7814 5014
rect 7750 4981 7814 4987
rect 7086 4979 7119 4981
rect 6681 4973 7119 4979
rect 6681 4956 6687 4973
rect 7113 4956 7119 4973
rect 6681 4950 7119 4956
rect 7229 4979 7671 4981
rect 7231 4973 7669 4979
rect 7231 4956 7237 4973
rect 7663 4956 7669 4973
rect 7231 4950 7669 4956
rect 7781 4979 7814 4981
rect 8186 4987 8227 5014
rect 8244 4987 8250 5413
rect 8186 4981 8250 4987
rect 8300 5413 8800 5419
rect 8300 4987 8306 5413
rect 8323 5365 8777 5413
rect 8323 5035 8385 5365
rect 8715 5035 8777 5365
rect 8323 4987 8777 5035
rect 8794 4987 8800 5413
rect 8300 4981 8800 4987
rect 8850 5413 8914 5419
rect 8850 4987 8856 5413
rect 8873 5386 8914 5413
rect 9286 5419 9319 5421
rect 9431 5444 9869 5450
rect 9431 5427 9437 5444
rect 9863 5427 9869 5444
rect 9431 5421 9869 5427
rect 9429 5419 9871 5421
rect 9981 5444 10419 5450
rect 9981 5427 9987 5444
rect 10413 5427 10419 5444
rect 9981 5421 10419 5427
rect 9981 5419 10014 5421
rect 9286 5413 9350 5419
rect 9286 5386 9327 5413
rect 8873 5014 8879 5386
rect 9321 5014 9327 5386
rect 8873 4987 8914 5014
rect 8850 4981 8914 4987
rect 8186 4979 8219 4981
rect 7781 4973 8219 4979
rect 7781 4956 7787 4973
rect 8213 4956 8219 4973
rect 7781 4950 8219 4956
rect 8329 4979 8771 4981
rect 8331 4973 8769 4979
rect 8331 4956 8337 4973
rect 8763 4956 8769 4973
rect 8331 4950 8769 4956
rect 8881 4979 8914 4981
rect 9286 4987 9327 5014
rect 9344 4987 9350 5413
rect 9286 4981 9350 4987
rect 9400 5413 9900 5419
rect 9400 4987 9406 5413
rect 9423 5365 9877 5413
rect 9423 5035 9485 5365
rect 9815 5035 9877 5365
rect 9423 4987 9877 5035
rect 9894 4987 9900 5413
rect 9400 4981 9900 4987
rect 9950 5413 10014 5419
rect 9950 4987 9956 5413
rect 9973 5386 10014 5413
rect 10386 5419 10419 5421
rect 10531 5444 10969 5450
rect 10531 5427 10537 5444
rect 10963 5427 10969 5444
rect 10531 5421 10969 5427
rect 10529 5419 10971 5421
rect 11081 5444 11519 5450
rect 11081 5427 11087 5444
rect 11513 5427 11519 5444
rect 11081 5421 11519 5427
rect 11081 5419 11114 5421
rect 10386 5413 10450 5419
rect 10386 5386 10427 5413
rect 9973 5014 9979 5386
rect 10421 5014 10427 5386
rect 9973 4987 10014 5014
rect 9950 4981 10014 4987
rect 9286 4979 9319 4981
rect 8881 4973 9319 4979
rect 8881 4956 8887 4973
rect 9313 4956 9319 4973
rect 8881 4950 9319 4956
rect 9429 4979 9871 4981
rect 9431 4973 9869 4979
rect 9431 4956 9437 4973
rect 9863 4956 9869 4973
rect 9431 4950 9869 4956
rect 9981 4979 10014 4981
rect 10386 4987 10427 5014
rect 10444 4987 10450 5413
rect 10386 4981 10450 4987
rect 10500 5413 11000 5419
rect 10500 4987 10506 5413
rect 10523 5365 10977 5413
rect 10523 5035 10585 5365
rect 10915 5035 10977 5365
rect 10523 4987 10977 5035
rect 10994 4987 11000 5413
rect 10500 4981 11000 4987
rect 11050 5413 11114 5419
rect 11050 4987 11056 5413
rect 11073 5386 11114 5413
rect 11486 5419 11519 5421
rect 11631 5444 12069 5450
rect 11631 5427 11637 5444
rect 12063 5427 12069 5444
rect 11631 5421 12069 5427
rect 11629 5419 12071 5421
rect 12181 5444 12619 5450
rect 12181 5427 12187 5444
rect 12613 5427 12619 5444
rect 12181 5421 12619 5427
rect 12181 5419 12214 5421
rect 11486 5413 11550 5419
rect 11486 5386 11527 5413
rect 11073 5014 11079 5386
rect 11521 5014 11527 5386
rect 11073 4987 11114 5014
rect 11050 4981 11114 4987
rect 10386 4979 10419 4981
rect 9981 4973 10419 4979
rect 9981 4956 9987 4973
rect 10413 4956 10419 4973
rect 9981 4950 10419 4956
rect 10529 4979 10971 4981
rect 10531 4973 10969 4979
rect 10531 4956 10537 4973
rect 10963 4956 10969 4973
rect 10531 4950 10969 4956
rect 11081 4979 11114 4981
rect 11486 4987 11527 5014
rect 11544 4987 11550 5413
rect 11486 4981 11550 4987
rect 11600 5413 12100 5419
rect 11600 4987 11606 5413
rect 11623 5365 12077 5413
rect 11623 5035 11685 5365
rect 12015 5035 12077 5365
rect 11623 4987 12077 5035
rect 12094 4987 12100 5413
rect 11600 4981 12100 4987
rect 12150 5413 12214 5419
rect 12150 4987 12156 5413
rect 12173 5386 12214 5413
rect 12586 5419 12619 5421
rect 12731 5444 13169 5450
rect 12731 5427 12737 5444
rect 13163 5427 13169 5444
rect 12731 5421 13169 5427
rect 12729 5419 13171 5421
rect 13281 5444 13719 5450
rect 13281 5427 13287 5444
rect 13713 5427 13719 5444
rect 13281 5421 13719 5427
rect 13281 5419 13314 5421
rect 12586 5413 12650 5419
rect 12586 5386 12627 5413
rect 12173 5014 12179 5386
rect 12621 5014 12627 5386
rect 12173 4987 12214 5014
rect 12150 4981 12214 4987
rect 11486 4979 11519 4981
rect 11081 4973 11519 4979
rect 11081 4956 11087 4973
rect 11513 4956 11519 4973
rect 11081 4950 11519 4956
rect 11629 4979 12071 4981
rect 11631 4973 12069 4979
rect 11631 4956 11637 4973
rect 12063 4956 12069 4973
rect 11631 4950 12069 4956
rect 12181 4979 12214 4981
rect 12586 4987 12627 5014
rect 12644 4987 12650 5413
rect 12586 4981 12650 4987
rect 12700 5413 13200 5419
rect 12700 4987 12706 5413
rect 12723 5365 13177 5413
rect 12723 5035 12785 5365
rect 13115 5035 13177 5365
rect 12723 4987 13177 5035
rect 13194 4987 13200 5413
rect 12700 4981 13200 4987
rect 13250 5413 13314 5419
rect 13250 4987 13256 5413
rect 13273 5386 13314 5413
rect 13273 5014 13279 5386
rect 13273 4987 13314 5014
rect 13250 4981 13314 4987
rect 12586 4979 12619 4981
rect 12181 4973 12619 4979
rect 12181 4956 12187 4973
rect 12613 4956 12619 4973
rect 12181 4950 12619 4956
rect 12729 4979 13171 4981
rect 12731 4973 13169 4979
rect 12731 4956 12737 4973
rect 13163 4956 13169 4973
rect 12731 4950 13169 4956
rect 13281 4979 13314 4981
rect 13281 4973 13719 4979
rect 13281 4956 13287 4973
rect 13713 4956 13719 4973
rect 13281 4950 13719 4956
rect -469 4894 -31 4900
rect -469 4877 -463 4894
rect -37 4877 -31 4894
rect -469 4871 -31 4877
rect -64 4869 -31 4871
rect 81 4894 519 4900
rect 81 4877 87 4894
rect 513 4877 519 4894
rect 81 4871 519 4877
rect 79 4869 521 4871
rect 631 4894 1069 4900
rect 631 4877 637 4894
rect 1063 4877 1069 4894
rect 631 4871 1069 4877
rect 631 4869 664 4871
rect -64 4863 0 4869
rect -64 4836 -23 4863
rect -29 4464 -23 4836
rect -64 4437 -23 4464
rect -6 4437 0 4863
rect -64 4431 0 4437
rect 50 4863 550 4869
rect 50 4437 56 4863
rect 73 4815 527 4863
rect 73 4485 135 4815
rect 465 4485 527 4815
rect 73 4437 527 4485
rect 544 4437 550 4863
rect 50 4431 550 4437
rect 600 4863 664 4869
rect 600 4437 606 4863
rect 623 4836 664 4863
rect 1036 4869 1069 4871
rect 1181 4894 1619 4900
rect 1181 4877 1187 4894
rect 1613 4877 1619 4894
rect 1181 4871 1619 4877
rect 1179 4869 1621 4871
rect 1731 4894 2169 4900
rect 1731 4877 1737 4894
rect 2163 4877 2169 4894
rect 1731 4871 2169 4877
rect 1731 4869 1764 4871
rect 1036 4863 1100 4869
rect 1036 4836 1077 4863
rect 623 4464 629 4836
rect 1071 4464 1077 4836
rect 623 4437 664 4464
rect 600 4431 664 4437
rect -64 4429 -31 4431
rect -469 4423 -31 4429
rect -469 4406 -463 4423
rect -37 4406 -31 4423
rect -469 4400 -31 4406
rect 79 4429 521 4431
rect 81 4423 519 4429
rect 81 4406 87 4423
rect 513 4406 519 4423
rect 81 4400 519 4406
rect 631 4429 664 4431
rect 1036 4437 1077 4464
rect 1094 4437 1100 4863
rect 1036 4431 1100 4437
rect 1150 4863 1650 4869
rect 1150 4437 1156 4863
rect 1173 4815 1627 4863
rect 1173 4485 1235 4815
rect 1565 4485 1627 4815
rect 1173 4437 1627 4485
rect 1644 4437 1650 4863
rect 1150 4431 1650 4437
rect 1700 4863 1764 4869
rect 1700 4437 1706 4863
rect 1723 4836 1764 4863
rect 2136 4869 2169 4871
rect 2281 4894 2719 4900
rect 2281 4877 2287 4894
rect 2713 4877 2719 4894
rect 2281 4871 2719 4877
rect 2279 4869 2721 4871
rect 2831 4894 3269 4900
rect 2831 4877 2837 4894
rect 3263 4877 3269 4894
rect 2831 4871 3269 4877
rect 2831 4869 2864 4871
rect 2136 4863 2200 4869
rect 2136 4836 2177 4863
rect 1723 4464 1729 4836
rect 2171 4464 2177 4836
rect 1723 4437 1764 4464
rect 1700 4431 1764 4437
rect 1036 4429 1069 4431
rect 631 4423 1069 4429
rect 631 4406 637 4423
rect 1063 4406 1069 4423
rect 631 4400 1069 4406
rect 1179 4429 1621 4431
rect 1181 4423 1619 4429
rect 1181 4406 1187 4423
rect 1613 4406 1619 4423
rect 1181 4400 1619 4406
rect 1731 4429 1764 4431
rect 2136 4437 2177 4464
rect 2194 4437 2200 4863
rect 2136 4431 2200 4437
rect 2250 4863 2750 4869
rect 2250 4437 2256 4863
rect 2273 4815 2727 4863
rect 2273 4485 2335 4815
rect 2665 4485 2727 4815
rect 2273 4437 2727 4485
rect 2744 4437 2750 4863
rect 2250 4431 2750 4437
rect 2800 4863 2864 4869
rect 2800 4437 2806 4863
rect 2823 4836 2864 4863
rect 3236 4869 3269 4871
rect 3381 4894 3819 4900
rect 3381 4877 3387 4894
rect 3813 4877 3819 4894
rect 3381 4871 3819 4877
rect 3379 4869 3821 4871
rect 3931 4894 4369 4900
rect 3931 4877 3937 4894
rect 4363 4877 4369 4894
rect 3931 4871 4369 4877
rect 3931 4869 3964 4871
rect 3236 4863 3300 4869
rect 3236 4836 3277 4863
rect 2823 4464 2829 4836
rect 3271 4464 3277 4836
rect 2823 4437 2864 4464
rect 2800 4431 2864 4437
rect 2136 4429 2169 4431
rect 1731 4423 2169 4429
rect 1731 4406 1737 4423
rect 2163 4406 2169 4423
rect 1731 4400 2169 4406
rect 2279 4429 2721 4431
rect 2281 4423 2719 4429
rect 2281 4406 2287 4423
rect 2713 4406 2719 4423
rect 2281 4400 2719 4406
rect 2831 4429 2864 4431
rect 3236 4437 3277 4464
rect 3294 4437 3300 4863
rect 3236 4431 3300 4437
rect 3350 4863 3850 4869
rect 3350 4437 3356 4863
rect 3373 4815 3827 4863
rect 3373 4485 3435 4815
rect 3765 4485 3827 4815
rect 3373 4437 3827 4485
rect 3844 4437 3850 4863
rect 3350 4431 3850 4437
rect 3900 4863 3964 4869
rect 3900 4437 3906 4863
rect 3923 4836 3964 4863
rect 4336 4869 4369 4871
rect 4481 4894 4919 4900
rect 4481 4877 4487 4894
rect 4913 4877 4919 4894
rect 4481 4871 4919 4877
rect 4479 4869 4921 4871
rect 5031 4894 5469 4900
rect 5031 4877 5037 4894
rect 5463 4877 5469 4894
rect 5031 4871 5469 4877
rect 5031 4869 5064 4871
rect 4336 4863 4400 4869
rect 4336 4836 4377 4863
rect 3923 4464 3929 4836
rect 4371 4464 4377 4836
rect 3923 4437 3964 4464
rect 3900 4431 3964 4437
rect 3236 4429 3269 4431
rect 2831 4423 3269 4429
rect 2831 4406 2837 4423
rect 3263 4406 3269 4423
rect 2831 4400 3269 4406
rect 3379 4429 3821 4431
rect 3381 4423 3819 4429
rect 3381 4406 3387 4423
rect 3813 4406 3819 4423
rect 3381 4400 3819 4406
rect 3931 4429 3964 4431
rect 4336 4437 4377 4464
rect 4394 4437 4400 4863
rect 4336 4431 4400 4437
rect 4450 4863 4950 4869
rect 4450 4437 4456 4863
rect 4473 4815 4927 4863
rect 4473 4485 4535 4815
rect 4865 4485 4927 4815
rect 4473 4437 4927 4485
rect 4944 4437 4950 4863
rect 4450 4431 4950 4437
rect 5000 4863 5064 4869
rect 5000 4437 5006 4863
rect 5023 4836 5064 4863
rect 5436 4869 5469 4871
rect 5581 4894 6019 4900
rect 5581 4877 5587 4894
rect 6013 4877 6019 4894
rect 5581 4871 6019 4877
rect 5579 4869 6021 4871
rect 6131 4894 6569 4900
rect 6131 4877 6137 4894
rect 6563 4877 6569 4894
rect 6131 4871 6569 4877
rect 6131 4869 6164 4871
rect 5436 4863 5500 4869
rect 5436 4836 5477 4863
rect 5023 4464 5029 4836
rect 5471 4464 5477 4836
rect 5023 4437 5064 4464
rect 5000 4431 5064 4437
rect 4336 4429 4369 4431
rect 3931 4423 4369 4429
rect 3931 4406 3937 4423
rect 4363 4406 4369 4423
rect 3931 4400 4369 4406
rect 4479 4429 4921 4431
rect 4481 4423 4919 4429
rect 4481 4406 4487 4423
rect 4913 4406 4919 4423
rect 4481 4400 4919 4406
rect 5031 4429 5064 4431
rect 5436 4437 5477 4464
rect 5494 4437 5500 4863
rect 5436 4431 5500 4437
rect 5550 4863 6050 4869
rect 5550 4437 5556 4863
rect 5573 4815 6027 4863
rect 5573 4485 5635 4815
rect 5965 4485 6027 4815
rect 5573 4437 6027 4485
rect 6044 4437 6050 4863
rect 5550 4431 6050 4437
rect 6100 4863 6164 4869
rect 6100 4437 6106 4863
rect 6123 4836 6164 4863
rect 6536 4869 6569 4871
rect 6681 4894 7119 4900
rect 6681 4877 6687 4894
rect 7113 4877 7119 4894
rect 6681 4871 7119 4877
rect 6679 4869 7121 4871
rect 7231 4894 7669 4900
rect 7231 4877 7237 4894
rect 7663 4877 7669 4894
rect 7231 4871 7669 4877
rect 7231 4869 7264 4871
rect 6536 4863 6600 4869
rect 6536 4836 6577 4863
rect 6123 4464 6129 4836
rect 6571 4464 6577 4836
rect 6123 4437 6164 4464
rect 6100 4431 6164 4437
rect 5436 4429 5469 4431
rect 5031 4423 5469 4429
rect 5031 4406 5037 4423
rect 5463 4406 5469 4423
rect 5031 4400 5469 4406
rect 5579 4429 6021 4431
rect 5581 4423 6019 4429
rect 5581 4406 5587 4423
rect 6013 4406 6019 4423
rect 5581 4400 6019 4406
rect 6131 4429 6164 4431
rect 6536 4437 6577 4464
rect 6594 4437 6600 4863
rect 6536 4431 6600 4437
rect 6650 4863 7150 4869
rect 6650 4437 6656 4863
rect 6673 4815 7127 4863
rect 6673 4485 6735 4815
rect 7065 4485 7127 4815
rect 6673 4437 7127 4485
rect 7144 4437 7150 4863
rect 6650 4431 7150 4437
rect 7200 4863 7264 4869
rect 7200 4437 7206 4863
rect 7223 4836 7264 4863
rect 7636 4869 7669 4871
rect 7781 4894 8219 4900
rect 7781 4877 7787 4894
rect 8213 4877 8219 4894
rect 7781 4871 8219 4877
rect 7779 4869 8221 4871
rect 8331 4894 8769 4900
rect 8331 4877 8337 4894
rect 8763 4877 8769 4894
rect 8331 4871 8769 4877
rect 8331 4869 8364 4871
rect 7636 4863 7700 4869
rect 7636 4836 7677 4863
rect 7223 4464 7229 4836
rect 7671 4464 7677 4836
rect 7223 4437 7264 4464
rect 7200 4431 7264 4437
rect 6536 4429 6569 4431
rect 6131 4423 6569 4429
rect 6131 4406 6137 4423
rect 6563 4406 6569 4423
rect 6131 4400 6569 4406
rect 6679 4429 7121 4431
rect 6681 4423 7119 4429
rect 6681 4406 6687 4423
rect 7113 4406 7119 4423
rect 6681 4400 7119 4406
rect 7231 4429 7264 4431
rect 7636 4437 7677 4464
rect 7694 4437 7700 4863
rect 7636 4431 7700 4437
rect 7750 4863 8250 4869
rect 7750 4437 7756 4863
rect 7773 4815 8227 4863
rect 7773 4485 7835 4815
rect 8165 4485 8227 4815
rect 7773 4437 8227 4485
rect 8244 4437 8250 4863
rect 7750 4431 8250 4437
rect 8300 4863 8364 4869
rect 8300 4437 8306 4863
rect 8323 4836 8364 4863
rect 8736 4869 8769 4871
rect 8881 4894 9319 4900
rect 8881 4877 8887 4894
rect 9313 4877 9319 4894
rect 8881 4871 9319 4877
rect 8879 4869 9321 4871
rect 9431 4894 9869 4900
rect 9431 4877 9437 4894
rect 9863 4877 9869 4894
rect 9431 4871 9869 4877
rect 9431 4869 9464 4871
rect 8736 4863 8800 4869
rect 8736 4836 8777 4863
rect 8323 4464 8329 4836
rect 8771 4464 8777 4836
rect 8323 4437 8364 4464
rect 8300 4431 8364 4437
rect 7636 4429 7669 4431
rect 7231 4423 7669 4429
rect 7231 4406 7237 4423
rect 7663 4406 7669 4423
rect 7231 4400 7669 4406
rect 7779 4429 8221 4431
rect 7781 4423 8219 4429
rect 7781 4406 7787 4423
rect 8213 4406 8219 4423
rect 7781 4400 8219 4406
rect 8331 4429 8364 4431
rect 8736 4437 8777 4464
rect 8794 4437 8800 4863
rect 8736 4431 8800 4437
rect 8850 4863 9350 4869
rect 8850 4437 8856 4863
rect 8873 4815 9327 4863
rect 8873 4485 8935 4815
rect 9265 4485 9327 4815
rect 8873 4437 9327 4485
rect 9344 4437 9350 4863
rect 8850 4431 9350 4437
rect 9400 4863 9464 4869
rect 9400 4437 9406 4863
rect 9423 4836 9464 4863
rect 9836 4869 9869 4871
rect 9981 4894 10419 4900
rect 9981 4877 9987 4894
rect 10413 4877 10419 4894
rect 9981 4871 10419 4877
rect 9979 4869 10421 4871
rect 10531 4894 10969 4900
rect 10531 4877 10537 4894
rect 10963 4877 10969 4894
rect 10531 4871 10969 4877
rect 10531 4869 10564 4871
rect 9836 4863 9900 4869
rect 9836 4836 9877 4863
rect 9423 4464 9429 4836
rect 9871 4464 9877 4836
rect 9423 4437 9464 4464
rect 9400 4431 9464 4437
rect 8736 4429 8769 4431
rect 8331 4423 8769 4429
rect 8331 4406 8337 4423
rect 8763 4406 8769 4423
rect 8331 4400 8769 4406
rect 8879 4429 9321 4431
rect 8881 4423 9319 4429
rect 8881 4406 8887 4423
rect 9313 4406 9319 4423
rect 8881 4400 9319 4406
rect 9431 4429 9464 4431
rect 9836 4437 9877 4464
rect 9894 4437 9900 4863
rect 9836 4431 9900 4437
rect 9950 4863 10450 4869
rect 9950 4437 9956 4863
rect 9973 4815 10427 4863
rect 9973 4485 10035 4815
rect 10365 4485 10427 4815
rect 9973 4437 10427 4485
rect 10444 4437 10450 4863
rect 9950 4431 10450 4437
rect 10500 4863 10564 4869
rect 10500 4437 10506 4863
rect 10523 4836 10564 4863
rect 10936 4869 10969 4871
rect 11081 4894 11519 4900
rect 11081 4877 11087 4894
rect 11513 4877 11519 4894
rect 11081 4871 11519 4877
rect 11079 4869 11521 4871
rect 11631 4894 12069 4900
rect 11631 4877 11637 4894
rect 12063 4877 12069 4894
rect 11631 4871 12069 4877
rect 11631 4869 11664 4871
rect 10936 4863 11000 4869
rect 10936 4836 10977 4863
rect 10523 4464 10529 4836
rect 10971 4464 10977 4836
rect 10523 4437 10564 4464
rect 10500 4431 10564 4437
rect 9836 4429 9869 4431
rect 9431 4423 9869 4429
rect 9431 4406 9437 4423
rect 9863 4406 9869 4423
rect 9431 4400 9869 4406
rect 9979 4429 10421 4431
rect 9981 4423 10419 4429
rect 9981 4406 9987 4423
rect 10413 4406 10419 4423
rect 9981 4400 10419 4406
rect 10531 4429 10564 4431
rect 10936 4437 10977 4464
rect 10994 4437 11000 4863
rect 10936 4431 11000 4437
rect 11050 4863 11550 4869
rect 11050 4437 11056 4863
rect 11073 4815 11527 4863
rect 11073 4485 11135 4815
rect 11465 4485 11527 4815
rect 11073 4437 11527 4485
rect 11544 4437 11550 4863
rect 11050 4431 11550 4437
rect 11600 4863 11664 4869
rect 11600 4437 11606 4863
rect 11623 4836 11664 4863
rect 12036 4869 12069 4871
rect 12181 4894 12619 4900
rect 12181 4877 12187 4894
rect 12613 4877 12619 4894
rect 12181 4871 12619 4877
rect 12179 4869 12621 4871
rect 12731 4894 13169 4900
rect 12731 4877 12737 4894
rect 13163 4877 13169 4894
rect 12731 4871 13169 4877
rect 12731 4869 12764 4871
rect 12036 4863 12100 4869
rect 12036 4836 12077 4863
rect 11623 4464 11629 4836
rect 12071 4464 12077 4836
rect 11623 4437 11664 4464
rect 11600 4431 11664 4437
rect 10936 4429 10969 4431
rect 10531 4423 10969 4429
rect 10531 4406 10537 4423
rect 10963 4406 10969 4423
rect 10531 4400 10969 4406
rect 11079 4429 11521 4431
rect 11081 4423 11519 4429
rect 11081 4406 11087 4423
rect 11513 4406 11519 4423
rect 11081 4400 11519 4406
rect 11631 4429 11664 4431
rect 12036 4437 12077 4464
rect 12094 4437 12100 4863
rect 12036 4431 12100 4437
rect 12150 4863 12650 4869
rect 12150 4437 12156 4863
rect 12173 4815 12627 4863
rect 12173 4485 12235 4815
rect 12565 4485 12627 4815
rect 12173 4437 12627 4485
rect 12644 4437 12650 4863
rect 12150 4431 12650 4437
rect 12700 4863 12764 4869
rect 12700 4437 12706 4863
rect 12723 4836 12764 4863
rect 13136 4869 13169 4871
rect 13281 4894 13719 4900
rect 13281 4877 13287 4894
rect 13713 4877 13719 4894
rect 13281 4871 13719 4877
rect 13279 4869 13721 4871
rect 13136 4863 13200 4869
rect 13136 4836 13177 4863
rect 12723 4464 12729 4836
rect 13171 4464 13177 4836
rect 12723 4437 12764 4464
rect 12700 4431 12764 4437
rect 12036 4429 12069 4431
rect 11631 4423 12069 4429
rect 11631 4406 11637 4423
rect 12063 4406 12069 4423
rect 11631 4400 12069 4406
rect 12179 4429 12621 4431
rect 12181 4423 12619 4429
rect 12181 4406 12187 4423
rect 12613 4406 12619 4423
rect 12181 4400 12619 4406
rect 12731 4429 12764 4431
rect 13136 4437 13177 4464
rect 13194 4437 13200 4863
rect 13136 4431 13200 4437
rect 13250 4863 13721 4869
rect 13250 4437 13256 4863
rect 13273 4815 13721 4863
rect 13273 4485 13335 4815
rect 13665 4485 13721 4815
rect 13273 4437 13721 4485
rect 13250 4431 13721 4437
rect 13136 4429 13169 4431
rect 12731 4423 13169 4429
rect 12731 4406 12737 4423
rect 13163 4406 13169 4423
rect 12731 4400 13169 4406
rect 13279 4429 13721 4431
rect 13281 4423 13719 4429
rect 13281 4406 13287 4423
rect 13713 4406 13719 4423
rect 13281 4400 13719 4406
rect -469 4344 -31 4350
rect -469 4327 -463 4344
rect -37 4327 -31 4344
rect -469 4321 -31 4327
rect -471 4319 -29 4321
rect 81 4344 519 4350
rect 81 4327 87 4344
rect 513 4327 519 4344
rect 81 4321 519 4327
rect 81 4319 114 4321
rect -471 4313 0 4319
rect -471 4265 -23 4313
rect -471 3935 -415 4265
rect -85 3935 -23 4265
rect -471 3887 -23 3935
rect -6 3887 0 4313
rect -471 3881 0 3887
rect 50 4313 114 4319
rect 50 3887 56 4313
rect 73 4286 114 4313
rect 486 4319 519 4321
rect 631 4344 1069 4350
rect 631 4327 637 4344
rect 1063 4327 1069 4344
rect 631 4321 1069 4327
rect 629 4319 1071 4321
rect 1181 4344 1619 4350
rect 1181 4327 1187 4344
rect 1613 4327 1619 4344
rect 1181 4321 1619 4327
rect 1181 4319 1214 4321
rect 486 4313 550 4319
rect 486 4286 527 4313
rect 73 3914 79 4286
rect 521 3914 527 4286
rect 73 3887 114 3914
rect 50 3881 114 3887
rect -471 3879 -29 3881
rect -469 3873 -31 3879
rect -469 3856 -463 3873
rect -37 3856 -31 3873
rect -469 3850 -31 3856
rect 81 3879 114 3881
rect 486 3887 527 3914
rect 544 3887 550 4313
rect 486 3881 550 3887
rect 600 4313 1100 4319
rect 600 3887 606 4313
rect 623 4265 1077 4313
rect 623 3935 685 4265
rect 1015 3935 1077 4265
rect 623 3887 1077 3935
rect 1094 3887 1100 4313
rect 600 3881 1100 3887
rect 1150 4313 1214 4319
rect 1150 3887 1156 4313
rect 1173 4286 1214 4313
rect 1586 4319 1619 4321
rect 1731 4344 2169 4350
rect 1731 4327 1737 4344
rect 2163 4327 2169 4344
rect 1731 4321 2169 4327
rect 1729 4319 2171 4321
rect 2281 4344 2719 4350
rect 2281 4327 2287 4344
rect 2713 4327 2719 4344
rect 2281 4321 2719 4327
rect 2281 4319 2314 4321
rect 1586 4313 1650 4319
rect 1586 4286 1627 4313
rect 1173 3914 1179 4286
rect 1621 3914 1627 4286
rect 1173 3887 1214 3914
rect 1150 3881 1214 3887
rect 486 3879 519 3881
rect 81 3873 519 3879
rect 81 3856 87 3873
rect 513 3856 519 3873
rect 81 3850 519 3856
rect 629 3879 1071 3881
rect 631 3873 1069 3879
rect 631 3856 637 3873
rect 1063 3856 1069 3873
rect 631 3850 1069 3856
rect 1181 3879 1214 3881
rect 1586 3887 1627 3914
rect 1644 3887 1650 4313
rect 1586 3881 1650 3887
rect 1700 4313 2200 4319
rect 1700 3887 1706 4313
rect 1723 4265 2177 4313
rect 1723 3935 1785 4265
rect 2115 3935 2177 4265
rect 1723 3887 2177 3935
rect 2194 3887 2200 4313
rect 1700 3881 2200 3887
rect 2250 4313 2314 4319
rect 2250 3887 2256 4313
rect 2273 4286 2314 4313
rect 2686 4319 2719 4321
rect 2831 4344 3269 4350
rect 2831 4327 2837 4344
rect 3263 4327 3269 4344
rect 2831 4321 3269 4327
rect 2829 4319 3271 4321
rect 3381 4344 3819 4350
rect 3381 4327 3387 4344
rect 3813 4327 3819 4344
rect 3381 4321 3819 4327
rect 3381 4319 3414 4321
rect 2686 4313 2750 4319
rect 2686 4286 2727 4313
rect 2273 3914 2279 4286
rect 2721 3914 2727 4286
rect 2273 3887 2314 3914
rect 2250 3881 2314 3887
rect 1586 3879 1619 3881
rect 1181 3873 1619 3879
rect 1181 3856 1187 3873
rect 1613 3856 1619 3873
rect 1181 3850 1619 3856
rect 1729 3879 2171 3881
rect 1731 3873 2169 3879
rect 1731 3856 1737 3873
rect 2163 3856 2169 3873
rect 1731 3850 2169 3856
rect 2281 3879 2314 3881
rect 2686 3887 2727 3914
rect 2744 3887 2750 4313
rect 2686 3881 2750 3887
rect 2800 4313 3300 4319
rect 2800 3887 2806 4313
rect 2823 4265 3277 4313
rect 2823 3935 2885 4265
rect 3215 3935 3277 4265
rect 2823 3887 3277 3935
rect 3294 3887 3300 4313
rect 2800 3881 3300 3887
rect 3350 4313 3414 4319
rect 3350 3887 3356 4313
rect 3373 4286 3414 4313
rect 3786 4319 3819 4321
rect 3931 4344 4369 4350
rect 3931 4327 3937 4344
rect 4363 4327 4369 4344
rect 3931 4321 4369 4327
rect 3929 4319 4371 4321
rect 4481 4344 4919 4350
rect 4481 4327 4487 4344
rect 4913 4327 4919 4344
rect 4481 4321 4919 4327
rect 4481 4319 4514 4321
rect 3786 4313 3850 4319
rect 3786 4286 3827 4313
rect 3373 3914 3379 4286
rect 3821 3914 3827 4286
rect 3373 3887 3414 3914
rect 3350 3881 3414 3887
rect 2686 3879 2719 3881
rect 2281 3873 2719 3879
rect 2281 3856 2287 3873
rect 2713 3856 2719 3873
rect 2281 3850 2719 3856
rect 2829 3879 3271 3881
rect 2831 3873 3269 3879
rect 2831 3856 2837 3873
rect 3263 3856 3269 3873
rect 2831 3850 3269 3856
rect 3381 3879 3414 3881
rect 3786 3887 3827 3914
rect 3844 3887 3850 4313
rect 3786 3881 3850 3887
rect 3900 4313 4400 4319
rect 3900 3887 3906 4313
rect 3923 4265 4377 4313
rect 3923 3935 3985 4265
rect 4315 3935 4377 4265
rect 3923 3887 4377 3935
rect 4394 3887 4400 4313
rect 3900 3881 4400 3887
rect 4450 4313 4514 4319
rect 4450 3887 4456 4313
rect 4473 4286 4514 4313
rect 4886 4319 4919 4321
rect 5031 4344 5469 4350
rect 5031 4327 5037 4344
rect 5463 4327 5469 4344
rect 5031 4321 5469 4327
rect 5029 4319 5471 4321
rect 5581 4344 6019 4350
rect 5581 4327 5587 4344
rect 6013 4327 6019 4344
rect 5581 4321 6019 4327
rect 5581 4319 5614 4321
rect 4886 4313 4950 4319
rect 4886 4286 4927 4313
rect 4473 3914 4479 4286
rect 4921 3914 4927 4286
rect 4473 3887 4514 3914
rect 4450 3881 4514 3887
rect 3786 3879 3819 3881
rect 3381 3873 3819 3879
rect 3381 3856 3387 3873
rect 3813 3856 3819 3873
rect 3381 3850 3819 3856
rect 3929 3879 4371 3881
rect 3931 3873 4369 3879
rect 3931 3856 3937 3873
rect 4363 3856 4369 3873
rect 3931 3850 4369 3856
rect 4481 3879 4514 3881
rect 4886 3887 4927 3914
rect 4944 3887 4950 4313
rect 4886 3881 4950 3887
rect 5000 4313 5500 4319
rect 5000 3887 5006 4313
rect 5023 4265 5477 4313
rect 5023 3935 5085 4265
rect 5415 3935 5477 4265
rect 5023 3887 5477 3935
rect 5494 3887 5500 4313
rect 5000 3881 5500 3887
rect 5550 4313 5614 4319
rect 5550 3887 5556 4313
rect 5573 4286 5614 4313
rect 5986 4319 6019 4321
rect 6131 4344 6569 4350
rect 6131 4327 6137 4344
rect 6563 4327 6569 4344
rect 6131 4321 6569 4327
rect 6129 4319 6571 4321
rect 6681 4344 7119 4350
rect 6681 4327 6687 4344
rect 7113 4327 7119 4344
rect 6681 4321 7119 4327
rect 6681 4319 6714 4321
rect 5986 4313 6050 4319
rect 5986 4286 6027 4313
rect 5573 3914 5579 4286
rect 6021 3914 6027 4286
rect 5573 3887 5614 3914
rect 5550 3881 5614 3887
rect 4886 3879 4919 3881
rect 4481 3873 4919 3879
rect 4481 3856 4487 3873
rect 4913 3856 4919 3873
rect 4481 3850 4919 3856
rect 5029 3879 5471 3881
rect 5031 3873 5469 3879
rect 5031 3856 5037 3873
rect 5463 3856 5469 3873
rect 5031 3850 5469 3856
rect 5581 3879 5614 3881
rect 5986 3887 6027 3914
rect 6044 3887 6050 4313
rect 5986 3881 6050 3887
rect 6100 4313 6600 4319
rect 6100 3887 6106 4313
rect 6123 4265 6577 4313
rect 6123 3935 6185 4265
rect 6515 3935 6577 4265
rect 6123 3887 6577 3935
rect 6594 3887 6600 4313
rect 6100 3881 6600 3887
rect 6650 4313 6714 4319
rect 6650 3887 6656 4313
rect 6673 4286 6714 4313
rect 7086 4319 7119 4321
rect 7231 4344 7669 4350
rect 7231 4327 7237 4344
rect 7663 4327 7669 4344
rect 7231 4321 7669 4327
rect 7229 4319 7671 4321
rect 7781 4344 8219 4350
rect 7781 4327 7787 4344
rect 8213 4327 8219 4344
rect 7781 4321 8219 4327
rect 7781 4319 7814 4321
rect 7086 4313 7150 4319
rect 7086 4286 7127 4313
rect 6673 3914 6679 4286
rect 7121 3914 7127 4286
rect 6673 3887 6714 3914
rect 6650 3881 6714 3887
rect 5986 3879 6019 3881
rect 5581 3873 6019 3879
rect 5581 3856 5587 3873
rect 6013 3856 6019 3873
rect 5581 3850 6019 3856
rect 6129 3879 6571 3881
rect 6131 3873 6569 3879
rect 6131 3856 6137 3873
rect 6563 3856 6569 3873
rect 6131 3850 6569 3856
rect 6681 3879 6714 3881
rect 7086 3887 7127 3914
rect 7144 3887 7150 4313
rect 7086 3881 7150 3887
rect 7200 4313 7700 4319
rect 7200 3887 7206 4313
rect 7223 4265 7677 4313
rect 7223 3935 7285 4265
rect 7615 3935 7677 4265
rect 7223 3887 7677 3935
rect 7694 3887 7700 4313
rect 7200 3881 7700 3887
rect 7750 4313 7814 4319
rect 7750 3887 7756 4313
rect 7773 4286 7814 4313
rect 8186 4319 8219 4321
rect 8331 4344 8769 4350
rect 8331 4327 8337 4344
rect 8763 4327 8769 4344
rect 8331 4321 8769 4327
rect 8329 4319 8771 4321
rect 8881 4344 9319 4350
rect 8881 4327 8887 4344
rect 9313 4327 9319 4344
rect 8881 4321 9319 4327
rect 8881 4319 8914 4321
rect 8186 4313 8250 4319
rect 8186 4286 8227 4313
rect 7773 3914 7779 4286
rect 8221 3914 8227 4286
rect 7773 3887 7814 3914
rect 7750 3881 7814 3887
rect 7086 3879 7119 3881
rect 6681 3873 7119 3879
rect 6681 3856 6687 3873
rect 7113 3856 7119 3873
rect 6681 3850 7119 3856
rect 7229 3879 7671 3881
rect 7231 3873 7669 3879
rect 7231 3856 7237 3873
rect 7663 3856 7669 3873
rect 7231 3850 7669 3856
rect 7781 3879 7814 3881
rect 8186 3887 8227 3914
rect 8244 3887 8250 4313
rect 8186 3881 8250 3887
rect 8300 4313 8800 4319
rect 8300 3887 8306 4313
rect 8323 4265 8777 4313
rect 8323 3935 8385 4265
rect 8715 3935 8777 4265
rect 8323 3887 8777 3935
rect 8794 3887 8800 4313
rect 8300 3881 8800 3887
rect 8850 4313 8914 4319
rect 8850 3887 8856 4313
rect 8873 4286 8914 4313
rect 9286 4319 9319 4321
rect 9431 4344 9869 4350
rect 9431 4327 9437 4344
rect 9863 4327 9869 4344
rect 9431 4321 9869 4327
rect 9429 4319 9871 4321
rect 9981 4344 10419 4350
rect 9981 4327 9987 4344
rect 10413 4327 10419 4344
rect 9981 4321 10419 4327
rect 9981 4319 10014 4321
rect 9286 4313 9350 4319
rect 9286 4286 9327 4313
rect 8873 3914 8879 4286
rect 9321 3914 9327 4286
rect 8873 3887 8914 3914
rect 8850 3881 8914 3887
rect 8186 3879 8219 3881
rect 7781 3873 8219 3879
rect 7781 3856 7787 3873
rect 8213 3856 8219 3873
rect 7781 3850 8219 3856
rect 8329 3879 8771 3881
rect 8331 3873 8769 3879
rect 8331 3856 8337 3873
rect 8763 3856 8769 3873
rect 8331 3850 8769 3856
rect 8881 3879 8914 3881
rect 9286 3887 9327 3914
rect 9344 3887 9350 4313
rect 9286 3881 9350 3887
rect 9400 4313 9900 4319
rect 9400 3887 9406 4313
rect 9423 4265 9877 4313
rect 9423 3935 9485 4265
rect 9815 3935 9877 4265
rect 9423 3887 9877 3935
rect 9894 3887 9900 4313
rect 9400 3881 9900 3887
rect 9950 4313 10014 4319
rect 9950 3887 9956 4313
rect 9973 4286 10014 4313
rect 10386 4319 10419 4321
rect 10531 4344 10969 4350
rect 10531 4327 10537 4344
rect 10963 4327 10969 4344
rect 10531 4321 10969 4327
rect 10529 4319 10971 4321
rect 11081 4344 11519 4350
rect 11081 4327 11087 4344
rect 11513 4327 11519 4344
rect 11081 4321 11519 4327
rect 11081 4319 11114 4321
rect 10386 4313 10450 4319
rect 10386 4286 10427 4313
rect 9973 3914 9979 4286
rect 10421 3914 10427 4286
rect 9973 3887 10014 3914
rect 9950 3881 10014 3887
rect 9286 3879 9319 3881
rect 8881 3873 9319 3879
rect 8881 3856 8887 3873
rect 9313 3856 9319 3873
rect 8881 3850 9319 3856
rect 9429 3879 9871 3881
rect 9431 3873 9869 3879
rect 9431 3856 9437 3873
rect 9863 3856 9869 3873
rect 9431 3850 9869 3856
rect 9981 3879 10014 3881
rect 10386 3887 10427 3914
rect 10444 3887 10450 4313
rect 10386 3881 10450 3887
rect 10500 4313 11000 4319
rect 10500 3887 10506 4313
rect 10523 4265 10977 4313
rect 10523 3935 10585 4265
rect 10915 3935 10977 4265
rect 10523 3887 10977 3935
rect 10994 3887 11000 4313
rect 10500 3881 11000 3887
rect 11050 4313 11114 4319
rect 11050 3887 11056 4313
rect 11073 4286 11114 4313
rect 11486 4319 11519 4321
rect 11631 4344 12069 4350
rect 11631 4327 11637 4344
rect 12063 4327 12069 4344
rect 11631 4321 12069 4327
rect 11629 4319 12071 4321
rect 12181 4344 12619 4350
rect 12181 4327 12187 4344
rect 12613 4327 12619 4344
rect 12181 4321 12619 4327
rect 12181 4319 12214 4321
rect 11486 4313 11550 4319
rect 11486 4286 11527 4313
rect 11073 3914 11079 4286
rect 11521 3914 11527 4286
rect 11073 3887 11114 3914
rect 11050 3881 11114 3887
rect 10386 3879 10419 3881
rect 9981 3873 10419 3879
rect 9981 3856 9987 3873
rect 10413 3856 10419 3873
rect 9981 3850 10419 3856
rect 10529 3879 10971 3881
rect 10531 3873 10969 3879
rect 10531 3856 10537 3873
rect 10963 3856 10969 3873
rect 10531 3850 10969 3856
rect 11081 3879 11114 3881
rect 11486 3887 11527 3914
rect 11544 3887 11550 4313
rect 11486 3881 11550 3887
rect 11600 4313 12100 4319
rect 11600 3887 11606 4313
rect 11623 4265 12077 4313
rect 11623 3935 11685 4265
rect 12015 3935 12077 4265
rect 11623 3887 12077 3935
rect 12094 3887 12100 4313
rect 11600 3881 12100 3887
rect 12150 4313 12214 4319
rect 12150 3887 12156 4313
rect 12173 4286 12214 4313
rect 12586 4319 12619 4321
rect 12731 4344 13169 4350
rect 12731 4327 12737 4344
rect 13163 4327 13169 4344
rect 12731 4321 13169 4327
rect 12729 4319 13171 4321
rect 13281 4344 13719 4350
rect 13281 4327 13287 4344
rect 13713 4327 13719 4344
rect 13281 4321 13719 4327
rect 13281 4319 13314 4321
rect 12586 4313 12650 4319
rect 12586 4286 12627 4313
rect 12173 3914 12179 4286
rect 12621 3914 12627 4286
rect 12173 3887 12214 3914
rect 12150 3881 12214 3887
rect 11486 3879 11519 3881
rect 11081 3873 11519 3879
rect 11081 3856 11087 3873
rect 11513 3856 11519 3873
rect 11081 3850 11519 3856
rect 11629 3879 12071 3881
rect 11631 3873 12069 3879
rect 11631 3856 11637 3873
rect 12063 3856 12069 3873
rect 11631 3850 12069 3856
rect 12181 3879 12214 3881
rect 12586 3887 12627 3914
rect 12644 3887 12650 4313
rect 12586 3881 12650 3887
rect 12700 4313 13200 4319
rect 12700 3887 12706 4313
rect 12723 4265 13177 4313
rect 12723 3935 12785 4265
rect 13115 3935 13177 4265
rect 12723 3887 13177 3935
rect 13194 3887 13200 4313
rect 12700 3881 13200 3887
rect 13250 4313 13314 4319
rect 13250 3887 13256 4313
rect 13273 4286 13314 4313
rect 13273 3914 13279 4286
rect 13273 3887 13314 3914
rect 13250 3881 13314 3887
rect 12586 3879 12619 3881
rect 12181 3873 12619 3879
rect 12181 3856 12187 3873
rect 12613 3856 12619 3873
rect 12181 3850 12619 3856
rect 12729 3879 13171 3881
rect 12731 3873 13169 3879
rect 12731 3856 12737 3873
rect 13163 3856 13169 3873
rect 12731 3850 13169 3856
rect 13281 3879 13314 3881
rect 13281 3873 13719 3879
rect 13281 3856 13287 3873
rect 13713 3856 13719 3873
rect 13281 3850 13719 3856
rect -469 3794 -31 3800
rect -469 3777 -463 3794
rect -37 3777 -31 3794
rect -469 3771 -31 3777
rect -64 3769 -31 3771
rect 81 3794 519 3800
rect 81 3777 87 3794
rect 513 3777 519 3794
rect 81 3771 519 3777
rect 79 3769 521 3771
rect 631 3794 1069 3800
rect 631 3777 637 3794
rect 1063 3777 1069 3794
rect 631 3771 1069 3777
rect 631 3769 664 3771
rect -64 3763 0 3769
rect -64 3736 -23 3763
rect -29 3364 -23 3736
rect -64 3337 -23 3364
rect -6 3337 0 3763
rect -64 3331 0 3337
rect 50 3763 550 3769
rect 50 3337 56 3763
rect 73 3715 527 3763
rect 73 3385 135 3715
rect 465 3385 527 3715
rect 73 3337 527 3385
rect 544 3337 550 3763
rect 50 3331 550 3337
rect 600 3763 664 3769
rect 600 3337 606 3763
rect 623 3736 664 3763
rect 1036 3769 1069 3771
rect 1181 3794 1619 3800
rect 1181 3777 1187 3794
rect 1613 3777 1619 3794
rect 1181 3771 1619 3777
rect 1179 3769 1621 3771
rect 1731 3794 2169 3800
rect 1731 3777 1737 3794
rect 2163 3777 2169 3794
rect 1731 3771 2169 3777
rect 1731 3769 1764 3771
rect 1036 3763 1100 3769
rect 1036 3736 1077 3763
rect 623 3364 629 3736
rect 1071 3364 1077 3736
rect 623 3337 664 3364
rect 600 3331 664 3337
rect -64 3329 -31 3331
rect -469 3323 -31 3329
rect -469 3306 -463 3323
rect -37 3306 -31 3323
rect -469 3300 -31 3306
rect 79 3329 521 3331
rect 81 3323 519 3329
rect 81 3306 87 3323
rect 513 3306 519 3323
rect 81 3300 519 3306
rect 631 3329 664 3331
rect 1036 3337 1077 3364
rect 1094 3337 1100 3763
rect 1036 3331 1100 3337
rect 1150 3763 1650 3769
rect 1150 3337 1156 3763
rect 1173 3715 1627 3763
rect 1173 3385 1235 3715
rect 1565 3385 1627 3715
rect 1173 3337 1627 3385
rect 1644 3337 1650 3763
rect 1150 3331 1650 3337
rect 1700 3763 1764 3769
rect 1700 3337 1706 3763
rect 1723 3736 1764 3763
rect 2136 3769 2169 3771
rect 2281 3794 2719 3800
rect 2281 3777 2287 3794
rect 2713 3777 2719 3794
rect 2281 3771 2719 3777
rect 2279 3769 2721 3771
rect 2831 3794 3269 3800
rect 2831 3777 2837 3794
rect 3263 3777 3269 3794
rect 2831 3771 3269 3777
rect 2831 3769 2864 3771
rect 2136 3763 2200 3769
rect 2136 3736 2177 3763
rect 1723 3364 1729 3736
rect 2171 3364 2177 3736
rect 1723 3337 1764 3364
rect 1700 3331 1764 3337
rect 1036 3329 1069 3331
rect 631 3323 1069 3329
rect 631 3306 637 3323
rect 1063 3306 1069 3323
rect 631 3300 1069 3306
rect 1179 3329 1621 3331
rect 1181 3323 1619 3329
rect 1181 3306 1187 3323
rect 1613 3306 1619 3323
rect 1181 3300 1619 3306
rect 1731 3329 1764 3331
rect 2136 3337 2177 3364
rect 2194 3337 2200 3763
rect 2136 3331 2200 3337
rect 2250 3763 2750 3769
rect 2250 3337 2256 3763
rect 2273 3715 2727 3763
rect 2273 3385 2335 3715
rect 2665 3385 2727 3715
rect 2273 3337 2727 3385
rect 2744 3337 2750 3763
rect 2250 3331 2750 3337
rect 2800 3763 2864 3769
rect 2800 3337 2806 3763
rect 2823 3736 2864 3763
rect 3236 3769 3269 3771
rect 3381 3794 3819 3800
rect 3381 3777 3387 3794
rect 3813 3777 3819 3794
rect 3381 3771 3819 3777
rect 3379 3769 3821 3771
rect 3931 3794 4369 3800
rect 3931 3777 3937 3794
rect 4363 3777 4369 3794
rect 3931 3771 4369 3777
rect 3931 3769 3964 3771
rect 3236 3763 3300 3769
rect 3236 3736 3277 3763
rect 2823 3364 2829 3736
rect 3271 3364 3277 3736
rect 2823 3337 2864 3364
rect 2800 3331 2864 3337
rect 2136 3329 2169 3331
rect 1731 3323 2169 3329
rect 1731 3306 1737 3323
rect 2163 3306 2169 3323
rect 1731 3300 2169 3306
rect 2279 3329 2721 3331
rect 2281 3323 2719 3329
rect 2281 3306 2287 3323
rect 2713 3306 2719 3323
rect 2281 3300 2719 3306
rect 2831 3329 2864 3331
rect 3236 3337 3277 3364
rect 3294 3337 3300 3763
rect 3236 3331 3300 3337
rect 3350 3763 3850 3769
rect 3350 3337 3356 3763
rect 3373 3715 3827 3763
rect 3373 3385 3435 3715
rect 3765 3385 3827 3715
rect 3373 3337 3827 3385
rect 3844 3337 3850 3763
rect 3350 3331 3850 3337
rect 3900 3763 3964 3769
rect 3900 3337 3906 3763
rect 3923 3736 3964 3763
rect 4336 3769 4369 3771
rect 4481 3794 4919 3800
rect 4481 3777 4487 3794
rect 4913 3777 4919 3794
rect 4481 3771 4919 3777
rect 4479 3769 4921 3771
rect 5031 3794 5469 3800
rect 5031 3777 5037 3794
rect 5463 3777 5469 3794
rect 5031 3771 5469 3777
rect 5031 3769 5064 3771
rect 4336 3763 4400 3769
rect 4336 3736 4377 3763
rect 3923 3364 3929 3736
rect 4371 3364 4377 3736
rect 3923 3337 3964 3364
rect 3900 3331 3964 3337
rect 3236 3329 3269 3331
rect 2831 3323 3269 3329
rect 2831 3306 2837 3323
rect 3263 3306 3269 3323
rect 2831 3300 3269 3306
rect 3379 3329 3821 3331
rect 3381 3323 3819 3329
rect 3381 3306 3387 3323
rect 3813 3306 3819 3323
rect 3381 3300 3819 3306
rect 3931 3329 3964 3331
rect 4336 3337 4377 3364
rect 4394 3337 4400 3763
rect 4336 3331 4400 3337
rect 4450 3763 4950 3769
rect 4450 3337 4456 3763
rect 4473 3715 4927 3763
rect 4473 3385 4535 3715
rect 4865 3385 4927 3715
rect 4473 3337 4927 3385
rect 4944 3337 4950 3763
rect 4450 3331 4950 3337
rect 5000 3763 5064 3769
rect 5000 3337 5006 3763
rect 5023 3736 5064 3763
rect 5436 3769 5469 3771
rect 5581 3794 6019 3800
rect 5581 3777 5587 3794
rect 6013 3777 6019 3794
rect 5581 3771 6019 3777
rect 5579 3769 6021 3771
rect 6131 3794 6569 3800
rect 6131 3777 6137 3794
rect 6563 3777 6569 3794
rect 6131 3771 6569 3777
rect 6131 3769 6164 3771
rect 5436 3763 5500 3769
rect 5436 3736 5477 3763
rect 5023 3364 5029 3736
rect 5471 3364 5477 3736
rect 5023 3337 5064 3364
rect 5000 3331 5064 3337
rect 4336 3329 4369 3331
rect 3931 3323 4369 3329
rect 3931 3306 3937 3323
rect 4363 3306 4369 3323
rect 3931 3300 4369 3306
rect 4479 3329 4921 3331
rect 4481 3323 4919 3329
rect 4481 3306 4487 3323
rect 4913 3306 4919 3323
rect 4481 3300 4919 3306
rect 5031 3329 5064 3331
rect 5436 3337 5477 3364
rect 5494 3337 5500 3763
rect 5436 3331 5500 3337
rect 5550 3763 6050 3769
rect 5550 3337 5556 3763
rect 5573 3715 6027 3763
rect 5573 3385 5635 3715
rect 5965 3385 6027 3715
rect 5573 3337 6027 3385
rect 6044 3337 6050 3763
rect 5550 3331 6050 3337
rect 6100 3763 6164 3769
rect 6100 3337 6106 3763
rect 6123 3736 6164 3763
rect 6536 3769 6569 3771
rect 6681 3794 7119 3800
rect 6681 3777 6687 3794
rect 7113 3777 7119 3794
rect 6681 3771 7119 3777
rect 6679 3769 7121 3771
rect 7231 3794 7669 3800
rect 7231 3777 7237 3794
rect 7663 3777 7669 3794
rect 7231 3771 7669 3777
rect 7231 3769 7264 3771
rect 6536 3763 6600 3769
rect 6536 3736 6577 3763
rect 6123 3364 6129 3736
rect 6571 3364 6577 3736
rect 6123 3337 6164 3364
rect 6100 3331 6164 3337
rect 5436 3329 5469 3331
rect 5031 3323 5469 3329
rect 5031 3306 5037 3323
rect 5463 3306 5469 3323
rect 5031 3300 5469 3306
rect 5579 3329 6021 3331
rect 5581 3323 6019 3329
rect 5581 3306 5587 3323
rect 6013 3306 6019 3323
rect 5581 3300 6019 3306
rect 6131 3329 6164 3331
rect 6536 3337 6577 3364
rect 6594 3337 6600 3763
rect 6536 3331 6600 3337
rect 6650 3763 7150 3769
rect 6650 3337 6656 3763
rect 6673 3715 7127 3763
rect 6673 3385 6735 3715
rect 7065 3385 7127 3715
rect 6673 3337 7127 3385
rect 7144 3337 7150 3763
rect 6650 3331 7150 3337
rect 7200 3763 7264 3769
rect 7200 3337 7206 3763
rect 7223 3736 7264 3763
rect 7636 3769 7669 3771
rect 7781 3794 8219 3800
rect 7781 3777 7787 3794
rect 8213 3777 8219 3794
rect 7781 3771 8219 3777
rect 7779 3769 8221 3771
rect 8331 3794 8769 3800
rect 8331 3777 8337 3794
rect 8763 3777 8769 3794
rect 8331 3771 8769 3777
rect 8331 3769 8364 3771
rect 7636 3763 7700 3769
rect 7636 3736 7677 3763
rect 7223 3364 7229 3736
rect 7671 3364 7677 3736
rect 7223 3337 7264 3364
rect 7200 3331 7264 3337
rect 6536 3329 6569 3331
rect 6131 3323 6569 3329
rect 6131 3306 6137 3323
rect 6563 3306 6569 3323
rect 6131 3300 6569 3306
rect 6679 3329 7121 3331
rect 6681 3323 7119 3329
rect 6681 3306 6687 3323
rect 7113 3306 7119 3323
rect 6681 3300 7119 3306
rect 7231 3329 7264 3331
rect 7636 3337 7677 3364
rect 7694 3337 7700 3763
rect 7636 3331 7700 3337
rect 7750 3763 8250 3769
rect 7750 3337 7756 3763
rect 7773 3715 8227 3763
rect 7773 3385 7835 3715
rect 8165 3385 8227 3715
rect 7773 3337 8227 3385
rect 8244 3337 8250 3763
rect 7750 3331 8250 3337
rect 8300 3763 8364 3769
rect 8300 3337 8306 3763
rect 8323 3736 8364 3763
rect 8736 3769 8769 3771
rect 8881 3794 9319 3800
rect 8881 3777 8887 3794
rect 9313 3777 9319 3794
rect 8881 3771 9319 3777
rect 8879 3769 9321 3771
rect 9431 3794 9869 3800
rect 9431 3777 9437 3794
rect 9863 3777 9869 3794
rect 9431 3771 9869 3777
rect 9431 3769 9464 3771
rect 8736 3763 8800 3769
rect 8736 3736 8777 3763
rect 8323 3364 8329 3736
rect 8771 3364 8777 3736
rect 8323 3337 8364 3364
rect 8300 3331 8364 3337
rect 7636 3329 7669 3331
rect 7231 3323 7669 3329
rect 7231 3306 7237 3323
rect 7663 3306 7669 3323
rect 7231 3300 7669 3306
rect 7779 3329 8221 3331
rect 7781 3323 8219 3329
rect 7781 3306 7787 3323
rect 8213 3306 8219 3323
rect 7781 3300 8219 3306
rect 8331 3329 8364 3331
rect 8736 3337 8777 3364
rect 8794 3337 8800 3763
rect 8736 3331 8800 3337
rect 8850 3763 9350 3769
rect 8850 3337 8856 3763
rect 8873 3715 9327 3763
rect 8873 3385 8935 3715
rect 9265 3385 9327 3715
rect 8873 3337 9327 3385
rect 9344 3337 9350 3763
rect 8850 3331 9350 3337
rect 9400 3763 9464 3769
rect 9400 3337 9406 3763
rect 9423 3736 9464 3763
rect 9836 3769 9869 3771
rect 9981 3794 10419 3800
rect 9981 3777 9987 3794
rect 10413 3777 10419 3794
rect 9981 3771 10419 3777
rect 9979 3769 10421 3771
rect 10531 3794 10969 3800
rect 10531 3777 10537 3794
rect 10963 3777 10969 3794
rect 10531 3771 10969 3777
rect 10531 3769 10564 3771
rect 9836 3763 9900 3769
rect 9836 3736 9877 3763
rect 9423 3364 9429 3736
rect 9871 3364 9877 3736
rect 9423 3337 9464 3364
rect 9400 3331 9464 3337
rect 8736 3329 8769 3331
rect 8331 3323 8769 3329
rect 8331 3306 8337 3323
rect 8763 3306 8769 3323
rect 8331 3300 8769 3306
rect 8879 3329 9321 3331
rect 8881 3323 9319 3329
rect 8881 3306 8887 3323
rect 9313 3306 9319 3323
rect 8881 3300 9319 3306
rect 9431 3329 9464 3331
rect 9836 3337 9877 3364
rect 9894 3337 9900 3763
rect 9836 3331 9900 3337
rect 9950 3763 10450 3769
rect 9950 3337 9956 3763
rect 9973 3715 10427 3763
rect 9973 3385 10035 3715
rect 10365 3385 10427 3715
rect 9973 3337 10427 3385
rect 10444 3337 10450 3763
rect 9950 3331 10450 3337
rect 10500 3763 10564 3769
rect 10500 3337 10506 3763
rect 10523 3736 10564 3763
rect 10936 3769 10969 3771
rect 11081 3794 11519 3800
rect 11081 3777 11087 3794
rect 11513 3777 11519 3794
rect 11081 3771 11519 3777
rect 11079 3769 11521 3771
rect 11631 3794 12069 3800
rect 11631 3777 11637 3794
rect 12063 3777 12069 3794
rect 11631 3771 12069 3777
rect 11631 3769 11664 3771
rect 10936 3763 11000 3769
rect 10936 3736 10977 3763
rect 10523 3364 10529 3736
rect 10971 3364 10977 3736
rect 10523 3337 10564 3364
rect 10500 3331 10564 3337
rect 9836 3329 9869 3331
rect 9431 3323 9869 3329
rect 9431 3306 9437 3323
rect 9863 3306 9869 3323
rect 9431 3300 9869 3306
rect 9979 3329 10421 3331
rect 9981 3323 10419 3329
rect 9981 3306 9987 3323
rect 10413 3306 10419 3323
rect 9981 3300 10419 3306
rect 10531 3329 10564 3331
rect 10936 3337 10977 3364
rect 10994 3337 11000 3763
rect 10936 3331 11000 3337
rect 11050 3763 11550 3769
rect 11050 3337 11056 3763
rect 11073 3715 11527 3763
rect 11073 3385 11135 3715
rect 11465 3385 11527 3715
rect 11073 3337 11527 3385
rect 11544 3337 11550 3763
rect 11050 3331 11550 3337
rect 11600 3763 11664 3769
rect 11600 3337 11606 3763
rect 11623 3736 11664 3763
rect 12036 3769 12069 3771
rect 12181 3794 12619 3800
rect 12181 3777 12187 3794
rect 12613 3777 12619 3794
rect 12181 3771 12619 3777
rect 12179 3769 12621 3771
rect 12731 3794 13169 3800
rect 12731 3777 12737 3794
rect 13163 3777 13169 3794
rect 12731 3771 13169 3777
rect 12731 3769 12764 3771
rect 12036 3763 12100 3769
rect 12036 3736 12077 3763
rect 11623 3364 11629 3736
rect 12071 3364 12077 3736
rect 11623 3337 11664 3364
rect 11600 3331 11664 3337
rect 10936 3329 10969 3331
rect 10531 3323 10969 3329
rect 10531 3306 10537 3323
rect 10963 3306 10969 3323
rect 10531 3300 10969 3306
rect 11079 3329 11521 3331
rect 11081 3323 11519 3329
rect 11081 3306 11087 3323
rect 11513 3306 11519 3323
rect 11081 3300 11519 3306
rect 11631 3329 11664 3331
rect 12036 3337 12077 3364
rect 12094 3337 12100 3763
rect 12036 3331 12100 3337
rect 12150 3763 12650 3769
rect 12150 3337 12156 3763
rect 12173 3715 12627 3763
rect 12173 3385 12235 3715
rect 12565 3385 12627 3715
rect 12173 3337 12627 3385
rect 12644 3337 12650 3763
rect 12150 3331 12650 3337
rect 12700 3763 12764 3769
rect 12700 3337 12706 3763
rect 12723 3736 12764 3763
rect 13136 3769 13169 3771
rect 13281 3794 13719 3800
rect 13281 3777 13287 3794
rect 13713 3777 13719 3794
rect 13281 3771 13719 3777
rect 13279 3769 13721 3771
rect 13136 3763 13200 3769
rect 13136 3736 13177 3763
rect 12723 3364 12729 3736
rect 13171 3364 13177 3736
rect 12723 3337 12764 3364
rect 12700 3331 12764 3337
rect 12036 3329 12069 3331
rect 11631 3323 12069 3329
rect 11631 3306 11637 3323
rect 12063 3306 12069 3323
rect 11631 3300 12069 3306
rect 12179 3329 12621 3331
rect 12181 3323 12619 3329
rect 12181 3306 12187 3323
rect 12613 3306 12619 3323
rect 12181 3300 12619 3306
rect 12731 3329 12764 3331
rect 13136 3337 13177 3364
rect 13194 3337 13200 3763
rect 13136 3331 13200 3337
rect 13250 3763 13721 3769
rect 13250 3337 13256 3763
rect 13273 3715 13721 3763
rect 13273 3385 13335 3715
rect 13665 3385 13721 3715
rect 13273 3337 13721 3385
rect 13250 3331 13721 3337
rect 13136 3329 13169 3331
rect 12731 3323 13169 3329
rect 12731 3306 12737 3323
rect 13163 3306 13169 3323
rect 12731 3300 13169 3306
rect 13279 3329 13721 3331
rect 13281 3323 13719 3329
rect 13281 3306 13287 3323
rect 13713 3306 13719 3323
rect 13281 3300 13719 3306
rect -469 3244 -31 3250
rect -469 3227 -463 3244
rect -37 3227 -31 3244
rect -469 3221 -31 3227
rect -471 3219 -29 3221
rect 81 3244 519 3250
rect 81 3227 87 3244
rect 513 3227 519 3244
rect 81 3221 519 3227
rect 81 3219 114 3221
rect -471 3213 0 3219
rect -471 3165 -23 3213
rect -471 2835 -415 3165
rect -85 2835 -23 3165
rect -471 2787 -23 2835
rect -6 2787 0 3213
rect -471 2781 0 2787
rect 50 3213 114 3219
rect 50 2787 56 3213
rect 73 3186 114 3213
rect 486 3219 519 3221
rect 631 3244 1069 3250
rect 631 3227 637 3244
rect 1063 3227 1069 3244
rect 631 3221 1069 3227
rect 629 3219 1071 3221
rect 1181 3244 1619 3250
rect 1181 3227 1187 3244
rect 1613 3227 1619 3244
rect 1181 3221 1619 3227
rect 1181 3219 1214 3221
rect 486 3213 550 3219
rect 486 3186 527 3213
rect 73 2814 79 3186
rect 521 2814 527 3186
rect 73 2787 114 2814
rect 50 2781 114 2787
rect -471 2779 -29 2781
rect -469 2773 -31 2779
rect -469 2756 -463 2773
rect -37 2756 -31 2773
rect -469 2750 -31 2756
rect 81 2779 114 2781
rect 486 2787 527 2814
rect 544 2787 550 3213
rect 486 2781 550 2787
rect 600 3213 1100 3219
rect 600 2787 606 3213
rect 623 3165 1077 3213
rect 623 2835 685 3165
rect 1015 2835 1077 3165
rect 623 2787 1077 2835
rect 1094 2787 1100 3213
rect 600 2781 1100 2787
rect 1150 3213 1214 3219
rect 1150 2787 1156 3213
rect 1173 3186 1214 3213
rect 1586 3219 1619 3221
rect 1731 3244 2169 3250
rect 1731 3227 1737 3244
rect 2163 3227 2169 3244
rect 1731 3221 2169 3227
rect 1729 3219 2171 3221
rect 2281 3244 2719 3250
rect 2281 3227 2287 3244
rect 2713 3227 2719 3244
rect 2281 3221 2719 3227
rect 2281 3219 2314 3221
rect 1586 3213 1650 3219
rect 1586 3186 1627 3213
rect 1173 2814 1179 3186
rect 1621 2814 1627 3186
rect 1173 2787 1214 2814
rect 1150 2781 1214 2787
rect 486 2779 519 2781
rect 81 2773 519 2779
rect 81 2756 87 2773
rect 513 2756 519 2773
rect 81 2750 519 2756
rect 629 2779 1071 2781
rect 631 2773 1069 2779
rect 631 2756 637 2773
rect 1063 2756 1069 2773
rect 631 2750 1069 2756
rect 1181 2779 1214 2781
rect 1586 2787 1627 2814
rect 1644 2787 1650 3213
rect 1586 2781 1650 2787
rect 1700 3213 2200 3219
rect 1700 2787 1706 3213
rect 1723 3165 2177 3213
rect 1723 2835 1785 3165
rect 2115 2835 2177 3165
rect 1723 2787 2177 2835
rect 2194 2787 2200 3213
rect 1700 2781 2200 2787
rect 2250 3213 2314 3219
rect 2250 2787 2256 3213
rect 2273 3186 2314 3213
rect 2686 3219 2719 3221
rect 2831 3244 3269 3250
rect 2831 3227 2837 3244
rect 3263 3227 3269 3244
rect 2831 3221 3269 3227
rect 2829 3219 3271 3221
rect 3381 3244 3819 3250
rect 3381 3227 3387 3244
rect 3813 3227 3819 3244
rect 3381 3221 3819 3227
rect 3381 3219 3414 3221
rect 2686 3213 2750 3219
rect 2686 3186 2727 3213
rect 2273 2814 2279 3186
rect 2721 2814 2727 3186
rect 2273 2787 2314 2814
rect 2250 2781 2314 2787
rect 1586 2779 1619 2781
rect 1181 2773 1619 2779
rect 1181 2756 1187 2773
rect 1613 2756 1619 2773
rect 1181 2750 1619 2756
rect 1729 2779 2171 2781
rect 1731 2773 2169 2779
rect 1731 2756 1737 2773
rect 2163 2756 2169 2773
rect 1731 2750 2169 2756
rect 2281 2779 2314 2781
rect 2686 2787 2727 2814
rect 2744 2787 2750 3213
rect 2686 2781 2750 2787
rect 2800 3213 3300 3219
rect 2800 2787 2806 3213
rect 2823 3165 3277 3213
rect 2823 2835 2885 3165
rect 3215 2835 3277 3165
rect 2823 2787 3277 2835
rect 3294 2787 3300 3213
rect 2800 2781 3300 2787
rect 3350 3213 3414 3219
rect 3350 2787 3356 3213
rect 3373 3186 3414 3213
rect 3786 3219 3819 3221
rect 3931 3244 4369 3250
rect 3931 3227 3937 3244
rect 4363 3227 4369 3244
rect 3931 3221 4369 3227
rect 3929 3219 4371 3221
rect 4481 3244 4919 3250
rect 4481 3227 4487 3244
rect 4913 3227 4919 3244
rect 4481 3221 4919 3227
rect 4481 3219 4514 3221
rect 3786 3213 3850 3219
rect 3786 3186 3827 3213
rect 3373 2814 3379 3186
rect 3821 2814 3827 3186
rect 3373 2787 3414 2814
rect 3350 2781 3414 2787
rect 2686 2779 2719 2781
rect 2281 2773 2719 2779
rect 2281 2756 2287 2773
rect 2713 2756 2719 2773
rect 2281 2750 2719 2756
rect 2829 2779 3271 2781
rect 2831 2773 3269 2779
rect 2831 2756 2837 2773
rect 3263 2756 3269 2773
rect 2831 2750 3269 2756
rect 3381 2779 3414 2781
rect 3786 2787 3827 2814
rect 3844 2787 3850 3213
rect 3786 2781 3850 2787
rect 3900 3213 4400 3219
rect 3900 2787 3906 3213
rect 3923 3165 4377 3213
rect 3923 2835 3985 3165
rect 4315 2835 4377 3165
rect 3923 2787 4377 2835
rect 4394 2787 4400 3213
rect 3900 2781 4400 2787
rect 4450 3213 4514 3219
rect 4450 2787 4456 3213
rect 4473 3186 4514 3213
rect 4886 3219 4919 3221
rect 5031 3244 5469 3250
rect 5031 3227 5037 3244
rect 5463 3227 5469 3244
rect 5031 3221 5469 3227
rect 5029 3219 5471 3221
rect 5581 3244 6019 3250
rect 5581 3227 5587 3244
rect 6013 3227 6019 3244
rect 5581 3221 6019 3227
rect 5581 3219 5614 3221
rect 4886 3213 4950 3219
rect 4886 3186 4927 3213
rect 4473 2814 4479 3186
rect 4921 2814 4927 3186
rect 4473 2787 4514 2814
rect 4450 2781 4514 2787
rect 3786 2779 3819 2781
rect 3381 2773 3819 2779
rect 3381 2756 3387 2773
rect 3813 2756 3819 2773
rect 3381 2750 3819 2756
rect 3929 2779 4371 2781
rect 3931 2773 4369 2779
rect 3931 2756 3937 2773
rect 4363 2756 4369 2773
rect 3931 2750 4369 2756
rect 4481 2779 4514 2781
rect 4886 2787 4927 2814
rect 4944 2787 4950 3213
rect 4886 2781 4950 2787
rect 5000 3213 5500 3219
rect 5000 2787 5006 3213
rect 5023 3165 5477 3213
rect 5023 2835 5085 3165
rect 5415 2835 5477 3165
rect 5023 2787 5477 2835
rect 5494 2787 5500 3213
rect 5000 2781 5500 2787
rect 5550 3213 5614 3219
rect 5550 2787 5556 3213
rect 5573 3186 5614 3213
rect 5986 3219 6019 3221
rect 6131 3244 6569 3250
rect 6131 3227 6137 3244
rect 6563 3227 6569 3244
rect 6131 3221 6569 3227
rect 6129 3219 6571 3221
rect 6681 3244 7119 3250
rect 6681 3227 6687 3244
rect 7113 3227 7119 3244
rect 6681 3221 7119 3227
rect 6681 3219 6714 3221
rect 5986 3213 6050 3219
rect 5986 3186 6027 3213
rect 5573 2814 5579 3186
rect 6021 2814 6027 3186
rect 5573 2787 5614 2814
rect 5550 2781 5614 2787
rect 4886 2779 4919 2781
rect 4481 2773 4919 2779
rect 4481 2756 4487 2773
rect 4913 2756 4919 2773
rect 4481 2750 4919 2756
rect 5029 2779 5471 2781
rect 5031 2773 5469 2779
rect 5031 2756 5037 2773
rect 5463 2756 5469 2773
rect 5031 2750 5469 2756
rect 5581 2779 5614 2781
rect 5986 2787 6027 2814
rect 6044 2787 6050 3213
rect 5986 2781 6050 2787
rect 6100 3213 6600 3219
rect 6100 2787 6106 3213
rect 6123 3165 6577 3213
rect 6123 2835 6185 3165
rect 6515 2835 6577 3165
rect 6123 2787 6577 2835
rect 6594 2787 6600 3213
rect 6100 2781 6600 2787
rect 6650 3213 6714 3219
rect 6650 2787 6656 3213
rect 6673 3186 6714 3213
rect 7086 3219 7119 3221
rect 7231 3244 7669 3250
rect 7231 3227 7237 3244
rect 7663 3227 7669 3244
rect 7231 3221 7669 3227
rect 7229 3219 7671 3221
rect 7781 3244 8219 3250
rect 7781 3227 7787 3244
rect 8213 3227 8219 3244
rect 7781 3221 8219 3227
rect 7781 3219 7814 3221
rect 7086 3213 7150 3219
rect 7086 3186 7127 3213
rect 6673 2814 6679 3186
rect 7121 2814 7127 3186
rect 6673 2787 6714 2814
rect 6650 2781 6714 2787
rect 5986 2779 6019 2781
rect 5581 2773 6019 2779
rect 5581 2756 5587 2773
rect 6013 2756 6019 2773
rect 5581 2750 6019 2756
rect 6129 2779 6571 2781
rect 6131 2773 6569 2779
rect 6131 2756 6137 2773
rect 6563 2756 6569 2773
rect 6131 2750 6569 2756
rect 6681 2779 6714 2781
rect 7086 2787 7127 2814
rect 7144 2787 7150 3213
rect 7086 2781 7150 2787
rect 7200 3213 7700 3219
rect 7200 2787 7206 3213
rect 7223 3165 7677 3213
rect 7223 2835 7285 3165
rect 7615 2835 7677 3165
rect 7223 2787 7677 2835
rect 7694 2787 7700 3213
rect 7200 2781 7700 2787
rect 7750 3213 7814 3219
rect 7750 2787 7756 3213
rect 7773 3186 7814 3213
rect 8186 3219 8219 3221
rect 8331 3244 8769 3250
rect 8331 3227 8337 3244
rect 8763 3227 8769 3244
rect 8331 3221 8769 3227
rect 8329 3219 8771 3221
rect 8881 3244 9319 3250
rect 8881 3227 8887 3244
rect 9313 3227 9319 3244
rect 8881 3221 9319 3227
rect 8881 3219 8914 3221
rect 8186 3213 8250 3219
rect 8186 3186 8227 3213
rect 7773 2814 7779 3186
rect 8221 2814 8227 3186
rect 7773 2787 7814 2814
rect 7750 2781 7814 2787
rect 7086 2779 7119 2781
rect 6681 2773 7119 2779
rect 6681 2756 6687 2773
rect 7113 2756 7119 2773
rect 6681 2750 7119 2756
rect 7229 2779 7671 2781
rect 7231 2773 7669 2779
rect 7231 2756 7237 2773
rect 7663 2756 7669 2773
rect 7231 2750 7669 2756
rect 7781 2779 7814 2781
rect 8186 2787 8227 2814
rect 8244 2787 8250 3213
rect 8186 2781 8250 2787
rect 8300 3213 8800 3219
rect 8300 2787 8306 3213
rect 8323 3165 8777 3213
rect 8323 2835 8385 3165
rect 8715 2835 8777 3165
rect 8323 2787 8777 2835
rect 8794 2787 8800 3213
rect 8300 2781 8800 2787
rect 8850 3213 8914 3219
rect 8850 2787 8856 3213
rect 8873 3186 8914 3213
rect 9286 3219 9319 3221
rect 9431 3244 9869 3250
rect 9431 3227 9437 3244
rect 9863 3227 9869 3244
rect 9431 3221 9869 3227
rect 9429 3219 9871 3221
rect 9981 3244 10419 3250
rect 9981 3227 9987 3244
rect 10413 3227 10419 3244
rect 9981 3221 10419 3227
rect 9981 3219 10014 3221
rect 9286 3213 9350 3219
rect 9286 3186 9327 3213
rect 8873 2814 8879 3186
rect 9321 2814 9327 3186
rect 8873 2787 8914 2814
rect 8850 2781 8914 2787
rect 8186 2779 8219 2781
rect 7781 2773 8219 2779
rect 7781 2756 7787 2773
rect 8213 2756 8219 2773
rect 7781 2750 8219 2756
rect 8329 2779 8771 2781
rect 8331 2773 8769 2779
rect 8331 2756 8337 2773
rect 8763 2756 8769 2773
rect 8331 2750 8769 2756
rect 8881 2779 8914 2781
rect 9286 2787 9327 2814
rect 9344 2787 9350 3213
rect 9286 2781 9350 2787
rect 9400 3213 9900 3219
rect 9400 2787 9406 3213
rect 9423 3165 9877 3213
rect 9423 2835 9485 3165
rect 9815 2835 9877 3165
rect 9423 2787 9877 2835
rect 9894 2787 9900 3213
rect 9400 2781 9900 2787
rect 9950 3213 10014 3219
rect 9950 2787 9956 3213
rect 9973 3186 10014 3213
rect 10386 3219 10419 3221
rect 10531 3244 10969 3250
rect 10531 3227 10537 3244
rect 10963 3227 10969 3244
rect 10531 3221 10969 3227
rect 10529 3219 10971 3221
rect 11081 3244 11519 3250
rect 11081 3227 11087 3244
rect 11513 3227 11519 3244
rect 11081 3221 11519 3227
rect 11081 3219 11114 3221
rect 10386 3213 10450 3219
rect 10386 3186 10427 3213
rect 9973 2814 9979 3186
rect 10421 2814 10427 3186
rect 9973 2787 10014 2814
rect 9950 2781 10014 2787
rect 9286 2779 9319 2781
rect 8881 2773 9319 2779
rect 8881 2756 8887 2773
rect 9313 2756 9319 2773
rect 8881 2750 9319 2756
rect 9429 2779 9871 2781
rect 9431 2773 9869 2779
rect 9431 2756 9437 2773
rect 9863 2756 9869 2773
rect 9431 2750 9869 2756
rect 9981 2779 10014 2781
rect 10386 2787 10427 2814
rect 10444 2787 10450 3213
rect 10386 2781 10450 2787
rect 10500 3213 11000 3219
rect 10500 2787 10506 3213
rect 10523 3165 10977 3213
rect 10523 2835 10585 3165
rect 10915 2835 10977 3165
rect 10523 2787 10977 2835
rect 10994 2787 11000 3213
rect 10500 2781 11000 2787
rect 11050 3213 11114 3219
rect 11050 2787 11056 3213
rect 11073 3186 11114 3213
rect 11486 3219 11519 3221
rect 11631 3244 12069 3250
rect 11631 3227 11637 3244
rect 12063 3227 12069 3244
rect 11631 3221 12069 3227
rect 11629 3219 12071 3221
rect 12181 3244 12619 3250
rect 12181 3227 12187 3244
rect 12613 3227 12619 3244
rect 12181 3221 12619 3227
rect 12181 3219 12214 3221
rect 11486 3213 11550 3219
rect 11486 3186 11527 3213
rect 11073 2814 11079 3186
rect 11521 2814 11527 3186
rect 11073 2787 11114 2814
rect 11050 2781 11114 2787
rect 10386 2779 10419 2781
rect 9981 2773 10419 2779
rect 9981 2756 9987 2773
rect 10413 2756 10419 2773
rect 9981 2750 10419 2756
rect 10529 2779 10971 2781
rect 10531 2773 10969 2779
rect 10531 2756 10537 2773
rect 10963 2756 10969 2773
rect 10531 2750 10969 2756
rect 11081 2779 11114 2781
rect 11486 2787 11527 2814
rect 11544 2787 11550 3213
rect 11486 2781 11550 2787
rect 11600 3213 12100 3219
rect 11600 2787 11606 3213
rect 11623 3165 12077 3213
rect 11623 2835 11685 3165
rect 12015 2835 12077 3165
rect 11623 2787 12077 2835
rect 12094 2787 12100 3213
rect 11600 2781 12100 2787
rect 12150 3213 12214 3219
rect 12150 2787 12156 3213
rect 12173 3186 12214 3213
rect 12586 3219 12619 3221
rect 12731 3244 13169 3250
rect 12731 3227 12737 3244
rect 13163 3227 13169 3244
rect 12731 3221 13169 3227
rect 12729 3219 13171 3221
rect 13281 3244 13719 3250
rect 13281 3227 13287 3244
rect 13713 3227 13719 3244
rect 13281 3221 13719 3227
rect 13281 3219 13314 3221
rect 12586 3213 12650 3219
rect 12586 3186 12627 3213
rect 12173 2814 12179 3186
rect 12621 2814 12627 3186
rect 12173 2787 12214 2814
rect 12150 2781 12214 2787
rect 11486 2779 11519 2781
rect 11081 2773 11519 2779
rect 11081 2756 11087 2773
rect 11513 2756 11519 2773
rect 11081 2750 11519 2756
rect 11629 2779 12071 2781
rect 11631 2773 12069 2779
rect 11631 2756 11637 2773
rect 12063 2756 12069 2773
rect 11631 2750 12069 2756
rect 12181 2779 12214 2781
rect 12586 2787 12627 2814
rect 12644 2787 12650 3213
rect 12586 2781 12650 2787
rect 12700 3213 13200 3219
rect 12700 2787 12706 3213
rect 12723 3165 13177 3213
rect 12723 2835 12785 3165
rect 13115 2835 13177 3165
rect 12723 2787 13177 2835
rect 13194 2787 13200 3213
rect 12700 2781 13200 2787
rect 13250 3213 13314 3219
rect 13250 2787 13256 3213
rect 13273 3186 13314 3213
rect 13273 2814 13279 3186
rect 13273 2787 13314 2814
rect 13250 2781 13314 2787
rect 12586 2779 12619 2781
rect 12181 2773 12619 2779
rect 12181 2756 12187 2773
rect 12613 2756 12619 2773
rect 12181 2750 12619 2756
rect 12729 2779 13171 2781
rect 12731 2773 13169 2779
rect 12731 2756 12737 2773
rect 13163 2756 13169 2773
rect 12731 2750 13169 2756
rect 13281 2779 13314 2781
rect 13281 2773 13719 2779
rect 13281 2756 13287 2773
rect 13713 2756 13719 2773
rect 13281 2750 13719 2756
rect -469 2694 -31 2700
rect -469 2677 -463 2694
rect -37 2677 -31 2694
rect -469 2671 -31 2677
rect -64 2669 -31 2671
rect 81 2694 519 2700
rect 81 2677 87 2694
rect 513 2677 519 2694
rect 81 2671 519 2677
rect 79 2669 521 2671
rect 631 2694 1069 2700
rect 631 2677 637 2694
rect 1063 2677 1069 2694
rect 631 2671 1069 2677
rect 631 2669 664 2671
rect -64 2663 0 2669
rect -64 2636 -23 2663
rect -29 2264 -23 2636
rect -64 2237 -23 2264
rect -6 2237 0 2663
rect -64 2231 0 2237
rect 50 2663 550 2669
rect 50 2237 56 2663
rect 73 2615 527 2663
rect 73 2285 135 2615
rect 465 2285 527 2615
rect 73 2237 527 2285
rect 544 2237 550 2663
rect 50 2231 550 2237
rect 600 2663 664 2669
rect 600 2237 606 2663
rect 623 2636 664 2663
rect 1036 2669 1069 2671
rect 1181 2694 1619 2700
rect 1181 2677 1187 2694
rect 1613 2677 1619 2694
rect 1181 2671 1619 2677
rect 1179 2669 1621 2671
rect 1731 2694 2169 2700
rect 1731 2677 1737 2694
rect 2163 2677 2169 2694
rect 1731 2671 2169 2677
rect 1731 2669 1764 2671
rect 1036 2663 1100 2669
rect 1036 2636 1077 2663
rect 623 2264 629 2636
rect 1071 2264 1077 2636
rect 623 2237 664 2264
rect 600 2231 664 2237
rect -64 2229 -31 2231
rect -469 2223 -31 2229
rect -469 2206 -463 2223
rect -37 2206 -31 2223
rect -469 2200 -31 2206
rect 79 2229 521 2231
rect 81 2223 519 2229
rect 81 2206 87 2223
rect 513 2206 519 2223
rect 81 2200 519 2206
rect 631 2229 664 2231
rect 1036 2237 1077 2264
rect 1094 2237 1100 2663
rect 1036 2231 1100 2237
rect 1150 2663 1650 2669
rect 1150 2237 1156 2663
rect 1173 2615 1627 2663
rect 1173 2285 1235 2615
rect 1565 2285 1627 2615
rect 1173 2237 1627 2285
rect 1644 2237 1650 2663
rect 1150 2231 1650 2237
rect 1700 2663 1764 2669
rect 1700 2237 1706 2663
rect 1723 2636 1764 2663
rect 2136 2669 2169 2671
rect 2281 2694 2719 2700
rect 2281 2677 2287 2694
rect 2713 2677 2719 2694
rect 2281 2671 2719 2677
rect 2279 2669 2721 2671
rect 2831 2694 3269 2700
rect 2831 2677 2837 2694
rect 3263 2677 3269 2694
rect 2831 2671 3269 2677
rect 2831 2669 2864 2671
rect 2136 2663 2200 2669
rect 2136 2636 2177 2663
rect 1723 2264 1729 2636
rect 2171 2264 2177 2636
rect 1723 2237 1764 2264
rect 1700 2231 1764 2237
rect 1036 2229 1069 2231
rect 631 2223 1069 2229
rect 631 2206 637 2223
rect 1063 2206 1069 2223
rect 631 2200 1069 2206
rect 1179 2229 1621 2231
rect 1181 2223 1619 2229
rect 1181 2206 1187 2223
rect 1613 2206 1619 2223
rect 1181 2200 1619 2206
rect 1731 2229 1764 2231
rect 2136 2237 2177 2264
rect 2194 2237 2200 2663
rect 2136 2231 2200 2237
rect 2250 2663 2750 2669
rect 2250 2237 2256 2663
rect 2273 2615 2727 2663
rect 2273 2285 2335 2615
rect 2665 2285 2727 2615
rect 2273 2237 2727 2285
rect 2744 2237 2750 2663
rect 2250 2231 2750 2237
rect 2800 2663 2864 2669
rect 2800 2237 2806 2663
rect 2823 2636 2864 2663
rect 3236 2669 3269 2671
rect 3381 2694 3819 2700
rect 3381 2677 3387 2694
rect 3813 2677 3819 2694
rect 3381 2671 3819 2677
rect 3379 2669 3821 2671
rect 3931 2694 4369 2700
rect 3931 2677 3937 2694
rect 4363 2677 4369 2694
rect 3931 2671 4369 2677
rect 3931 2669 3964 2671
rect 3236 2663 3300 2669
rect 3236 2636 3277 2663
rect 2823 2264 2829 2636
rect 3271 2264 3277 2636
rect 2823 2237 2864 2264
rect 2800 2231 2864 2237
rect 2136 2229 2169 2231
rect 1731 2223 2169 2229
rect 1731 2206 1737 2223
rect 2163 2206 2169 2223
rect 1731 2200 2169 2206
rect 2279 2229 2721 2231
rect 2281 2223 2719 2229
rect 2281 2206 2287 2223
rect 2713 2206 2719 2223
rect 2281 2200 2719 2206
rect 2831 2229 2864 2231
rect 3236 2237 3277 2264
rect 3294 2237 3300 2663
rect 3236 2231 3300 2237
rect 3350 2663 3850 2669
rect 3350 2237 3356 2663
rect 3373 2615 3827 2663
rect 3373 2285 3435 2615
rect 3765 2285 3827 2615
rect 3373 2237 3827 2285
rect 3844 2237 3850 2663
rect 3350 2231 3850 2237
rect 3900 2663 3964 2669
rect 3900 2237 3906 2663
rect 3923 2636 3964 2663
rect 4336 2669 4369 2671
rect 4481 2694 4919 2700
rect 4481 2677 4487 2694
rect 4913 2677 4919 2694
rect 4481 2671 4919 2677
rect 4479 2669 4921 2671
rect 5031 2694 5469 2700
rect 5031 2677 5037 2694
rect 5463 2677 5469 2694
rect 5031 2671 5469 2677
rect 5031 2669 5064 2671
rect 4336 2663 4400 2669
rect 4336 2636 4377 2663
rect 3923 2264 3929 2636
rect 4371 2264 4377 2636
rect 3923 2237 3964 2264
rect 3900 2231 3964 2237
rect 3236 2229 3269 2231
rect 2831 2223 3269 2229
rect 2831 2206 2837 2223
rect 3263 2206 3269 2223
rect 2831 2200 3269 2206
rect 3379 2229 3821 2231
rect 3381 2223 3819 2229
rect 3381 2206 3387 2223
rect 3813 2206 3819 2223
rect 3381 2200 3819 2206
rect 3931 2229 3964 2231
rect 4336 2237 4377 2264
rect 4394 2237 4400 2663
rect 4336 2231 4400 2237
rect 4450 2663 4950 2669
rect 4450 2237 4456 2663
rect 4473 2615 4927 2663
rect 4473 2285 4535 2615
rect 4865 2285 4927 2615
rect 4473 2237 4927 2285
rect 4944 2237 4950 2663
rect 4450 2231 4950 2237
rect 5000 2663 5064 2669
rect 5000 2237 5006 2663
rect 5023 2636 5064 2663
rect 5436 2669 5469 2671
rect 5581 2694 6019 2700
rect 5581 2677 5587 2694
rect 6013 2677 6019 2694
rect 5581 2671 6019 2677
rect 5579 2669 6021 2671
rect 6131 2694 6569 2700
rect 6131 2677 6137 2694
rect 6563 2677 6569 2694
rect 6131 2671 6569 2677
rect 6131 2669 6164 2671
rect 5436 2663 5500 2669
rect 5436 2636 5477 2663
rect 5023 2264 5029 2636
rect 5471 2264 5477 2636
rect 5023 2237 5064 2264
rect 5000 2231 5064 2237
rect 4336 2229 4369 2231
rect 3931 2223 4369 2229
rect 3931 2206 3937 2223
rect 4363 2206 4369 2223
rect 3931 2200 4369 2206
rect 4479 2229 4921 2231
rect 4481 2223 4919 2229
rect 4481 2206 4487 2223
rect 4913 2206 4919 2223
rect 4481 2200 4919 2206
rect 5031 2229 5064 2231
rect 5436 2237 5477 2264
rect 5494 2237 5500 2663
rect 5436 2231 5500 2237
rect 5550 2663 6050 2669
rect 5550 2237 5556 2663
rect 5573 2615 6027 2663
rect 5573 2285 5635 2615
rect 5965 2285 6027 2615
rect 5573 2237 6027 2285
rect 6044 2237 6050 2663
rect 5550 2231 6050 2237
rect 6100 2663 6164 2669
rect 6100 2237 6106 2663
rect 6123 2636 6164 2663
rect 6536 2669 6569 2671
rect 6681 2694 7119 2700
rect 6681 2677 6687 2694
rect 7113 2677 7119 2694
rect 6681 2671 7119 2677
rect 6679 2669 7121 2671
rect 7231 2694 7669 2700
rect 7231 2677 7237 2694
rect 7663 2677 7669 2694
rect 7231 2671 7669 2677
rect 7231 2669 7264 2671
rect 6536 2663 6600 2669
rect 6536 2636 6577 2663
rect 6123 2264 6129 2636
rect 6571 2264 6577 2636
rect 6123 2237 6164 2264
rect 6100 2231 6164 2237
rect 5436 2229 5469 2231
rect 5031 2223 5469 2229
rect 5031 2206 5037 2223
rect 5463 2206 5469 2223
rect 5031 2200 5469 2206
rect 5579 2229 6021 2231
rect 5581 2223 6019 2229
rect 5581 2206 5587 2223
rect 6013 2206 6019 2223
rect 5581 2200 6019 2206
rect 6131 2229 6164 2231
rect 6536 2237 6577 2264
rect 6594 2237 6600 2663
rect 6536 2231 6600 2237
rect 6650 2663 7150 2669
rect 6650 2237 6656 2663
rect 6673 2615 7127 2663
rect 6673 2285 6735 2615
rect 7065 2285 7127 2615
rect 6673 2237 7127 2285
rect 7144 2237 7150 2663
rect 6650 2231 7150 2237
rect 7200 2663 7264 2669
rect 7200 2237 7206 2663
rect 7223 2636 7264 2663
rect 7636 2669 7669 2671
rect 7781 2694 8219 2700
rect 7781 2677 7787 2694
rect 8213 2677 8219 2694
rect 7781 2671 8219 2677
rect 7779 2669 8221 2671
rect 8331 2694 8769 2700
rect 8331 2677 8337 2694
rect 8763 2677 8769 2694
rect 8331 2671 8769 2677
rect 8331 2669 8364 2671
rect 7636 2663 7700 2669
rect 7636 2636 7677 2663
rect 7223 2264 7229 2636
rect 7671 2264 7677 2636
rect 7223 2237 7264 2264
rect 7200 2231 7264 2237
rect 6536 2229 6569 2231
rect 6131 2223 6569 2229
rect 6131 2206 6137 2223
rect 6563 2206 6569 2223
rect 6131 2200 6569 2206
rect 6679 2229 7121 2231
rect 6681 2223 7119 2229
rect 6681 2206 6687 2223
rect 7113 2206 7119 2223
rect 6681 2200 7119 2206
rect 7231 2229 7264 2231
rect 7636 2237 7677 2264
rect 7694 2237 7700 2663
rect 7636 2231 7700 2237
rect 7750 2663 8250 2669
rect 7750 2237 7756 2663
rect 7773 2615 8227 2663
rect 7773 2285 7835 2615
rect 8165 2285 8227 2615
rect 7773 2237 8227 2285
rect 8244 2237 8250 2663
rect 7750 2231 8250 2237
rect 8300 2663 8364 2669
rect 8300 2237 8306 2663
rect 8323 2636 8364 2663
rect 8736 2669 8769 2671
rect 8881 2694 9319 2700
rect 8881 2677 8887 2694
rect 9313 2677 9319 2694
rect 8881 2671 9319 2677
rect 8879 2669 9321 2671
rect 9431 2694 9869 2700
rect 9431 2677 9437 2694
rect 9863 2677 9869 2694
rect 9431 2671 9869 2677
rect 9431 2669 9464 2671
rect 8736 2663 8800 2669
rect 8736 2636 8777 2663
rect 8323 2264 8329 2636
rect 8771 2264 8777 2636
rect 8323 2237 8364 2264
rect 8300 2231 8364 2237
rect 7636 2229 7669 2231
rect 7231 2223 7669 2229
rect 7231 2206 7237 2223
rect 7663 2206 7669 2223
rect 7231 2200 7669 2206
rect 7779 2229 8221 2231
rect 7781 2223 8219 2229
rect 7781 2206 7787 2223
rect 8213 2206 8219 2223
rect 7781 2200 8219 2206
rect 8331 2229 8364 2231
rect 8736 2237 8777 2264
rect 8794 2237 8800 2663
rect 8736 2231 8800 2237
rect 8850 2663 9350 2669
rect 8850 2237 8856 2663
rect 8873 2615 9327 2663
rect 8873 2285 8935 2615
rect 9265 2285 9327 2615
rect 8873 2237 9327 2285
rect 9344 2237 9350 2663
rect 8850 2231 9350 2237
rect 9400 2663 9464 2669
rect 9400 2237 9406 2663
rect 9423 2636 9464 2663
rect 9836 2669 9869 2671
rect 9981 2694 10419 2700
rect 9981 2677 9987 2694
rect 10413 2677 10419 2694
rect 9981 2671 10419 2677
rect 9979 2669 10421 2671
rect 10531 2694 10969 2700
rect 10531 2677 10537 2694
rect 10963 2677 10969 2694
rect 10531 2671 10969 2677
rect 10531 2669 10564 2671
rect 9836 2663 9900 2669
rect 9836 2636 9877 2663
rect 9423 2264 9429 2636
rect 9871 2264 9877 2636
rect 9423 2237 9464 2264
rect 9400 2231 9464 2237
rect 8736 2229 8769 2231
rect 8331 2223 8769 2229
rect 8331 2206 8337 2223
rect 8763 2206 8769 2223
rect 8331 2200 8769 2206
rect 8879 2229 9321 2231
rect 8881 2223 9319 2229
rect 8881 2206 8887 2223
rect 9313 2206 9319 2223
rect 8881 2200 9319 2206
rect 9431 2229 9464 2231
rect 9836 2237 9877 2264
rect 9894 2237 9900 2663
rect 9836 2231 9900 2237
rect 9950 2663 10450 2669
rect 9950 2237 9956 2663
rect 9973 2615 10427 2663
rect 9973 2285 10035 2615
rect 10365 2285 10427 2615
rect 9973 2237 10427 2285
rect 10444 2237 10450 2663
rect 9950 2231 10450 2237
rect 10500 2663 10564 2669
rect 10500 2237 10506 2663
rect 10523 2636 10564 2663
rect 10936 2669 10969 2671
rect 11081 2694 11519 2700
rect 11081 2677 11087 2694
rect 11513 2677 11519 2694
rect 11081 2671 11519 2677
rect 11079 2669 11521 2671
rect 11631 2694 12069 2700
rect 11631 2677 11637 2694
rect 12063 2677 12069 2694
rect 11631 2671 12069 2677
rect 11631 2669 11664 2671
rect 10936 2663 11000 2669
rect 10936 2636 10977 2663
rect 10523 2264 10529 2636
rect 10971 2264 10977 2636
rect 10523 2237 10564 2264
rect 10500 2231 10564 2237
rect 9836 2229 9869 2231
rect 9431 2223 9869 2229
rect 9431 2206 9437 2223
rect 9863 2206 9869 2223
rect 9431 2200 9869 2206
rect 9979 2229 10421 2231
rect 9981 2223 10419 2229
rect 9981 2206 9987 2223
rect 10413 2206 10419 2223
rect 9981 2200 10419 2206
rect 10531 2229 10564 2231
rect 10936 2237 10977 2264
rect 10994 2237 11000 2663
rect 10936 2231 11000 2237
rect 11050 2663 11550 2669
rect 11050 2237 11056 2663
rect 11073 2615 11527 2663
rect 11073 2285 11135 2615
rect 11465 2285 11527 2615
rect 11073 2237 11527 2285
rect 11544 2237 11550 2663
rect 11050 2231 11550 2237
rect 11600 2663 11664 2669
rect 11600 2237 11606 2663
rect 11623 2636 11664 2663
rect 12036 2669 12069 2671
rect 12181 2694 12619 2700
rect 12181 2677 12187 2694
rect 12613 2677 12619 2694
rect 12181 2671 12619 2677
rect 12179 2669 12621 2671
rect 12731 2694 13169 2700
rect 12731 2677 12737 2694
rect 13163 2677 13169 2694
rect 12731 2671 13169 2677
rect 12731 2669 12764 2671
rect 12036 2663 12100 2669
rect 12036 2636 12077 2663
rect 11623 2264 11629 2636
rect 12071 2264 12077 2636
rect 11623 2237 11664 2264
rect 11600 2231 11664 2237
rect 10936 2229 10969 2231
rect 10531 2223 10969 2229
rect 10531 2206 10537 2223
rect 10963 2206 10969 2223
rect 10531 2200 10969 2206
rect 11079 2229 11521 2231
rect 11081 2223 11519 2229
rect 11081 2206 11087 2223
rect 11513 2206 11519 2223
rect 11081 2200 11519 2206
rect 11631 2229 11664 2231
rect 12036 2237 12077 2264
rect 12094 2237 12100 2663
rect 12036 2231 12100 2237
rect 12150 2663 12650 2669
rect 12150 2237 12156 2663
rect 12173 2615 12627 2663
rect 12173 2285 12235 2615
rect 12565 2285 12627 2615
rect 12173 2237 12627 2285
rect 12644 2237 12650 2663
rect 12150 2231 12650 2237
rect 12700 2663 12764 2669
rect 12700 2237 12706 2663
rect 12723 2636 12764 2663
rect 13136 2669 13169 2671
rect 13281 2694 13719 2700
rect 13281 2677 13287 2694
rect 13713 2677 13719 2694
rect 13281 2671 13719 2677
rect 13279 2669 13721 2671
rect 13136 2663 13200 2669
rect 13136 2636 13177 2663
rect 12723 2264 12729 2636
rect 13171 2264 13177 2636
rect 12723 2237 12764 2264
rect 12700 2231 12764 2237
rect 12036 2229 12069 2231
rect 11631 2223 12069 2229
rect 11631 2206 11637 2223
rect 12063 2206 12069 2223
rect 11631 2200 12069 2206
rect 12179 2229 12621 2231
rect 12181 2223 12619 2229
rect 12181 2206 12187 2223
rect 12613 2206 12619 2223
rect 12181 2200 12619 2206
rect 12731 2229 12764 2231
rect 13136 2237 13177 2264
rect 13194 2237 13200 2663
rect 13136 2231 13200 2237
rect 13250 2663 13721 2669
rect 13250 2237 13256 2663
rect 13273 2615 13721 2663
rect 13273 2285 13335 2615
rect 13665 2285 13721 2615
rect 13273 2237 13721 2285
rect 13250 2231 13721 2237
rect 13136 2229 13169 2231
rect 12731 2223 13169 2229
rect 12731 2206 12737 2223
rect 13163 2206 13169 2223
rect 12731 2200 13169 2206
rect 13279 2229 13721 2231
rect 13281 2223 13719 2229
rect 13281 2206 13287 2223
rect 13713 2206 13719 2223
rect 13281 2200 13719 2206
rect -469 2144 -31 2150
rect -469 2127 -463 2144
rect -37 2127 -31 2144
rect -469 2121 -31 2127
rect -471 2119 -29 2121
rect 81 2144 519 2150
rect 81 2127 87 2144
rect 513 2127 519 2144
rect 81 2121 519 2127
rect 81 2119 114 2121
rect -471 2113 0 2119
rect -471 2065 -23 2113
rect -471 1735 -415 2065
rect -85 1735 -23 2065
rect -471 1687 -23 1735
rect -6 1687 0 2113
rect -471 1681 0 1687
rect 50 2113 114 2119
rect 50 1687 56 2113
rect 73 2086 114 2113
rect 486 2119 519 2121
rect 631 2144 1069 2150
rect 631 2127 637 2144
rect 1063 2127 1069 2144
rect 631 2121 1069 2127
rect 629 2119 1071 2121
rect 1181 2144 1619 2150
rect 1181 2127 1187 2144
rect 1613 2127 1619 2144
rect 1181 2121 1619 2127
rect 1181 2119 1214 2121
rect 486 2113 550 2119
rect 486 2086 527 2113
rect 73 1714 79 2086
rect 521 1714 527 2086
rect 73 1687 114 1714
rect 50 1681 114 1687
rect -471 1679 -29 1681
rect -469 1673 -31 1679
rect -469 1656 -463 1673
rect -37 1656 -31 1673
rect -469 1650 -31 1656
rect 81 1679 114 1681
rect 486 1687 527 1714
rect 544 1687 550 2113
rect 486 1681 550 1687
rect 600 2113 1100 2119
rect 600 1687 606 2113
rect 623 2065 1077 2113
rect 623 1735 685 2065
rect 1015 1735 1077 2065
rect 623 1687 1077 1735
rect 1094 1687 1100 2113
rect 600 1681 1100 1687
rect 1150 2113 1214 2119
rect 1150 1687 1156 2113
rect 1173 2086 1214 2113
rect 1586 2119 1619 2121
rect 1731 2144 2169 2150
rect 1731 2127 1737 2144
rect 2163 2127 2169 2144
rect 1731 2121 2169 2127
rect 1729 2119 2171 2121
rect 2281 2144 2719 2150
rect 2281 2127 2287 2144
rect 2713 2127 2719 2144
rect 2281 2121 2719 2127
rect 2281 2119 2314 2121
rect 1586 2113 1650 2119
rect 1586 2086 1627 2113
rect 1173 1714 1179 2086
rect 1621 1714 1627 2086
rect 1173 1687 1214 1714
rect 1150 1681 1214 1687
rect 486 1679 519 1681
rect 81 1673 519 1679
rect 81 1656 87 1673
rect 513 1656 519 1673
rect 81 1650 519 1656
rect 629 1679 1071 1681
rect 631 1673 1069 1679
rect 631 1656 637 1673
rect 1063 1656 1069 1673
rect 631 1650 1069 1656
rect 1181 1679 1214 1681
rect 1586 1687 1627 1714
rect 1644 1687 1650 2113
rect 1586 1681 1650 1687
rect 1700 2113 2200 2119
rect 1700 1687 1706 2113
rect 1723 2065 2177 2113
rect 1723 1735 1785 2065
rect 2115 1735 2177 2065
rect 1723 1687 2177 1735
rect 2194 1687 2200 2113
rect 1700 1681 2200 1687
rect 2250 2113 2314 2119
rect 2250 1687 2256 2113
rect 2273 2086 2314 2113
rect 2686 2119 2719 2121
rect 2831 2144 3269 2150
rect 2831 2127 2837 2144
rect 3263 2127 3269 2144
rect 2831 2121 3269 2127
rect 2829 2119 3271 2121
rect 3381 2144 3819 2150
rect 3381 2127 3387 2144
rect 3813 2127 3819 2144
rect 3381 2121 3819 2127
rect 3381 2119 3414 2121
rect 2686 2113 2750 2119
rect 2686 2086 2727 2113
rect 2273 1714 2279 2086
rect 2721 1714 2727 2086
rect 2273 1687 2314 1714
rect 2250 1681 2314 1687
rect 1586 1679 1619 1681
rect 1181 1673 1619 1679
rect 1181 1656 1187 1673
rect 1613 1656 1619 1673
rect 1181 1650 1619 1656
rect 1729 1679 2171 1681
rect 1731 1673 2169 1679
rect 1731 1656 1737 1673
rect 2163 1656 2169 1673
rect 1731 1650 2169 1656
rect 2281 1679 2314 1681
rect 2686 1687 2727 1714
rect 2744 1687 2750 2113
rect 2686 1681 2750 1687
rect 2800 2113 3300 2119
rect 2800 1687 2806 2113
rect 2823 2065 3277 2113
rect 2823 1735 2885 2065
rect 3215 1735 3277 2065
rect 2823 1687 3277 1735
rect 3294 1687 3300 2113
rect 2800 1681 3300 1687
rect 3350 2113 3414 2119
rect 3350 1687 3356 2113
rect 3373 2086 3414 2113
rect 3786 2119 3819 2121
rect 3931 2144 4369 2150
rect 3931 2127 3937 2144
rect 4363 2127 4369 2144
rect 3931 2121 4369 2127
rect 3929 2119 4371 2121
rect 4481 2144 4919 2150
rect 4481 2127 4487 2144
rect 4913 2127 4919 2144
rect 4481 2121 4919 2127
rect 4481 2119 4514 2121
rect 3786 2113 3850 2119
rect 3786 2086 3827 2113
rect 3373 1714 3379 2086
rect 3821 1714 3827 2086
rect 3373 1687 3414 1714
rect 3350 1681 3414 1687
rect 2686 1679 2719 1681
rect 2281 1673 2719 1679
rect 2281 1656 2287 1673
rect 2713 1656 2719 1673
rect 2281 1650 2719 1656
rect 2829 1679 3271 1681
rect 2831 1673 3269 1679
rect 2831 1656 2837 1673
rect 3263 1656 3269 1673
rect 2831 1650 3269 1656
rect 3381 1679 3414 1681
rect 3786 1687 3827 1714
rect 3844 1687 3850 2113
rect 3786 1681 3850 1687
rect 3900 2113 4400 2119
rect 3900 1687 3906 2113
rect 3923 2065 4377 2113
rect 3923 1735 3985 2065
rect 4315 1735 4377 2065
rect 3923 1687 4377 1735
rect 4394 1687 4400 2113
rect 3900 1681 4400 1687
rect 4450 2113 4514 2119
rect 4450 1687 4456 2113
rect 4473 2086 4514 2113
rect 4886 2119 4919 2121
rect 5031 2144 5469 2150
rect 5031 2127 5037 2144
rect 5463 2127 5469 2144
rect 5031 2121 5469 2127
rect 5029 2119 5471 2121
rect 5581 2144 6019 2150
rect 5581 2127 5587 2144
rect 6013 2127 6019 2144
rect 5581 2121 6019 2127
rect 5581 2119 5614 2121
rect 4886 2113 4950 2119
rect 4886 2086 4927 2113
rect 4473 1714 4479 2086
rect 4921 1714 4927 2086
rect 4473 1687 4514 1714
rect 4450 1681 4514 1687
rect 3786 1679 3819 1681
rect 3381 1673 3819 1679
rect 3381 1656 3387 1673
rect 3813 1656 3819 1673
rect 3381 1650 3819 1656
rect 3929 1679 4371 1681
rect 3931 1673 4369 1679
rect 3931 1656 3937 1673
rect 4363 1656 4369 1673
rect 3931 1650 4369 1656
rect 4481 1679 4514 1681
rect 4886 1687 4927 1714
rect 4944 1687 4950 2113
rect 4886 1681 4950 1687
rect 5000 2113 5500 2119
rect 5000 1687 5006 2113
rect 5023 2065 5477 2113
rect 5023 1735 5085 2065
rect 5415 1735 5477 2065
rect 5023 1687 5477 1735
rect 5494 1687 5500 2113
rect 5000 1681 5500 1687
rect 5550 2113 5614 2119
rect 5550 1687 5556 2113
rect 5573 2086 5614 2113
rect 5986 2119 6019 2121
rect 6131 2144 6569 2150
rect 6131 2127 6137 2144
rect 6563 2127 6569 2144
rect 6131 2121 6569 2127
rect 6129 2119 6571 2121
rect 6681 2144 7119 2150
rect 6681 2127 6687 2144
rect 7113 2127 7119 2144
rect 6681 2121 7119 2127
rect 6681 2119 6714 2121
rect 5986 2113 6050 2119
rect 5986 2086 6027 2113
rect 5573 1714 5579 2086
rect 6021 1714 6027 2086
rect 5573 1687 5614 1714
rect 5550 1681 5614 1687
rect 4886 1679 4919 1681
rect 4481 1673 4919 1679
rect 4481 1656 4487 1673
rect 4913 1656 4919 1673
rect 4481 1650 4919 1656
rect 5029 1679 5471 1681
rect 5031 1673 5469 1679
rect 5031 1656 5037 1673
rect 5463 1656 5469 1673
rect 5031 1650 5469 1656
rect 5581 1679 5614 1681
rect 5986 1687 6027 1714
rect 6044 1687 6050 2113
rect 5986 1681 6050 1687
rect 6100 2113 6600 2119
rect 6100 1687 6106 2113
rect 6123 2065 6577 2113
rect 6123 1735 6185 2065
rect 6515 1735 6577 2065
rect 6123 1687 6577 1735
rect 6594 1687 6600 2113
rect 6100 1681 6600 1687
rect 6650 2113 6714 2119
rect 6650 1687 6656 2113
rect 6673 2086 6714 2113
rect 7086 2119 7119 2121
rect 7231 2144 7669 2150
rect 7231 2127 7237 2144
rect 7663 2127 7669 2144
rect 7231 2121 7669 2127
rect 7229 2119 7671 2121
rect 7781 2144 8219 2150
rect 7781 2127 7787 2144
rect 8213 2127 8219 2144
rect 7781 2121 8219 2127
rect 7781 2119 7814 2121
rect 7086 2113 7150 2119
rect 7086 2086 7127 2113
rect 6673 1714 6679 2086
rect 7121 1714 7127 2086
rect 6673 1687 6714 1714
rect 6650 1681 6714 1687
rect 5986 1679 6019 1681
rect 5581 1673 6019 1679
rect 5581 1656 5587 1673
rect 6013 1656 6019 1673
rect 5581 1650 6019 1656
rect 6129 1679 6571 1681
rect 6131 1673 6569 1679
rect 6131 1656 6137 1673
rect 6563 1656 6569 1673
rect 6131 1650 6569 1656
rect 6681 1679 6714 1681
rect 7086 1687 7127 1714
rect 7144 1687 7150 2113
rect 7086 1681 7150 1687
rect 7200 2113 7700 2119
rect 7200 1687 7206 2113
rect 7223 2065 7677 2113
rect 7223 1735 7285 2065
rect 7615 1735 7677 2065
rect 7223 1687 7677 1735
rect 7694 1687 7700 2113
rect 7200 1681 7700 1687
rect 7750 2113 7814 2119
rect 7750 1687 7756 2113
rect 7773 2086 7814 2113
rect 8186 2119 8219 2121
rect 8331 2144 8769 2150
rect 8331 2127 8337 2144
rect 8763 2127 8769 2144
rect 8331 2121 8769 2127
rect 8329 2119 8771 2121
rect 8881 2144 9319 2150
rect 8881 2127 8887 2144
rect 9313 2127 9319 2144
rect 8881 2121 9319 2127
rect 8881 2119 8914 2121
rect 8186 2113 8250 2119
rect 8186 2086 8227 2113
rect 7773 1714 7779 2086
rect 8221 1714 8227 2086
rect 7773 1687 7814 1714
rect 7750 1681 7814 1687
rect 7086 1679 7119 1681
rect 6681 1673 7119 1679
rect 6681 1656 6687 1673
rect 7113 1656 7119 1673
rect 6681 1650 7119 1656
rect 7229 1679 7671 1681
rect 7231 1673 7669 1679
rect 7231 1656 7237 1673
rect 7663 1656 7669 1673
rect 7231 1650 7669 1656
rect 7781 1679 7814 1681
rect 8186 1687 8227 1714
rect 8244 1687 8250 2113
rect 8186 1681 8250 1687
rect 8300 2113 8800 2119
rect 8300 1687 8306 2113
rect 8323 2065 8777 2113
rect 8323 1735 8385 2065
rect 8715 1735 8777 2065
rect 8323 1687 8777 1735
rect 8794 1687 8800 2113
rect 8300 1681 8800 1687
rect 8850 2113 8914 2119
rect 8850 1687 8856 2113
rect 8873 2086 8914 2113
rect 9286 2119 9319 2121
rect 9431 2144 9869 2150
rect 9431 2127 9437 2144
rect 9863 2127 9869 2144
rect 9431 2121 9869 2127
rect 9429 2119 9871 2121
rect 9981 2144 10419 2150
rect 9981 2127 9987 2144
rect 10413 2127 10419 2144
rect 9981 2121 10419 2127
rect 9981 2119 10014 2121
rect 9286 2113 9350 2119
rect 9286 2086 9327 2113
rect 8873 1714 8879 2086
rect 9321 1714 9327 2086
rect 8873 1687 8914 1714
rect 8850 1681 8914 1687
rect 8186 1679 8219 1681
rect 7781 1673 8219 1679
rect 7781 1656 7787 1673
rect 8213 1656 8219 1673
rect 7781 1650 8219 1656
rect 8329 1679 8771 1681
rect 8331 1673 8769 1679
rect 8331 1656 8337 1673
rect 8763 1656 8769 1673
rect 8331 1650 8769 1656
rect 8881 1679 8914 1681
rect 9286 1687 9327 1714
rect 9344 1687 9350 2113
rect 9286 1681 9350 1687
rect 9400 2113 9900 2119
rect 9400 1687 9406 2113
rect 9423 2065 9877 2113
rect 9423 1735 9485 2065
rect 9815 1735 9877 2065
rect 9423 1687 9877 1735
rect 9894 1687 9900 2113
rect 9400 1681 9900 1687
rect 9950 2113 10014 2119
rect 9950 1687 9956 2113
rect 9973 2086 10014 2113
rect 10386 2119 10419 2121
rect 10531 2144 10969 2150
rect 10531 2127 10537 2144
rect 10963 2127 10969 2144
rect 10531 2121 10969 2127
rect 10529 2119 10971 2121
rect 11081 2144 11519 2150
rect 11081 2127 11087 2144
rect 11513 2127 11519 2144
rect 11081 2121 11519 2127
rect 11081 2119 11114 2121
rect 10386 2113 10450 2119
rect 10386 2086 10427 2113
rect 9973 1714 9979 2086
rect 10421 1714 10427 2086
rect 9973 1687 10014 1714
rect 9950 1681 10014 1687
rect 9286 1679 9319 1681
rect 8881 1673 9319 1679
rect 8881 1656 8887 1673
rect 9313 1656 9319 1673
rect 8881 1650 9319 1656
rect 9429 1679 9871 1681
rect 9431 1673 9869 1679
rect 9431 1656 9437 1673
rect 9863 1656 9869 1673
rect 9431 1650 9869 1656
rect 9981 1679 10014 1681
rect 10386 1687 10427 1714
rect 10444 1687 10450 2113
rect 10386 1681 10450 1687
rect 10500 2113 11000 2119
rect 10500 1687 10506 2113
rect 10523 2065 10977 2113
rect 10523 1735 10585 2065
rect 10915 1735 10977 2065
rect 10523 1687 10977 1735
rect 10994 1687 11000 2113
rect 10500 1681 11000 1687
rect 11050 2113 11114 2119
rect 11050 1687 11056 2113
rect 11073 2086 11114 2113
rect 11486 2119 11519 2121
rect 11631 2144 12069 2150
rect 11631 2127 11637 2144
rect 12063 2127 12069 2144
rect 11631 2121 12069 2127
rect 11629 2119 12071 2121
rect 12181 2144 12619 2150
rect 12181 2127 12187 2144
rect 12613 2127 12619 2144
rect 12181 2121 12619 2127
rect 12181 2119 12214 2121
rect 11486 2113 11550 2119
rect 11486 2086 11527 2113
rect 11073 1714 11079 2086
rect 11521 1714 11527 2086
rect 11073 1687 11114 1714
rect 11050 1681 11114 1687
rect 10386 1679 10419 1681
rect 9981 1673 10419 1679
rect 9981 1656 9987 1673
rect 10413 1656 10419 1673
rect 9981 1650 10419 1656
rect 10529 1679 10971 1681
rect 10531 1673 10969 1679
rect 10531 1656 10537 1673
rect 10963 1656 10969 1673
rect 10531 1650 10969 1656
rect 11081 1679 11114 1681
rect 11486 1687 11527 1714
rect 11544 1687 11550 2113
rect 11486 1681 11550 1687
rect 11600 2113 12100 2119
rect 11600 1687 11606 2113
rect 11623 2065 12077 2113
rect 11623 1735 11685 2065
rect 12015 1735 12077 2065
rect 11623 1687 12077 1735
rect 12094 1687 12100 2113
rect 11600 1681 12100 1687
rect 12150 2113 12214 2119
rect 12150 1687 12156 2113
rect 12173 2086 12214 2113
rect 12586 2119 12619 2121
rect 12731 2144 13169 2150
rect 12731 2127 12737 2144
rect 13163 2127 13169 2144
rect 12731 2121 13169 2127
rect 12729 2119 13171 2121
rect 13281 2144 13719 2150
rect 13281 2127 13287 2144
rect 13713 2127 13719 2144
rect 13281 2121 13719 2127
rect 13281 2119 13314 2121
rect 12586 2113 12650 2119
rect 12586 2086 12627 2113
rect 12173 1714 12179 2086
rect 12621 1714 12627 2086
rect 12173 1687 12214 1714
rect 12150 1681 12214 1687
rect 11486 1679 11519 1681
rect 11081 1673 11519 1679
rect 11081 1656 11087 1673
rect 11513 1656 11519 1673
rect 11081 1650 11519 1656
rect 11629 1679 12071 1681
rect 11631 1673 12069 1679
rect 11631 1656 11637 1673
rect 12063 1656 12069 1673
rect 11631 1650 12069 1656
rect 12181 1679 12214 1681
rect 12586 1687 12627 1714
rect 12644 1687 12650 2113
rect 12586 1681 12650 1687
rect 12700 2113 13200 2119
rect 12700 1687 12706 2113
rect 12723 2065 13177 2113
rect 12723 1735 12785 2065
rect 13115 1735 13177 2065
rect 12723 1687 13177 1735
rect 13194 1687 13200 2113
rect 12700 1681 13200 1687
rect 13250 2113 13314 2119
rect 13250 1687 13256 2113
rect 13273 2086 13314 2113
rect 13273 1714 13279 2086
rect 13273 1687 13314 1714
rect 13250 1681 13314 1687
rect 12586 1679 12619 1681
rect 12181 1673 12619 1679
rect 12181 1656 12187 1673
rect 12613 1656 12619 1673
rect 12181 1650 12619 1656
rect 12729 1679 13171 1681
rect 12731 1673 13169 1679
rect 12731 1656 12737 1673
rect 13163 1656 13169 1673
rect 12731 1650 13169 1656
rect 13281 1679 13314 1681
rect 13281 1673 13719 1679
rect 13281 1656 13287 1673
rect 13713 1656 13719 1673
rect 13281 1650 13719 1656
rect -469 1594 -31 1600
rect -469 1577 -463 1594
rect -37 1577 -31 1594
rect -469 1571 -31 1577
rect -64 1569 -31 1571
rect 81 1594 519 1600
rect 81 1577 87 1594
rect 513 1577 519 1594
rect 81 1571 519 1577
rect 79 1569 521 1571
rect 631 1594 1069 1600
rect 631 1577 637 1594
rect 1063 1577 1069 1594
rect 631 1571 1069 1577
rect 631 1569 664 1571
rect -64 1563 0 1569
rect -64 1536 -23 1563
rect -29 1164 -23 1536
rect -64 1137 -23 1164
rect -6 1137 0 1563
rect -64 1131 0 1137
rect 50 1563 550 1569
rect 50 1137 56 1563
rect 73 1515 527 1563
rect 73 1185 135 1515
rect 465 1185 527 1515
rect 73 1137 527 1185
rect 544 1137 550 1563
rect 50 1131 550 1137
rect 600 1563 664 1569
rect 600 1137 606 1563
rect 623 1536 664 1563
rect 1036 1569 1069 1571
rect 1181 1594 1619 1600
rect 1181 1577 1187 1594
rect 1613 1577 1619 1594
rect 1181 1571 1619 1577
rect 1179 1569 1621 1571
rect 1731 1594 2169 1600
rect 1731 1577 1737 1594
rect 2163 1577 2169 1594
rect 1731 1571 2169 1577
rect 1731 1569 1764 1571
rect 1036 1563 1100 1569
rect 1036 1536 1077 1563
rect 623 1164 629 1536
rect 1071 1164 1077 1536
rect 623 1137 664 1164
rect 600 1131 664 1137
rect -64 1129 -31 1131
rect -469 1123 -31 1129
rect -469 1106 -463 1123
rect -37 1106 -31 1123
rect -469 1100 -31 1106
rect 79 1129 521 1131
rect 81 1123 519 1129
rect 81 1106 87 1123
rect 513 1106 519 1123
rect 81 1100 519 1106
rect 631 1129 664 1131
rect 1036 1137 1077 1164
rect 1094 1137 1100 1563
rect 1036 1131 1100 1137
rect 1150 1563 1650 1569
rect 1150 1137 1156 1563
rect 1173 1515 1627 1563
rect 1173 1185 1235 1515
rect 1565 1185 1627 1515
rect 1173 1137 1627 1185
rect 1644 1137 1650 1563
rect 1150 1131 1650 1137
rect 1700 1563 1764 1569
rect 1700 1137 1706 1563
rect 1723 1536 1764 1563
rect 2136 1569 2169 1571
rect 2281 1594 2719 1600
rect 2281 1577 2287 1594
rect 2713 1577 2719 1594
rect 2281 1571 2719 1577
rect 2279 1569 2721 1571
rect 2831 1594 3269 1600
rect 2831 1577 2837 1594
rect 3263 1577 3269 1594
rect 2831 1571 3269 1577
rect 2831 1569 2864 1571
rect 2136 1563 2200 1569
rect 2136 1536 2177 1563
rect 1723 1164 1729 1536
rect 2171 1164 2177 1536
rect 1723 1137 1764 1164
rect 1700 1131 1764 1137
rect 1036 1129 1069 1131
rect 631 1123 1069 1129
rect 631 1106 637 1123
rect 1063 1106 1069 1123
rect 631 1100 1069 1106
rect 1179 1129 1621 1131
rect 1181 1123 1619 1129
rect 1181 1106 1187 1123
rect 1613 1106 1619 1123
rect 1181 1100 1619 1106
rect 1731 1129 1764 1131
rect 2136 1137 2177 1164
rect 2194 1137 2200 1563
rect 2136 1131 2200 1137
rect 2250 1563 2750 1569
rect 2250 1137 2256 1563
rect 2273 1515 2727 1563
rect 2273 1185 2335 1515
rect 2665 1185 2727 1515
rect 2273 1137 2727 1185
rect 2744 1137 2750 1563
rect 2250 1131 2750 1137
rect 2800 1563 2864 1569
rect 2800 1137 2806 1563
rect 2823 1536 2864 1563
rect 3236 1569 3269 1571
rect 3381 1594 3819 1600
rect 3381 1577 3387 1594
rect 3813 1577 3819 1594
rect 3381 1571 3819 1577
rect 3379 1569 3821 1571
rect 3931 1594 4369 1600
rect 3931 1577 3937 1594
rect 4363 1577 4369 1594
rect 3931 1571 4369 1577
rect 3931 1569 3964 1571
rect 3236 1563 3300 1569
rect 3236 1536 3277 1563
rect 2823 1164 2829 1536
rect 3271 1164 3277 1536
rect 2823 1137 2864 1164
rect 2800 1131 2864 1137
rect 2136 1129 2169 1131
rect 1731 1123 2169 1129
rect 1731 1106 1737 1123
rect 2163 1106 2169 1123
rect 1731 1100 2169 1106
rect 2279 1129 2721 1131
rect 2281 1123 2719 1129
rect 2281 1106 2287 1123
rect 2713 1106 2719 1123
rect 2281 1100 2719 1106
rect 2831 1129 2864 1131
rect 3236 1137 3277 1164
rect 3294 1137 3300 1563
rect 3236 1131 3300 1137
rect 3350 1563 3850 1569
rect 3350 1137 3356 1563
rect 3373 1515 3827 1563
rect 3373 1185 3435 1515
rect 3765 1185 3827 1515
rect 3373 1137 3827 1185
rect 3844 1137 3850 1563
rect 3350 1131 3850 1137
rect 3900 1563 3964 1569
rect 3900 1137 3906 1563
rect 3923 1536 3964 1563
rect 4336 1569 4369 1571
rect 4481 1594 4919 1600
rect 4481 1577 4487 1594
rect 4913 1577 4919 1594
rect 4481 1571 4919 1577
rect 4479 1569 4921 1571
rect 5031 1594 5469 1600
rect 5031 1577 5037 1594
rect 5463 1577 5469 1594
rect 5031 1571 5469 1577
rect 5031 1569 5064 1571
rect 4336 1563 4400 1569
rect 4336 1536 4377 1563
rect 3923 1164 3929 1536
rect 4371 1164 4377 1536
rect 3923 1137 3964 1164
rect 3900 1131 3964 1137
rect 3236 1129 3269 1131
rect 2831 1123 3269 1129
rect 2831 1106 2837 1123
rect 3263 1106 3269 1123
rect 2831 1100 3269 1106
rect 3379 1129 3821 1131
rect 3381 1123 3819 1129
rect 3381 1106 3387 1123
rect 3813 1106 3819 1123
rect 3381 1100 3819 1106
rect 3931 1129 3964 1131
rect 4336 1137 4377 1164
rect 4394 1137 4400 1563
rect 4336 1131 4400 1137
rect 4450 1563 4950 1569
rect 4450 1137 4456 1563
rect 4473 1515 4927 1563
rect 4473 1185 4535 1515
rect 4865 1185 4927 1515
rect 4473 1137 4927 1185
rect 4944 1137 4950 1563
rect 4450 1131 4950 1137
rect 5000 1563 5064 1569
rect 5000 1137 5006 1563
rect 5023 1536 5064 1563
rect 5436 1569 5469 1571
rect 5581 1594 6019 1600
rect 5581 1577 5587 1594
rect 6013 1577 6019 1594
rect 5581 1571 6019 1577
rect 5579 1569 6021 1571
rect 6131 1594 6569 1600
rect 6131 1577 6137 1594
rect 6563 1577 6569 1594
rect 6131 1571 6569 1577
rect 6131 1569 6164 1571
rect 5436 1563 5500 1569
rect 5436 1536 5477 1563
rect 5023 1164 5029 1536
rect 5471 1164 5477 1536
rect 5023 1137 5064 1164
rect 5000 1131 5064 1137
rect 4336 1129 4369 1131
rect 3931 1123 4369 1129
rect 3931 1106 3937 1123
rect 4363 1106 4369 1123
rect 3931 1100 4369 1106
rect 4479 1129 4921 1131
rect 4481 1123 4919 1129
rect 4481 1106 4487 1123
rect 4913 1106 4919 1123
rect 4481 1100 4919 1106
rect 5031 1129 5064 1131
rect 5436 1137 5477 1164
rect 5494 1137 5500 1563
rect 5436 1131 5500 1137
rect 5550 1563 6050 1569
rect 5550 1137 5556 1563
rect 5573 1515 6027 1563
rect 5573 1185 5635 1515
rect 5965 1185 6027 1515
rect 5573 1137 6027 1185
rect 6044 1137 6050 1563
rect 5550 1131 6050 1137
rect 6100 1563 6164 1569
rect 6100 1137 6106 1563
rect 6123 1536 6164 1563
rect 6536 1569 6569 1571
rect 6681 1594 7119 1600
rect 6681 1577 6687 1594
rect 7113 1577 7119 1594
rect 6681 1571 7119 1577
rect 6679 1569 7121 1571
rect 7231 1594 7669 1600
rect 7231 1577 7237 1594
rect 7663 1577 7669 1594
rect 7231 1571 7669 1577
rect 7231 1569 7264 1571
rect 6536 1563 6600 1569
rect 6536 1536 6577 1563
rect 6123 1164 6129 1536
rect 6571 1164 6577 1536
rect 6123 1137 6164 1164
rect 6100 1131 6164 1137
rect 5436 1129 5469 1131
rect 5031 1123 5469 1129
rect 5031 1106 5037 1123
rect 5463 1106 5469 1123
rect 5031 1100 5469 1106
rect 5579 1129 6021 1131
rect 5581 1123 6019 1129
rect 5581 1106 5587 1123
rect 6013 1106 6019 1123
rect 5581 1100 6019 1106
rect 6131 1129 6164 1131
rect 6536 1137 6577 1164
rect 6594 1137 6600 1563
rect 6536 1131 6600 1137
rect 6650 1563 7150 1569
rect 6650 1137 6656 1563
rect 6673 1515 7127 1563
rect 6673 1185 6735 1515
rect 7065 1185 7127 1515
rect 6673 1137 7127 1185
rect 7144 1137 7150 1563
rect 6650 1131 7150 1137
rect 7200 1563 7264 1569
rect 7200 1137 7206 1563
rect 7223 1536 7264 1563
rect 7636 1569 7669 1571
rect 7781 1594 8219 1600
rect 7781 1577 7787 1594
rect 8213 1577 8219 1594
rect 7781 1571 8219 1577
rect 7779 1569 8221 1571
rect 8331 1594 8769 1600
rect 8331 1577 8337 1594
rect 8763 1577 8769 1594
rect 8331 1571 8769 1577
rect 8331 1569 8364 1571
rect 7636 1563 7700 1569
rect 7636 1536 7677 1563
rect 7223 1164 7229 1536
rect 7671 1164 7677 1536
rect 7223 1137 7264 1164
rect 7200 1131 7264 1137
rect 6536 1129 6569 1131
rect 6131 1123 6569 1129
rect 6131 1106 6137 1123
rect 6563 1106 6569 1123
rect 6131 1100 6569 1106
rect 6679 1129 7121 1131
rect 6681 1123 7119 1129
rect 6681 1106 6687 1123
rect 7113 1106 7119 1123
rect 6681 1100 7119 1106
rect 7231 1129 7264 1131
rect 7636 1137 7677 1164
rect 7694 1137 7700 1563
rect 7636 1131 7700 1137
rect 7750 1563 8250 1569
rect 7750 1137 7756 1563
rect 7773 1515 8227 1563
rect 7773 1185 7835 1515
rect 8165 1185 8227 1515
rect 7773 1137 8227 1185
rect 8244 1137 8250 1563
rect 7750 1131 8250 1137
rect 8300 1563 8364 1569
rect 8300 1137 8306 1563
rect 8323 1536 8364 1563
rect 8736 1569 8769 1571
rect 8881 1594 9319 1600
rect 8881 1577 8887 1594
rect 9313 1577 9319 1594
rect 8881 1571 9319 1577
rect 8879 1569 9321 1571
rect 9431 1594 9869 1600
rect 9431 1577 9437 1594
rect 9863 1577 9869 1594
rect 9431 1571 9869 1577
rect 9431 1569 9464 1571
rect 8736 1563 8800 1569
rect 8736 1536 8777 1563
rect 8323 1164 8329 1536
rect 8771 1164 8777 1536
rect 8323 1137 8364 1164
rect 8300 1131 8364 1137
rect 7636 1129 7669 1131
rect 7231 1123 7669 1129
rect 7231 1106 7237 1123
rect 7663 1106 7669 1123
rect 7231 1100 7669 1106
rect 7779 1129 8221 1131
rect 7781 1123 8219 1129
rect 7781 1106 7787 1123
rect 8213 1106 8219 1123
rect 7781 1100 8219 1106
rect 8331 1129 8364 1131
rect 8736 1137 8777 1164
rect 8794 1137 8800 1563
rect 8736 1131 8800 1137
rect 8850 1563 9350 1569
rect 8850 1137 8856 1563
rect 8873 1515 9327 1563
rect 8873 1185 8935 1515
rect 9265 1185 9327 1515
rect 8873 1137 9327 1185
rect 9344 1137 9350 1563
rect 8850 1131 9350 1137
rect 9400 1563 9464 1569
rect 9400 1137 9406 1563
rect 9423 1536 9464 1563
rect 9836 1569 9869 1571
rect 9981 1594 10419 1600
rect 9981 1577 9987 1594
rect 10413 1577 10419 1594
rect 9981 1571 10419 1577
rect 9979 1569 10421 1571
rect 10531 1594 10969 1600
rect 10531 1577 10537 1594
rect 10963 1577 10969 1594
rect 10531 1571 10969 1577
rect 10531 1569 10564 1571
rect 9836 1563 9900 1569
rect 9836 1536 9877 1563
rect 9423 1164 9429 1536
rect 9871 1164 9877 1536
rect 9423 1137 9464 1164
rect 9400 1131 9464 1137
rect 8736 1129 8769 1131
rect 8331 1123 8769 1129
rect 8331 1106 8337 1123
rect 8763 1106 8769 1123
rect 8331 1100 8769 1106
rect 8879 1129 9321 1131
rect 8881 1123 9319 1129
rect 8881 1106 8887 1123
rect 9313 1106 9319 1123
rect 8881 1100 9319 1106
rect 9431 1129 9464 1131
rect 9836 1137 9877 1164
rect 9894 1137 9900 1563
rect 9836 1131 9900 1137
rect 9950 1563 10450 1569
rect 9950 1137 9956 1563
rect 9973 1515 10427 1563
rect 9973 1185 10035 1515
rect 10365 1185 10427 1515
rect 9973 1137 10427 1185
rect 10444 1137 10450 1563
rect 9950 1131 10450 1137
rect 10500 1563 10564 1569
rect 10500 1137 10506 1563
rect 10523 1536 10564 1563
rect 10936 1569 10969 1571
rect 11081 1594 11519 1600
rect 11081 1577 11087 1594
rect 11513 1577 11519 1594
rect 11081 1571 11519 1577
rect 11079 1569 11521 1571
rect 11631 1594 12069 1600
rect 11631 1577 11637 1594
rect 12063 1577 12069 1594
rect 11631 1571 12069 1577
rect 11631 1569 11664 1571
rect 10936 1563 11000 1569
rect 10936 1536 10977 1563
rect 10523 1164 10529 1536
rect 10971 1164 10977 1536
rect 10523 1137 10564 1164
rect 10500 1131 10564 1137
rect 9836 1129 9869 1131
rect 9431 1123 9869 1129
rect 9431 1106 9437 1123
rect 9863 1106 9869 1123
rect 9431 1100 9869 1106
rect 9979 1129 10421 1131
rect 9981 1123 10419 1129
rect 9981 1106 9987 1123
rect 10413 1106 10419 1123
rect 9981 1100 10419 1106
rect 10531 1129 10564 1131
rect 10936 1137 10977 1164
rect 10994 1137 11000 1563
rect 10936 1131 11000 1137
rect 11050 1563 11550 1569
rect 11050 1137 11056 1563
rect 11073 1515 11527 1563
rect 11073 1185 11135 1515
rect 11465 1185 11527 1515
rect 11073 1137 11527 1185
rect 11544 1137 11550 1563
rect 11050 1131 11550 1137
rect 11600 1563 11664 1569
rect 11600 1137 11606 1563
rect 11623 1536 11664 1563
rect 12036 1569 12069 1571
rect 12181 1594 12619 1600
rect 12181 1577 12187 1594
rect 12613 1577 12619 1594
rect 12181 1571 12619 1577
rect 12179 1569 12621 1571
rect 12731 1594 13169 1600
rect 12731 1577 12737 1594
rect 13163 1577 13169 1594
rect 12731 1571 13169 1577
rect 12731 1569 12764 1571
rect 12036 1563 12100 1569
rect 12036 1536 12077 1563
rect 11623 1164 11629 1536
rect 12071 1164 12077 1536
rect 11623 1137 11664 1164
rect 11600 1131 11664 1137
rect 10936 1129 10969 1131
rect 10531 1123 10969 1129
rect 10531 1106 10537 1123
rect 10963 1106 10969 1123
rect 10531 1100 10969 1106
rect 11079 1129 11521 1131
rect 11081 1123 11519 1129
rect 11081 1106 11087 1123
rect 11513 1106 11519 1123
rect 11081 1100 11519 1106
rect 11631 1129 11664 1131
rect 12036 1137 12077 1164
rect 12094 1137 12100 1563
rect 12036 1131 12100 1137
rect 12150 1563 12650 1569
rect 12150 1137 12156 1563
rect 12173 1515 12627 1563
rect 12173 1185 12235 1515
rect 12565 1185 12627 1515
rect 12173 1137 12627 1185
rect 12644 1137 12650 1563
rect 12150 1131 12650 1137
rect 12700 1563 12764 1569
rect 12700 1137 12706 1563
rect 12723 1536 12764 1563
rect 13136 1569 13169 1571
rect 13281 1594 13719 1600
rect 13281 1577 13287 1594
rect 13713 1577 13719 1594
rect 13281 1571 13719 1577
rect 13279 1569 13721 1571
rect 13136 1563 13200 1569
rect 13136 1536 13177 1563
rect 12723 1164 12729 1536
rect 13171 1164 13177 1536
rect 12723 1137 12764 1164
rect 12700 1131 12764 1137
rect 12036 1129 12069 1131
rect 11631 1123 12069 1129
rect 11631 1106 11637 1123
rect 12063 1106 12069 1123
rect 11631 1100 12069 1106
rect 12179 1129 12621 1131
rect 12181 1123 12619 1129
rect 12181 1106 12187 1123
rect 12613 1106 12619 1123
rect 12181 1100 12619 1106
rect 12731 1129 12764 1131
rect 13136 1137 13177 1164
rect 13194 1137 13200 1563
rect 13136 1131 13200 1137
rect 13250 1563 13721 1569
rect 13250 1137 13256 1563
rect 13273 1515 13721 1563
rect 13273 1185 13335 1515
rect 13665 1185 13721 1515
rect 13273 1137 13721 1185
rect 13250 1131 13721 1137
rect 13136 1129 13169 1131
rect 12731 1123 13169 1129
rect 12731 1106 12737 1123
rect 13163 1106 13169 1123
rect 12731 1100 13169 1106
rect 13279 1129 13721 1131
rect 13281 1123 13719 1129
rect 13281 1106 13287 1123
rect 13713 1106 13719 1123
rect 13281 1100 13719 1106
rect -469 1044 -31 1050
rect -469 1027 -463 1044
rect -37 1027 -31 1044
rect -469 1021 -31 1027
rect -471 1019 -29 1021
rect 81 1044 519 1050
rect 81 1027 87 1044
rect 513 1027 519 1044
rect 81 1021 519 1027
rect 81 1019 114 1021
rect -471 1013 0 1019
rect -471 965 -23 1013
rect -471 635 -415 965
rect -85 635 -23 965
rect -471 587 -23 635
rect -6 587 0 1013
rect -471 581 0 587
rect 50 1013 114 1019
rect 50 587 56 1013
rect 73 986 114 1013
rect 486 1019 519 1021
rect 631 1044 1069 1050
rect 631 1027 637 1044
rect 1063 1027 1069 1044
rect 631 1021 1069 1027
rect 629 1019 1071 1021
rect 1181 1044 1619 1050
rect 1181 1027 1187 1044
rect 1613 1027 1619 1044
rect 1181 1021 1619 1027
rect 1181 1019 1214 1021
rect 486 1013 550 1019
rect 486 986 527 1013
rect 73 614 79 986
rect 521 614 527 986
rect 73 587 114 614
rect 50 581 114 587
rect -471 579 -29 581
rect -469 573 -31 579
rect -469 556 -463 573
rect -37 556 -31 573
rect -469 550 -31 556
rect 81 579 114 581
rect 486 587 527 614
rect 544 587 550 1013
rect 486 581 550 587
rect 600 1013 1100 1019
rect 600 587 606 1013
rect 623 965 1077 1013
rect 623 635 685 965
rect 1015 635 1077 965
rect 623 587 1077 635
rect 1094 587 1100 1013
rect 600 581 1100 587
rect 1150 1013 1214 1019
rect 1150 587 1156 1013
rect 1173 986 1214 1013
rect 1586 1019 1619 1021
rect 1731 1044 2169 1050
rect 1731 1027 1737 1044
rect 2163 1027 2169 1044
rect 1731 1021 2169 1027
rect 1729 1019 2171 1021
rect 2281 1044 2719 1050
rect 2281 1027 2287 1044
rect 2713 1027 2719 1044
rect 2281 1021 2719 1027
rect 2281 1019 2314 1021
rect 1586 1013 1650 1019
rect 1586 986 1627 1013
rect 1173 614 1179 986
rect 1621 614 1627 986
rect 1173 587 1214 614
rect 1150 581 1214 587
rect 486 579 519 581
rect 81 573 519 579
rect 81 556 87 573
rect 513 556 519 573
rect 81 550 519 556
rect 629 579 1071 581
rect 631 573 1069 579
rect 631 556 637 573
rect 1063 556 1069 573
rect 631 550 1069 556
rect 1181 579 1214 581
rect 1586 587 1627 614
rect 1644 587 1650 1013
rect 1586 581 1650 587
rect 1700 1013 2200 1019
rect 1700 587 1706 1013
rect 1723 965 2177 1013
rect 1723 635 1785 965
rect 2115 635 2177 965
rect 1723 587 2177 635
rect 2194 587 2200 1013
rect 1700 581 2200 587
rect 2250 1013 2314 1019
rect 2250 587 2256 1013
rect 2273 986 2314 1013
rect 2686 1019 2719 1021
rect 2831 1044 3269 1050
rect 2831 1027 2837 1044
rect 3263 1027 3269 1044
rect 2831 1021 3269 1027
rect 2829 1019 3271 1021
rect 3381 1044 3819 1050
rect 3381 1027 3387 1044
rect 3813 1027 3819 1044
rect 3381 1021 3819 1027
rect 3381 1019 3414 1021
rect 2686 1013 2750 1019
rect 2686 986 2727 1013
rect 2273 614 2279 986
rect 2721 614 2727 986
rect 2273 587 2314 614
rect 2250 581 2314 587
rect 1586 579 1619 581
rect 1181 573 1619 579
rect 1181 556 1187 573
rect 1613 556 1619 573
rect 1181 550 1619 556
rect 1729 579 2171 581
rect 1731 573 2169 579
rect 1731 556 1737 573
rect 2163 556 2169 573
rect 1731 550 2169 556
rect 2281 579 2314 581
rect 2686 587 2727 614
rect 2744 587 2750 1013
rect 2686 581 2750 587
rect 2800 1013 3300 1019
rect 2800 587 2806 1013
rect 2823 965 3277 1013
rect 2823 635 2885 965
rect 3215 635 3277 965
rect 2823 587 3277 635
rect 3294 587 3300 1013
rect 2800 581 3300 587
rect 3350 1013 3414 1019
rect 3350 587 3356 1013
rect 3373 986 3414 1013
rect 3786 1019 3819 1021
rect 3931 1044 4369 1050
rect 3931 1027 3937 1044
rect 4363 1027 4369 1044
rect 3931 1021 4369 1027
rect 3929 1019 4371 1021
rect 4481 1044 4919 1050
rect 4481 1027 4487 1044
rect 4913 1027 4919 1044
rect 4481 1021 4919 1027
rect 4481 1019 4514 1021
rect 3786 1013 3850 1019
rect 3786 986 3827 1013
rect 3373 614 3379 986
rect 3821 614 3827 986
rect 3373 587 3414 614
rect 3350 581 3414 587
rect 2686 579 2719 581
rect 2281 573 2719 579
rect 2281 556 2287 573
rect 2713 556 2719 573
rect 2281 550 2719 556
rect 2829 579 3271 581
rect 2831 573 3269 579
rect 2831 556 2837 573
rect 3263 556 3269 573
rect 2831 550 3269 556
rect 3381 579 3414 581
rect 3786 587 3827 614
rect 3844 587 3850 1013
rect 3786 581 3850 587
rect 3900 1013 4400 1019
rect 3900 587 3906 1013
rect 3923 965 4377 1013
rect 3923 635 3985 965
rect 4315 635 4377 965
rect 3923 587 4377 635
rect 4394 587 4400 1013
rect 3900 581 4400 587
rect 4450 1013 4514 1019
rect 4450 587 4456 1013
rect 4473 986 4514 1013
rect 4886 1019 4919 1021
rect 5031 1044 5469 1050
rect 5031 1027 5037 1044
rect 5463 1027 5469 1044
rect 5031 1021 5469 1027
rect 5029 1019 5471 1021
rect 5581 1044 6019 1050
rect 5581 1027 5587 1044
rect 6013 1027 6019 1044
rect 5581 1021 6019 1027
rect 5581 1019 5614 1021
rect 4886 1013 4950 1019
rect 4886 986 4927 1013
rect 4473 614 4479 986
rect 4921 614 4927 986
rect 4473 587 4514 614
rect 4450 581 4514 587
rect 3786 579 3819 581
rect 3381 573 3819 579
rect 3381 556 3387 573
rect 3813 556 3819 573
rect 3381 550 3819 556
rect 3929 579 4371 581
rect 3931 573 4369 579
rect 3931 556 3937 573
rect 4363 556 4369 573
rect 3931 550 4369 556
rect 4481 579 4514 581
rect 4886 587 4927 614
rect 4944 587 4950 1013
rect 4886 581 4950 587
rect 5000 1013 5500 1019
rect 5000 587 5006 1013
rect 5023 965 5477 1013
rect 5023 635 5085 965
rect 5415 635 5477 965
rect 5023 587 5477 635
rect 5494 587 5500 1013
rect 5000 581 5500 587
rect 5550 1013 5614 1019
rect 5550 587 5556 1013
rect 5573 986 5614 1013
rect 5986 1019 6019 1021
rect 6131 1044 6569 1050
rect 6131 1027 6137 1044
rect 6563 1027 6569 1044
rect 6131 1021 6569 1027
rect 6129 1019 6571 1021
rect 6681 1044 7119 1050
rect 6681 1027 6687 1044
rect 7113 1027 7119 1044
rect 6681 1021 7119 1027
rect 6681 1019 6714 1021
rect 5986 1013 6050 1019
rect 5986 986 6027 1013
rect 5573 614 5579 986
rect 6021 614 6027 986
rect 5573 587 5614 614
rect 5550 581 5614 587
rect 4886 579 4919 581
rect 4481 573 4919 579
rect 4481 556 4487 573
rect 4913 556 4919 573
rect 4481 550 4919 556
rect 5029 579 5471 581
rect 5031 573 5469 579
rect 5031 556 5037 573
rect 5463 556 5469 573
rect 5031 550 5469 556
rect 5581 579 5614 581
rect 5986 587 6027 614
rect 6044 587 6050 1013
rect 5986 581 6050 587
rect 6100 1013 6600 1019
rect 6100 587 6106 1013
rect 6123 965 6577 1013
rect 6123 635 6185 965
rect 6515 635 6577 965
rect 6123 587 6577 635
rect 6594 587 6600 1013
rect 6100 581 6600 587
rect 6650 1013 6714 1019
rect 6650 587 6656 1013
rect 6673 986 6714 1013
rect 7086 1019 7119 1021
rect 7231 1044 7669 1050
rect 7231 1027 7237 1044
rect 7663 1027 7669 1044
rect 7231 1021 7669 1027
rect 7229 1019 7671 1021
rect 7781 1044 8219 1050
rect 7781 1027 7787 1044
rect 8213 1027 8219 1044
rect 7781 1021 8219 1027
rect 7781 1019 7814 1021
rect 7086 1013 7150 1019
rect 7086 986 7127 1013
rect 6673 614 6679 986
rect 7121 614 7127 986
rect 6673 587 6714 614
rect 6650 581 6714 587
rect 5986 579 6019 581
rect 5581 573 6019 579
rect 5581 556 5587 573
rect 6013 556 6019 573
rect 5581 550 6019 556
rect 6129 579 6571 581
rect 6131 573 6569 579
rect 6131 556 6137 573
rect 6563 556 6569 573
rect 6131 550 6569 556
rect 6681 579 6714 581
rect 7086 587 7127 614
rect 7144 587 7150 1013
rect 7086 581 7150 587
rect 7200 1013 7700 1019
rect 7200 587 7206 1013
rect 7223 965 7677 1013
rect 7223 635 7285 965
rect 7615 635 7677 965
rect 7223 587 7677 635
rect 7694 587 7700 1013
rect 7200 581 7700 587
rect 7750 1013 7814 1019
rect 7750 587 7756 1013
rect 7773 986 7814 1013
rect 8186 1019 8219 1021
rect 8331 1044 8769 1050
rect 8331 1027 8337 1044
rect 8763 1027 8769 1044
rect 8331 1021 8769 1027
rect 8329 1019 8771 1021
rect 8881 1044 9319 1050
rect 8881 1027 8887 1044
rect 9313 1027 9319 1044
rect 8881 1021 9319 1027
rect 8881 1019 8914 1021
rect 8186 1013 8250 1019
rect 8186 986 8227 1013
rect 7773 614 7779 986
rect 8221 614 8227 986
rect 7773 587 7814 614
rect 7750 581 7814 587
rect 7086 579 7119 581
rect 6681 573 7119 579
rect 6681 556 6687 573
rect 7113 556 7119 573
rect 6681 550 7119 556
rect 7229 579 7671 581
rect 7231 573 7669 579
rect 7231 556 7237 573
rect 7663 556 7669 573
rect 7231 550 7669 556
rect 7781 579 7814 581
rect 8186 587 8227 614
rect 8244 587 8250 1013
rect 8186 581 8250 587
rect 8300 1013 8800 1019
rect 8300 587 8306 1013
rect 8323 965 8777 1013
rect 8323 635 8385 965
rect 8715 635 8777 965
rect 8323 587 8777 635
rect 8794 587 8800 1013
rect 8300 581 8800 587
rect 8850 1013 8914 1019
rect 8850 587 8856 1013
rect 8873 986 8914 1013
rect 9286 1019 9319 1021
rect 9431 1044 9869 1050
rect 9431 1027 9437 1044
rect 9863 1027 9869 1044
rect 9431 1021 9869 1027
rect 9429 1019 9871 1021
rect 9981 1044 10419 1050
rect 9981 1027 9987 1044
rect 10413 1027 10419 1044
rect 9981 1021 10419 1027
rect 9981 1019 10014 1021
rect 9286 1013 9350 1019
rect 9286 986 9327 1013
rect 8873 614 8879 986
rect 9321 614 9327 986
rect 8873 587 8914 614
rect 8850 581 8914 587
rect 8186 579 8219 581
rect 7781 573 8219 579
rect 7781 556 7787 573
rect 8213 556 8219 573
rect 7781 550 8219 556
rect 8329 579 8771 581
rect 8331 573 8769 579
rect 8331 556 8337 573
rect 8763 556 8769 573
rect 8331 550 8769 556
rect 8881 579 8914 581
rect 9286 587 9327 614
rect 9344 587 9350 1013
rect 9286 581 9350 587
rect 9400 1013 9900 1019
rect 9400 587 9406 1013
rect 9423 965 9877 1013
rect 9423 635 9485 965
rect 9815 635 9877 965
rect 9423 587 9877 635
rect 9894 587 9900 1013
rect 9400 581 9900 587
rect 9950 1013 10014 1019
rect 9950 587 9956 1013
rect 9973 986 10014 1013
rect 10386 1019 10419 1021
rect 10531 1044 10969 1050
rect 10531 1027 10537 1044
rect 10963 1027 10969 1044
rect 10531 1021 10969 1027
rect 10529 1019 10971 1021
rect 11081 1044 11519 1050
rect 11081 1027 11087 1044
rect 11513 1027 11519 1044
rect 11081 1021 11519 1027
rect 11081 1019 11114 1021
rect 10386 1013 10450 1019
rect 10386 986 10427 1013
rect 9973 614 9979 986
rect 10421 614 10427 986
rect 9973 587 10014 614
rect 9950 581 10014 587
rect 9286 579 9319 581
rect 8881 573 9319 579
rect 8881 556 8887 573
rect 9313 556 9319 573
rect 8881 550 9319 556
rect 9429 579 9871 581
rect 9431 573 9869 579
rect 9431 556 9437 573
rect 9863 556 9869 573
rect 9431 550 9869 556
rect 9981 579 10014 581
rect 10386 587 10427 614
rect 10444 587 10450 1013
rect 10386 581 10450 587
rect 10500 1013 11000 1019
rect 10500 587 10506 1013
rect 10523 965 10977 1013
rect 10523 635 10585 965
rect 10915 635 10977 965
rect 10523 587 10977 635
rect 10994 587 11000 1013
rect 10500 581 11000 587
rect 11050 1013 11114 1019
rect 11050 587 11056 1013
rect 11073 986 11114 1013
rect 11486 1019 11519 1021
rect 11631 1044 12069 1050
rect 11631 1027 11637 1044
rect 12063 1027 12069 1044
rect 11631 1021 12069 1027
rect 11629 1019 12071 1021
rect 12181 1044 12619 1050
rect 12181 1027 12187 1044
rect 12613 1027 12619 1044
rect 12181 1021 12619 1027
rect 12181 1019 12214 1021
rect 11486 1013 11550 1019
rect 11486 986 11527 1013
rect 11073 614 11079 986
rect 11521 614 11527 986
rect 11073 587 11114 614
rect 11050 581 11114 587
rect 10386 579 10419 581
rect 9981 573 10419 579
rect 9981 556 9987 573
rect 10413 556 10419 573
rect 9981 550 10419 556
rect 10529 579 10971 581
rect 10531 573 10969 579
rect 10531 556 10537 573
rect 10963 556 10969 573
rect 10531 550 10969 556
rect 11081 579 11114 581
rect 11486 587 11527 614
rect 11544 587 11550 1013
rect 11486 581 11550 587
rect 11600 1013 12100 1019
rect 11600 587 11606 1013
rect 11623 965 12077 1013
rect 11623 635 11685 965
rect 12015 635 12077 965
rect 11623 587 12077 635
rect 12094 587 12100 1013
rect 11600 581 12100 587
rect 12150 1013 12214 1019
rect 12150 587 12156 1013
rect 12173 986 12214 1013
rect 12586 1019 12619 1021
rect 12731 1044 13169 1050
rect 12731 1027 12737 1044
rect 13163 1027 13169 1044
rect 12731 1021 13169 1027
rect 12729 1019 13171 1021
rect 13281 1044 13719 1050
rect 13281 1027 13287 1044
rect 13713 1027 13719 1044
rect 13281 1021 13719 1027
rect 13281 1019 13314 1021
rect 12586 1013 12650 1019
rect 12586 986 12627 1013
rect 12173 614 12179 986
rect 12621 614 12627 986
rect 12173 587 12214 614
rect 12150 581 12214 587
rect 11486 579 11519 581
rect 11081 573 11519 579
rect 11081 556 11087 573
rect 11513 556 11519 573
rect 11081 550 11519 556
rect 11629 579 12071 581
rect 11631 573 12069 579
rect 11631 556 11637 573
rect 12063 556 12069 573
rect 11631 550 12069 556
rect 12181 579 12214 581
rect 12586 587 12627 614
rect 12644 587 12650 1013
rect 12586 581 12650 587
rect 12700 1013 13200 1019
rect 12700 587 12706 1013
rect 12723 965 13177 1013
rect 12723 635 12785 965
rect 13115 635 13177 965
rect 12723 587 13177 635
rect 13194 587 13200 1013
rect 12700 581 13200 587
rect 13250 1013 13314 1019
rect 13250 587 13256 1013
rect 13273 986 13314 1013
rect 13273 614 13279 986
rect 13273 587 13314 614
rect 13250 581 13314 587
rect 12586 579 12619 581
rect 12181 573 12619 579
rect 12181 556 12187 573
rect 12613 556 12619 573
rect 12181 550 12619 556
rect 12729 579 13171 581
rect 12731 573 13169 579
rect 12731 556 12737 573
rect 13163 556 13169 573
rect 12731 550 13169 556
rect 13281 579 13314 581
rect 13281 573 13719 579
rect 13281 556 13287 573
rect 13713 556 13719 573
rect 13281 550 13719 556
rect -469 494 -31 500
rect -469 477 -463 494
rect -37 477 -31 494
rect -469 471 -31 477
rect -64 469 -31 471
rect 81 494 519 500
rect 81 477 87 494
rect 513 477 519 494
rect 81 471 519 477
rect 79 469 521 471
rect 631 494 1069 500
rect 631 477 637 494
rect 1063 477 1069 494
rect 631 471 1069 477
rect 631 469 664 471
rect -64 463 0 469
rect -64 436 -23 463
rect -29 64 -23 436
rect -64 37 -23 64
rect -6 37 0 463
rect -64 31 0 37
rect 50 463 550 469
rect 50 37 56 463
rect 73 415 527 463
rect 73 85 135 415
rect 465 85 527 415
rect 73 37 527 85
rect 544 37 550 463
rect 50 31 550 37
rect 600 463 664 469
rect 600 37 606 463
rect 623 436 664 463
rect 1036 469 1069 471
rect 1181 494 1619 500
rect 1181 477 1187 494
rect 1613 477 1619 494
rect 1181 471 1619 477
rect 1179 469 1621 471
rect 1731 494 2169 500
rect 1731 477 1737 494
rect 2163 477 2169 494
rect 1731 471 2169 477
rect 1731 469 1764 471
rect 1036 463 1100 469
rect 1036 436 1077 463
rect 623 64 629 436
rect 1071 64 1077 436
rect 623 37 664 64
rect 600 31 664 37
rect -64 29 -31 31
rect -469 23 -31 29
rect -469 6 -463 23
rect -37 6 -31 23
rect -469 0 -31 6
rect 79 29 521 31
rect 81 23 519 29
rect 81 6 87 23
rect 513 6 519 23
rect 81 0 519 6
rect 631 29 664 31
rect 1036 37 1077 64
rect 1094 37 1100 463
rect 1036 31 1100 37
rect 1150 463 1650 469
rect 1150 37 1156 463
rect 1173 415 1627 463
rect 1173 85 1235 415
rect 1565 85 1627 415
rect 1173 37 1627 85
rect 1644 37 1650 463
rect 1150 31 1650 37
rect 1700 463 1764 469
rect 1700 37 1706 463
rect 1723 436 1764 463
rect 2136 469 2169 471
rect 2281 494 2719 500
rect 2281 477 2287 494
rect 2713 477 2719 494
rect 2281 471 2719 477
rect 2279 469 2721 471
rect 2831 494 3269 500
rect 2831 477 2837 494
rect 3263 477 3269 494
rect 2831 471 3269 477
rect 2831 469 2864 471
rect 2136 463 2200 469
rect 2136 436 2177 463
rect 1723 64 1729 436
rect 2171 64 2177 436
rect 1723 37 1764 64
rect 1700 31 1764 37
rect 1036 29 1069 31
rect 631 23 1069 29
rect 631 6 637 23
rect 1063 6 1069 23
rect 631 0 1069 6
rect 1179 29 1621 31
rect 1181 23 1619 29
rect 1181 6 1187 23
rect 1613 6 1619 23
rect 1181 0 1619 6
rect 1731 29 1764 31
rect 2136 37 2177 64
rect 2194 37 2200 463
rect 2136 31 2200 37
rect 2250 463 2750 469
rect 2250 37 2256 463
rect 2273 415 2727 463
rect 2273 85 2335 415
rect 2665 85 2727 415
rect 2273 37 2727 85
rect 2744 37 2750 463
rect 2250 31 2750 37
rect 2800 463 2864 469
rect 2800 37 2806 463
rect 2823 436 2864 463
rect 3236 469 3269 471
rect 3381 494 3819 500
rect 3381 477 3387 494
rect 3813 477 3819 494
rect 3381 471 3819 477
rect 3379 469 3821 471
rect 3931 494 4369 500
rect 3931 477 3937 494
rect 4363 477 4369 494
rect 3931 471 4369 477
rect 3931 469 3964 471
rect 3236 463 3300 469
rect 3236 436 3277 463
rect 2823 64 2829 436
rect 3271 64 3277 436
rect 2823 37 2864 64
rect 2800 31 2864 37
rect 2136 29 2169 31
rect 1731 23 2169 29
rect 1731 6 1737 23
rect 2163 6 2169 23
rect 1731 0 2169 6
rect 2279 29 2721 31
rect 2281 23 2719 29
rect 2281 6 2287 23
rect 2713 6 2719 23
rect 2281 0 2719 6
rect 2831 29 2864 31
rect 3236 37 3277 64
rect 3294 37 3300 463
rect 3236 31 3300 37
rect 3350 463 3850 469
rect 3350 37 3356 463
rect 3373 415 3827 463
rect 3373 85 3435 415
rect 3765 85 3827 415
rect 3373 37 3827 85
rect 3844 37 3850 463
rect 3350 31 3850 37
rect 3900 463 3964 469
rect 3900 37 3906 463
rect 3923 436 3964 463
rect 4336 469 4369 471
rect 4481 494 4919 500
rect 4481 477 4487 494
rect 4913 477 4919 494
rect 4481 471 4919 477
rect 4479 469 4921 471
rect 5031 494 5469 500
rect 5031 477 5037 494
rect 5463 477 5469 494
rect 5031 471 5469 477
rect 5031 469 5064 471
rect 4336 463 4400 469
rect 4336 436 4377 463
rect 3923 64 3929 436
rect 4371 64 4377 436
rect 3923 37 3964 64
rect 3900 31 3964 37
rect 3236 29 3269 31
rect 2831 23 3269 29
rect 2831 6 2837 23
rect 3263 6 3269 23
rect 2831 0 3269 6
rect 3379 29 3821 31
rect 3381 23 3819 29
rect 3381 6 3387 23
rect 3813 6 3819 23
rect 3381 0 3819 6
rect 3931 29 3964 31
rect 4336 37 4377 64
rect 4394 37 4400 463
rect 4336 31 4400 37
rect 4450 463 4950 469
rect 4450 37 4456 463
rect 4473 415 4927 463
rect 4473 85 4535 415
rect 4865 85 4927 415
rect 4473 37 4927 85
rect 4944 37 4950 463
rect 4450 31 4950 37
rect 5000 463 5064 469
rect 5000 37 5006 463
rect 5023 436 5064 463
rect 5436 469 5469 471
rect 5581 494 6019 500
rect 5581 477 5587 494
rect 6013 477 6019 494
rect 5581 471 6019 477
rect 5579 469 6021 471
rect 6131 494 6569 500
rect 6131 477 6137 494
rect 6563 477 6569 494
rect 6131 471 6569 477
rect 6131 469 6164 471
rect 5436 463 5500 469
rect 5436 436 5477 463
rect 5023 64 5029 436
rect 5471 64 5477 436
rect 5023 37 5064 64
rect 5000 31 5064 37
rect 4336 29 4369 31
rect 3931 23 4369 29
rect 3931 6 3937 23
rect 4363 6 4369 23
rect 3931 0 4369 6
rect 4479 29 4921 31
rect 4481 23 4919 29
rect 4481 6 4487 23
rect 4913 6 4919 23
rect 4481 0 4919 6
rect 5031 29 5064 31
rect 5436 37 5477 64
rect 5494 37 5500 463
rect 5436 31 5500 37
rect 5550 463 6050 469
rect 5550 37 5556 463
rect 5573 415 6027 463
rect 5573 85 5635 415
rect 5965 85 6027 415
rect 5573 37 6027 85
rect 6044 37 6050 463
rect 5550 31 6050 37
rect 6100 463 6164 469
rect 6100 37 6106 463
rect 6123 436 6164 463
rect 6536 469 6569 471
rect 6681 494 7119 500
rect 6681 477 6687 494
rect 7113 477 7119 494
rect 6681 471 7119 477
rect 6679 469 7121 471
rect 7231 494 7669 500
rect 7231 477 7237 494
rect 7663 477 7669 494
rect 7231 471 7669 477
rect 7231 469 7264 471
rect 6536 463 6600 469
rect 6536 436 6577 463
rect 6123 64 6129 436
rect 6571 64 6577 436
rect 6123 37 6164 64
rect 6100 31 6164 37
rect 5436 29 5469 31
rect 5031 23 5469 29
rect 5031 6 5037 23
rect 5463 6 5469 23
rect 5031 0 5469 6
rect 5579 29 6021 31
rect 5581 23 6019 29
rect 5581 6 5587 23
rect 6013 6 6019 23
rect 5581 0 6019 6
rect 6131 29 6164 31
rect 6536 37 6577 64
rect 6594 37 6600 463
rect 6536 31 6600 37
rect 6650 463 7150 469
rect 6650 37 6656 463
rect 6673 415 7127 463
rect 6673 85 6735 415
rect 7065 85 7127 415
rect 6673 37 7127 85
rect 7144 37 7150 463
rect 6650 31 7150 37
rect 7200 463 7264 469
rect 7200 37 7206 463
rect 7223 436 7264 463
rect 7636 469 7669 471
rect 7781 494 8219 500
rect 7781 477 7787 494
rect 8213 477 8219 494
rect 7781 471 8219 477
rect 7779 469 8221 471
rect 8331 494 8769 500
rect 8331 477 8337 494
rect 8763 477 8769 494
rect 8331 471 8769 477
rect 8331 469 8364 471
rect 7636 463 7700 469
rect 7636 436 7677 463
rect 7223 64 7229 436
rect 7671 64 7677 436
rect 7223 37 7264 64
rect 7200 31 7264 37
rect 6536 29 6569 31
rect 6131 23 6569 29
rect 6131 6 6137 23
rect 6563 6 6569 23
rect 6131 0 6569 6
rect 6679 29 7121 31
rect 6681 23 7119 29
rect 6681 6 6687 23
rect 7113 6 7119 23
rect 6681 0 7119 6
rect 7231 29 7264 31
rect 7636 37 7677 64
rect 7694 37 7700 463
rect 7636 31 7700 37
rect 7750 463 8250 469
rect 7750 37 7756 463
rect 7773 415 8227 463
rect 7773 85 7835 415
rect 8165 85 8227 415
rect 7773 37 8227 85
rect 8244 37 8250 463
rect 7750 31 8250 37
rect 8300 463 8364 469
rect 8300 37 8306 463
rect 8323 436 8364 463
rect 8736 469 8769 471
rect 8881 494 9319 500
rect 8881 477 8887 494
rect 9313 477 9319 494
rect 8881 471 9319 477
rect 8879 469 9321 471
rect 9431 494 9869 500
rect 9431 477 9437 494
rect 9863 477 9869 494
rect 9431 471 9869 477
rect 9431 469 9464 471
rect 8736 463 8800 469
rect 8736 436 8777 463
rect 8323 64 8329 436
rect 8771 64 8777 436
rect 8323 37 8364 64
rect 8300 31 8364 37
rect 7636 29 7669 31
rect 7231 23 7669 29
rect 7231 6 7237 23
rect 7663 6 7669 23
rect 7231 0 7669 6
rect 7779 29 8221 31
rect 7781 23 8219 29
rect 7781 6 7787 23
rect 8213 6 8219 23
rect 7781 0 8219 6
rect 8331 29 8364 31
rect 8736 37 8777 64
rect 8794 37 8800 463
rect 8736 31 8800 37
rect 8850 463 9350 469
rect 8850 37 8856 463
rect 8873 415 9327 463
rect 8873 85 8935 415
rect 9265 85 9327 415
rect 8873 37 9327 85
rect 9344 37 9350 463
rect 8850 31 9350 37
rect 9400 463 9464 469
rect 9400 37 9406 463
rect 9423 436 9464 463
rect 9836 469 9869 471
rect 9981 494 10419 500
rect 9981 477 9987 494
rect 10413 477 10419 494
rect 9981 471 10419 477
rect 9979 469 10421 471
rect 10531 494 10969 500
rect 10531 477 10537 494
rect 10963 477 10969 494
rect 10531 471 10969 477
rect 10531 469 10564 471
rect 9836 463 9900 469
rect 9836 436 9877 463
rect 9423 64 9429 436
rect 9871 64 9877 436
rect 9423 37 9464 64
rect 9400 31 9464 37
rect 8736 29 8769 31
rect 8331 23 8769 29
rect 8331 6 8337 23
rect 8763 6 8769 23
rect 8331 0 8769 6
rect 8879 29 9321 31
rect 8881 23 9319 29
rect 8881 6 8887 23
rect 9313 6 9319 23
rect 8881 0 9319 6
rect 9431 29 9464 31
rect 9836 37 9877 64
rect 9894 37 9900 463
rect 9836 31 9900 37
rect 9950 463 10450 469
rect 9950 37 9956 463
rect 9973 415 10427 463
rect 9973 85 10035 415
rect 10365 85 10427 415
rect 9973 37 10427 85
rect 10444 37 10450 463
rect 9950 31 10450 37
rect 10500 463 10564 469
rect 10500 37 10506 463
rect 10523 436 10564 463
rect 10936 469 10969 471
rect 11081 494 11519 500
rect 11081 477 11087 494
rect 11513 477 11519 494
rect 11081 471 11519 477
rect 11079 469 11521 471
rect 11631 494 12069 500
rect 11631 477 11637 494
rect 12063 477 12069 494
rect 11631 471 12069 477
rect 11631 469 11664 471
rect 10936 463 11000 469
rect 10936 436 10977 463
rect 10523 64 10529 436
rect 10971 64 10977 436
rect 10523 37 10564 64
rect 10500 31 10564 37
rect 9836 29 9869 31
rect 9431 23 9869 29
rect 9431 6 9437 23
rect 9863 6 9869 23
rect 9431 0 9869 6
rect 9979 29 10421 31
rect 9981 23 10419 29
rect 9981 6 9987 23
rect 10413 6 10419 23
rect 9981 0 10419 6
rect 10531 29 10564 31
rect 10936 37 10977 64
rect 10994 37 11000 463
rect 10936 31 11000 37
rect 11050 463 11550 469
rect 11050 37 11056 463
rect 11073 415 11527 463
rect 11073 85 11135 415
rect 11465 85 11527 415
rect 11073 37 11527 85
rect 11544 37 11550 463
rect 11050 31 11550 37
rect 11600 463 11664 469
rect 11600 37 11606 463
rect 11623 436 11664 463
rect 12036 469 12069 471
rect 12181 494 12619 500
rect 12181 477 12187 494
rect 12613 477 12619 494
rect 12181 471 12619 477
rect 12179 469 12621 471
rect 12731 494 13169 500
rect 12731 477 12737 494
rect 13163 477 13169 494
rect 12731 471 13169 477
rect 12731 469 12764 471
rect 12036 463 12100 469
rect 12036 436 12077 463
rect 11623 64 11629 436
rect 12071 64 12077 436
rect 11623 37 11664 64
rect 11600 31 11664 37
rect 10936 29 10969 31
rect 10531 23 10969 29
rect 10531 6 10537 23
rect 10963 6 10969 23
rect 10531 0 10969 6
rect 11079 29 11521 31
rect 11081 23 11519 29
rect 11081 6 11087 23
rect 11513 6 11519 23
rect 11081 0 11519 6
rect 11631 29 11664 31
rect 12036 37 12077 64
rect 12094 37 12100 463
rect 12036 31 12100 37
rect 12150 463 12650 469
rect 12150 37 12156 463
rect 12173 415 12627 463
rect 12173 85 12235 415
rect 12565 85 12627 415
rect 12173 37 12627 85
rect 12644 37 12650 463
rect 12150 31 12650 37
rect 12700 463 12764 469
rect 12700 37 12706 463
rect 12723 436 12764 463
rect 13136 469 13169 471
rect 13281 494 13719 500
rect 13281 477 13287 494
rect 13713 477 13719 494
rect 13281 471 13719 477
rect 13279 469 13721 471
rect 13136 463 13200 469
rect 13136 436 13177 463
rect 12723 64 12729 436
rect 13171 64 13177 436
rect 12723 37 12764 64
rect 12700 31 12764 37
rect 12036 29 12069 31
rect 11631 23 12069 29
rect 11631 6 11637 23
rect 12063 6 12069 23
rect 11631 0 12069 6
rect 12179 29 12621 31
rect 12181 23 12619 29
rect 12181 6 12187 23
rect 12613 6 12619 23
rect 12181 0 12619 6
rect 12731 29 12764 31
rect 13136 37 13177 64
rect 13194 37 13200 463
rect 13136 31 13200 37
rect 13250 463 13721 469
rect 13250 37 13256 463
rect 13273 415 13721 463
rect 13273 85 13335 415
rect 13665 85 13721 415
rect 13273 37 13721 85
rect 13250 31 13721 37
rect 13136 29 13169 31
rect 12731 23 13169 29
rect 12731 6 12737 23
rect 13163 6 13169 23
rect 12731 0 13169 6
rect 13279 29 13721 31
rect 13281 23 13719 29
rect 13281 6 13287 23
rect 13713 6 13719 23
rect 13281 0 13719 6
rect -469 -56 -31 -50
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -79 -31 -73
rect -471 -81 -29 -79
rect 81 -56 519 -50
rect 81 -73 87 -56
rect 513 -73 519 -56
rect 81 -79 519 -73
rect 81 -81 114 -79
rect -471 -87 0 -81
rect -471 -135 -23 -87
rect -471 -465 -415 -135
rect -85 -465 -23 -135
rect -471 -513 -23 -465
rect -6 -513 0 -87
rect -471 -519 0 -513
rect 50 -87 114 -81
rect 50 -513 56 -87
rect 73 -114 114 -87
rect 486 -81 519 -79
rect 631 -56 1069 -50
rect 631 -73 637 -56
rect 1063 -73 1069 -56
rect 631 -79 1069 -73
rect 629 -81 1071 -79
rect 1181 -56 1619 -50
rect 1181 -73 1187 -56
rect 1613 -73 1619 -56
rect 1181 -79 1619 -73
rect 1181 -81 1214 -79
rect 486 -87 550 -81
rect 486 -114 527 -87
rect 73 -513 79 -114
rect 50 -519 79 -513
rect 521 -513 527 -114
rect 544 -513 550 -87
rect 521 -519 550 -513
rect 600 -87 1100 -81
rect 600 -513 606 -87
rect 623 -135 1077 -87
rect 623 -465 685 -135
rect 1015 -465 1077 -135
rect 623 -513 1077 -465
rect 1094 -513 1100 -87
rect 600 -519 1100 -513
rect 1150 -87 1214 -81
rect 1150 -513 1156 -87
rect 1173 -114 1214 -87
rect 1586 -81 1619 -79
rect 1731 -56 2169 -50
rect 1731 -73 1737 -56
rect 2163 -73 2169 -56
rect 1731 -79 2169 -73
rect 1729 -81 2171 -79
rect 2281 -56 2719 -50
rect 2281 -73 2287 -56
rect 2713 -73 2719 -56
rect 2281 -79 2719 -73
rect 2281 -81 2314 -79
rect 1586 -87 1650 -81
rect 1586 -114 1627 -87
rect 1173 -513 1179 -114
rect 1150 -519 1179 -513
rect 1621 -513 1627 -114
rect 1644 -513 1650 -87
rect 1621 -519 1650 -513
rect 1700 -87 2200 -81
rect 1700 -513 1706 -87
rect 1723 -135 2177 -87
rect 1723 -465 1785 -135
rect 2115 -465 2177 -135
rect 1723 -513 2177 -465
rect 2194 -513 2200 -87
rect 1700 -519 2200 -513
rect 2250 -87 2314 -81
rect 2250 -513 2256 -87
rect 2273 -114 2314 -87
rect 2686 -81 2719 -79
rect 2831 -56 3269 -50
rect 2831 -73 2837 -56
rect 3263 -73 3269 -56
rect 2831 -79 3269 -73
rect 2829 -81 3271 -79
rect 3381 -56 3819 -50
rect 3381 -73 3387 -56
rect 3813 -73 3819 -56
rect 3381 -79 3819 -73
rect 3381 -81 3414 -79
rect 2686 -87 2750 -81
rect 2686 -114 2727 -87
rect 2273 -513 2279 -114
rect 2250 -519 2279 -513
rect 2721 -513 2727 -114
rect 2744 -513 2750 -87
rect 2721 -519 2750 -513
rect 2800 -87 3300 -81
rect 2800 -513 2806 -87
rect 2823 -135 3277 -87
rect 2823 -465 2885 -135
rect 3215 -465 3277 -135
rect 2823 -513 3277 -465
rect 3294 -513 3300 -87
rect 2800 -519 3300 -513
rect 3350 -87 3414 -81
rect 3350 -513 3356 -87
rect 3373 -114 3414 -87
rect 3786 -81 3819 -79
rect 3931 -56 4369 -50
rect 3931 -73 3937 -56
rect 4363 -73 4369 -56
rect 3931 -79 4369 -73
rect 3929 -81 4371 -79
rect 4481 -56 4919 -50
rect 4481 -73 4487 -56
rect 4913 -73 4919 -56
rect 4481 -79 4919 -73
rect 4481 -81 4514 -79
rect 3786 -87 3850 -81
rect 3786 -114 3827 -87
rect 3373 -513 3379 -114
rect 3350 -519 3379 -513
rect 3821 -513 3827 -114
rect 3844 -513 3850 -87
rect 3821 -519 3850 -513
rect 3900 -87 4400 -81
rect 3900 -513 3906 -87
rect 3923 -135 4377 -87
rect 3923 -465 3985 -135
rect 4315 -465 4377 -135
rect 3923 -513 4377 -465
rect 4394 -513 4400 -87
rect 3900 -519 4400 -513
rect 4450 -87 4514 -81
rect 4450 -513 4456 -87
rect 4473 -114 4514 -87
rect 4886 -81 4919 -79
rect 5031 -56 5469 -50
rect 5031 -73 5037 -56
rect 5463 -73 5469 -56
rect 5031 -79 5469 -73
rect 5029 -81 5471 -79
rect 5581 -56 6019 -50
rect 5581 -73 5587 -56
rect 6013 -73 6019 -56
rect 5581 -79 6019 -73
rect 5581 -81 5614 -79
rect 4886 -87 4950 -81
rect 4886 -114 4927 -87
rect 4473 -513 4479 -114
rect 4450 -519 4479 -513
rect 4921 -513 4927 -114
rect 4944 -513 4950 -87
rect 4921 -519 4950 -513
rect 5000 -87 5500 -81
rect 5000 -513 5006 -87
rect 5023 -135 5477 -87
rect 5023 -465 5085 -135
rect 5415 -465 5477 -135
rect 5023 -513 5477 -465
rect 5494 -513 5500 -87
rect 5000 -519 5500 -513
rect 5550 -87 5614 -81
rect 5550 -513 5556 -87
rect 5573 -114 5614 -87
rect 5986 -81 6019 -79
rect 6131 -56 6569 -50
rect 6131 -73 6137 -56
rect 6563 -73 6569 -56
rect 6131 -79 6569 -73
rect 6129 -81 6571 -79
rect 6681 -56 7119 -50
rect 6681 -73 6687 -56
rect 7113 -73 7119 -56
rect 6681 -79 7119 -73
rect 6681 -81 6714 -79
rect 5986 -87 6050 -81
rect 5986 -114 6027 -87
rect 5573 -513 5579 -114
rect 5550 -519 5579 -513
rect 6021 -513 6027 -114
rect 6044 -513 6050 -87
rect 6021 -519 6050 -513
rect 6100 -87 6600 -81
rect 6100 -513 6106 -87
rect 6123 -135 6577 -87
rect 6123 -465 6185 -135
rect 6515 -465 6577 -135
rect 6123 -513 6577 -465
rect 6594 -513 6600 -87
rect 6100 -519 6600 -513
rect 6650 -87 6714 -81
rect 6650 -513 6656 -87
rect 6673 -114 6714 -87
rect 7086 -81 7119 -79
rect 7231 -56 7669 -50
rect 7231 -73 7237 -56
rect 7663 -73 7669 -56
rect 7231 -79 7669 -73
rect 7229 -81 7671 -79
rect 7781 -56 8219 -50
rect 7781 -73 7787 -56
rect 8213 -73 8219 -56
rect 7781 -79 8219 -73
rect 7781 -81 7814 -79
rect 7086 -87 7150 -81
rect 7086 -114 7127 -87
rect 6673 -513 6679 -114
rect 6650 -519 6679 -513
rect 7121 -513 7127 -114
rect 7144 -513 7150 -87
rect 7121 -519 7150 -513
rect 7200 -87 7700 -81
rect 7200 -513 7206 -87
rect 7223 -135 7677 -87
rect 7223 -465 7285 -135
rect 7615 -465 7677 -135
rect 7223 -513 7677 -465
rect 7694 -513 7700 -87
rect 7200 -519 7700 -513
rect 7750 -87 7814 -81
rect 7750 -513 7756 -87
rect 7773 -114 7814 -87
rect 8186 -81 8219 -79
rect 8331 -56 8769 -50
rect 8331 -73 8337 -56
rect 8763 -73 8769 -56
rect 8331 -79 8769 -73
rect 8329 -81 8771 -79
rect 8881 -56 9319 -50
rect 8881 -73 8887 -56
rect 9313 -73 9319 -56
rect 8881 -79 9319 -73
rect 8881 -81 8914 -79
rect 8186 -87 8250 -81
rect 8186 -114 8227 -87
rect 7773 -513 7779 -114
rect 7750 -519 7779 -513
rect 8221 -513 8227 -114
rect 8244 -513 8250 -87
rect 8221 -519 8250 -513
rect 8300 -87 8800 -81
rect 8300 -513 8306 -87
rect 8323 -135 8777 -87
rect 8323 -465 8385 -135
rect 8715 -465 8777 -135
rect 8323 -513 8777 -465
rect 8794 -513 8800 -87
rect 8300 -519 8800 -513
rect 8850 -87 8914 -81
rect 8850 -513 8856 -87
rect 8873 -114 8914 -87
rect 9286 -81 9319 -79
rect 9431 -56 9869 -50
rect 9431 -73 9437 -56
rect 9863 -73 9869 -56
rect 9431 -79 9869 -73
rect 9429 -81 9871 -79
rect 9981 -56 10419 -50
rect 9981 -73 9987 -56
rect 10413 -73 10419 -56
rect 9981 -79 10419 -73
rect 9981 -81 10014 -79
rect 9286 -87 9350 -81
rect 9286 -114 9327 -87
rect 8873 -513 8879 -114
rect 8850 -519 8879 -513
rect 9321 -513 9327 -114
rect 9344 -513 9350 -87
rect 9321 -519 9350 -513
rect 9400 -87 9900 -81
rect 9400 -513 9406 -87
rect 9423 -135 9877 -87
rect 9423 -465 9485 -135
rect 9815 -465 9877 -135
rect 9423 -513 9877 -465
rect 9894 -513 9900 -87
rect 9400 -519 9900 -513
rect 9950 -87 10014 -81
rect 9950 -513 9956 -87
rect 9973 -114 10014 -87
rect 10386 -81 10419 -79
rect 10531 -56 10969 -50
rect 10531 -73 10537 -56
rect 10963 -73 10969 -56
rect 10531 -79 10969 -73
rect 10529 -81 10971 -79
rect 11081 -56 11519 -50
rect 11081 -73 11087 -56
rect 11513 -73 11519 -56
rect 11081 -79 11519 -73
rect 11081 -81 11114 -79
rect 10386 -87 10450 -81
rect 10386 -114 10427 -87
rect 9973 -513 9979 -114
rect 9950 -519 9979 -513
rect 10421 -513 10427 -114
rect 10444 -513 10450 -87
rect 10421 -519 10450 -513
rect 10500 -87 11000 -81
rect 10500 -513 10506 -87
rect 10523 -135 10977 -87
rect 10523 -465 10585 -135
rect 10915 -465 10977 -135
rect 10523 -513 10977 -465
rect 10994 -513 11000 -87
rect 10500 -519 11000 -513
rect 11050 -87 11114 -81
rect 11050 -513 11056 -87
rect 11073 -114 11114 -87
rect 11486 -81 11519 -79
rect 11631 -56 12069 -50
rect 11631 -73 11637 -56
rect 12063 -73 12069 -56
rect 11631 -79 12069 -73
rect 11629 -81 12071 -79
rect 12181 -56 12619 -50
rect 12181 -73 12187 -56
rect 12613 -73 12619 -56
rect 12181 -79 12619 -73
rect 12181 -81 12214 -79
rect 11486 -87 11550 -81
rect 11486 -114 11527 -87
rect 11073 -513 11079 -114
rect 11050 -519 11079 -513
rect 11521 -513 11527 -114
rect 11544 -513 11550 -87
rect 11521 -519 11550 -513
rect 11600 -87 12100 -81
rect 11600 -513 11606 -87
rect 11623 -135 12077 -87
rect 11623 -465 11685 -135
rect 12015 -465 12077 -135
rect 11623 -513 12077 -465
rect 12094 -513 12100 -87
rect 11600 -519 12100 -513
rect 12150 -87 12214 -81
rect 12150 -513 12156 -87
rect 12173 -114 12214 -87
rect 12586 -81 12619 -79
rect 12731 -56 13169 -50
rect 12731 -73 12737 -56
rect 13163 -73 13169 -56
rect 12731 -79 13169 -73
rect 12729 -81 13171 -79
rect 13281 -56 13719 -50
rect 13281 -73 13287 -56
rect 13713 -73 13719 -56
rect 13281 -79 13719 -73
rect 13281 -81 13314 -79
rect 12586 -87 12650 -81
rect 12586 -114 12627 -87
rect 12173 -513 12179 -114
rect 12150 -519 12179 -513
rect 12621 -513 12627 -114
rect 12644 -513 12650 -87
rect 12621 -519 12650 -513
rect 12700 -87 13200 -81
rect 12700 -513 12706 -87
rect 12723 -135 13177 -87
rect 12723 -465 12785 -135
rect 13115 -465 13177 -135
rect 12723 -513 13177 -465
rect 13194 -513 13200 -87
rect 12700 -519 13200 -513
rect 13250 -87 13314 -81
rect 13250 -513 13256 -87
rect 13273 -114 13314 -87
rect 13273 -513 13279 -114
rect 13250 -519 13279 -513
rect -471 -521 -29 -519
rect 629 -521 1071 -519
rect 1729 -521 2171 -519
rect 2829 -521 3271 -519
rect 3929 -521 4371 -519
rect 5029 -521 5471 -519
rect 6129 -521 6571 -519
rect 7229 -521 7671 -519
rect 8329 -521 8771 -519
rect 9429 -521 9871 -519
rect 10529 -521 10971 -519
rect 11629 -521 12071 -519
rect 12729 -521 13171 -519
<< mvpdiffc >>
rect -23 13237 -6 13663
rect 56 13237 73 13663
rect 527 13237 544 13663
rect 606 13237 623 13663
rect -463 13206 -37 13223
rect 87 13206 513 13223
rect 1077 13237 1094 13663
rect 1156 13237 1173 13663
rect 1627 13237 1644 13663
rect 1706 13237 1723 13663
rect 637 13206 1063 13223
rect 1187 13206 1613 13223
rect 2177 13237 2194 13663
rect 2256 13237 2273 13663
rect 2727 13237 2744 13663
rect 2806 13237 2823 13663
rect 1737 13206 2163 13223
rect 2287 13206 2713 13223
rect 3277 13237 3294 13663
rect 3356 13237 3373 13663
rect 3827 13237 3844 13663
rect 3906 13237 3923 13663
rect 2837 13206 3263 13223
rect 3387 13206 3813 13223
rect 4377 13237 4394 13663
rect 4456 13237 4473 13663
rect 4927 13237 4944 13663
rect 5006 13237 5023 13663
rect 3937 13206 4363 13223
rect 4487 13206 4913 13223
rect 5477 13237 5494 13663
rect 5556 13237 5573 13663
rect 6027 13237 6044 13663
rect 6106 13237 6123 13663
rect 5037 13206 5463 13223
rect 5587 13206 6013 13223
rect 6577 13237 6594 13663
rect 6656 13237 6673 13663
rect 7127 13237 7144 13663
rect 7206 13237 7223 13663
rect 6137 13206 6563 13223
rect 6687 13206 7113 13223
rect 7677 13237 7694 13663
rect 7756 13237 7773 13663
rect 8227 13237 8244 13663
rect 8306 13237 8323 13663
rect 7237 13206 7663 13223
rect 7787 13206 8213 13223
rect 8777 13237 8794 13663
rect 8856 13237 8873 13663
rect 9327 13237 9344 13663
rect 9406 13237 9423 13663
rect 8337 13206 8763 13223
rect 8887 13206 9313 13223
rect 9877 13237 9894 13663
rect 9956 13237 9973 13663
rect 10427 13237 10444 13663
rect 10506 13237 10523 13663
rect 9437 13206 9863 13223
rect 9987 13206 10413 13223
rect 10977 13237 10994 13663
rect 11056 13237 11073 13663
rect 11527 13237 11544 13663
rect 11606 13237 11623 13663
rect 10537 13206 10963 13223
rect 11087 13206 11513 13223
rect 12077 13237 12094 13663
rect 12156 13237 12173 13663
rect 12627 13237 12644 13663
rect 12706 13237 12723 13663
rect 11637 13206 12063 13223
rect 12187 13206 12613 13223
rect 13177 13237 13194 13663
rect 13256 13237 13273 13663
rect 12737 13206 13163 13223
rect 13287 13206 13713 13223
rect -463 13127 -37 13144
rect 87 13127 513 13144
rect -23 12687 -6 13113
rect 56 12687 73 13113
rect 637 13127 1063 13144
rect 1187 13127 1613 13144
rect -463 12656 -37 12673
rect 527 12687 544 13113
rect 606 12687 623 13113
rect 1077 12687 1094 13113
rect 1156 12687 1173 13113
rect 1737 13127 2163 13144
rect 2287 13127 2713 13144
rect 87 12656 513 12673
rect 637 12656 1063 12673
rect 1627 12687 1644 13113
rect 1706 12687 1723 13113
rect 2177 12687 2194 13113
rect 2256 12687 2273 13113
rect 2837 13127 3263 13144
rect 3387 13127 3813 13144
rect 1187 12656 1613 12673
rect 1737 12656 2163 12673
rect 2727 12687 2744 13113
rect 2806 12687 2823 13113
rect 3277 12687 3294 13113
rect 3356 12687 3373 13113
rect 3937 13127 4363 13144
rect 4487 13127 4913 13144
rect 2287 12656 2713 12673
rect 2837 12656 3263 12673
rect 3827 12687 3844 13113
rect 3906 12687 3923 13113
rect 4377 12687 4394 13113
rect 4456 12687 4473 13113
rect 5037 13127 5463 13144
rect 5587 13127 6013 13144
rect 3387 12656 3813 12673
rect 3937 12656 4363 12673
rect 4927 12687 4944 13113
rect 5006 12687 5023 13113
rect 5477 12687 5494 13113
rect 5556 12687 5573 13113
rect 6137 13127 6563 13144
rect 6687 13127 7113 13144
rect 4487 12656 4913 12673
rect 5037 12656 5463 12673
rect 6027 12687 6044 13113
rect 6106 12687 6123 13113
rect 6577 12687 6594 13113
rect 6656 12687 6673 13113
rect 7237 13127 7663 13144
rect 7787 13127 8213 13144
rect 5587 12656 6013 12673
rect 6137 12656 6563 12673
rect 7127 12687 7144 13113
rect 7206 12687 7223 13113
rect 7677 12687 7694 13113
rect 7756 12687 7773 13113
rect 8337 13127 8763 13144
rect 8887 13127 9313 13144
rect 6687 12656 7113 12673
rect 7237 12656 7663 12673
rect 8227 12687 8244 13113
rect 8306 12687 8323 13113
rect 8777 12687 8794 13113
rect 8856 12687 8873 13113
rect 9437 13127 9863 13144
rect 9987 13127 10413 13144
rect 7787 12656 8213 12673
rect 8337 12656 8763 12673
rect 9327 12687 9344 13113
rect 9406 12687 9423 13113
rect 9877 12687 9894 13113
rect 9956 12687 9973 13113
rect 10537 13127 10963 13144
rect 11087 13127 11513 13144
rect 8887 12656 9313 12673
rect 9437 12656 9863 12673
rect 10427 12687 10444 13113
rect 10506 12687 10523 13113
rect 10977 12687 10994 13113
rect 11056 12687 11073 13113
rect 11637 13127 12063 13144
rect 12187 13127 12613 13144
rect 9987 12656 10413 12673
rect 10537 12656 10963 12673
rect 11527 12687 11544 13113
rect 11606 12687 11623 13113
rect 12077 12687 12094 13113
rect 12156 12687 12173 13113
rect 12737 13127 13163 13144
rect 13287 13127 13713 13144
rect 11087 12656 11513 12673
rect 11637 12656 12063 12673
rect 12627 12687 12644 13113
rect 12706 12687 12723 13113
rect 13177 12687 13194 13113
rect 13256 12687 13273 13113
rect 12187 12656 12613 12673
rect 12737 12656 13163 12673
rect 13287 12656 13713 12673
rect -463 12577 -37 12594
rect 87 12577 513 12594
rect 637 12577 1063 12594
rect -23 12137 -6 12563
rect 56 12137 73 12563
rect 527 12137 544 12563
rect 606 12137 623 12563
rect 1187 12577 1613 12594
rect 1737 12577 2163 12594
rect -463 12106 -37 12123
rect 87 12106 513 12123
rect 1077 12137 1094 12563
rect 1156 12137 1173 12563
rect 1627 12137 1644 12563
rect 1706 12137 1723 12563
rect 2287 12577 2713 12594
rect 2837 12577 3263 12594
rect 637 12106 1063 12123
rect 1187 12106 1613 12123
rect 2177 12137 2194 12563
rect 2256 12137 2273 12563
rect 2727 12137 2744 12563
rect 2806 12137 2823 12563
rect 3387 12577 3813 12594
rect 3937 12577 4363 12594
rect 1737 12106 2163 12123
rect 2287 12106 2713 12123
rect 3277 12137 3294 12563
rect 3356 12137 3373 12563
rect 3827 12137 3844 12563
rect 3906 12137 3923 12563
rect 4487 12577 4913 12594
rect 5037 12577 5463 12594
rect 2837 12106 3263 12123
rect 3387 12106 3813 12123
rect 4377 12137 4394 12563
rect 4456 12137 4473 12563
rect 4927 12137 4944 12563
rect 5006 12137 5023 12563
rect 5587 12577 6013 12594
rect 6137 12577 6563 12594
rect 3937 12106 4363 12123
rect 4487 12106 4913 12123
rect 5477 12137 5494 12563
rect 5556 12137 5573 12563
rect 6027 12137 6044 12563
rect 6106 12137 6123 12563
rect 6687 12577 7113 12594
rect 7237 12577 7663 12594
rect 5037 12106 5463 12123
rect 5587 12106 6013 12123
rect 6577 12137 6594 12563
rect 6656 12137 6673 12563
rect 7127 12137 7144 12563
rect 7206 12137 7223 12563
rect 7787 12577 8213 12594
rect 8337 12577 8763 12594
rect 6137 12106 6563 12123
rect 6687 12106 7113 12123
rect 7677 12137 7694 12563
rect 7756 12137 7773 12563
rect 8227 12137 8244 12563
rect 8306 12137 8323 12563
rect 8887 12577 9313 12594
rect 9437 12577 9863 12594
rect 7237 12106 7663 12123
rect 7787 12106 8213 12123
rect 8777 12137 8794 12563
rect 8856 12137 8873 12563
rect 9327 12137 9344 12563
rect 9406 12137 9423 12563
rect 9987 12577 10413 12594
rect 10537 12577 10963 12594
rect 8337 12106 8763 12123
rect 8887 12106 9313 12123
rect 9877 12137 9894 12563
rect 9956 12137 9973 12563
rect 10427 12137 10444 12563
rect 10506 12137 10523 12563
rect 11087 12577 11513 12594
rect 11637 12577 12063 12594
rect 9437 12106 9863 12123
rect 9987 12106 10413 12123
rect 10977 12137 10994 12563
rect 11056 12137 11073 12563
rect 11527 12137 11544 12563
rect 11606 12137 11623 12563
rect 12187 12577 12613 12594
rect 12737 12577 13163 12594
rect 10537 12106 10963 12123
rect 11087 12106 11513 12123
rect 12077 12137 12094 12563
rect 12156 12137 12173 12563
rect 12627 12137 12644 12563
rect 12706 12137 12723 12563
rect 13287 12577 13713 12594
rect 11637 12106 12063 12123
rect 12187 12106 12613 12123
rect 13177 12137 13194 12563
rect 13256 12137 13273 12563
rect 12737 12106 13163 12123
rect 13287 12106 13713 12123
rect -463 12027 -37 12044
rect 87 12027 513 12044
rect -23 11587 -6 12013
rect 56 11587 73 12013
rect 637 12027 1063 12044
rect 1187 12027 1613 12044
rect -463 11556 -37 11573
rect 527 11587 544 12013
rect 606 11587 623 12013
rect 1077 11587 1094 12013
rect 1156 11587 1173 12013
rect 1737 12027 2163 12044
rect 2287 12027 2713 12044
rect 87 11556 513 11573
rect 637 11556 1063 11573
rect 1627 11587 1644 12013
rect 1706 11587 1723 12013
rect 2177 11587 2194 12013
rect 2256 11587 2273 12013
rect 2837 12027 3263 12044
rect 3387 12027 3813 12044
rect 1187 11556 1613 11573
rect 1737 11556 2163 11573
rect 2727 11587 2744 12013
rect 2806 11587 2823 12013
rect 3277 11587 3294 12013
rect 3356 11587 3373 12013
rect 3937 12027 4363 12044
rect 4487 12027 4913 12044
rect 2287 11556 2713 11573
rect 2837 11556 3263 11573
rect 3827 11587 3844 12013
rect 3906 11587 3923 12013
rect 4377 11587 4394 12013
rect 4456 11587 4473 12013
rect 5037 12027 5463 12044
rect 5587 12027 6013 12044
rect 3387 11556 3813 11573
rect 3937 11556 4363 11573
rect 4927 11587 4944 12013
rect 5006 11587 5023 12013
rect 5477 11587 5494 12013
rect 5556 11587 5573 12013
rect 6137 12027 6563 12044
rect 6687 12027 7113 12044
rect 4487 11556 4913 11573
rect 5037 11556 5463 11573
rect 6027 11587 6044 12013
rect 6106 11587 6123 12013
rect 6577 11587 6594 12013
rect 6656 11587 6673 12013
rect 7237 12027 7663 12044
rect 7787 12027 8213 12044
rect 5587 11556 6013 11573
rect 6137 11556 6563 11573
rect 7127 11587 7144 12013
rect 7206 11587 7223 12013
rect 7677 11587 7694 12013
rect 7756 11587 7773 12013
rect 8337 12027 8763 12044
rect 8887 12027 9313 12044
rect 6687 11556 7113 11573
rect 7237 11556 7663 11573
rect 8227 11587 8244 12013
rect 8306 11587 8323 12013
rect 8777 11587 8794 12013
rect 8856 11587 8873 12013
rect 9437 12027 9863 12044
rect 9987 12027 10413 12044
rect 7787 11556 8213 11573
rect 8337 11556 8763 11573
rect 9327 11587 9344 12013
rect 9406 11587 9423 12013
rect 9877 11587 9894 12013
rect 9956 11587 9973 12013
rect 10537 12027 10963 12044
rect 11087 12027 11513 12044
rect 8887 11556 9313 11573
rect 9437 11556 9863 11573
rect 10427 11587 10444 12013
rect 10506 11587 10523 12013
rect 10977 11587 10994 12013
rect 11056 11587 11073 12013
rect 11637 12027 12063 12044
rect 12187 12027 12613 12044
rect 9987 11556 10413 11573
rect 10537 11556 10963 11573
rect 11527 11587 11544 12013
rect 11606 11587 11623 12013
rect 12077 11587 12094 12013
rect 12156 11587 12173 12013
rect 12737 12027 13163 12044
rect 13287 12027 13713 12044
rect 11087 11556 11513 11573
rect 11637 11556 12063 11573
rect 12627 11587 12644 12013
rect 12706 11587 12723 12013
rect 13177 11587 13194 12013
rect 13256 11587 13273 12013
rect 12187 11556 12613 11573
rect 12737 11556 13163 11573
rect 13287 11556 13713 11573
rect -463 11477 -37 11494
rect 87 11477 513 11494
rect 637 11477 1063 11494
rect -23 11037 -6 11463
rect 56 11037 73 11463
rect 527 11037 544 11463
rect 606 11037 623 11463
rect 1187 11477 1613 11494
rect 1737 11477 2163 11494
rect -463 11006 -37 11023
rect 87 11006 513 11023
rect 1077 11037 1094 11463
rect 1156 11037 1173 11463
rect 1627 11037 1644 11463
rect 1706 11037 1723 11463
rect 2287 11477 2713 11494
rect 2837 11477 3263 11494
rect 637 11006 1063 11023
rect 1187 11006 1613 11023
rect 2177 11037 2194 11463
rect 2256 11037 2273 11463
rect 2727 11037 2744 11463
rect 2806 11037 2823 11463
rect 3387 11477 3813 11494
rect 3937 11477 4363 11494
rect 1737 11006 2163 11023
rect 2287 11006 2713 11023
rect 3277 11037 3294 11463
rect 3356 11037 3373 11463
rect 3827 11037 3844 11463
rect 3906 11037 3923 11463
rect 4487 11477 4913 11494
rect 5037 11477 5463 11494
rect 2837 11006 3263 11023
rect 3387 11006 3813 11023
rect 4377 11037 4394 11463
rect 4456 11037 4473 11463
rect 4927 11037 4944 11463
rect 5006 11037 5023 11463
rect 5587 11477 6013 11494
rect 6137 11477 6563 11494
rect 3937 11006 4363 11023
rect 4487 11006 4913 11023
rect 5477 11037 5494 11463
rect 5556 11037 5573 11463
rect 6027 11037 6044 11463
rect 6106 11037 6123 11463
rect 6687 11477 7113 11494
rect 7237 11477 7663 11494
rect 5037 11006 5463 11023
rect 5587 11006 6013 11023
rect 6577 11037 6594 11463
rect 6656 11037 6673 11463
rect 7127 11037 7144 11463
rect 7206 11037 7223 11463
rect 7787 11477 8213 11494
rect 8337 11477 8763 11494
rect 6137 11006 6563 11023
rect 6687 11006 7113 11023
rect 7677 11037 7694 11463
rect 7756 11037 7773 11463
rect 8227 11037 8244 11463
rect 8306 11037 8323 11463
rect 8887 11477 9313 11494
rect 9437 11477 9863 11494
rect 7237 11006 7663 11023
rect 7787 11006 8213 11023
rect 8777 11037 8794 11463
rect 8856 11037 8873 11463
rect 9327 11037 9344 11463
rect 9406 11037 9423 11463
rect 9987 11477 10413 11494
rect 10537 11477 10963 11494
rect 8337 11006 8763 11023
rect 8887 11006 9313 11023
rect 9877 11037 9894 11463
rect 9956 11037 9973 11463
rect 10427 11037 10444 11463
rect 10506 11037 10523 11463
rect 11087 11477 11513 11494
rect 11637 11477 12063 11494
rect 9437 11006 9863 11023
rect 9987 11006 10413 11023
rect 10977 11037 10994 11463
rect 11056 11037 11073 11463
rect 11527 11037 11544 11463
rect 11606 11037 11623 11463
rect 12187 11477 12613 11494
rect 12737 11477 13163 11494
rect 10537 11006 10963 11023
rect 11087 11006 11513 11023
rect 12077 11037 12094 11463
rect 12156 11037 12173 11463
rect 12627 11037 12644 11463
rect 12706 11037 12723 11463
rect 13287 11477 13713 11494
rect 11637 11006 12063 11023
rect 12187 11006 12613 11023
rect 13177 11037 13194 11463
rect 13256 11037 13273 11463
rect 12737 11006 13163 11023
rect 13287 11006 13713 11023
rect -463 10927 -37 10944
rect 87 10927 513 10944
rect -23 10487 -6 10913
rect 56 10487 73 10913
rect 637 10927 1063 10944
rect 1187 10927 1613 10944
rect -463 10456 -37 10473
rect 527 10487 544 10913
rect 606 10487 623 10913
rect 1077 10487 1094 10913
rect 1156 10487 1173 10913
rect 1737 10927 2163 10944
rect 2287 10927 2713 10944
rect 87 10456 513 10473
rect 637 10456 1063 10473
rect 1627 10487 1644 10913
rect 1706 10487 1723 10913
rect 2177 10487 2194 10913
rect 2256 10487 2273 10913
rect 2837 10927 3263 10944
rect 3387 10927 3813 10944
rect 1187 10456 1613 10473
rect 1737 10456 2163 10473
rect 2727 10487 2744 10913
rect 2806 10487 2823 10913
rect 3277 10487 3294 10913
rect 3356 10487 3373 10913
rect 3937 10927 4363 10944
rect 4487 10927 4913 10944
rect 2287 10456 2713 10473
rect 2837 10456 3263 10473
rect 3827 10487 3844 10913
rect 3906 10487 3923 10913
rect 4377 10487 4394 10913
rect 4456 10487 4473 10913
rect 5037 10927 5463 10944
rect 5587 10927 6013 10944
rect 3387 10456 3813 10473
rect 3937 10456 4363 10473
rect 4927 10487 4944 10913
rect 5006 10487 5023 10913
rect 5477 10487 5494 10913
rect 5556 10487 5573 10913
rect 6137 10927 6563 10944
rect 6687 10927 7113 10944
rect 4487 10456 4913 10473
rect 5037 10456 5463 10473
rect 6027 10487 6044 10913
rect 6106 10487 6123 10913
rect 6577 10487 6594 10913
rect 6656 10487 6673 10913
rect 7237 10927 7663 10944
rect 7787 10927 8213 10944
rect 5587 10456 6013 10473
rect 6137 10456 6563 10473
rect 7127 10487 7144 10913
rect 7206 10487 7223 10913
rect 7677 10487 7694 10913
rect 7756 10487 7773 10913
rect 8337 10927 8763 10944
rect 8887 10927 9313 10944
rect 6687 10456 7113 10473
rect 7237 10456 7663 10473
rect 8227 10487 8244 10913
rect 8306 10487 8323 10913
rect 8777 10487 8794 10913
rect 8856 10487 8873 10913
rect 9437 10927 9863 10944
rect 9987 10927 10413 10944
rect 7787 10456 8213 10473
rect 8337 10456 8763 10473
rect 9327 10487 9344 10913
rect 9406 10487 9423 10913
rect 9877 10487 9894 10913
rect 9956 10487 9973 10913
rect 10537 10927 10963 10944
rect 11087 10927 11513 10944
rect 8887 10456 9313 10473
rect 9437 10456 9863 10473
rect 10427 10487 10444 10913
rect 10506 10487 10523 10913
rect 10977 10487 10994 10913
rect 11056 10487 11073 10913
rect 11637 10927 12063 10944
rect 12187 10927 12613 10944
rect 9987 10456 10413 10473
rect 10537 10456 10963 10473
rect 11527 10487 11544 10913
rect 11606 10487 11623 10913
rect 12077 10487 12094 10913
rect 12156 10487 12173 10913
rect 12737 10927 13163 10944
rect 13287 10927 13713 10944
rect 11087 10456 11513 10473
rect 11637 10456 12063 10473
rect 12627 10487 12644 10913
rect 12706 10487 12723 10913
rect 13177 10487 13194 10913
rect 13256 10487 13273 10913
rect 12187 10456 12613 10473
rect 12737 10456 13163 10473
rect 13287 10456 13713 10473
rect -463 10377 -37 10394
rect 87 10377 513 10394
rect 637 10377 1063 10394
rect -23 9937 -6 10363
rect 56 9937 73 10363
rect 527 9937 544 10363
rect 606 9937 623 10363
rect 1187 10377 1613 10394
rect 1737 10377 2163 10394
rect -463 9906 -37 9923
rect 87 9906 513 9923
rect 1077 9937 1094 10363
rect 1156 9937 1173 10363
rect 1627 9937 1644 10363
rect 1706 9937 1723 10363
rect 2287 10377 2713 10394
rect 2837 10377 3263 10394
rect 637 9906 1063 9923
rect 1187 9906 1613 9923
rect 2177 9937 2194 10363
rect 2256 9937 2273 10363
rect 2727 9937 2744 10363
rect 2806 9937 2823 10363
rect 3387 10377 3813 10394
rect 3937 10377 4363 10394
rect 1737 9906 2163 9923
rect 2287 9906 2713 9923
rect 3277 9937 3294 10363
rect 3356 9937 3373 10363
rect 3827 9937 3844 10363
rect 3906 9937 3923 10363
rect 4487 10377 4913 10394
rect 5037 10377 5463 10394
rect 2837 9906 3263 9923
rect 3387 9906 3813 9923
rect 4377 9937 4394 10363
rect 4456 9937 4473 10363
rect 4927 9937 4944 10363
rect 5006 9937 5023 10363
rect 5587 10377 6013 10394
rect 6137 10377 6563 10394
rect 3937 9906 4363 9923
rect 4487 9906 4913 9923
rect 5477 9937 5494 10363
rect 5556 9937 5573 10363
rect 6027 9937 6044 10363
rect 6106 9937 6123 10363
rect 6687 10377 7113 10394
rect 7237 10377 7663 10394
rect 5037 9906 5463 9923
rect 5587 9906 6013 9923
rect 6577 9937 6594 10363
rect 6656 9937 6673 10363
rect 7127 9937 7144 10363
rect 7206 9937 7223 10363
rect 7787 10377 8213 10394
rect 8337 10377 8763 10394
rect 6137 9906 6563 9923
rect 6687 9906 7113 9923
rect 7677 9937 7694 10363
rect 7756 9937 7773 10363
rect 8227 9937 8244 10363
rect 8306 9937 8323 10363
rect 8887 10377 9313 10394
rect 9437 10377 9863 10394
rect 7237 9906 7663 9923
rect 7787 9906 8213 9923
rect 8777 9937 8794 10363
rect 8856 9937 8873 10363
rect 9327 9937 9344 10363
rect 9406 9937 9423 10363
rect 9987 10377 10413 10394
rect 10537 10377 10963 10394
rect 8337 9906 8763 9923
rect 8887 9906 9313 9923
rect 9877 9937 9894 10363
rect 9956 9937 9973 10363
rect 10427 9937 10444 10363
rect 10506 9937 10523 10363
rect 11087 10377 11513 10394
rect 11637 10377 12063 10394
rect 9437 9906 9863 9923
rect 9987 9906 10413 9923
rect 10977 9937 10994 10363
rect 11056 9937 11073 10363
rect 11527 9937 11544 10363
rect 11606 9937 11623 10363
rect 12187 10377 12613 10394
rect 12737 10377 13163 10394
rect 10537 9906 10963 9923
rect 11087 9906 11513 9923
rect 12077 9937 12094 10363
rect 12156 9937 12173 10363
rect 12627 9937 12644 10363
rect 12706 9937 12723 10363
rect 13287 10377 13713 10394
rect 11637 9906 12063 9923
rect 12187 9906 12613 9923
rect 13177 9937 13194 10363
rect 13256 9937 13273 10363
rect 12737 9906 13163 9923
rect 13287 9906 13713 9923
rect -463 9827 -37 9844
rect 87 9827 513 9844
rect -23 9387 -6 9813
rect 56 9387 73 9813
rect 637 9827 1063 9844
rect 1187 9827 1613 9844
rect -463 9356 -37 9373
rect 527 9387 544 9813
rect 606 9387 623 9813
rect 1077 9387 1094 9813
rect 1156 9387 1173 9813
rect 1737 9827 2163 9844
rect 2287 9827 2713 9844
rect 87 9356 513 9373
rect 637 9356 1063 9373
rect 1627 9387 1644 9813
rect 1706 9387 1723 9813
rect 2177 9387 2194 9813
rect 2256 9387 2273 9813
rect 2837 9827 3263 9844
rect 3387 9827 3813 9844
rect 1187 9356 1613 9373
rect 1737 9356 2163 9373
rect 2727 9387 2744 9813
rect 2806 9387 2823 9813
rect 3277 9387 3294 9813
rect 3356 9387 3373 9813
rect 3937 9827 4363 9844
rect 4487 9827 4913 9844
rect 2287 9356 2713 9373
rect 2837 9356 3263 9373
rect 3827 9387 3844 9813
rect 3906 9387 3923 9813
rect 4377 9387 4394 9813
rect 4456 9387 4473 9813
rect 5037 9827 5463 9844
rect 5587 9827 6013 9844
rect 3387 9356 3813 9373
rect 3937 9356 4363 9373
rect 4927 9387 4944 9813
rect 5006 9387 5023 9813
rect 5477 9387 5494 9813
rect 5556 9387 5573 9813
rect 6137 9827 6563 9844
rect 6687 9827 7113 9844
rect 4487 9356 4913 9373
rect 5037 9356 5463 9373
rect 6027 9387 6044 9813
rect 6106 9387 6123 9813
rect 6577 9387 6594 9813
rect 6656 9387 6673 9813
rect 7237 9827 7663 9844
rect 7787 9827 8213 9844
rect 5587 9356 6013 9373
rect 6137 9356 6563 9373
rect 7127 9387 7144 9813
rect 7206 9387 7223 9813
rect 7677 9387 7694 9813
rect 7756 9387 7773 9813
rect 8337 9827 8763 9844
rect 8887 9827 9313 9844
rect 6687 9356 7113 9373
rect 7237 9356 7663 9373
rect 8227 9387 8244 9813
rect 8306 9387 8323 9813
rect 8777 9387 8794 9813
rect 8856 9387 8873 9813
rect 9437 9827 9863 9844
rect 9987 9827 10413 9844
rect 7787 9356 8213 9373
rect 8337 9356 8763 9373
rect 9327 9387 9344 9813
rect 9406 9387 9423 9813
rect 9877 9387 9894 9813
rect 9956 9387 9973 9813
rect 10537 9827 10963 9844
rect 11087 9827 11513 9844
rect 8887 9356 9313 9373
rect 9437 9356 9863 9373
rect 10427 9387 10444 9813
rect 10506 9387 10523 9813
rect 10977 9387 10994 9813
rect 11056 9387 11073 9813
rect 11637 9827 12063 9844
rect 12187 9827 12613 9844
rect 9987 9356 10413 9373
rect 10537 9356 10963 9373
rect 11527 9387 11544 9813
rect 11606 9387 11623 9813
rect 12077 9387 12094 9813
rect 12156 9387 12173 9813
rect 12737 9827 13163 9844
rect 13287 9827 13713 9844
rect 11087 9356 11513 9373
rect 11637 9356 12063 9373
rect 12627 9387 12644 9813
rect 12706 9387 12723 9813
rect 13177 9387 13194 9813
rect 13256 9387 13273 9813
rect 12187 9356 12613 9373
rect 12737 9356 13163 9373
rect 13287 9356 13713 9373
rect -463 9277 -37 9294
rect 87 9277 513 9294
rect 637 9277 1063 9294
rect -23 8837 -6 9263
rect 56 8837 73 9263
rect 527 8837 544 9263
rect 606 8837 623 9263
rect 1187 9277 1613 9294
rect 1737 9277 2163 9294
rect -463 8806 -37 8823
rect 87 8806 513 8823
rect 1077 8837 1094 9263
rect 1156 8837 1173 9263
rect 1627 8837 1644 9263
rect 1706 8837 1723 9263
rect 2287 9277 2713 9294
rect 2837 9277 3263 9294
rect 637 8806 1063 8823
rect 1187 8806 1613 8823
rect 2177 8837 2194 9263
rect 2256 8837 2273 9263
rect 2727 8837 2744 9263
rect 2806 8837 2823 9263
rect 3387 9277 3813 9294
rect 3937 9277 4363 9294
rect 1737 8806 2163 8823
rect 2287 8806 2713 8823
rect 3277 8837 3294 9263
rect 3356 8837 3373 9263
rect 3827 8837 3844 9263
rect 3906 8837 3923 9263
rect 4487 9277 4913 9294
rect 5037 9277 5463 9294
rect 2837 8806 3263 8823
rect 3387 8806 3813 8823
rect 4377 8837 4394 9263
rect 4456 8837 4473 9263
rect 4927 8837 4944 9263
rect 5006 8837 5023 9263
rect 5587 9277 6013 9294
rect 6137 9277 6563 9294
rect 3937 8806 4363 8823
rect 4487 8806 4913 8823
rect 5477 8837 5494 9263
rect 5556 8837 5573 9263
rect 6027 8837 6044 9263
rect 6106 8837 6123 9263
rect 6687 9277 7113 9294
rect 7237 9277 7663 9294
rect 5037 8806 5463 8823
rect 5587 8806 6013 8823
rect 6577 8837 6594 9263
rect 6656 8837 6673 9263
rect 7127 8837 7144 9263
rect 7206 8837 7223 9263
rect 7787 9277 8213 9294
rect 8337 9277 8763 9294
rect 6137 8806 6563 8823
rect 6687 8806 7113 8823
rect 7677 8837 7694 9263
rect 7756 8837 7773 9263
rect 8227 8837 8244 9263
rect 8306 8837 8323 9263
rect 8887 9277 9313 9294
rect 9437 9277 9863 9294
rect 7237 8806 7663 8823
rect 7787 8806 8213 8823
rect 8777 8837 8794 9263
rect 8856 8837 8873 9263
rect 9327 8837 9344 9263
rect 9406 8837 9423 9263
rect 9987 9277 10413 9294
rect 10537 9277 10963 9294
rect 8337 8806 8763 8823
rect 8887 8806 9313 8823
rect 9877 8837 9894 9263
rect 9956 8837 9973 9263
rect 10427 8837 10444 9263
rect 10506 8837 10523 9263
rect 11087 9277 11513 9294
rect 11637 9277 12063 9294
rect 9437 8806 9863 8823
rect 9987 8806 10413 8823
rect 10977 8837 10994 9263
rect 11056 8837 11073 9263
rect 11527 8837 11544 9263
rect 11606 8837 11623 9263
rect 12187 9277 12613 9294
rect 12737 9277 13163 9294
rect 10537 8806 10963 8823
rect 11087 8806 11513 8823
rect 12077 8837 12094 9263
rect 12156 8837 12173 9263
rect 12627 8837 12644 9263
rect 12706 8837 12723 9263
rect 13287 9277 13713 9294
rect 11637 8806 12063 8823
rect 12187 8806 12613 8823
rect 13177 8837 13194 9263
rect 13256 8837 13273 9263
rect 12737 8806 13163 8823
rect 13287 8806 13713 8823
rect -463 8727 -37 8744
rect 87 8727 513 8744
rect -23 8287 -6 8713
rect 56 8287 73 8713
rect 637 8727 1063 8744
rect 1187 8727 1613 8744
rect -463 8256 -37 8273
rect 527 8287 544 8713
rect 606 8287 623 8713
rect 1077 8287 1094 8713
rect 1156 8287 1173 8713
rect 1737 8727 2163 8744
rect 2287 8727 2713 8744
rect 87 8256 513 8273
rect 637 8256 1063 8273
rect 1627 8287 1644 8713
rect 1706 8287 1723 8713
rect 2177 8287 2194 8713
rect 2256 8287 2273 8713
rect 2837 8727 3263 8744
rect 3387 8727 3813 8744
rect 1187 8256 1613 8273
rect 1737 8256 2163 8273
rect 2727 8287 2744 8713
rect 2806 8287 2823 8713
rect 3277 8287 3294 8713
rect 3356 8287 3373 8713
rect 3937 8727 4363 8744
rect 4487 8727 4913 8744
rect 2287 8256 2713 8273
rect 2837 8256 3263 8273
rect 3827 8287 3844 8713
rect 3906 8287 3923 8713
rect 4377 8287 4394 8713
rect 4456 8287 4473 8713
rect 5037 8727 5463 8744
rect 5587 8727 6013 8744
rect 3387 8256 3813 8273
rect 3937 8256 4363 8273
rect 4927 8287 4944 8713
rect 5006 8287 5023 8713
rect 5477 8287 5494 8713
rect 5556 8287 5573 8713
rect 6137 8727 6563 8744
rect 6687 8727 7113 8744
rect 4487 8256 4913 8273
rect 5037 8256 5463 8273
rect 6027 8287 6044 8713
rect 6106 8287 6123 8713
rect 6577 8287 6594 8713
rect 6656 8287 6673 8713
rect 7237 8727 7663 8744
rect 7787 8727 8213 8744
rect 5587 8256 6013 8273
rect 6137 8256 6563 8273
rect 7127 8287 7144 8713
rect 7206 8287 7223 8713
rect 7677 8287 7694 8713
rect 7756 8287 7773 8713
rect 8337 8727 8763 8744
rect 8887 8727 9313 8744
rect 6687 8256 7113 8273
rect 7237 8256 7663 8273
rect 8227 8287 8244 8713
rect 8306 8287 8323 8713
rect 8777 8287 8794 8713
rect 8856 8287 8873 8713
rect 9437 8727 9863 8744
rect 9987 8727 10413 8744
rect 7787 8256 8213 8273
rect 8337 8256 8763 8273
rect 9327 8287 9344 8713
rect 9406 8287 9423 8713
rect 9877 8287 9894 8713
rect 9956 8287 9973 8713
rect 10537 8727 10963 8744
rect 11087 8727 11513 8744
rect 8887 8256 9313 8273
rect 9437 8256 9863 8273
rect 10427 8287 10444 8713
rect 10506 8287 10523 8713
rect 10977 8287 10994 8713
rect 11056 8287 11073 8713
rect 11637 8727 12063 8744
rect 12187 8727 12613 8744
rect 9987 8256 10413 8273
rect 10537 8256 10963 8273
rect 11527 8287 11544 8713
rect 11606 8287 11623 8713
rect 12077 8287 12094 8713
rect 12156 8287 12173 8713
rect 12737 8727 13163 8744
rect 13287 8727 13713 8744
rect 11087 8256 11513 8273
rect 11637 8256 12063 8273
rect 12627 8287 12644 8713
rect 12706 8287 12723 8713
rect 13177 8287 13194 8713
rect 13256 8287 13273 8713
rect 12187 8256 12613 8273
rect 12737 8256 13163 8273
rect 13287 8256 13713 8273
rect -463 8177 -37 8194
rect 87 8177 513 8194
rect 637 8177 1063 8194
rect -23 7737 -6 8163
rect 56 7737 73 8163
rect 527 7737 544 8163
rect 606 7737 623 8163
rect 1187 8177 1613 8194
rect 1737 8177 2163 8194
rect -463 7706 -37 7723
rect 87 7706 513 7723
rect 1077 7737 1094 8163
rect 1156 7737 1173 8163
rect 1627 7737 1644 8163
rect 1706 7737 1723 8163
rect 2287 8177 2713 8194
rect 2837 8177 3263 8194
rect 637 7706 1063 7723
rect 1187 7706 1613 7723
rect 2177 7737 2194 8163
rect 2256 7737 2273 8163
rect 2727 7737 2744 8163
rect 2806 7737 2823 8163
rect 3387 8177 3813 8194
rect 3937 8177 4363 8194
rect 1737 7706 2163 7723
rect 2287 7706 2713 7723
rect 3277 7737 3294 8163
rect 3356 7737 3373 8163
rect 3827 7737 3844 8163
rect 3906 7737 3923 8163
rect 4487 8177 4913 8194
rect 5037 8177 5463 8194
rect 2837 7706 3263 7723
rect 3387 7706 3813 7723
rect 4377 7737 4394 8163
rect 4456 7737 4473 8163
rect 4927 7737 4944 8163
rect 5006 7737 5023 8163
rect 5587 8177 6013 8194
rect 6137 8177 6563 8194
rect 3937 7706 4363 7723
rect 4487 7706 4913 7723
rect 5477 7737 5494 8163
rect 5556 7737 5573 8163
rect 6027 7737 6044 8163
rect 6106 7737 6123 8163
rect 6687 8177 7113 8194
rect 7237 8177 7663 8194
rect 5037 7706 5463 7723
rect 5587 7706 6013 7723
rect 6577 7737 6594 8163
rect 6656 7737 6673 8163
rect 7127 7737 7144 8163
rect 7206 7737 7223 8163
rect 7787 8177 8213 8194
rect 8337 8177 8763 8194
rect 6137 7706 6563 7723
rect 6687 7706 7113 7723
rect 7677 7737 7694 8163
rect 7756 7737 7773 8163
rect 8227 7737 8244 8163
rect 8306 7737 8323 8163
rect 8887 8177 9313 8194
rect 9437 8177 9863 8194
rect 7237 7706 7663 7723
rect 7787 7706 8213 7723
rect 8777 7737 8794 8163
rect 8856 7737 8873 8163
rect 9327 7737 9344 8163
rect 9406 7737 9423 8163
rect 9987 8177 10413 8194
rect 10537 8177 10963 8194
rect 8337 7706 8763 7723
rect 8887 7706 9313 7723
rect 9877 7737 9894 8163
rect 9956 7737 9973 8163
rect 10427 7737 10444 8163
rect 10506 7737 10523 8163
rect 11087 8177 11513 8194
rect 11637 8177 12063 8194
rect 9437 7706 9863 7723
rect 9987 7706 10413 7723
rect 10977 7737 10994 8163
rect 11056 7737 11073 8163
rect 11527 7737 11544 8163
rect 11606 7737 11623 8163
rect 12187 8177 12613 8194
rect 12737 8177 13163 8194
rect 10537 7706 10963 7723
rect 11087 7706 11513 7723
rect 12077 7737 12094 8163
rect 12156 7737 12173 8163
rect 12627 7737 12644 8163
rect 12706 7737 12723 8163
rect 13287 8177 13713 8194
rect 11637 7706 12063 7723
rect 12187 7706 12613 7723
rect 13177 7737 13194 8163
rect 13256 7737 13273 8163
rect 12737 7706 13163 7723
rect 13287 7706 13713 7723
rect -463 7627 -37 7644
rect 87 7627 513 7644
rect -23 7187 -6 7613
rect 56 7187 73 7613
rect 637 7627 1063 7644
rect 1187 7627 1613 7644
rect -463 7156 -37 7173
rect 527 7187 544 7613
rect 606 7187 623 7613
rect 1077 7187 1094 7613
rect 1156 7187 1173 7613
rect 1737 7627 2163 7644
rect 2287 7627 2713 7644
rect 87 7156 513 7173
rect 637 7156 1063 7173
rect 1627 7187 1644 7613
rect 1706 7187 1723 7613
rect 2177 7187 2194 7613
rect 2256 7187 2273 7613
rect 2837 7627 3263 7644
rect 3387 7627 3813 7644
rect 1187 7156 1613 7173
rect 1737 7156 2163 7173
rect 2727 7187 2744 7613
rect 2806 7187 2823 7613
rect 3277 7187 3294 7613
rect 3356 7187 3373 7613
rect 3937 7627 4363 7644
rect 4487 7627 4913 7644
rect 2287 7156 2713 7173
rect 2837 7156 3263 7173
rect 3827 7187 3844 7613
rect 3906 7187 3923 7613
rect 4377 7187 4394 7613
rect 4456 7187 4473 7613
rect 5037 7627 5463 7644
rect 5587 7627 6013 7644
rect 3387 7156 3813 7173
rect 3937 7156 4363 7173
rect 4927 7187 4944 7613
rect 5006 7187 5023 7613
rect 5477 7187 5494 7613
rect 5556 7187 5573 7613
rect 6137 7627 6563 7644
rect 6687 7627 7113 7644
rect 4487 7156 4913 7173
rect 5037 7156 5463 7173
rect 6027 7187 6044 7613
rect 6106 7187 6123 7613
rect 6577 7187 6594 7613
rect 6656 7187 6673 7613
rect 7237 7627 7663 7644
rect 7787 7627 8213 7644
rect 5587 7156 6013 7173
rect 6137 7156 6563 7173
rect 7127 7187 7144 7613
rect 7206 7187 7223 7613
rect 7677 7187 7694 7613
rect 7756 7187 7773 7613
rect 8337 7627 8763 7644
rect 8887 7627 9313 7644
rect 6687 7156 7113 7173
rect 7237 7156 7663 7173
rect 8227 7187 8244 7613
rect 8306 7187 8323 7613
rect 8777 7187 8794 7613
rect 8856 7187 8873 7613
rect 9437 7627 9863 7644
rect 9987 7627 10413 7644
rect 7787 7156 8213 7173
rect 8337 7156 8763 7173
rect 9327 7187 9344 7613
rect 9406 7187 9423 7613
rect 9877 7187 9894 7613
rect 9956 7187 9973 7613
rect 10537 7627 10963 7644
rect 11087 7627 11513 7644
rect 8887 7156 9313 7173
rect 9437 7156 9863 7173
rect 10427 7187 10444 7613
rect 10506 7187 10523 7613
rect 10977 7187 10994 7613
rect 11056 7187 11073 7613
rect 11637 7627 12063 7644
rect 12187 7627 12613 7644
rect 9987 7156 10413 7173
rect 10537 7156 10963 7173
rect 11527 7187 11544 7613
rect 11606 7187 11623 7613
rect 12077 7187 12094 7613
rect 12156 7187 12173 7613
rect 12737 7627 13163 7644
rect 13287 7627 13713 7644
rect 11087 7156 11513 7173
rect 11637 7156 12063 7173
rect 12627 7187 12644 7613
rect 12706 7187 12723 7613
rect 13177 7187 13194 7613
rect 13256 7187 13273 7613
rect 12187 7156 12613 7173
rect 12737 7156 13163 7173
rect 13287 7156 13713 7173
rect -463 7077 -37 7094
rect 87 7077 513 7094
rect 637 7077 1063 7094
rect -23 6637 -6 7063
rect 56 6637 73 7063
rect 527 6637 544 7063
rect 606 6637 623 7063
rect 1187 7077 1613 7094
rect 1737 7077 2163 7094
rect -463 6606 -37 6623
rect 87 6606 513 6623
rect 1077 6637 1094 7063
rect 1156 6637 1173 7063
rect 1627 6637 1644 7063
rect 1706 6637 1723 7063
rect 2287 7077 2713 7094
rect 2837 7077 3263 7094
rect 637 6606 1063 6623
rect 1187 6606 1613 6623
rect 2177 6637 2194 7063
rect 2256 6637 2273 7063
rect 2727 6637 2744 7063
rect 2806 6637 2823 7063
rect 3387 7077 3813 7094
rect 3937 7077 4363 7094
rect 1737 6606 2163 6623
rect 2287 6606 2713 6623
rect 3277 6637 3294 7063
rect 3356 6637 3373 7063
rect 3827 6637 3844 7063
rect 3906 6637 3923 7063
rect 4487 7077 4913 7094
rect 5037 7077 5463 7094
rect 2837 6606 3263 6623
rect 3387 6606 3813 6623
rect 4377 6637 4394 7063
rect 4456 6637 4473 7063
rect 4927 6637 4944 7063
rect 5006 6637 5023 7063
rect 5587 7077 6013 7094
rect 6137 7077 6563 7094
rect 3937 6606 4363 6623
rect 4487 6606 4913 6623
rect 5477 6637 5494 7063
rect 5556 6637 5573 7063
rect 6027 6637 6044 7063
rect 6106 6637 6123 7063
rect 6687 7077 7113 7094
rect 7237 7077 7663 7094
rect 5037 6606 5463 6623
rect 5587 6606 6013 6623
rect 6577 6637 6594 7063
rect 6656 6637 6673 7063
rect 7127 6637 7144 7063
rect 7206 6637 7223 7063
rect 7787 7077 8213 7094
rect 8337 7077 8763 7094
rect 6137 6606 6563 6623
rect 6687 6606 7113 6623
rect 7677 6637 7694 7063
rect 7756 6637 7773 7063
rect 8227 6637 8244 7063
rect 8306 6637 8323 7063
rect 8887 7077 9313 7094
rect 9437 7077 9863 7094
rect 7237 6606 7663 6623
rect 7787 6606 8213 6623
rect 8777 6637 8794 7063
rect 8856 6637 8873 7063
rect 9327 6637 9344 7063
rect 9406 6637 9423 7063
rect 9987 7077 10413 7094
rect 10537 7077 10963 7094
rect 8337 6606 8763 6623
rect 8887 6606 9313 6623
rect 9877 6637 9894 7063
rect 9956 6637 9973 7063
rect 10427 6637 10444 7063
rect 10506 6637 10523 7063
rect 11087 7077 11513 7094
rect 11637 7077 12063 7094
rect 9437 6606 9863 6623
rect 9987 6606 10413 6623
rect 10977 6637 10994 7063
rect 11056 6637 11073 7063
rect 11527 6637 11544 7063
rect 11606 6637 11623 7063
rect 12187 7077 12613 7094
rect 12737 7077 13163 7094
rect 10537 6606 10963 6623
rect 11087 6606 11513 6623
rect 12077 6637 12094 7063
rect 12156 6637 12173 7063
rect 12627 6637 12644 7063
rect 12706 6637 12723 7063
rect 13287 7077 13713 7094
rect 11637 6606 12063 6623
rect 12187 6606 12613 6623
rect 13177 6637 13194 7063
rect 13256 6637 13273 7063
rect 12737 6606 13163 6623
rect 13287 6606 13713 6623
rect -463 6527 -37 6544
rect 87 6527 513 6544
rect -23 6087 -6 6513
rect 56 6087 73 6513
rect 637 6527 1063 6544
rect 1187 6527 1613 6544
rect -463 6056 -37 6073
rect 527 6087 544 6513
rect 606 6087 623 6513
rect 1077 6087 1094 6513
rect 1156 6087 1173 6513
rect 1737 6527 2163 6544
rect 2287 6527 2713 6544
rect 87 6056 513 6073
rect 637 6056 1063 6073
rect 1627 6087 1644 6513
rect 1706 6087 1723 6513
rect 2177 6087 2194 6513
rect 2256 6087 2273 6513
rect 2837 6527 3263 6544
rect 3387 6527 3813 6544
rect 1187 6056 1613 6073
rect 1737 6056 2163 6073
rect 2727 6087 2744 6513
rect 2806 6087 2823 6513
rect 3277 6087 3294 6513
rect 3356 6087 3373 6513
rect 3937 6527 4363 6544
rect 4487 6527 4913 6544
rect 2287 6056 2713 6073
rect 2837 6056 3263 6073
rect 3827 6087 3844 6513
rect 3906 6087 3923 6513
rect 4377 6087 4394 6513
rect 4456 6087 4473 6513
rect 5037 6527 5463 6544
rect 5587 6527 6013 6544
rect 3387 6056 3813 6073
rect 3937 6056 4363 6073
rect 4927 6087 4944 6513
rect 5006 6087 5023 6513
rect 5477 6087 5494 6513
rect 5556 6087 5573 6513
rect 6137 6527 6563 6544
rect 6687 6527 7113 6544
rect 4487 6056 4913 6073
rect 5037 6056 5463 6073
rect 6027 6087 6044 6513
rect 6106 6087 6123 6513
rect 6577 6087 6594 6513
rect 6656 6087 6673 6513
rect 7237 6527 7663 6544
rect 7787 6527 8213 6544
rect 5587 6056 6013 6073
rect 6137 6056 6563 6073
rect 7127 6087 7144 6513
rect 7206 6087 7223 6513
rect 7677 6087 7694 6513
rect 7756 6087 7773 6513
rect 8337 6527 8763 6544
rect 8887 6527 9313 6544
rect 6687 6056 7113 6073
rect 7237 6056 7663 6073
rect 8227 6087 8244 6513
rect 8306 6087 8323 6513
rect 8777 6087 8794 6513
rect 8856 6087 8873 6513
rect 9437 6527 9863 6544
rect 9987 6527 10413 6544
rect 7787 6056 8213 6073
rect 8337 6056 8763 6073
rect 9327 6087 9344 6513
rect 9406 6087 9423 6513
rect 9877 6087 9894 6513
rect 9956 6087 9973 6513
rect 10537 6527 10963 6544
rect 11087 6527 11513 6544
rect 8887 6056 9313 6073
rect 9437 6056 9863 6073
rect 10427 6087 10444 6513
rect 10506 6087 10523 6513
rect 10977 6087 10994 6513
rect 11056 6087 11073 6513
rect 11637 6527 12063 6544
rect 12187 6527 12613 6544
rect 9987 6056 10413 6073
rect 10537 6056 10963 6073
rect 11527 6087 11544 6513
rect 11606 6087 11623 6513
rect 12077 6087 12094 6513
rect 12156 6087 12173 6513
rect 12737 6527 13163 6544
rect 13287 6527 13713 6544
rect 11087 6056 11513 6073
rect 11637 6056 12063 6073
rect 12627 6087 12644 6513
rect 12706 6087 12723 6513
rect 13177 6087 13194 6513
rect 13256 6087 13273 6513
rect 12187 6056 12613 6073
rect 12737 6056 13163 6073
rect 13287 6056 13713 6073
rect -463 5977 -37 5994
rect 87 5977 513 5994
rect 637 5977 1063 5994
rect -23 5537 -6 5963
rect 56 5537 73 5963
rect 527 5537 544 5963
rect 606 5537 623 5963
rect 1187 5977 1613 5994
rect 1737 5977 2163 5994
rect -463 5506 -37 5523
rect 87 5506 513 5523
rect 1077 5537 1094 5963
rect 1156 5537 1173 5963
rect 1627 5537 1644 5963
rect 1706 5537 1723 5963
rect 2287 5977 2713 5994
rect 2837 5977 3263 5994
rect 637 5506 1063 5523
rect 1187 5506 1613 5523
rect 2177 5537 2194 5963
rect 2256 5537 2273 5963
rect 2727 5537 2744 5963
rect 2806 5537 2823 5963
rect 3387 5977 3813 5994
rect 3937 5977 4363 5994
rect 1737 5506 2163 5523
rect 2287 5506 2713 5523
rect 3277 5537 3294 5963
rect 3356 5537 3373 5963
rect 3827 5537 3844 5963
rect 3906 5537 3923 5963
rect 4487 5977 4913 5994
rect 5037 5977 5463 5994
rect 2837 5506 3263 5523
rect 3387 5506 3813 5523
rect 4377 5537 4394 5963
rect 4456 5537 4473 5963
rect 4927 5537 4944 5963
rect 5006 5537 5023 5963
rect 5587 5977 6013 5994
rect 6137 5977 6563 5994
rect 3937 5506 4363 5523
rect 4487 5506 4913 5523
rect 5477 5537 5494 5963
rect 5556 5537 5573 5963
rect 6027 5537 6044 5963
rect 6106 5537 6123 5963
rect 6687 5977 7113 5994
rect 7237 5977 7663 5994
rect 5037 5506 5463 5523
rect 5587 5506 6013 5523
rect 6577 5537 6594 5963
rect 6656 5537 6673 5963
rect 7127 5537 7144 5963
rect 7206 5537 7223 5963
rect 7787 5977 8213 5994
rect 8337 5977 8763 5994
rect 6137 5506 6563 5523
rect 6687 5506 7113 5523
rect 7677 5537 7694 5963
rect 7756 5537 7773 5963
rect 8227 5537 8244 5963
rect 8306 5537 8323 5963
rect 8887 5977 9313 5994
rect 9437 5977 9863 5994
rect 7237 5506 7663 5523
rect 7787 5506 8213 5523
rect 8777 5537 8794 5963
rect 8856 5537 8873 5963
rect 9327 5537 9344 5963
rect 9406 5537 9423 5963
rect 9987 5977 10413 5994
rect 10537 5977 10963 5994
rect 8337 5506 8763 5523
rect 8887 5506 9313 5523
rect 9877 5537 9894 5963
rect 9956 5537 9973 5963
rect 10427 5537 10444 5963
rect 10506 5537 10523 5963
rect 11087 5977 11513 5994
rect 11637 5977 12063 5994
rect 9437 5506 9863 5523
rect 9987 5506 10413 5523
rect 10977 5537 10994 5963
rect 11056 5537 11073 5963
rect 11527 5537 11544 5963
rect 11606 5537 11623 5963
rect 12187 5977 12613 5994
rect 12737 5977 13163 5994
rect 10537 5506 10963 5523
rect 11087 5506 11513 5523
rect 12077 5537 12094 5963
rect 12156 5537 12173 5963
rect 12627 5537 12644 5963
rect 12706 5537 12723 5963
rect 13287 5977 13713 5994
rect 11637 5506 12063 5523
rect 12187 5506 12613 5523
rect 13177 5537 13194 5963
rect 13256 5537 13273 5963
rect 12737 5506 13163 5523
rect 13287 5506 13713 5523
rect -463 5427 -37 5444
rect 87 5427 513 5444
rect -23 4987 -6 5413
rect 56 4987 73 5413
rect 637 5427 1063 5444
rect 1187 5427 1613 5444
rect -463 4956 -37 4973
rect 527 4987 544 5413
rect 606 4987 623 5413
rect 1077 4987 1094 5413
rect 1156 4987 1173 5413
rect 1737 5427 2163 5444
rect 2287 5427 2713 5444
rect 87 4956 513 4973
rect 637 4956 1063 4973
rect 1627 4987 1644 5413
rect 1706 4987 1723 5413
rect 2177 4987 2194 5413
rect 2256 4987 2273 5413
rect 2837 5427 3263 5444
rect 3387 5427 3813 5444
rect 1187 4956 1613 4973
rect 1737 4956 2163 4973
rect 2727 4987 2744 5413
rect 2806 4987 2823 5413
rect 3277 4987 3294 5413
rect 3356 4987 3373 5413
rect 3937 5427 4363 5444
rect 4487 5427 4913 5444
rect 2287 4956 2713 4973
rect 2837 4956 3263 4973
rect 3827 4987 3844 5413
rect 3906 4987 3923 5413
rect 4377 4987 4394 5413
rect 4456 4987 4473 5413
rect 5037 5427 5463 5444
rect 5587 5427 6013 5444
rect 3387 4956 3813 4973
rect 3937 4956 4363 4973
rect 4927 4987 4944 5413
rect 5006 4987 5023 5413
rect 5477 4987 5494 5413
rect 5556 4987 5573 5413
rect 6137 5427 6563 5444
rect 6687 5427 7113 5444
rect 4487 4956 4913 4973
rect 5037 4956 5463 4973
rect 6027 4987 6044 5413
rect 6106 4987 6123 5413
rect 6577 4987 6594 5413
rect 6656 4987 6673 5413
rect 7237 5427 7663 5444
rect 7787 5427 8213 5444
rect 5587 4956 6013 4973
rect 6137 4956 6563 4973
rect 7127 4987 7144 5413
rect 7206 4987 7223 5413
rect 7677 4987 7694 5413
rect 7756 4987 7773 5413
rect 8337 5427 8763 5444
rect 8887 5427 9313 5444
rect 6687 4956 7113 4973
rect 7237 4956 7663 4973
rect 8227 4987 8244 5413
rect 8306 4987 8323 5413
rect 8777 4987 8794 5413
rect 8856 4987 8873 5413
rect 9437 5427 9863 5444
rect 9987 5427 10413 5444
rect 7787 4956 8213 4973
rect 8337 4956 8763 4973
rect 9327 4987 9344 5413
rect 9406 4987 9423 5413
rect 9877 4987 9894 5413
rect 9956 4987 9973 5413
rect 10537 5427 10963 5444
rect 11087 5427 11513 5444
rect 8887 4956 9313 4973
rect 9437 4956 9863 4973
rect 10427 4987 10444 5413
rect 10506 4987 10523 5413
rect 10977 4987 10994 5413
rect 11056 4987 11073 5413
rect 11637 5427 12063 5444
rect 12187 5427 12613 5444
rect 9987 4956 10413 4973
rect 10537 4956 10963 4973
rect 11527 4987 11544 5413
rect 11606 4987 11623 5413
rect 12077 4987 12094 5413
rect 12156 4987 12173 5413
rect 12737 5427 13163 5444
rect 13287 5427 13713 5444
rect 11087 4956 11513 4973
rect 11637 4956 12063 4973
rect 12627 4987 12644 5413
rect 12706 4987 12723 5413
rect 13177 4987 13194 5413
rect 13256 4987 13273 5413
rect 12187 4956 12613 4973
rect 12737 4956 13163 4973
rect 13287 4956 13713 4973
rect -463 4877 -37 4894
rect 87 4877 513 4894
rect 637 4877 1063 4894
rect -23 4437 -6 4863
rect 56 4437 73 4863
rect 527 4437 544 4863
rect 606 4437 623 4863
rect 1187 4877 1613 4894
rect 1737 4877 2163 4894
rect -463 4406 -37 4423
rect 87 4406 513 4423
rect 1077 4437 1094 4863
rect 1156 4437 1173 4863
rect 1627 4437 1644 4863
rect 1706 4437 1723 4863
rect 2287 4877 2713 4894
rect 2837 4877 3263 4894
rect 637 4406 1063 4423
rect 1187 4406 1613 4423
rect 2177 4437 2194 4863
rect 2256 4437 2273 4863
rect 2727 4437 2744 4863
rect 2806 4437 2823 4863
rect 3387 4877 3813 4894
rect 3937 4877 4363 4894
rect 1737 4406 2163 4423
rect 2287 4406 2713 4423
rect 3277 4437 3294 4863
rect 3356 4437 3373 4863
rect 3827 4437 3844 4863
rect 3906 4437 3923 4863
rect 4487 4877 4913 4894
rect 5037 4877 5463 4894
rect 2837 4406 3263 4423
rect 3387 4406 3813 4423
rect 4377 4437 4394 4863
rect 4456 4437 4473 4863
rect 4927 4437 4944 4863
rect 5006 4437 5023 4863
rect 5587 4877 6013 4894
rect 6137 4877 6563 4894
rect 3937 4406 4363 4423
rect 4487 4406 4913 4423
rect 5477 4437 5494 4863
rect 5556 4437 5573 4863
rect 6027 4437 6044 4863
rect 6106 4437 6123 4863
rect 6687 4877 7113 4894
rect 7237 4877 7663 4894
rect 5037 4406 5463 4423
rect 5587 4406 6013 4423
rect 6577 4437 6594 4863
rect 6656 4437 6673 4863
rect 7127 4437 7144 4863
rect 7206 4437 7223 4863
rect 7787 4877 8213 4894
rect 8337 4877 8763 4894
rect 6137 4406 6563 4423
rect 6687 4406 7113 4423
rect 7677 4437 7694 4863
rect 7756 4437 7773 4863
rect 8227 4437 8244 4863
rect 8306 4437 8323 4863
rect 8887 4877 9313 4894
rect 9437 4877 9863 4894
rect 7237 4406 7663 4423
rect 7787 4406 8213 4423
rect 8777 4437 8794 4863
rect 8856 4437 8873 4863
rect 9327 4437 9344 4863
rect 9406 4437 9423 4863
rect 9987 4877 10413 4894
rect 10537 4877 10963 4894
rect 8337 4406 8763 4423
rect 8887 4406 9313 4423
rect 9877 4437 9894 4863
rect 9956 4437 9973 4863
rect 10427 4437 10444 4863
rect 10506 4437 10523 4863
rect 11087 4877 11513 4894
rect 11637 4877 12063 4894
rect 9437 4406 9863 4423
rect 9987 4406 10413 4423
rect 10977 4437 10994 4863
rect 11056 4437 11073 4863
rect 11527 4437 11544 4863
rect 11606 4437 11623 4863
rect 12187 4877 12613 4894
rect 12737 4877 13163 4894
rect 10537 4406 10963 4423
rect 11087 4406 11513 4423
rect 12077 4437 12094 4863
rect 12156 4437 12173 4863
rect 12627 4437 12644 4863
rect 12706 4437 12723 4863
rect 13287 4877 13713 4894
rect 11637 4406 12063 4423
rect 12187 4406 12613 4423
rect 13177 4437 13194 4863
rect 13256 4437 13273 4863
rect 12737 4406 13163 4423
rect 13287 4406 13713 4423
rect -463 4327 -37 4344
rect 87 4327 513 4344
rect -23 3887 -6 4313
rect 56 3887 73 4313
rect 637 4327 1063 4344
rect 1187 4327 1613 4344
rect -463 3856 -37 3873
rect 527 3887 544 4313
rect 606 3887 623 4313
rect 1077 3887 1094 4313
rect 1156 3887 1173 4313
rect 1737 4327 2163 4344
rect 2287 4327 2713 4344
rect 87 3856 513 3873
rect 637 3856 1063 3873
rect 1627 3887 1644 4313
rect 1706 3887 1723 4313
rect 2177 3887 2194 4313
rect 2256 3887 2273 4313
rect 2837 4327 3263 4344
rect 3387 4327 3813 4344
rect 1187 3856 1613 3873
rect 1737 3856 2163 3873
rect 2727 3887 2744 4313
rect 2806 3887 2823 4313
rect 3277 3887 3294 4313
rect 3356 3887 3373 4313
rect 3937 4327 4363 4344
rect 4487 4327 4913 4344
rect 2287 3856 2713 3873
rect 2837 3856 3263 3873
rect 3827 3887 3844 4313
rect 3906 3887 3923 4313
rect 4377 3887 4394 4313
rect 4456 3887 4473 4313
rect 5037 4327 5463 4344
rect 5587 4327 6013 4344
rect 3387 3856 3813 3873
rect 3937 3856 4363 3873
rect 4927 3887 4944 4313
rect 5006 3887 5023 4313
rect 5477 3887 5494 4313
rect 5556 3887 5573 4313
rect 6137 4327 6563 4344
rect 6687 4327 7113 4344
rect 4487 3856 4913 3873
rect 5037 3856 5463 3873
rect 6027 3887 6044 4313
rect 6106 3887 6123 4313
rect 6577 3887 6594 4313
rect 6656 3887 6673 4313
rect 7237 4327 7663 4344
rect 7787 4327 8213 4344
rect 5587 3856 6013 3873
rect 6137 3856 6563 3873
rect 7127 3887 7144 4313
rect 7206 3887 7223 4313
rect 7677 3887 7694 4313
rect 7756 3887 7773 4313
rect 8337 4327 8763 4344
rect 8887 4327 9313 4344
rect 6687 3856 7113 3873
rect 7237 3856 7663 3873
rect 8227 3887 8244 4313
rect 8306 3887 8323 4313
rect 8777 3887 8794 4313
rect 8856 3887 8873 4313
rect 9437 4327 9863 4344
rect 9987 4327 10413 4344
rect 7787 3856 8213 3873
rect 8337 3856 8763 3873
rect 9327 3887 9344 4313
rect 9406 3887 9423 4313
rect 9877 3887 9894 4313
rect 9956 3887 9973 4313
rect 10537 4327 10963 4344
rect 11087 4327 11513 4344
rect 8887 3856 9313 3873
rect 9437 3856 9863 3873
rect 10427 3887 10444 4313
rect 10506 3887 10523 4313
rect 10977 3887 10994 4313
rect 11056 3887 11073 4313
rect 11637 4327 12063 4344
rect 12187 4327 12613 4344
rect 9987 3856 10413 3873
rect 10537 3856 10963 3873
rect 11527 3887 11544 4313
rect 11606 3887 11623 4313
rect 12077 3887 12094 4313
rect 12156 3887 12173 4313
rect 12737 4327 13163 4344
rect 13287 4327 13713 4344
rect 11087 3856 11513 3873
rect 11637 3856 12063 3873
rect 12627 3887 12644 4313
rect 12706 3887 12723 4313
rect 13177 3887 13194 4313
rect 13256 3887 13273 4313
rect 12187 3856 12613 3873
rect 12737 3856 13163 3873
rect 13287 3856 13713 3873
rect -463 3777 -37 3794
rect 87 3777 513 3794
rect 637 3777 1063 3794
rect -23 3337 -6 3763
rect 56 3337 73 3763
rect 527 3337 544 3763
rect 606 3337 623 3763
rect 1187 3777 1613 3794
rect 1737 3777 2163 3794
rect -463 3306 -37 3323
rect 87 3306 513 3323
rect 1077 3337 1094 3763
rect 1156 3337 1173 3763
rect 1627 3337 1644 3763
rect 1706 3337 1723 3763
rect 2287 3777 2713 3794
rect 2837 3777 3263 3794
rect 637 3306 1063 3323
rect 1187 3306 1613 3323
rect 2177 3337 2194 3763
rect 2256 3337 2273 3763
rect 2727 3337 2744 3763
rect 2806 3337 2823 3763
rect 3387 3777 3813 3794
rect 3937 3777 4363 3794
rect 1737 3306 2163 3323
rect 2287 3306 2713 3323
rect 3277 3337 3294 3763
rect 3356 3337 3373 3763
rect 3827 3337 3844 3763
rect 3906 3337 3923 3763
rect 4487 3777 4913 3794
rect 5037 3777 5463 3794
rect 2837 3306 3263 3323
rect 3387 3306 3813 3323
rect 4377 3337 4394 3763
rect 4456 3337 4473 3763
rect 4927 3337 4944 3763
rect 5006 3337 5023 3763
rect 5587 3777 6013 3794
rect 6137 3777 6563 3794
rect 3937 3306 4363 3323
rect 4487 3306 4913 3323
rect 5477 3337 5494 3763
rect 5556 3337 5573 3763
rect 6027 3337 6044 3763
rect 6106 3337 6123 3763
rect 6687 3777 7113 3794
rect 7237 3777 7663 3794
rect 5037 3306 5463 3323
rect 5587 3306 6013 3323
rect 6577 3337 6594 3763
rect 6656 3337 6673 3763
rect 7127 3337 7144 3763
rect 7206 3337 7223 3763
rect 7787 3777 8213 3794
rect 8337 3777 8763 3794
rect 6137 3306 6563 3323
rect 6687 3306 7113 3323
rect 7677 3337 7694 3763
rect 7756 3337 7773 3763
rect 8227 3337 8244 3763
rect 8306 3337 8323 3763
rect 8887 3777 9313 3794
rect 9437 3777 9863 3794
rect 7237 3306 7663 3323
rect 7787 3306 8213 3323
rect 8777 3337 8794 3763
rect 8856 3337 8873 3763
rect 9327 3337 9344 3763
rect 9406 3337 9423 3763
rect 9987 3777 10413 3794
rect 10537 3777 10963 3794
rect 8337 3306 8763 3323
rect 8887 3306 9313 3323
rect 9877 3337 9894 3763
rect 9956 3337 9973 3763
rect 10427 3337 10444 3763
rect 10506 3337 10523 3763
rect 11087 3777 11513 3794
rect 11637 3777 12063 3794
rect 9437 3306 9863 3323
rect 9987 3306 10413 3323
rect 10977 3337 10994 3763
rect 11056 3337 11073 3763
rect 11527 3337 11544 3763
rect 11606 3337 11623 3763
rect 12187 3777 12613 3794
rect 12737 3777 13163 3794
rect 10537 3306 10963 3323
rect 11087 3306 11513 3323
rect 12077 3337 12094 3763
rect 12156 3337 12173 3763
rect 12627 3337 12644 3763
rect 12706 3337 12723 3763
rect 13287 3777 13713 3794
rect 11637 3306 12063 3323
rect 12187 3306 12613 3323
rect 13177 3337 13194 3763
rect 13256 3337 13273 3763
rect 12737 3306 13163 3323
rect 13287 3306 13713 3323
rect -463 3227 -37 3244
rect 87 3227 513 3244
rect -23 2787 -6 3213
rect 56 2787 73 3213
rect 637 3227 1063 3244
rect 1187 3227 1613 3244
rect -463 2756 -37 2773
rect 527 2787 544 3213
rect 606 2787 623 3213
rect 1077 2787 1094 3213
rect 1156 2787 1173 3213
rect 1737 3227 2163 3244
rect 2287 3227 2713 3244
rect 87 2756 513 2773
rect 637 2756 1063 2773
rect 1627 2787 1644 3213
rect 1706 2787 1723 3213
rect 2177 2787 2194 3213
rect 2256 2787 2273 3213
rect 2837 3227 3263 3244
rect 3387 3227 3813 3244
rect 1187 2756 1613 2773
rect 1737 2756 2163 2773
rect 2727 2787 2744 3213
rect 2806 2787 2823 3213
rect 3277 2787 3294 3213
rect 3356 2787 3373 3213
rect 3937 3227 4363 3244
rect 4487 3227 4913 3244
rect 2287 2756 2713 2773
rect 2837 2756 3263 2773
rect 3827 2787 3844 3213
rect 3906 2787 3923 3213
rect 4377 2787 4394 3213
rect 4456 2787 4473 3213
rect 5037 3227 5463 3244
rect 5587 3227 6013 3244
rect 3387 2756 3813 2773
rect 3937 2756 4363 2773
rect 4927 2787 4944 3213
rect 5006 2787 5023 3213
rect 5477 2787 5494 3213
rect 5556 2787 5573 3213
rect 6137 3227 6563 3244
rect 6687 3227 7113 3244
rect 4487 2756 4913 2773
rect 5037 2756 5463 2773
rect 6027 2787 6044 3213
rect 6106 2787 6123 3213
rect 6577 2787 6594 3213
rect 6656 2787 6673 3213
rect 7237 3227 7663 3244
rect 7787 3227 8213 3244
rect 5587 2756 6013 2773
rect 6137 2756 6563 2773
rect 7127 2787 7144 3213
rect 7206 2787 7223 3213
rect 7677 2787 7694 3213
rect 7756 2787 7773 3213
rect 8337 3227 8763 3244
rect 8887 3227 9313 3244
rect 6687 2756 7113 2773
rect 7237 2756 7663 2773
rect 8227 2787 8244 3213
rect 8306 2787 8323 3213
rect 8777 2787 8794 3213
rect 8856 2787 8873 3213
rect 9437 3227 9863 3244
rect 9987 3227 10413 3244
rect 7787 2756 8213 2773
rect 8337 2756 8763 2773
rect 9327 2787 9344 3213
rect 9406 2787 9423 3213
rect 9877 2787 9894 3213
rect 9956 2787 9973 3213
rect 10537 3227 10963 3244
rect 11087 3227 11513 3244
rect 8887 2756 9313 2773
rect 9437 2756 9863 2773
rect 10427 2787 10444 3213
rect 10506 2787 10523 3213
rect 10977 2787 10994 3213
rect 11056 2787 11073 3213
rect 11637 3227 12063 3244
rect 12187 3227 12613 3244
rect 9987 2756 10413 2773
rect 10537 2756 10963 2773
rect 11527 2787 11544 3213
rect 11606 2787 11623 3213
rect 12077 2787 12094 3213
rect 12156 2787 12173 3213
rect 12737 3227 13163 3244
rect 13287 3227 13713 3244
rect 11087 2756 11513 2773
rect 11637 2756 12063 2773
rect 12627 2787 12644 3213
rect 12706 2787 12723 3213
rect 13177 2787 13194 3213
rect 13256 2787 13273 3213
rect 12187 2756 12613 2773
rect 12737 2756 13163 2773
rect 13287 2756 13713 2773
rect -463 2677 -37 2694
rect 87 2677 513 2694
rect 637 2677 1063 2694
rect -23 2237 -6 2663
rect 56 2237 73 2663
rect 527 2237 544 2663
rect 606 2237 623 2663
rect 1187 2677 1613 2694
rect 1737 2677 2163 2694
rect -463 2206 -37 2223
rect 87 2206 513 2223
rect 1077 2237 1094 2663
rect 1156 2237 1173 2663
rect 1627 2237 1644 2663
rect 1706 2237 1723 2663
rect 2287 2677 2713 2694
rect 2837 2677 3263 2694
rect 637 2206 1063 2223
rect 1187 2206 1613 2223
rect 2177 2237 2194 2663
rect 2256 2237 2273 2663
rect 2727 2237 2744 2663
rect 2806 2237 2823 2663
rect 3387 2677 3813 2694
rect 3937 2677 4363 2694
rect 1737 2206 2163 2223
rect 2287 2206 2713 2223
rect 3277 2237 3294 2663
rect 3356 2237 3373 2663
rect 3827 2237 3844 2663
rect 3906 2237 3923 2663
rect 4487 2677 4913 2694
rect 5037 2677 5463 2694
rect 2837 2206 3263 2223
rect 3387 2206 3813 2223
rect 4377 2237 4394 2663
rect 4456 2237 4473 2663
rect 4927 2237 4944 2663
rect 5006 2237 5023 2663
rect 5587 2677 6013 2694
rect 6137 2677 6563 2694
rect 3937 2206 4363 2223
rect 4487 2206 4913 2223
rect 5477 2237 5494 2663
rect 5556 2237 5573 2663
rect 6027 2237 6044 2663
rect 6106 2237 6123 2663
rect 6687 2677 7113 2694
rect 7237 2677 7663 2694
rect 5037 2206 5463 2223
rect 5587 2206 6013 2223
rect 6577 2237 6594 2663
rect 6656 2237 6673 2663
rect 7127 2237 7144 2663
rect 7206 2237 7223 2663
rect 7787 2677 8213 2694
rect 8337 2677 8763 2694
rect 6137 2206 6563 2223
rect 6687 2206 7113 2223
rect 7677 2237 7694 2663
rect 7756 2237 7773 2663
rect 8227 2237 8244 2663
rect 8306 2237 8323 2663
rect 8887 2677 9313 2694
rect 9437 2677 9863 2694
rect 7237 2206 7663 2223
rect 7787 2206 8213 2223
rect 8777 2237 8794 2663
rect 8856 2237 8873 2663
rect 9327 2237 9344 2663
rect 9406 2237 9423 2663
rect 9987 2677 10413 2694
rect 10537 2677 10963 2694
rect 8337 2206 8763 2223
rect 8887 2206 9313 2223
rect 9877 2237 9894 2663
rect 9956 2237 9973 2663
rect 10427 2237 10444 2663
rect 10506 2237 10523 2663
rect 11087 2677 11513 2694
rect 11637 2677 12063 2694
rect 9437 2206 9863 2223
rect 9987 2206 10413 2223
rect 10977 2237 10994 2663
rect 11056 2237 11073 2663
rect 11527 2237 11544 2663
rect 11606 2237 11623 2663
rect 12187 2677 12613 2694
rect 12737 2677 13163 2694
rect 10537 2206 10963 2223
rect 11087 2206 11513 2223
rect 12077 2237 12094 2663
rect 12156 2237 12173 2663
rect 12627 2237 12644 2663
rect 12706 2237 12723 2663
rect 13287 2677 13713 2694
rect 11637 2206 12063 2223
rect 12187 2206 12613 2223
rect 13177 2237 13194 2663
rect 13256 2237 13273 2663
rect 12737 2206 13163 2223
rect 13287 2206 13713 2223
rect -463 2127 -37 2144
rect 87 2127 513 2144
rect -23 1687 -6 2113
rect 56 1687 73 2113
rect 637 2127 1063 2144
rect 1187 2127 1613 2144
rect -463 1656 -37 1673
rect 527 1687 544 2113
rect 606 1687 623 2113
rect 1077 1687 1094 2113
rect 1156 1687 1173 2113
rect 1737 2127 2163 2144
rect 2287 2127 2713 2144
rect 87 1656 513 1673
rect 637 1656 1063 1673
rect 1627 1687 1644 2113
rect 1706 1687 1723 2113
rect 2177 1687 2194 2113
rect 2256 1687 2273 2113
rect 2837 2127 3263 2144
rect 3387 2127 3813 2144
rect 1187 1656 1613 1673
rect 1737 1656 2163 1673
rect 2727 1687 2744 2113
rect 2806 1687 2823 2113
rect 3277 1687 3294 2113
rect 3356 1687 3373 2113
rect 3937 2127 4363 2144
rect 4487 2127 4913 2144
rect 2287 1656 2713 1673
rect 2837 1656 3263 1673
rect 3827 1687 3844 2113
rect 3906 1687 3923 2113
rect 4377 1687 4394 2113
rect 4456 1687 4473 2113
rect 5037 2127 5463 2144
rect 5587 2127 6013 2144
rect 3387 1656 3813 1673
rect 3937 1656 4363 1673
rect 4927 1687 4944 2113
rect 5006 1687 5023 2113
rect 5477 1687 5494 2113
rect 5556 1687 5573 2113
rect 6137 2127 6563 2144
rect 6687 2127 7113 2144
rect 4487 1656 4913 1673
rect 5037 1656 5463 1673
rect 6027 1687 6044 2113
rect 6106 1687 6123 2113
rect 6577 1687 6594 2113
rect 6656 1687 6673 2113
rect 7237 2127 7663 2144
rect 7787 2127 8213 2144
rect 5587 1656 6013 1673
rect 6137 1656 6563 1673
rect 7127 1687 7144 2113
rect 7206 1687 7223 2113
rect 7677 1687 7694 2113
rect 7756 1687 7773 2113
rect 8337 2127 8763 2144
rect 8887 2127 9313 2144
rect 6687 1656 7113 1673
rect 7237 1656 7663 1673
rect 8227 1687 8244 2113
rect 8306 1687 8323 2113
rect 8777 1687 8794 2113
rect 8856 1687 8873 2113
rect 9437 2127 9863 2144
rect 9987 2127 10413 2144
rect 7787 1656 8213 1673
rect 8337 1656 8763 1673
rect 9327 1687 9344 2113
rect 9406 1687 9423 2113
rect 9877 1687 9894 2113
rect 9956 1687 9973 2113
rect 10537 2127 10963 2144
rect 11087 2127 11513 2144
rect 8887 1656 9313 1673
rect 9437 1656 9863 1673
rect 10427 1687 10444 2113
rect 10506 1687 10523 2113
rect 10977 1687 10994 2113
rect 11056 1687 11073 2113
rect 11637 2127 12063 2144
rect 12187 2127 12613 2144
rect 9987 1656 10413 1673
rect 10537 1656 10963 1673
rect 11527 1687 11544 2113
rect 11606 1687 11623 2113
rect 12077 1687 12094 2113
rect 12156 1687 12173 2113
rect 12737 2127 13163 2144
rect 13287 2127 13713 2144
rect 11087 1656 11513 1673
rect 11637 1656 12063 1673
rect 12627 1687 12644 2113
rect 12706 1687 12723 2113
rect 13177 1687 13194 2113
rect 13256 1687 13273 2113
rect 12187 1656 12613 1673
rect 12737 1656 13163 1673
rect 13287 1656 13713 1673
rect -463 1577 -37 1594
rect 87 1577 513 1594
rect 637 1577 1063 1594
rect -23 1137 -6 1563
rect 56 1137 73 1563
rect 527 1137 544 1563
rect 606 1137 623 1563
rect 1187 1577 1613 1594
rect 1737 1577 2163 1594
rect -463 1106 -37 1123
rect 87 1106 513 1123
rect 1077 1137 1094 1563
rect 1156 1137 1173 1563
rect 1627 1137 1644 1563
rect 1706 1137 1723 1563
rect 2287 1577 2713 1594
rect 2837 1577 3263 1594
rect 637 1106 1063 1123
rect 1187 1106 1613 1123
rect 2177 1137 2194 1563
rect 2256 1137 2273 1563
rect 2727 1137 2744 1563
rect 2806 1137 2823 1563
rect 3387 1577 3813 1594
rect 3937 1577 4363 1594
rect 1737 1106 2163 1123
rect 2287 1106 2713 1123
rect 3277 1137 3294 1563
rect 3356 1137 3373 1563
rect 3827 1137 3844 1563
rect 3906 1137 3923 1563
rect 4487 1577 4913 1594
rect 5037 1577 5463 1594
rect 2837 1106 3263 1123
rect 3387 1106 3813 1123
rect 4377 1137 4394 1563
rect 4456 1137 4473 1563
rect 4927 1137 4944 1563
rect 5006 1137 5023 1563
rect 5587 1577 6013 1594
rect 6137 1577 6563 1594
rect 3937 1106 4363 1123
rect 4487 1106 4913 1123
rect 5477 1137 5494 1563
rect 5556 1137 5573 1563
rect 6027 1137 6044 1563
rect 6106 1137 6123 1563
rect 6687 1577 7113 1594
rect 7237 1577 7663 1594
rect 5037 1106 5463 1123
rect 5587 1106 6013 1123
rect 6577 1137 6594 1563
rect 6656 1137 6673 1563
rect 7127 1137 7144 1563
rect 7206 1137 7223 1563
rect 7787 1577 8213 1594
rect 8337 1577 8763 1594
rect 6137 1106 6563 1123
rect 6687 1106 7113 1123
rect 7677 1137 7694 1563
rect 7756 1137 7773 1563
rect 8227 1137 8244 1563
rect 8306 1137 8323 1563
rect 8887 1577 9313 1594
rect 9437 1577 9863 1594
rect 7237 1106 7663 1123
rect 7787 1106 8213 1123
rect 8777 1137 8794 1563
rect 8856 1137 8873 1563
rect 9327 1137 9344 1563
rect 9406 1137 9423 1563
rect 9987 1577 10413 1594
rect 10537 1577 10963 1594
rect 8337 1106 8763 1123
rect 8887 1106 9313 1123
rect 9877 1137 9894 1563
rect 9956 1137 9973 1563
rect 10427 1137 10444 1563
rect 10506 1137 10523 1563
rect 11087 1577 11513 1594
rect 11637 1577 12063 1594
rect 9437 1106 9863 1123
rect 9987 1106 10413 1123
rect 10977 1137 10994 1563
rect 11056 1137 11073 1563
rect 11527 1137 11544 1563
rect 11606 1137 11623 1563
rect 12187 1577 12613 1594
rect 12737 1577 13163 1594
rect 10537 1106 10963 1123
rect 11087 1106 11513 1123
rect 12077 1137 12094 1563
rect 12156 1137 12173 1563
rect 12627 1137 12644 1563
rect 12706 1137 12723 1563
rect 13287 1577 13713 1594
rect 11637 1106 12063 1123
rect 12187 1106 12613 1123
rect 13177 1137 13194 1563
rect 13256 1137 13273 1563
rect 12737 1106 13163 1123
rect 13287 1106 13713 1123
rect -463 1027 -37 1044
rect 87 1027 513 1044
rect -23 587 -6 1013
rect 56 587 73 1013
rect 637 1027 1063 1044
rect 1187 1027 1613 1044
rect -463 556 -37 573
rect 527 587 544 1013
rect 606 587 623 1013
rect 1077 587 1094 1013
rect 1156 587 1173 1013
rect 1737 1027 2163 1044
rect 2287 1027 2713 1044
rect 87 556 513 573
rect 637 556 1063 573
rect 1627 587 1644 1013
rect 1706 587 1723 1013
rect 2177 587 2194 1013
rect 2256 587 2273 1013
rect 2837 1027 3263 1044
rect 3387 1027 3813 1044
rect 1187 556 1613 573
rect 1737 556 2163 573
rect 2727 587 2744 1013
rect 2806 587 2823 1013
rect 3277 587 3294 1013
rect 3356 587 3373 1013
rect 3937 1027 4363 1044
rect 4487 1027 4913 1044
rect 2287 556 2713 573
rect 2837 556 3263 573
rect 3827 587 3844 1013
rect 3906 587 3923 1013
rect 4377 587 4394 1013
rect 4456 587 4473 1013
rect 5037 1027 5463 1044
rect 5587 1027 6013 1044
rect 3387 556 3813 573
rect 3937 556 4363 573
rect 4927 587 4944 1013
rect 5006 587 5023 1013
rect 5477 587 5494 1013
rect 5556 587 5573 1013
rect 6137 1027 6563 1044
rect 6687 1027 7113 1044
rect 4487 556 4913 573
rect 5037 556 5463 573
rect 6027 587 6044 1013
rect 6106 587 6123 1013
rect 6577 587 6594 1013
rect 6656 587 6673 1013
rect 7237 1027 7663 1044
rect 7787 1027 8213 1044
rect 5587 556 6013 573
rect 6137 556 6563 573
rect 7127 587 7144 1013
rect 7206 587 7223 1013
rect 7677 587 7694 1013
rect 7756 587 7773 1013
rect 8337 1027 8763 1044
rect 8887 1027 9313 1044
rect 6687 556 7113 573
rect 7237 556 7663 573
rect 8227 587 8244 1013
rect 8306 587 8323 1013
rect 8777 587 8794 1013
rect 8856 587 8873 1013
rect 9437 1027 9863 1044
rect 9987 1027 10413 1044
rect 7787 556 8213 573
rect 8337 556 8763 573
rect 9327 587 9344 1013
rect 9406 587 9423 1013
rect 9877 587 9894 1013
rect 9956 587 9973 1013
rect 10537 1027 10963 1044
rect 11087 1027 11513 1044
rect 8887 556 9313 573
rect 9437 556 9863 573
rect 10427 587 10444 1013
rect 10506 587 10523 1013
rect 10977 587 10994 1013
rect 11056 587 11073 1013
rect 11637 1027 12063 1044
rect 12187 1027 12613 1044
rect 9987 556 10413 573
rect 10537 556 10963 573
rect 11527 587 11544 1013
rect 11606 587 11623 1013
rect 12077 587 12094 1013
rect 12156 587 12173 1013
rect 12737 1027 13163 1044
rect 13287 1027 13713 1044
rect 11087 556 11513 573
rect 11637 556 12063 573
rect 12627 587 12644 1013
rect 12706 587 12723 1013
rect 13177 587 13194 1013
rect 13256 587 13273 1013
rect 12187 556 12613 573
rect 12737 556 13163 573
rect 13287 556 13713 573
rect -463 477 -37 494
rect 87 477 513 494
rect 637 477 1063 494
rect -23 37 -6 463
rect 56 37 73 463
rect 527 37 544 463
rect 606 37 623 463
rect 1187 477 1613 494
rect 1737 477 2163 494
rect -463 6 -37 23
rect 87 6 513 23
rect 1077 37 1094 463
rect 1156 37 1173 463
rect 1627 37 1644 463
rect 1706 37 1723 463
rect 2287 477 2713 494
rect 2837 477 3263 494
rect 637 6 1063 23
rect 1187 6 1613 23
rect 2177 37 2194 463
rect 2256 37 2273 463
rect 2727 37 2744 463
rect 2806 37 2823 463
rect 3387 477 3813 494
rect 3937 477 4363 494
rect 1737 6 2163 23
rect 2287 6 2713 23
rect 3277 37 3294 463
rect 3356 37 3373 463
rect 3827 37 3844 463
rect 3906 37 3923 463
rect 4487 477 4913 494
rect 5037 477 5463 494
rect 2837 6 3263 23
rect 3387 6 3813 23
rect 4377 37 4394 463
rect 4456 37 4473 463
rect 4927 37 4944 463
rect 5006 37 5023 463
rect 5587 477 6013 494
rect 6137 477 6563 494
rect 3937 6 4363 23
rect 4487 6 4913 23
rect 5477 37 5494 463
rect 5556 37 5573 463
rect 6027 37 6044 463
rect 6106 37 6123 463
rect 6687 477 7113 494
rect 7237 477 7663 494
rect 5037 6 5463 23
rect 5587 6 6013 23
rect 6577 37 6594 463
rect 6656 37 6673 463
rect 7127 37 7144 463
rect 7206 37 7223 463
rect 7787 477 8213 494
rect 8337 477 8763 494
rect 6137 6 6563 23
rect 6687 6 7113 23
rect 7677 37 7694 463
rect 7756 37 7773 463
rect 8227 37 8244 463
rect 8306 37 8323 463
rect 8887 477 9313 494
rect 9437 477 9863 494
rect 7237 6 7663 23
rect 7787 6 8213 23
rect 8777 37 8794 463
rect 8856 37 8873 463
rect 9327 37 9344 463
rect 9406 37 9423 463
rect 9987 477 10413 494
rect 10537 477 10963 494
rect 8337 6 8763 23
rect 8887 6 9313 23
rect 9877 37 9894 463
rect 9956 37 9973 463
rect 10427 37 10444 463
rect 10506 37 10523 463
rect 11087 477 11513 494
rect 11637 477 12063 494
rect 9437 6 9863 23
rect 9987 6 10413 23
rect 10977 37 10994 463
rect 11056 37 11073 463
rect 11527 37 11544 463
rect 11606 37 11623 463
rect 12187 477 12613 494
rect 12737 477 13163 494
rect 10537 6 10963 23
rect 11087 6 11513 23
rect 12077 37 12094 463
rect 12156 37 12173 463
rect 12627 37 12644 463
rect 12706 37 12723 463
rect 13287 477 13713 494
rect 11637 6 12063 23
rect 12187 6 12613 23
rect 13177 37 13194 463
rect 13256 37 13273 463
rect 12737 6 13163 23
rect 13287 6 13713 23
rect -463 -73 -37 -56
rect 87 -73 513 -56
rect -23 -513 -6 -87
rect 56 -513 73 -87
rect 637 -73 1063 -56
rect 1187 -73 1613 -56
rect 527 -513 544 -87
rect 606 -513 623 -87
rect 1077 -513 1094 -87
rect 1156 -513 1173 -87
rect 1737 -73 2163 -56
rect 2287 -73 2713 -56
rect 1627 -513 1644 -87
rect 1706 -513 1723 -87
rect 2177 -513 2194 -87
rect 2256 -513 2273 -87
rect 2837 -73 3263 -56
rect 3387 -73 3813 -56
rect 2727 -513 2744 -87
rect 2806 -513 2823 -87
rect 3277 -513 3294 -87
rect 3356 -513 3373 -87
rect 3937 -73 4363 -56
rect 4487 -73 4913 -56
rect 3827 -513 3844 -87
rect 3906 -513 3923 -87
rect 4377 -513 4394 -87
rect 4456 -513 4473 -87
rect 5037 -73 5463 -56
rect 5587 -73 6013 -56
rect 4927 -513 4944 -87
rect 5006 -513 5023 -87
rect 5477 -513 5494 -87
rect 5556 -513 5573 -87
rect 6137 -73 6563 -56
rect 6687 -73 7113 -56
rect 6027 -513 6044 -87
rect 6106 -513 6123 -87
rect 6577 -513 6594 -87
rect 6656 -513 6673 -87
rect 7237 -73 7663 -56
rect 7787 -73 8213 -56
rect 7127 -513 7144 -87
rect 7206 -513 7223 -87
rect 7677 -513 7694 -87
rect 7756 -513 7773 -87
rect 8337 -73 8763 -56
rect 8887 -73 9313 -56
rect 8227 -513 8244 -87
rect 8306 -513 8323 -87
rect 8777 -513 8794 -87
rect 8856 -513 8873 -87
rect 9437 -73 9863 -56
rect 9987 -73 10413 -56
rect 9327 -513 9344 -87
rect 9406 -513 9423 -87
rect 9877 -513 9894 -87
rect 9956 -513 9973 -87
rect 10537 -73 10963 -56
rect 11087 -73 11513 -56
rect 10427 -513 10444 -87
rect 10506 -513 10523 -87
rect 10977 -513 10994 -87
rect 11056 -513 11073 -87
rect 11637 -73 12063 -56
rect 12187 -73 12613 -56
rect 11527 -513 11544 -87
rect 11606 -513 11623 -87
rect 12077 -513 12094 -87
rect 12156 -513 12173 -87
rect 12737 -73 13163 -56
rect 13287 -73 13713 -56
rect 12627 -513 12644 -87
rect 12706 -513 12723 -87
rect 13177 -513 13194 -87
rect 13256 -513 13273 -87
<< mvpsubdiff >>
rect -5525 18713 18775 18725
rect -5525 -5563 -5513 18713
rect -1537 14725 14787 14737
rect -1537 -1575 -1525 14725
rect 14775 -1575 14787 14725
rect -1537 -1587 14787 -1575
rect 18763 -5563 18775 18713
rect -5525 -5575 18775 -5563
<< mvnsubdiff >>
rect -1025 14213 14275 14225
rect -1025 13217 -1013 14213
rect -17 13937 0 14213
rect 533 13937 550 14213
rect 1083 13937 1100 14213
rect 1633 13937 1650 14213
rect 2183 13937 2200 14213
rect 2733 13937 2750 14213
rect 3283 13937 3300 14213
rect 3833 13937 3850 14213
rect 4383 13937 4400 14213
rect 4933 13937 4950 14213
rect 5483 13937 5500 14213
rect 6033 13937 6050 14213
rect 6583 13937 6600 14213
rect 7133 13937 7150 14213
rect 7683 13937 7700 14213
rect 8233 13937 8250 14213
rect 8783 13937 8800 14213
rect 9333 13937 9350 14213
rect 9883 13937 9900 14213
rect 10433 13937 10450 14213
rect 10983 13937 11000 14213
rect 11533 13937 11550 14213
rect 12083 13937 12100 14213
rect 12633 13937 12650 14213
rect 13183 13937 13200 14213
rect -737 13925 13987 13937
rect -737 13217 -725 13925
rect -1025 13200 -725 13217
rect -1025 12667 -1013 13200
rect -737 12667 -725 13200
rect -1025 12650 -725 12667
rect -1025 12117 -1013 12650
rect -737 12117 -725 12650
rect -1025 12100 -725 12117
rect -1025 11567 -1013 12100
rect -737 11567 -725 12100
rect -1025 11550 -725 11567
rect -1025 11017 -1013 11550
rect -737 11017 -725 11550
rect -1025 11000 -725 11017
rect -1025 10467 -1013 11000
rect -737 10467 -725 11000
rect -1025 10450 -725 10467
rect -1025 9917 -1013 10450
rect -737 9917 -725 10450
rect -1025 9900 -725 9917
rect -1025 9367 -1013 9900
rect -737 9367 -725 9900
rect -1025 9350 -725 9367
rect -1025 8817 -1013 9350
rect -737 8817 -725 9350
rect -1025 8800 -725 8817
rect -1025 8267 -1013 8800
rect -737 8267 -725 8800
rect -1025 8250 -725 8267
rect -1025 7717 -1013 8250
rect -737 7717 -725 8250
rect -1025 7700 -725 7717
rect -1025 7167 -1013 7700
rect -737 7167 -725 7700
rect -1025 7150 -725 7167
rect -1025 6617 -1013 7150
rect -737 6617 -725 7150
rect -1025 6600 -725 6617
rect -1025 6067 -1013 6600
rect -737 6067 -725 6600
rect -1025 6050 -725 6067
rect -1025 5517 -1013 6050
rect -737 5517 -725 6050
rect -1025 5500 -725 5517
rect -1025 4967 -1013 5500
rect -737 4967 -725 5500
rect -1025 4950 -725 4967
rect -1025 4417 -1013 4950
rect -737 4417 -725 4950
rect -1025 4400 -725 4417
rect -1025 3867 -1013 4400
rect -737 3867 -725 4400
rect -1025 3850 -725 3867
rect -1025 3317 -1013 3850
rect -737 3317 -725 3850
rect -1025 3300 -725 3317
rect -1025 2767 -1013 3300
rect -737 2767 -725 3300
rect -1025 2750 -725 2767
rect -1025 2217 -1013 2750
rect -737 2217 -725 2750
rect -1025 2200 -725 2217
rect -1025 1667 -1013 2200
rect -737 1667 -725 2200
rect -1025 1650 -725 1667
rect -1025 1117 -1013 1650
rect -737 1117 -725 1650
rect -1025 1100 -725 1117
rect -1025 567 -1013 1100
rect -737 567 -725 1100
rect -1025 550 -725 567
rect -1025 17 -1013 550
rect -737 17 -725 550
rect -1025 0 -725 17
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect 135 13603 465 13615
rect 135 13297 147 13603
rect 453 13297 465 13603
rect 135 13285 465 13297
rect 1235 13603 1565 13615
rect 1235 13297 1247 13603
rect 1553 13297 1565 13603
rect 1235 13285 1565 13297
rect 2335 13603 2665 13615
rect 2335 13297 2347 13603
rect 2653 13297 2665 13603
rect 2335 13285 2665 13297
rect 3435 13603 3765 13615
rect 3435 13297 3447 13603
rect 3753 13297 3765 13603
rect 3435 13285 3765 13297
rect 4535 13603 4865 13615
rect 4535 13297 4547 13603
rect 4853 13297 4865 13603
rect 4535 13285 4865 13297
rect 5635 13603 5965 13615
rect 5635 13297 5647 13603
rect 5953 13297 5965 13603
rect 5635 13285 5965 13297
rect 6735 13603 7065 13615
rect 6735 13297 6747 13603
rect 7053 13297 7065 13603
rect 6735 13285 7065 13297
rect 7835 13603 8165 13615
rect 7835 13297 7847 13603
rect 8153 13297 8165 13603
rect 7835 13285 8165 13297
rect 8935 13603 9265 13615
rect 8935 13297 8947 13603
rect 9253 13297 9265 13603
rect 8935 13285 9265 13297
rect 10035 13603 10365 13615
rect 10035 13297 10047 13603
rect 10353 13297 10365 13603
rect 10035 13285 10365 13297
rect 11135 13603 11465 13615
rect 11135 13297 11147 13603
rect 11453 13297 11465 13603
rect 11135 13285 11465 13297
rect 12235 13603 12565 13615
rect 12235 13297 12247 13603
rect 12553 13297 12565 13603
rect 12235 13285 12565 13297
rect 13335 13603 13665 13615
rect 13335 13297 13347 13603
rect 13653 13297 13665 13603
rect 13335 13285 13665 13297
rect -415 13053 -85 13065
rect -415 12747 -403 13053
rect -97 12747 -85 13053
rect -415 12735 -85 12747
rect 685 13053 1015 13065
rect 685 12747 697 13053
rect 1003 12747 1015 13053
rect 685 12735 1015 12747
rect 1785 13053 2115 13065
rect 1785 12747 1797 13053
rect 2103 12747 2115 13053
rect 1785 12735 2115 12747
rect 2885 13053 3215 13065
rect 2885 12747 2897 13053
rect 3203 12747 3215 13053
rect 2885 12735 3215 12747
rect 3985 13053 4315 13065
rect 3985 12747 3997 13053
rect 4303 12747 4315 13053
rect 3985 12735 4315 12747
rect 5085 13053 5415 13065
rect 5085 12747 5097 13053
rect 5403 12747 5415 13053
rect 5085 12735 5415 12747
rect 6185 13053 6515 13065
rect 6185 12747 6197 13053
rect 6503 12747 6515 13053
rect 6185 12735 6515 12747
rect 7285 13053 7615 13065
rect 7285 12747 7297 13053
rect 7603 12747 7615 13053
rect 7285 12735 7615 12747
rect 8385 13053 8715 13065
rect 8385 12747 8397 13053
rect 8703 12747 8715 13053
rect 8385 12735 8715 12747
rect 9485 13053 9815 13065
rect 9485 12747 9497 13053
rect 9803 12747 9815 13053
rect 9485 12735 9815 12747
rect 10585 13053 10915 13065
rect 10585 12747 10597 13053
rect 10903 12747 10915 13053
rect 10585 12735 10915 12747
rect 11685 13053 12015 13065
rect 11685 12747 11697 13053
rect 12003 12747 12015 13053
rect 11685 12735 12015 12747
rect 12785 13053 13115 13065
rect 12785 12747 12797 13053
rect 13103 12747 13115 13053
rect 12785 12735 13115 12747
rect 135 12503 465 12515
rect 135 12197 147 12503
rect 453 12197 465 12503
rect 135 12185 465 12197
rect 1235 12503 1565 12515
rect 1235 12197 1247 12503
rect 1553 12197 1565 12503
rect 1235 12185 1565 12197
rect 2335 12503 2665 12515
rect 2335 12197 2347 12503
rect 2653 12197 2665 12503
rect 2335 12185 2665 12197
rect 3435 12503 3765 12515
rect 3435 12197 3447 12503
rect 3753 12197 3765 12503
rect 3435 12185 3765 12197
rect 4535 12503 4865 12515
rect 4535 12197 4547 12503
rect 4853 12197 4865 12503
rect 4535 12185 4865 12197
rect 5635 12503 5965 12515
rect 5635 12197 5647 12503
rect 5953 12197 5965 12503
rect 5635 12185 5965 12197
rect 6735 12503 7065 12515
rect 6735 12197 6747 12503
rect 7053 12197 7065 12503
rect 6735 12185 7065 12197
rect 7835 12503 8165 12515
rect 7835 12197 7847 12503
rect 8153 12197 8165 12503
rect 7835 12185 8165 12197
rect 8935 12503 9265 12515
rect 8935 12197 8947 12503
rect 9253 12197 9265 12503
rect 8935 12185 9265 12197
rect 10035 12503 10365 12515
rect 10035 12197 10047 12503
rect 10353 12197 10365 12503
rect 10035 12185 10365 12197
rect 11135 12503 11465 12515
rect 11135 12197 11147 12503
rect 11453 12197 11465 12503
rect 11135 12185 11465 12197
rect 12235 12503 12565 12515
rect 12235 12197 12247 12503
rect 12553 12197 12565 12503
rect 12235 12185 12565 12197
rect 13335 12503 13665 12515
rect 13335 12197 13347 12503
rect 13653 12197 13665 12503
rect 13335 12185 13665 12197
rect -415 11953 -85 11965
rect -415 11647 -403 11953
rect -97 11647 -85 11953
rect -415 11635 -85 11647
rect 685 11953 1015 11965
rect 685 11647 697 11953
rect 1003 11647 1015 11953
rect 685 11635 1015 11647
rect 1785 11953 2115 11965
rect 1785 11647 1797 11953
rect 2103 11647 2115 11953
rect 1785 11635 2115 11647
rect 2885 11953 3215 11965
rect 2885 11647 2897 11953
rect 3203 11647 3215 11953
rect 2885 11635 3215 11647
rect 3985 11953 4315 11965
rect 3985 11647 3997 11953
rect 4303 11647 4315 11953
rect 3985 11635 4315 11647
rect 5085 11953 5415 11965
rect 5085 11647 5097 11953
rect 5403 11647 5415 11953
rect 5085 11635 5415 11647
rect 6185 11953 6515 11965
rect 6185 11647 6197 11953
rect 6503 11647 6515 11953
rect 6185 11635 6515 11647
rect 7285 11953 7615 11965
rect 7285 11647 7297 11953
rect 7603 11647 7615 11953
rect 7285 11635 7615 11647
rect 8385 11953 8715 11965
rect 8385 11647 8397 11953
rect 8703 11647 8715 11953
rect 8385 11635 8715 11647
rect 9485 11953 9815 11965
rect 9485 11647 9497 11953
rect 9803 11647 9815 11953
rect 9485 11635 9815 11647
rect 10585 11953 10915 11965
rect 10585 11647 10597 11953
rect 10903 11647 10915 11953
rect 10585 11635 10915 11647
rect 11685 11953 12015 11965
rect 11685 11647 11697 11953
rect 12003 11647 12015 11953
rect 11685 11635 12015 11647
rect 12785 11953 13115 11965
rect 12785 11647 12797 11953
rect 13103 11647 13115 11953
rect 12785 11635 13115 11647
rect 135 11403 465 11415
rect 135 11097 147 11403
rect 453 11097 465 11403
rect 135 11085 465 11097
rect 1235 11403 1565 11415
rect 1235 11097 1247 11403
rect 1553 11097 1565 11403
rect 1235 11085 1565 11097
rect 2335 11403 2665 11415
rect 2335 11097 2347 11403
rect 2653 11097 2665 11403
rect 2335 11085 2665 11097
rect 3435 11403 3765 11415
rect 3435 11097 3447 11403
rect 3753 11097 3765 11403
rect 3435 11085 3765 11097
rect 4535 11403 4865 11415
rect 4535 11097 4547 11403
rect 4853 11097 4865 11403
rect 4535 11085 4865 11097
rect 5635 11403 5965 11415
rect 5635 11097 5647 11403
rect 5953 11097 5965 11403
rect 5635 11085 5965 11097
rect 6735 11403 7065 11415
rect 6735 11097 6747 11403
rect 7053 11097 7065 11403
rect 6735 11085 7065 11097
rect 7835 11403 8165 11415
rect 7835 11097 7847 11403
rect 8153 11097 8165 11403
rect 7835 11085 8165 11097
rect 8935 11403 9265 11415
rect 8935 11097 8947 11403
rect 9253 11097 9265 11403
rect 8935 11085 9265 11097
rect 10035 11403 10365 11415
rect 10035 11097 10047 11403
rect 10353 11097 10365 11403
rect 10035 11085 10365 11097
rect 11135 11403 11465 11415
rect 11135 11097 11147 11403
rect 11453 11097 11465 11403
rect 11135 11085 11465 11097
rect 12235 11403 12565 11415
rect 12235 11097 12247 11403
rect 12553 11097 12565 11403
rect 12235 11085 12565 11097
rect 13335 11403 13665 11415
rect 13335 11097 13347 11403
rect 13653 11097 13665 11403
rect 13335 11085 13665 11097
rect -415 10853 -85 10865
rect -415 10547 -403 10853
rect -97 10547 -85 10853
rect -415 10535 -85 10547
rect 685 10853 1015 10865
rect 685 10547 697 10853
rect 1003 10547 1015 10853
rect 685 10535 1015 10547
rect 1785 10853 2115 10865
rect 1785 10547 1797 10853
rect 2103 10547 2115 10853
rect 1785 10535 2115 10547
rect 2885 10853 3215 10865
rect 2885 10547 2897 10853
rect 3203 10547 3215 10853
rect 2885 10535 3215 10547
rect 3985 10853 4315 10865
rect 3985 10547 3997 10853
rect 4303 10547 4315 10853
rect 3985 10535 4315 10547
rect 5085 10853 5415 10865
rect 5085 10547 5097 10853
rect 5403 10547 5415 10853
rect 5085 10535 5415 10547
rect 6185 10853 6515 10865
rect 6185 10547 6197 10853
rect 6503 10547 6515 10853
rect 6185 10535 6515 10547
rect 7285 10853 7615 10865
rect 7285 10547 7297 10853
rect 7603 10547 7615 10853
rect 7285 10535 7615 10547
rect 8385 10853 8715 10865
rect 8385 10547 8397 10853
rect 8703 10547 8715 10853
rect 8385 10535 8715 10547
rect 9485 10853 9815 10865
rect 9485 10547 9497 10853
rect 9803 10547 9815 10853
rect 9485 10535 9815 10547
rect 10585 10853 10915 10865
rect 10585 10547 10597 10853
rect 10903 10547 10915 10853
rect 10585 10535 10915 10547
rect 11685 10853 12015 10865
rect 11685 10547 11697 10853
rect 12003 10547 12015 10853
rect 11685 10535 12015 10547
rect 12785 10853 13115 10865
rect 12785 10547 12797 10853
rect 13103 10547 13115 10853
rect 12785 10535 13115 10547
rect 135 10303 465 10315
rect 135 9997 147 10303
rect 453 9997 465 10303
rect 135 9985 465 9997
rect 1235 10303 1565 10315
rect 1235 9997 1247 10303
rect 1553 9997 1565 10303
rect 1235 9985 1565 9997
rect 2335 10303 2665 10315
rect 2335 9997 2347 10303
rect 2653 9997 2665 10303
rect 2335 9985 2665 9997
rect 3435 10303 3765 10315
rect 3435 9997 3447 10303
rect 3753 9997 3765 10303
rect 3435 9985 3765 9997
rect 4535 10303 4865 10315
rect 4535 9997 4547 10303
rect 4853 9997 4865 10303
rect 4535 9985 4865 9997
rect 5635 10303 5965 10315
rect 5635 9997 5647 10303
rect 5953 9997 5965 10303
rect 5635 9985 5965 9997
rect 6735 10303 7065 10315
rect 6735 9997 6747 10303
rect 7053 9997 7065 10303
rect 6735 9985 7065 9997
rect 7835 10303 8165 10315
rect 7835 9997 7847 10303
rect 8153 9997 8165 10303
rect 7835 9985 8165 9997
rect 8935 10303 9265 10315
rect 8935 9997 8947 10303
rect 9253 9997 9265 10303
rect 8935 9985 9265 9997
rect 10035 10303 10365 10315
rect 10035 9997 10047 10303
rect 10353 9997 10365 10303
rect 10035 9985 10365 9997
rect 11135 10303 11465 10315
rect 11135 9997 11147 10303
rect 11453 9997 11465 10303
rect 11135 9985 11465 9997
rect 12235 10303 12565 10315
rect 12235 9997 12247 10303
rect 12553 9997 12565 10303
rect 12235 9985 12565 9997
rect 13335 10303 13665 10315
rect 13335 9997 13347 10303
rect 13653 9997 13665 10303
rect 13335 9985 13665 9997
rect -415 9753 -85 9765
rect -415 9447 -403 9753
rect -97 9447 -85 9753
rect -415 9435 -85 9447
rect 685 9753 1015 9765
rect 685 9447 697 9753
rect 1003 9447 1015 9753
rect 685 9435 1015 9447
rect 1785 9753 2115 9765
rect 1785 9447 1797 9753
rect 2103 9447 2115 9753
rect 1785 9435 2115 9447
rect 2885 9753 3215 9765
rect 2885 9447 2897 9753
rect 3203 9447 3215 9753
rect 2885 9435 3215 9447
rect 3985 9753 4315 9765
rect 3985 9447 3997 9753
rect 4303 9447 4315 9753
rect 3985 9435 4315 9447
rect 5085 9753 5415 9765
rect 5085 9447 5097 9753
rect 5403 9447 5415 9753
rect 5085 9435 5415 9447
rect 6185 9753 6515 9765
rect 6185 9447 6197 9753
rect 6503 9447 6515 9753
rect 6185 9435 6515 9447
rect 7285 9753 7615 9765
rect 7285 9447 7297 9753
rect 7603 9447 7615 9753
rect 7285 9435 7615 9447
rect 8385 9753 8715 9765
rect 8385 9447 8397 9753
rect 8703 9447 8715 9753
rect 8385 9435 8715 9447
rect 9485 9753 9815 9765
rect 9485 9447 9497 9753
rect 9803 9447 9815 9753
rect 9485 9435 9815 9447
rect 10585 9753 10915 9765
rect 10585 9447 10597 9753
rect 10903 9447 10915 9753
rect 10585 9435 10915 9447
rect 11685 9753 12015 9765
rect 11685 9447 11697 9753
rect 12003 9447 12015 9753
rect 11685 9435 12015 9447
rect 12785 9753 13115 9765
rect 12785 9447 12797 9753
rect 13103 9447 13115 9753
rect 12785 9435 13115 9447
rect 135 9203 465 9215
rect 135 8897 147 9203
rect 453 8897 465 9203
rect 135 8885 465 8897
rect 1235 9203 1565 9215
rect 1235 8897 1247 9203
rect 1553 8897 1565 9203
rect 1235 8885 1565 8897
rect 2335 9203 2665 9215
rect 2335 8897 2347 9203
rect 2653 8897 2665 9203
rect 2335 8885 2665 8897
rect 3435 9203 3765 9215
rect 3435 8897 3447 9203
rect 3753 8897 3765 9203
rect 3435 8885 3765 8897
rect 4535 9203 4865 9215
rect 4535 8897 4547 9203
rect 4853 8897 4865 9203
rect 4535 8885 4865 8897
rect 5635 9203 5965 9215
rect 5635 8897 5647 9203
rect 5953 8897 5965 9203
rect 5635 8885 5965 8897
rect 6735 9203 7065 9215
rect 6735 8897 6747 9203
rect 7053 8897 7065 9203
rect 6735 8885 7065 8897
rect 7835 9203 8165 9215
rect 7835 8897 7847 9203
rect 8153 8897 8165 9203
rect 7835 8885 8165 8897
rect 8935 9203 9265 9215
rect 8935 8897 8947 9203
rect 9253 8897 9265 9203
rect 8935 8885 9265 8897
rect 10035 9203 10365 9215
rect 10035 8897 10047 9203
rect 10353 8897 10365 9203
rect 10035 8885 10365 8897
rect 11135 9203 11465 9215
rect 11135 8897 11147 9203
rect 11453 8897 11465 9203
rect 11135 8885 11465 8897
rect 12235 9203 12565 9215
rect 12235 8897 12247 9203
rect 12553 8897 12565 9203
rect 12235 8885 12565 8897
rect 13335 9203 13665 9215
rect 13335 8897 13347 9203
rect 13653 8897 13665 9203
rect 13335 8885 13665 8897
rect -415 8653 -85 8665
rect -415 8347 -403 8653
rect -97 8347 -85 8653
rect -415 8335 -85 8347
rect 685 8653 1015 8665
rect 685 8347 697 8653
rect 1003 8347 1015 8653
rect 685 8335 1015 8347
rect 1785 8653 2115 8665
rect 1785 8347 1797 8653
rect 2103 8347 2115 8653
rect 1785 8335 2115 8347
rect 2885 8653 3215 8665
rect 2885 8347 2897 8653
rect 3203 8347 3215 8653
rect 2885 8335 3215 8347
rect 3985 8653 4315 8665
rect 3985 8347 3997 8653
rect 4303 8347 4315 8653
rect 3985 8335 4315 8347
rect 5085 8653 5415 8665
rect 5085 8347 5097 8653
rect 5403 8347 5415 8653
rect 5085 8335 5415 8347
rect 6185 8653 6515 8665
rect 6185 8347 6197 8653
rect 6503 8347 6515 8653
rect 6185 8335 6515 8347
rect 7285 8653 7615 8665
rect 7285 8347 7297 8653
rect 7603 8347 7615 8653
rect 7285 8335 7615 8347
rect 8385 8653 8715 8665
rect 8385 8347 8397 8653
rect 8703 8347 8715 8653
rect 8385 8335 8715 8347
rect 9485 8653 9815 8665
rect 9485 8347 9497 8653
rect 9803 8347 9815 8653
rect 9485 8335 9815 8347
rect 10585 8653 10915 8665
rect 10585 8347 10597 8653
rect 10903 8347 10915 8653
rect 10585 8335 10915 8347
rect 11685 8653 12015 8665
rect 11685 8347 11697 8653
rect 12003 8347 12015 8653
rect 11685 8335 12015 8347
rect 12785 8653 13115 8665
rect 12785 8347 12797 8653
rect 13103 8347 13115 8653
rect 12785 8335 13115 8347
rect 135 8103 465 8115
rect 135 7797 147 8103
rect 453 7797 465 8103
rect 135 7785 465 7797
rect 1235 8103 1565 8115
rect 1235 7797 1247 8103
rect 1553 7797 1565 8103
rect 1235 7785 1565 7797
rect 2335 8103 2665 8115
rect 2335 7797 2347 8103
rect 2653 7797 2665 8103
rect 2335 7785 2665 7797
rect 3435 8103 3765 8115
rect 3435 7797 3447 8103
rect 3753 7797 3765 8103
rect 3435 7785 3765 7797
rect 4535 8103 4865 8115
rect 4535 7797 4547 8103
rect 4853 7797 4865 8103
rect 4535 7785 4865 7797
rect 5635 8103 5965 8115
rect 5635 7797 5647 8103
rect 5953 7797 5965 8103
rect 5635 7785 5965 7797
rect 6735 8103 7065 8115
rect 6735 7797 6747 8103
rect 7053 7797 7065 8103
rect 6735 7785 7065 7797
rect 7835 8103 8165 8115
rect 7835 7797 7847 8103
rect 8153 7797 8165 8103
rect 7835 7785 8165 7797
rect 8935 8103 9265 8115
rect 8935 7797 8947 8103
rect 9253 7797 9265 8103
rect 8935 7785 9265 7797
rect 10035 8103 10365 8115
rect 10035 7797 10047 8103
rect 10353 7797 10365 8103
rect 10035 7785 10365 7797
rect 11135 8103 11465 8115
rect 11135 7797 11147 8103
rect 11453 7797 11465 8103
rect 11135 7785 11465 7797
rect 12235 8103 12565 8115
rect 12235 7797 12247 8103
rect 12553 7797 12565 8103
rect 12235 7785 12565 7797
rect 13335 8103 13665 8115
rect 13335 7797 13347 8103
rect 13653 7797 13665 8103
rect 13335 7785 13665 7797
rect -415 7553 -85 7565
rect -415 7247 -403 7553
rect -97 7247 -85 7553
rect -415 7235 -85 7247
rect 685 7553 1015 7565
rect 685 7247 697 7553
rect 1003 7247 1015 7553
rect 685 7235 1015 7247
rect 1785 7553 2115 7565
rect 1785 7247 1797 7553
rect 2103 7247 2115 7553
rect 1785 7235 2115 7247
rect 2885 7553 3215 7565
rect 2885 7247 2897 7553
rect 3203 7247 3215 7553
rect 2885 7235 3215 7247
rect 3985 7553 4315 7565
rect 3985 7247 3997 7553
rect 4303 7247 4315 7553
rect 3985 7235 4315 7247
rect 5085 7553 5415 7565
rect 5085 7247 5097 7553
rect 5403 7247 5415 7553
rect 5085 7235 5415 7247
rect 6185 7553 6515 7565
rect 6185 7247 6197 7553
rect 6503 7247 6515 7553
rect 6185 7235 6515 7247
rect 7285 7553 7615 7565
rect 7285 7247 7297 7553
rect 7603 7247 7615 7553
rect 7285 7235 7615 7247
rect 8385 7553 8715 7565
rect 8385 7247 8397 7553
rect 8703 7247 8715 7553
rect 8385 7235 8715 7247
rect 9485 7553 9815 7565
rect 9485 7247 9497 7553
rect 9803 7247 9815 7553
rect 9485 7235 9815 7247
rect 10585 7553 10915 7565
rect 10585 7247 10597 7553
rect 10903 7247 10915 7553
rect 10585 7235 10915 7247
rect 11685 7553 12015 7565
rect 11685 7247 11697 7553
rect 12003 7247 12015 7553
rect 11685 7235 12015 7247
rect 12785 7553 13115 7565
rect 12785 7247 12797 7553
rect 13103 7247 13115 7553
rect 12785 7235 13115 7247
rect 135 7003 465 7015
rect 135 6697 147 7003
rect 453 6697 465 7003
rect 135 6685 465 6697
rect 1235 7003 1565 7015
rect 1235 6697 1247 7003
rect 1553 6697 1565 7003
rect 1235 6685 1565 6697
rect 2335 7003 2665 7015
rect 2335 6697 2347 7003
rect 2653 6697 2665 7003
rect 2335 6685 2665 6697
rect 3435 7003 3765 7015
rect 3435 6697 3447 7003
rect 3753 6697 3765 7003
rect 3435 6685 3765 6697
rect 4535 7003 4865 7015
rect 4535 6697 4547 7003
rect 4853 6697 4865 7003
rect 4535 6685 4865 6697
rect 5635 7003 5965 7015
rect 5635 6697 5647 7003
rect 5953 6697 5965 7003
rect 5635 6685 5965 6697
rect 6735 7003 7065 7015
rect 6735 6697 6747 7003
rect 7053 6697 7065 7003
rect 6735 6685 7065 6697
rect 7835 7003 8165 7015
rect 7835 6697 7847 7003
rect 8153 6697 8165 7003
rect 7835 6685 8165 6697
rect 8935 7003 9265 7015
rect 8935 6697 8947 7003
rect 9253 6697 9265 7003
rect 8935 6685 9265 6697
rect 10035 7003 10365 7015
rect 10035 6697 10047 7003
rect 10353 6697 10365 7003
rect 10035 6685 10365 6697
rect 11135 7003 11465 7015
rect 11135 6697 11147 7003
rect 11453 6697 11465 7003
rect 11135 6685 11465 6697
rect 12235 7003 12565 7015
rect 12235 6697 12247 7003
rect 12553 6697 12565 7003
rect 12235 6685 12565 6697
rect 13335 7003 13665 7015
rect 13335 6697 13347 7003
rect 13653 6697 13665 7003
rect 13335 6685 13665 6697
rect -415 6453 -85 6465
rect -415 6147 -403 6453
rect -97 6147 -85 6453
rect -415 6135 -85 6147
rect 685 6453 1015 6465
rect 685 6147 697 6453
rect 1003 6147 1015 6453
rect 685 6135 1015 6147
rect 1785 6453 2115 6465
rect 1785 6147 1797 6453
rect 2103 6147 2115 6453
rect 1785 6135 2115 6147
rect 2885 6453 3215 6465
rect 2885 6147 2897 6453
rect 3203 6147 3215 6453
rect 2885 6135 3215 6147
rect 3985 6453 4315 6465
rect 3985 6147 3997 6453
rect 4303 6147 4315 6453
rect 3985 6135 4315 6147
rect 5085 6453 5415 6465
rect 5085 6147 5097 6453
rect 5403 6147 5415 6453
rect 5085 6135 5415 6147
rect 6185 6453 6515 6465
rect 6185 6147 6197 6453
rect 6503 6147 6515 6453
rect 6185 6135 6515 6147
rect 7285 6453 7615 6465
rect 7285 6147 7297 6453
rect 7603 6147 7615 6453
rect 7285 6135 7615 6147
rect 8385 6453 8715 6465
rect 8385 6147 8397 6453
rect 8703 6147 8715 6453
rect 8385 6135 8715 6147
rect 9485 6453 9815 6465
rect 9485 6147 9497 6453
rect 9803 6147 9815 6453
rect 9485 6135 9815 6147
rect 10585 6453 10915 6465
rect 10585 6147 10597 6453
rect 10903 6147 10915 6453
rect 10585 6135 10915 6147
rect 11685 6453 12015 6465
rect 11685 6147 11697 6453
rect 12003 6147 12015 6453
rect 11685 6135 12015 6147
rect 12785 6453 13115 6465
rect 12785 6147 12797 6453
rect 13103 6147 13115 6453
rect 12785 6135 13115 6147
rect 135 5903 465 5915
rect 135 5597 147 5903
rect 453 5597 465 5903
rect 135 5585 465 5597
rect 1235 5903 1565 5915
rect 1235 5597 1247 5903
rect 1553 5597 1565 5903
rect 1235 5585 1565 5597
rect 2335 5903 2665 5915
rect 2335 5597 2347 5903
rect 2653 5597 2665 5903
rect 2335 5585 2665 5597
rect 3435 5903 3765 5915
rect 3435 5597 3447 5903
rect 3753 5597 3765 5903
rect 3435 5585 3765 5597
rect 4535 5903 4865 5915
rect 4535 5597 4547 5903
rect 4853 5597 4865 5903
rect 4535 5585 4865 5597
rect 5635 5903 5965 5915
rect 5635 5597 5647 5903
rect 5953 5597 5965 5903
rect 5635 5585 5965 5597
rect 6735 5903 7065 5915
rect 6735 5597 6747 5903
rect 7053 5597 7065 5903
rect 6735 5585 7065 5597
rect 7835 5903 8165 5915
rect 7835 5597 7847 5903
rect 8153 5597 8165 5903
rect 7835 5585 8165 5597
rect 8935 5903 9265 5915
rect 8935 5597 8947 5903
rect 9253 5597 9265 5903
rect 8935 5585 9265 5597
rect 10035 5903 10365 5915
rect 10035 5597 10047 5903
rect 10353 5597 10365 5903
rect 10035 5585 10365 5597
rect 11135 5903 11465 5915
rect 11135 5597 11147 5903
rect 11453 5597 11465 5903
rect 11135 5585 11465 5597
rect 12235 5903 12565 5915
rect 12235 5597 12247 5903
rect 12553 5597 12565 5903
rect 12235 5585 12565 5597
rect 13335 5903 13665 5915
rect 13335 5597 13347 5903
rect 13653 5597 13665 5903
rect 13335 5585 13665 5597
rect -415 5353 -85 5365
rect -415 5047 -403 5353
rect -97 5047 -85 5353
rect -415 5035 -85 5047
rect 685 5353 1015 5365
rect 685 5047 697 5353
rect 1003 5047 1015 5353
rect 685 5035 1015 5047
rect 1785 5353 2115 5365
rect 1785 5047 1797 5353
rect 2103 5047 2115 5353
rect 1785 5035 2115 5047
rect 2885 5353 3215 5365
rect 2885 5047 2897 5353
rect 3203 5047 3215 5353
rect 2885 5035 3215 5047
rect 3985 5353 4315 5365
rect 3985 5047 3997 5353
rect 4303 5047 4315 5353
rect 3985 5035 4315 5047
rect 5085 5353 5415 5365
rect 5085 5047 5097 5353
rect 5403 5047 5415 5353
rect 5085 5035 5415 5047
rect 6185 5353 6515 5365
rect 6185 5047 6197 5353
rect 6503 5047 6515 5353
rect 6185 5035 6515 5047
rect 7285 5353 7615 5365
rect 7285 5047 7297 5353
rect 7603 5047 7615 5353
rect 7285 5035 7615 5047
rect 8385 5353 8715 5365
rect 8385 5047 8397 5353
rect 8703 5047 8715 5353
rect 8385 5035 8715 5047
rect 9485 5353 9815 5365
rect 9485 5047 9497 5353
rect 9803 5047 9815 5353
rect 9485 5035 9815 5047
rect 10585 5353 10915 5365
rect 10585 5047 10597 5353
rect 10903 5047 10915 5353
rect 10585 5035 10915 5047
rect 11685 5353 12015 5365
rect 11685 5047 11697 5353
rect 12003 5047 12015 5353
rect 11685 5035 12015 5047
rect 12785 5353 13115 5365
rect 12785 5047 12797 5353
rect 13103 5047 13115 5353
rect 12785 5035 13115 5047
rect 135 4803 465 4815
rect 135 4497 147 4803
rect 453 4497 465 4803
rect 135 4485 465 4497
rect 1235 4803 1565 4815
rect 1235 4497 1247 4803
rect 1553 4497 1565 4803
rect 1235 4485 1565 4497
rect 2335 4803 2665 4815
rect 2335 4497 2347 4803
rect 2653 4497 2665 4803
rect 2335 4485 2665 4497
rect 3435 4803 3765 4815
rect 3435 4497 3447 4803
rect 3753 4497 3765 4803
rect 3435 4485 3765 4497
rect 4535 4803 4865 4815
rect 4535 4497 4547 4803
rect 4853 4497 4865 4803
rect 4535 4485 4865 4497
rect 5635 4803 5965 4815
rect 5635 4497 5647 4803
rect 5953 4497 5965 4803
rect 5635 4485 5965 4497
rect 6735 4803 7065 4815
rect 6735 4497 6747 4803
rect 7053 4497 7065 4803
rect 6735 4485 7065 4497
rect 7835 4803 8165 4815
rect 7835 4497 7847 4803
rect 8153 4497 8165 4803
rect 7835 4485 8165 4497
rect 8935 4803 9265 4815
rect 8935 4497 8947 4803
rect 9253 4497 9265 4803
rect 8935 4485 9265 4497
rect 10035 4803 10365 4815
rect 10035 4497 10047 4803
rect 10353 4497 10365 4803
rect 10035 4485 10365 4497
rect 11135 4803 11465 4815
rect 11135 4497 11147 4803
rect 11453 4497 11465 4803
rect 11135 4485 11465 4497
rect 12235 4803 12565 4815
rect 12235 4497 12247 4803
rect 12553 4497 12565 4803
rect 12235 4485 12565 4497
rect 13335 4803 13665 4815
rect 13335 4497 13347 4803
rect 13653 4497 13665 4803
rect 13335 4485 13665 4497
rect -415 4253 -85 4265
rect -415 3947 -403 4253
rect -97 3947 -85 4253
rect -415 3935 -85 3947
rect 685 4253 1015 4265
rect 685 3947 697 4253
rect 1003 3947 1015 4253
rect 685 3935 1015 3947
rect 1785 4253 2115 4265
rect 1785 3947 1797 4253
rect 2103 3947 2115 4253
rect 1785 3935 2115 3947
rect 2885 4253 3215 4265
rect 2885 3947 2897 4253
rect 3203 3947 3215 4253
rect 2885 3935 3215 3947
rect 3985 4253 4315 4265
rect 3985 3947 3997 4253
rect 4303 3947 4315 4253
rect 3985 3935 4315 3947
rect 5085 4253 5415 4265
rect 5085 3947 5097 4253
rect 5403 3947 5415 4253
rect 5085 3935 5415 3947
rect 6185 4253 6515 4265
rect 6185 3947 6197 4253
rect 6503 3947 6515 4253
rect 6185 3935 6515 3947
rect 7285 4253 7615 4265
rect 7285 3947 7297 4253
rect 7603 3947 7615 4253
rect 7285 3935 7615 3947
rect 8385 4253 8715 4265
rect 8385 3947 8397 4253
rect 8703 3947 8715 4253
rect 8385 3935 8715 3947
rect 9485 4253 9815 4265
rect 9485 3947 9497 4253
rect 9803 3947 9815 4253
rect 9485 3935 9815 3947
rect 10585 4253 10915 4265
rect 10585 3947 10597 4253
rect 10903 3947 10915 4253
rect 10585 3935 10915 3947
rect 11685 4253 12015 4265
rect 11685 3947 11697 4253
rect 12003 3947 12015 4253
rect 11685 3935 12015 3947
rect 12785 4253 13115 4265
rect 12785 3947 12797 4253
rect 13103 3947 13115 4253
rect 12785 3935 13115 3947
rect 135 3703 465 3715
rect 135 3397 147 3703
rect 453 3397 465 3703
rect 135 3385 465 3397
rect 1235 3703 1565 3715
rect 1235 3397 1247 3703
rect 1553 3397 1565 3703
rect 1235 3385 1565 3397
rect 2335 3703 2665 3715
rect 2335 3397 2347 3703
rect 2653 3397 2665 3703
rect 2335 3385 2665 3397
rect 3435 3703 3765 3715
rect 3435 3397 3447 3703
rect 3753 3397 3765 3703
rect 3435 3385 3765 3397
rect 4535 3703 4865 3715
rect 4535 3397 4547 3703
rect 4853 3397 4865 3703
rect 4535 3385 4865 3397
rect 5635 3703 5965 3715
rect 5635 3397 5647 3703
rect 5953 3397 5965 3703
rect 5635 3385 5965 3397
rect 6735 3703 7065 3715
rect 6735 3397 6747 3703
rect 7053 3397 7065 3703
rect 6735 3385 7065 3397
rect 7835 3703 8165 3715
rect 7835 3397 7847 3703
rect 8153 3397 8165 3703
rect 7835 3385 8165 3397
rect 8935 3703 9265 3715
rect 8935 3397 8947 3703
rect 9253 3397 9265 3703
rect 8935 3385 9265 3397
rect 10035 3703 10365 3715
rect 10035 3397 10047 3703
rect 10353 3397 10365 3703
rect 10035 3385 10365 3397
rect 11135 3703 11465 3715
rect 11135 3397 11147 3703
rect 11453 3397 11465 3703
rect 11135 3385 11465 3397
rect 12235 3703 12565 3715
rect 12235 3397 12247 3703
rect 12553 3397 12565 3703
rect 12235 3385 12565 3397
rect 13335 3703 13665 3715
rect 13335 3397 13347 3703
rect 13653 3397 13665 3703
rect 13335 3385 13665 3397
rect -415 3153 -85 3165
rect -415 2847 -403 3153
rect -97 2847 -85 3153
rect -415 2835 -85 2847
rect 685 3153 1015 3165
rect 685 2847 697 3153
rect 1003 2847 1015 3153
rect 685 2835 1015 2847
rect 1785 3153 2115 3165
rect 1785 2847 1797 3153
rect 2103 2847 2115 3153
rect 1785 2835 2115 2847
rect 2885 3153 3215 3165
rect 2885 2847 2897 3153
rect 3203 2847 3215 3153
rect 2885 2835 3215 2847
rect 3985 3153 4315 3165
rect 3985 2847 3997 3153
rect 4303 2847 4315 3153
rect 3985 2835 4315 2847
rect 5085 3153 5415 3165
rect 5085 2847 5097 3153
rect 5403 2847 5415 3153
rect 5085 2835 5415 2847
rect 6185 3153 6515 3165
rect 6185 2847 6197 3153
rect 6503 2847 6515 3153
rect 6185 2835 6515 2847
rect 7285 3153 7615 3165
rect 7285 2847 7297 3153
rect 7603 2847 7615 3153
rect 7285 2835 7615 2847
rect 8385 3153 8715 3165
rect 8385 2847 8397 3153
rect 8703 2847 8715 3153
rect 8385 2835 8715 2847
rect 9485 3153 9815 3165
rect 9485 2847 9497 3153
rect 9803 2847 9815 3153
rect 9485 2835 9815 2847
rect 10585 3153 10915 3165
rect 10585 2847 10597 3153
rect 10903 2847 10915 3153
rect 10585 2835 10915 2847
rect 11685 3153 12015 3165
rect 11685 2847 11697 3153
rect 12003 2847 12015 3153
rect 11685 2835 12015 2847
rect 12785 3153 13115 3165
rect 12785 2847 12797 3153
rect 13103 2847 13115 3153
rect 12785 2835 13115 2847
rect 135 2603 465 2615
rect 135 2297 147 2603
rect 453 2297 465 2603
rect 135 2285 465 2297
rect 1235 2603 1565 2615
rect 1235 2297 1247 2603
rect 1553 2297 1565 2603
rect 1235 2285 1565 2297
rect 2335 2603 2665 2615
rect 2335 2297 2347 2603
rect 2653 2297 2665 2603
rect 2335 2285 2665 2297
rect 3435 2603 3765 2615
rect 3435 2297 3447 2603
rect 3753 2297 3765 2603
rect 3435 2285 3765 2297
rect 4535 2603 4865 2615
rect 4535 2297 4547 2603
rect 4853 2297 4865 2603
rect 4535 2285 4865 2297
rect 5635 2603 5965 2615
rect 5635 2297 5647 2603
rect 5953 2297 5965 2603
rect 5635 2285 5965 2297
rect 6735 2603 7065 2615
rect 6735 2297 6747 2603
rect 7053 2297 7065 2603
rect 6735 2285 7065 2297
rect 7835 2603 8165 2615
rect 7835 2297 7847 2603
rect 8153 2297 8165 2603
rect 7835 2285 8165 2297
rect 8935 2603 9265 2615
rect 8935 2297 8947 2603
rect 9253 2297 9265 2603
rect 8935 2285 9265 2297
rect 10035 2603 10365 2615
rect 10035 2297 10047 2603
rect 10353 2297 10365 2603
rect 10035 2285 10365 2297
rect 11135 2603 11465 2615
rect 11135 2297 11147 2603
rect 11453 2297 11465 2603
rect 11135 2285 11465 2297
rect 12235 2603 12565 2615
rect 12235 2297 12247 2603
rect 12553 2297 12565 2603
rect 12235 2285 12565 2297
rect 13335 2603 13665 2615
rect 13335 2297 13347 2603
rect 13653 2297 13665 2603
rect 13335 2285 13665 2297
rect -415 2053 -85 2065
rect -415 1747 -403 2053
rect -97 1747 -85 2053
rect -415 1735 -85 1747
rect 685 2053 1015 2065
rect 685 1747 697 2053
rect 1003 1747 1015 2053
rect 685 1735 1015 1747
rect 1785 2053 2115 2065
rect 1785 1747 1797 2053
rect 2103 1747 2115 2053
rect 1785 1735 2115 1747
rect 2885 2053 3215 2065
rect 2885 1747 2897 2053
rect 3203 1747 3215 2053
rect 2885 1735 3215 1747
rect 3985 2053 4315 2065
rect 3985 1747 3997 2053
rect 4303 1747 4315 2053
rect 3985 1735 4315 1747
rect 5085 2053 5415 2065
rect 5085 1747 5097 2053
rect 5403 1747 5415 2053
rect 5085 1735 5415 1747
rect 6185 2053 6515 2065
rect 6185 1747 6197 2053
rect 6503 1747 6515 2053
rect 6185 1735 6515 1747
rect 7285 2053 7615 2065
rect 7285 1747 7297 2053
rect 7603 1747 7615 2053
rect 7285 1735 7615 1747
rect 8385 2053 8715 2065
rect 8385 1747 8397 2053
rect 8703 1747 8715 2053
rect 8385 1735 8715 1747
rect 9485 2053 9815 2065
rect 9485 1747 9497 2053
rect 9803 1747 9815 2053
rect 9485 1735 9815 1747
rect 10585 2053 10915 2065
rect 10585 1747 10597 2053
rect 10903 1747 10915 2053
rect 10585 1735 10915 1747
rect 11685 2053 12015 2065
rect 11685 1747 11697 2053
rect 12003 1747 12015 2053
rect 11685 1735 12015 1747
rect 12785 2053 13115 2065
rect 12785 1747 12797 2053
rect 13103 1747 13115 2053
rect 12785 1735 13115 1747
rect 135 1503 465 1515
rect 135 1197 147 1503
rect 453 1197 465 1503
rect 135 1185 465 1197
rect 1235 1503 1565 1515
rect 1235 1197 1247 1503
rect 1553 1197 1565 1503
rect 1235 1185 1565 1197
rect 2335 1503 2665 1515
rect 2335 1197 2347 1503
rect 2653 1197 2665 1503
rect 2335 1185 2665 1197
rect 3435 1503 3765 1515
rect 3435 1197 3447 1503
rect 3753 1197 3765 1503
rect 3435 1185 3765 1197
rect 4535 1503 4865 1515
rect 4535 1197 4547 1503
rect 4853 1197 4865 1503
rect 4535 1185 4865 1197
rect 5635 1503 5965 1515
rect 5635 1197 5647 1503
rect 5953 1197 5965 1503
rect 5635 1185 5965 1197
rect 6735 1503 7065 1515
rect 6735 1197 6747 1503
rect 7053 1197 7065 1503
rect 6735 1185 7065 1197
rect 7835 1503 8165 1515
rect 7835 1197 7847 1503
rect 8153 1197 8165 1503
rect 7835 1185 8165 1197
rect 8935 1503 9265 1515
rect 8935 1197 8947 1503
rect 9253 1197 9265 1503
rect 8935 1185 9265 1197
rect 10035 1503 10365 1515
rect 10035 1197 10047 1503
rect 10353 1197 10365 1503
rect 10035 1185 10365 1197
rect 11135 1503 11465 1515
rect 11135 1197 11147 1503
rect 11453 1197 11465 1503
rect 11135 1185 11465 1197
rect 12235 1503 12565 1515
rect 12235 1197 12247 1503
rect 12553 1197 12565 1503
rect 12235 1185 12565 1197
rect 13335 1503 13665 1515
rect 13335 1197 13347 1503
rect 13653 1197 13665 1503
rect 13335 1185 13665 1197
rect -415 953 -85 965
rect -415 647 -403 953
rect -97 647 -85 953
rect -415 635 -85 647
rect 685 953 1015 965
rect 685 647 697 953
rect 1003 647 1015 953
rect 685 635 1015 647
rect 1785 953 2115 965
rect 1785 647 1797 953
rect 2103 647 2115 953
rect 1785 635 2115 647
rect 2885 953 3215 965
rect 2885 647 2897 953
rect 3203 647 3215 953
rect 2885 635 3215 647
rect 3985 953 4315 965
rect 3985 647 3997 953
rect 4303 647 4315 953
rect 3985 635 4315 647
rect 5085 953 5415 965
rect 5085 647 5097 953
rect 5403 647 5415 953
rect 5085 635 5415 647
rect 6185 953 6515 965
rect 6185 647 6197 953
rect 6503 647 6515 953
rect 6185 635 6515 647
rect 7285 953 7615 965
rect 7285 647 7297 953
rect 7603 647 7615 953
rect 7285 635 7615 647
rect 8385 953 8715 965
rect 8385 647 8397 953
rect 8703 647 8715 953
rect 8385 635 8715 647
rect 9485 953 9815 965
rect 9485 647 9497 953
rect 9803 647 9815 953
rect 9485 635 9815 647
rect 10585 953 10915 965
rect 10585 647 10597 953
rect 10903 647 10915 953
rect 10585 635 10915 647
rect 11685 953 12015 965
rect 11685 647 11697 953
rect 12003 647 12015 953
rect 11685 635 12015 647
rect 12785 953 13115 965
rect 12785 647 12797 953
rect 13103 647 13115 953
rect 12785 635 13115 647
rect 135 403 465 415
rect 135 97 147 403
rect 453 97 465 403
rect 135 85 465 97
rect 1235 403 1565 415
rect 1235 97 1247 403
rect 1553 97 1565 403
rect 1235 85 1565 97
rect 2335 403 2665 415
rect 2335 97 2347 403
rect 2653 97 2665 403
rect 2335 85 2665 97
rect 3435 403 3765 415
rect 3435 97 3447 403
rect 3753 97 3765 403
rect 3435 85 3765 97
rect 4535 403 4865 415
rect 4535 97 4547 403
rect 4853 97 4865 403
rect 4535 85 4865 97
rect 5635 403 5965 415
rect 5635 97 5647 403
rect 5953 97 5965 403
rect 5635 85 5965 97
rect 6735 403 7065 415
rect 6735 97 6747 403
rect 7053 97 7065 403
rect 6735 85 7065 97
rect 7835 403 8165 415
rect 7835 97 7847 403
rect 8153 97 8165 403
rect 7835 85 8165 97
rect 8935 403 9265 415
rect 8935 97 8947 403
rect 9253 97 9265 403
rect 8935 85 9265 97
rect 10035 403 10365 415
rect 10035 97 10047 403
rect 10353 97 10365 403
rect 10035 85 10365 97
rect 11135 403 11465 415
rect 11135 97 11147 403
rect 11453 97 11465 403
rect 11135 85 11465 97
rect 12235 403 12565 415
rect 12235 97 12247 403
rect 12553 97 12565 403
rect 12235 85 12565 97
rect 13335 403 13665 415
rect 13335 97 13347 403
rect 13653 97 13665 403
rect 13335 85 13665 97
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect 685 -147 1015 -135
rect 685 -453 697 -147
rect 1003 -453 1015 -147
rect 685 -465 1015 -453
rect 1785 -147 2115 -135
rect 1785 -453 1797 -147
rect 2103 -453 2115 -147
rect 1785 -465 2115 -453
rect 2885 -147 3215 -135
rect 2885 -453 2897 -147
rect 3203 -453 3215 -147
rect 2885 -465 3215 -453
rect 3985 -147 4315 -135
rect 3985 -453 3997 -147
rect 4303 -453 4315 -147
rect 3985 -465 4315 -453
rect 5085 -147 5415 -135
rect 5085 -453 5097 -147
rect 5403 -453 5415 -147
rect 5085 -465 5415 -453
rect 6185 -147 6515 -135
rect 6185 -453 6197 -147
rect 6503 -453 6515 -147
rect 6185 -465 6515 -453
rect 7285 -147 7615 -135
rect 7285 -453 7297 -147
rect 7603 -453 7615 -147
rect 7285 -465 7615 -453
rect 8385 -147 8715 -135
rect 8385 -453 8397 -147
rect 8703 -453 8715 -147
rect 8385 -465 8715 -453
rect 9485 -147 9815 -135
rect 9485 -453 9497 -147
rect 9803 -453 9815 -147
rect 9485 -465 9815 -453
rect 10585 -147 10915 -135
rect 10585 -453 10597 -147
rect 10903 -453 10915 -147
rect 10585 -465 10915 -453
rect 11685 -147 12015 -135
rect 11685 -453 11697 -147
rect 12003 -453 12015 -147
rect 11685 -465 12015 -453
rect 12785 -147 13115 -135
rect 12785 -453 12797 -147
rect 13103 -453 13115 -147
rect 12785 -465 13115 -453
rect 13975 13217 13987 13925
rect 14263 13217 14275 14213
rect 13975 13200 14275 13217
rect 13975 12669 13987 13200
rect 14263 12669 14275 13200
rect 13975 12650 14275 12669
rect 13975 12117 13987 12650
rect 14263 12117 14275 12650
rect 13975 12100 14275 12117
rect 13975 11569 13987 12100
rect 14263 11569 14275 12100
rect 13975 11550 14275 11569
rect 13975 11017 13987 11550
rect 14263 11017 14275 11550
rect 13975 11000 14275 11017
rect 13975 10469 13987 11000
rect 14263 10469 14275 11000
rect 13975 10450 14275 10469
rect 13975 9917 13987 10450
rect 14263 9917 14275 10450
rect 13975 9900 14275 9917
rect 13975 9369 13987 9900
rect 14263 9369 14275 9900
rect 13975 9350 14275 9369
rect 13975 8817 13987 9350
rect 14263 8817 14275 9350
rect 13975 8800 14275 8817
rect 13975 8269 13987 8800
rect 14263 8269 14275 8800
rect 13975 8250 14275 8269
rect 13975 7717 13987 8250
rect 14263 7717 14275 8250
rect 13975 7700 14275 7717
rect 13975 7169 13987 7700
rect 14263 7169 14275 7700
rect 13975 7150 14275 7169
rect 13975 6617 13987 7150
rect 14263 6617 14275 7150
rect 13975 6600 14275 6617
rect 13975 6069 13987 6600
rect 14263 6069 14275 6600
rect 13975 6050 14275 6069
rect 13975 5517 13987 6050
rect 14263 5517 14275 6050
rect 13975 5500 14275 5517
rect 13975 4969 13987 5500
rect 14263 4969 14275 5500
rect 13975 4950 14275 4969
rect 13975 4417 13987 4950
rect 14263 4417 14275 4950
rect 13975 4400 14275 4417
rect 13975 3869 13987 4400
rect 14263 3869 14275 4400
rect 13975 3850 14275 3869
rect 13975 3317 13987 3850
rect 14263 3317 14275 3850
rect 13975 3300 14275 3317
rect 13975 2769 13987 3300
rect 14263 2769 14275 3300
rect 13975 2750 14275 2769
rect 13975 2217 13987 2750
rect 14263 2217 14275 2750
rect 13975 2200 14275 2217
rect 13975 1669 13987 2200
rect 14263 1669 14275 2200
rect 13975 1650 14275 1669
rect 13975 1117 13987 1650
rect 14263 1117 14275 1650
rect 13975 1100 14275 1117
rect 13975 569 13987 1100
rect 14263 569 14275 1100
rect 13975 550 14275 569
rect 13975 17 13987 550
rect 14263 17 14275 550
rect 13975 0 14275 17
rect 13975 -775 13987 0
rect -737 -787 13987 -775
rect -17 -1063 0 -787
rect 531 -1063 550 -787
rect 1083 -1063 1100 -787
rect 1631 -1063 1650 -787
rect 2183 -1063 2200 -787
rect 2731 -1063 2750 -787
rect 3283 -1063 3300 -787
rect 3831 -1063 3850 -787
rect 4383 -1063 4400 -787
rect 4931 -1063 4950 -787
rect 5483 -1063 5500 -787
rect 6031 -1063 6050 -787
rect 6583 -1063 6600 -787
rect 7131 -1063 7150 -787
rect 7683 -1063 7700 -787
rect 8231 -1063 8250 -787
rect 8783 -1063 8800 -787
rect 9331 -1063 9350 -787
rect 9883 -1063 9900 -787
rect 10431 -1063 10450 -787
rect 10983 -1063 11000 -787
rect 11531 -1063 11550 -787
rect 12083 -1063 12100 -787
rect 12631 -1063 12650 -787
rect 13183 -1063 13200 -787
rect 14263 -1063 14275 0
rect -1025 -1075 14275 -1063
<< mvpsubdiffcont >>
rect -5513 14737 18763 18713
rect -5513 -1587 -1537 14737
rect 14787 -1587 18763 14737
rect -5513 -5563 18763 -1587
<< mvnsubdiffcont >>
rect -1013 13937 -17 14213
rect 0 13937 533 14213
rect 550 13937 1083 14213
rect 1100 13937 1633 14213
rect 1650 13937 2183 14213
rect 2200 13937 2733 14213
rect 2750 13937 3283 14213
rect 3300 13937 3833 14213
rect 3850 13937 4383 14213
rect 4400 13937 4933 14213
rect 4950 13937 5483 14213
rect 5500 13937 6033 14213
rect 6050 13937 6583 14213
rect 6600 13937 7133 14213
rect 7150 13937 7683 14213
rect 7700 13937 8233 14213
rect 8250 13937 8783 14213
rect 8800 13937 9333 14213
rect 9350 13937 9883 14213
rect 9900 13937 10433 14213
rect 10450 13937 10983 14213
rect 11000 13937 11533 14213
rect 11550 13937 12083 14213
rect 12100 13937 12633 14213
rect 12650 13937 13183 14213
rect 13200 13937 14263 14213
rect -1013 13217 -737 13937
rect -1013 12667 -737 13200
rect -1013 12117 -737 12650
rect -1013 11567 -737 12100
rect -1013 11017 -737 11550
rect -1013 10467 -737 11000
rect -1013 9917 -737 10450
rect -1013 9367 -737 9900
rect -1013 8817 -737 9350
rect -1013 8267 -737 8800
rect -1013 7717 -737 8250
rect -1013 7167 -737 7700
rect -1013 6617 -737 7150
rect -1013 6067 -737 6600
rect -1013 5517 -737 6050
rect -1013 4967 -737 5500
rect -1013 4417 -737 4950
rect -1013 3867 -737 4400
rect -1013 3317 -737 3850
rect -1013 2767 -737 3300
rect -1013 2217 -737 2750
rect -1013 1667 -737 2200
rect -1013 1117 -737 1650
rect -1013 567 -737 1100
rect -1013 17 -737 550
rect -1013 -787 -737 0
rect 147 13297 453 13603
rect 1247 13297 1553 13603
rect 2347 13297 2653 13603
rect 3447 13297 3753 13603
rect 4547 13297 4853 13603
rect 5647 13297 5953 13603
rect 6747 13297 7053 13603
rect 7847 13297 8153 13603
rect 8947 13297 9253 13603
rect 10047 13297 10353 13603
rect 11147 13297 11453 13603
rect 12247 13297 12553 13603
rect 13347 13297 13653 13603
rect -403 12747 -97 13053
rect 697 12747 1003 13053
rect 1797 12747 2103 13053
rect 2897 12747 3203 13053
rect 3997 12747 4303 13053
rect 5097 12747 5403 13053
rect 6197 12747 6503 13053
rect 7297 12747 7603 13053
rect 8397 12747 8703 13053
rect 9497 12747 9803 13053
rect 10597 12747 10903 13053
rect 11697 12747 12003 13053
rect 12797 12747 13103 13053
rect 147 12197 453 12503
rect 1247 12197 1553 12503
rect 2347 12197 2653 12503
rect 3447 12197 3753 12503
rect 4547 12197 4853 12503
rect 5647 12197 5953 12503
rect 6747 12197 7053 12503
rect 7847 12197 8153 12503
rect 8947 12197 9253 12503
rect 10047 12197 10353 12503
rect 11147 12197 11453 12503
rect 12247 12197 12553 12503
rect 13347 12197 13653 12503
rect -403 11647 -97 11953
rect 697 11647 1003 11953
rect 1797 11647 2103 11953
rect 2897 11647 3203 11953
rect 3997 11647 4303 11953
rect 5097 11647 5403 11953
rect 6197 11647 6503 11953
rect 7297 11647 7603 11953
rect 8397 11647 8703 11953
rect 9497 11647 9803 11953
rect 10597 11647 10903 11953
rect 11697 11647 12003 11953
rect 12797 11647 13103 11953
rect 147 11097 453 11403
rect 1247 11097 1553 11403
rect 2347 11097 2653 11403
rect 3447 11097 3753 11403
rect 4547 11097 4853 11403
rect 5647 11097 5953 11403
rect 6747 11097 7053 11403
rect 7847 11097 8153 11403
rect 8947 11097 9253 11403
rect 10047 11097 10353 11403
rect 11147 11097 11453 11403
rect 12247 11097 12553 11403
rect 13347 11097 13653 11403
rect -403 10547 -97 10853
rect 697 10547 1003 10853
rect 1797 10547 2103 10853
rect 2897 10547 3203 10853
rect 3997 10547 4303 10853
rect 5097 10547 5403 10853
rect 6197 10547 6503 10853
rect 7297 10547 7603 10853
rect 8397 10547 8703 10853
rect 9497 10547 9803 10853
rect 10597 10547 10903 10853
rect 11697 10547 12003 10853
rect 12797 10547 13103 10853
rect 147 9997 453 10303
rect 1247 9997 1553 10303
rect 2347 9997 2653 10303
rect 3447 9997 3753 10303
rect 4547 9997 4853 10303
rect 5647 9997 5953 10303
rect 6747 9997 7053 10303
rect 7847 9997 8153 10303
rect 8947 9997 9253 10303
rect 10047 9997 10353 10303
rect 11147 9997 11453 10303
rect 12247 9997 12553 10303
rect 13347 9997 13653 10303
rect -403 9447 -97 9753
rect 697 9447 1003 9753
rect 1797 9447 2103 9753
rect 2897 9447 3203 9753
rect 3997 9447 4303 9753
rect 5097 9447 5403 9753
rect 6197 9447 6503 9753
rect 7297 9447 7603 9753
rect 8397 9447 8703 9753
rect 9497 9447 9803 9753
rect 10597 9447 10903 9753
rect 11697 9447 12003 9753
rect 12797 9447 13103 9753
rect 147 8897 453 9203
rect 1247 8897 1553 9203
rect 2347 8897 2653 9203
rect 3447 8897 3753 9203
rect 4547 8897 4853 9203
rect 5647 8897 5953 9203
rect 6747 8897 7053 9203
rect 7847 8897 8153 9203
rect 8947 8897 9253 9203
rect 10047 8897 10353 9203
rect 11147 8897 11453 9203
rect 12247 8897 12553 9203
rect 13347 8897 13653 9203
rect -403 8347 -97 8653
rect 697 8347 1003 8653
rect 1797 8347 2103 8653
rect 2897 8347 3203 8653
rect 3997 8347 4303 8653
rect 5097 8347 5403 8653
rect 6197 8347 6503 8653
rect 7297 8347 7603 8653
rect 8397 8347 8703 8653
rect 9497 8347 9803 8653
rect 10597 8347 10903 8653
rect 11697 8347 12003 8653
rect 12797 8347 13103 8653
rect 147 7797 453 8103
rect 1247 7797 1553 8103
rect 2347 7797 2653 8103
rect 3447 7797 3753 8103
rect 4547 7797 4853 8103
rect 5647 7797 5953 8103
rect 6747 7797 7053 8103
rect 7847 7797 8153 8103
rect 8947 7797 9253 8103
rect 10047 7797 10353 8103
rect 11147 7797 11453 8103
rect 12247 7797 12553 8103
rect 13347 7797 13653 8103
rect -403 7247 -97 7553
rect 697 7247 1003 7553
rect 1797 7247 2103 7553
rect 2897 7247 3203 7553
rect 3997 7247 4303 7553
rect 5097 7247 5403 7553
rect 6197 7247 6503 7553
rect 7297 7247 7603 7553
rect 8397 7247 8703 7553
rect 9497 7247 9803 7553
rect 10597 7247 10903 7553
rect 11697 7247 12003 7553
rect 12797 7247 13103 7553
rect 147 6697 453 7003
rect 1247 6697 1553 7003
rect 2347 6697 2653 7003
rect 3447 6697 3753 7003
rect 4547 6697 4853 7003
rect 5647 6697 5953 7003
rect 6747 6697 7053 7003
rect 7847 6697 8153 7003
rect 8947 6697 9253 7003
rect 10047 6697 10353 7003
rect 11147 6697 11453 7003
rect 12247 6697 12553 7003
rect 13347 6697 13653 7003
rect -403 6147 -97 6453
rect 697 6147 1003 6453
rect 1797 6147 2103 6453
rect 2897 6147 3203 6453
rect 3997 6147 4303 6453
rect 5097 6147 5403 6453
rect 6197 6147 6503 6453
rect 7297 6147 7603 6453
rect 8397 6147 8703 6453
rect 9497 6147 9803 6453
rect 10597 6147 10903 6453
rect 11697 6147 12003 6453
rect 12797 6147 13103 6453
rect 147 5597 453 5903
rect 1247 5597 1553 5903
rect 2347 5597 2653 5903
rect 3447 5597 3753 5903
rect 4547 5597 4853 5903
rect 5647 5597 5953 5903
rect 6747 5597 7053 5903
rect 7847 5597 8153 5903
rect 8947 5597 9253 5903
rect 10047 5597 10353 5903
rect 11147 5597 11453 5903
rect 12247 5597 12553 5903
rect 13347 5597 13653 5903
rect -403 5047 -97 5353
rect 697 5047 1003 5353
rect 1797 5047 2103 5353
rect 2897 5047 3203 5353
rect 3997 5047 4303 5353
rect 5097 5047 5403 5353
rect 6197 5047 6503 5353
rect 7297 5047 7603 5353
rect 8397 5047 8703 5353
rect 9497 5047 9803 5353
rect 10597 5047 10903 5353
rect 11697 5047 12003 5353
rect 12797 5047 13103 5353
rect 147 4497 453 4803
rect 1247 4497 1553 4803
rect 2347 4497 2653 4803
rect 3447 4497 3753 4803
rect 4547 4497 4853 4803
rect 5647 4497 5953 4803
rect 6747 4497 7053 4803
rect 7847 4497 8153 4803
rect 8947 4497 9253 4803
rect 10047 4497 10353 4803
rect 11147 4497 11453 4803
rect 12247 4497 12553 4803
rect 13347 4497 13653 4803
rect -403 3947 -97 4253
rect 697 3947 1003 4253
rect 1797 3947 2103 4253
rect 2897 3947 3203 4253
rect 3997 3947 4303 4253
rect 5097 3947 5403 4253
rect 6197 3947 6503 4253
rect 7297 3947 7603 4253
rect 8397 3947 8703 4253
rect 9497 3947 9803 4253
rect 10597 3947 10903 4253
rect 11697 3947 12003 4253
rect 12797 3947 13103 4253
rect 147 3397 453 3703
rect 1247 3397 1553 3703
rect 2347 3397 2653 3703
rect 3447 3397 3753 3703
rect 4547 3397 4853 3703
rect 5647 3397 5953 3703
rect 6747 3397 7053 3703
rect 7847 3397 8153 3703
rect 8947 3397 9253 3703
rect 10047 3397 10353 3703
rect 11147 3397 11453 3703
rect 12247 3397 12553 3703
rect 13347 3397 13653 3703
rect -403 2847 -97 3153
rect 697 2847 1003 3153
rect 1797 2847 2103 3153
rect 2897 2847 3203 3153
rect 3997 2847 4303 3153
rect 5097 2847 5403 3153
rect 6197 2847 6503 3153
rect 7297 2847 7603 3153
rect 8397 2847 8703 3153
rect 9497 2847 9803 3153
rect 10597 2847 10903 3153
rect 11697 2847 12003 3153
rect 12797 2847 13103 3153
rect 147 2297 453 2603
rect 1247 2297 1553 2603
rect 2347 2297 2653 2603
rect 3447 2297 3753 2603
rect 4547 2297 4853 2603
rect 5647 2297 5953 2603
rect 6747 2297 7053 2603
rect 7847 2297 8153 2603
rect 8947 2297 9253 2603
rect 10047 2297 10353 2603
rect 11147 2297 11453 2603
rect 12247 2297 12553 2603
rect 13347 2297 13653 2603
rect -403 1747 -97 2053
rect 697 1747 1003 2053
rect 1797 1747 2103 2053
rect 2897 1747 3203 2053
rect 3997 1747 4303 2053
rect 5097 1747 5403 2053
rect 6197 1747 6503 2053
rect 7297 1747 7603 2053
rect 8397 1747 8703 2053
rect 9497 1747 9803 2053
rect 10597 1747 10903 2053
rect 11697 1747 12003 2053
rect 12797 1747 13103 2053
rect 147 1197 453 1503
rect 1247 1197 1553 1503
rect 2347 1197 2653 1503
rect 3447 1197 3753 1503
rect 4547 1197 4853 1503
rect 5647 1197 5953 1503
rect 6747 1197 7053 1503
rect 7847 1197 8153 1503
rect 8947 1197 9253 1503
rect 10047 1197 10353 1503
rect 11147 1197 11453 1503
rect 12247 1197 12553 1503
rect 13347 1197 13653 1503
rect -403 647 -97 953
rect 697 647 1003 953
rect 1797 647 2103 953
rect 2897 647 3203 953
rect 3997 647 4303 953
rect 5097 647 5403 953
rect 6197 647 6503 953
rect 7297 647 7603 953
rect 8397 647 8703 953
rect 9497 647 9803 953
rect 10597 647 10903 953
rect 11697 647 12003 953
rect 12797 647 13103 953
rect 147 97 453 403
rect 1247 97 1553 403
rect 2347 97 2653 403
rect 3447 97 3753 403
rect 4547 97 4853 403
rect 5647 97 5953 403
rect 6747 97 7053 403
rect 7847 97 8153 403
rect 8947 97 9253 403
rect 10047 97 10353 403
rect 11147 97 11453 403
rect 12247 97 12553 403
rect 13347 97 13653 403
rect -403 -453 -97 -147
rect 697 -453 1003 -147
rect 1797 -453 2103 -147
rect 2897 -453 3203 -147
rect 3997 -453 4303 -147
rect 5097 -453 5403 -147
rect 6197 -453 6503 -147
rect 7297 -453 7603 -147
rect 8397 -453 8703 -147
rect 9497 -453 9803 -147
rect 10597 -453 10903 -147
rect 11697 -453 12003 -147
rect 12797 -453 13103 -147
rect 13987 13217 14263 13937
rect 13987 12669 14263 13200
rect 13987 12117 14263 12650
rect 13987 11569 14263 12100
rect 13987 11017 14263 11550
rect 13987 10469 14263 11000
rect 13987 9917 14263 10450
rect 13987 9369 14263 9900
rect 13987 8817 14263 9350
rect 13987 8269 14263 8800
rect 13987 7717 14263 8250
rect 13987 7169 14263 7700
rect 13987 6617 14263 7150
rect 13987 6069 14263 6600
rect 13987 5517 14263 6050
rect 13987 4969 14263 5500
rect 13987 4417 14263 4950
rect 13987 3869 14263 4400
rect 13987 3317 14263 3850
rect 13987 2769 14263 3300
rect 13987 2217 14263 2750
rect 13987 1669 14263 2200
rect 13987 1117 14263 1650
rect 13987 569 14263 1100
rect 13987 17 14263 550
rect 13987 -787 14263 0
rect -1013 -1063 -17 -787
rect 0 -1063 531 -787
rect 550 -1063 1083 -787
rect 1100 -1063 1631 -787
rect 1650 -1063 2183 -787
rect 2200 -1063 2731 -787
rect 2750 -1063 3283 -787
rect 3300 -1063 3831 -787
rect 3850 -1063 4383 -787
rect 4400 -1063 4931 -787
rect 4950 -1063 5483 -787
rect 5500 -1063 6031 -787
rect 6050 -1063 6583 -787
rect 6600 -1063 7131 -787
rect 7150 -1063 7683 -787
rect 7700 -1063 8231 -787
rect 8250 -1063 8783 -787
rect 8800 -1063 9331 -787
rect 9350 -1063 9883 -787
rect 9900 -1063 10431 -787
rect 10450 -1063 10983 -787
rect 11000 -1063 11531 -787
rect 11550 -1063 12083 -787
rect 12100 -1063 12631 -787
rect 12650 -1063 13183 -787
rect 13200 -1063 14263 -787
<< poly >>
rect -550 13742 13800 13750
rect -550 13708 -542 13742
rect -508 13708 8 13742
rect 42 13708 558 13742
rect 592 13708 1108 13742
rect 1142 13708 1658 13742
rect 1692 13708 2208 13742
rect 2242 13708 2758 13742
rect 2792 13708 3308 13742
rect 3342 13708 3858 13742
rect 3892 13708 4408 13742
rect 4442 13708 4958 13742
rect 4992 13708 5508 13742
rect 5542 13708 6058 13742
rect 6092 13708 6608 13742
rect 6642 13708 7158 13742
rect 7192 13708 7708 13742
rect 7742 13708 8258 13742
rect 8292 13708 8808 13742
rect 8842 13708 9358 13742
rect 9392 13708 9908 13742
rect 9942 13708 10458 13742
rect 10492 13708 11008 13742
rect 11042 13708 11558 13742
rect 11592 13708 12108 13742
rect 12142 13708 12658 13742
rect 12692 13708 13208 13742
rect 13242 13708 13758 13742
rect 13792 13708 13800 13742
rect -550 13700 13800 13708
rect -550 13200 -500 13700
rect 0 13669 50 13700
rect 550 13669 600 13700
rect 1100 13669 1150 13700
rect 1650 13669 1700 13700
rect 2200 13669 2250 13700
rect 2750 13669 2800 13700
rect 3300 13669 3350 13700
rect 3850 13669 3900 13700
rect 4400 13669 4450 13700
rect 4950 13669 5000 13700
rect 5500 13669 5550 13700
rect 6050 13669 6100 13700
rect 6600 13669 6650 13700
rect 7150 13669 7200 13700
rect 7700 13669 7750 13700
rect 8250 13669 8300 13700
rect 8800 13669 8850 13700
rect 9350 13669 9400 13700
rect 9900 13669 9950 13700
rect 10450 13669 10500 13700
rect 11000 13669 11050 13700
rect 11550 13669 11600 13700
rect 12100 13669 12150 13700
rect 12650 13669 12700 13700
rect 13200 13669 13250 13700
rect 0 13200 50 13231
rect 550 13200 600 13231
rect 1100 13200 1150 13231
rect 1650 13200 1700 13231
rect 2200 13200 2250 13231
rect 2750 13200 2800 13231
rect 3300 13200 3350 13231
rect 3850 13200 3900 13231
rect 4400 13200 4450 13231
rect 4950 13200 5000 13231
rect 5500 13200 5550 13231
rect 6050 13200 6100 13231
rect 6600 13200 6650 13231
rect 7150 13200 7200 13231
rect 7700 13200 7750 13231
rect 8250 13200 8300 13231
rect 8800 13200 8850 13231
rect 9350 13200 9400 13231
rect 9900 13200 9950 13231
rect 10450 13200 10500 13231
rect 11000 13200 11050 13231
rect 11550 13200 11600 13231
rect 12100 13200 12150 13231
rect 12650 13200 12700 13231
rect 13200 13200 13250 13231
rect 13750 13200 13800 13700
rect -550 13192 -469 13200
rect -550 13158 -542 13192
rect -508 13158 -469 13192
rect -550 13150 -469 13158
rect -31 13192 81 13200
rect -31 13158 8 13192
rect 42 13158 81 13192
rect -31 13150 81 13158
rect 519 13192 631 13200
rect 519 13158 558 13192
rect 592 13158 631 13192
rect 519 13150 631 13158
rect 1069 13192 1181 13200
rect 1069 13158 1108 13192
rect 1142 13158 1181 13192
rect 1069 13150 1181 13158
rect 1619 13192 1731 13200
rect 1619 13158 1658 13192
rect 1692 13158 1731 13192
rect 1619 13150 1731 13158
rect 2169 13192 2281 13200
rect 2169 13158 2208 13192
rect 2242 13158 2281 13192
rect 2169 13150 2281 13158
rect 2719 13192 2831 13200
rect 2719 13158 2758 13192
rect 2792 13158 2831 13192
rect 2719 13150 2831 13158
rect 3269 13192 3381 13200
rect 3269 13158 3308 13192
rect 3342 13158 3381 13192
rect 3269 13150 3381 13158
rect 3819 13192 3931 13200
rect 3819 13158 3858 13192
rect 3892 13158 3931 13192
rect 3819 13150 3931 13158
rect 4369 13192 4481 13200
rect 4369 13158 4408 13192
rect 4442 13158 4481 13192
rect 4369 13150 4481 13158
rect 4919 13192 5031 13200
rect 4919 13158 4958 13192
rect 4992 13158 5031 13192
rect 4919 13150 5031 13158
rect 5469 13192 5581 13200
rect 5469 13158 5508 13192
rect 5542 13158 5581 13192
rect 5469 13150 5581 13158
rect 6019 13192 6131 13200
rect 6019 13158 6058 13192
rect 6092 13158 6131 13192
rect 6019 13150 6131 13158
rect 6569 13192 6681 13200
rect 6569 13158 6608 13192
rect 6642 13158 6681 13192
rect 6569 13150 6681 13158
rect 7119 13192 7231 13200
rect 7119 13158 7158 13192
rect 7192 13158 7231 13192
rect 7119 13150 7231 13158
rect 7669 13192 7781 13200
rect 7669 13158 7708 13192
rect 7742 13158 7781 13192
rect 7669 13150 7781 13158
rect 8219 13192 8331 13200
rect 8219 13158 8258 13192
rect 8292 13158 8331 13192
rect 8219 13150 8331 13158
rect 8769 13192 8881 13200
rect 8769 13158 8808 13192
rect 8842 13158 8881 13192
rect 8769 13150 8881 13158
rect 9319 13192 9431 13200
rect 9319 13158 9358 13192
rect 9392 13158 9431 13192
rect 9319 13150 9431 13158
rect 9869 13192 9981 13200
rect 9869 13158 9908 13192
rect 9942 13158 9981 13192
rect 9869 13150 9981 13158
rect 10419 13192 10531 13200
rect 10419 13158 10458 13192
rect 10492 13158 10531 13192
rect 10419 13150 10531 13158
rect 10969 13192 11081 13200
rect 10969 13158 11008 13192
rect 11042 13158 11081 13192
rect 10969 13150 11081 13158
rect 11519 13192 11631 13200
rect 11519 13158 11558 13192
rect 11592 13158 11631 13192
rect 11519 13150 11631 13158
rect 12069 13192 12181 13200
rect 12069 13158 12108 13192
rect 12142 13158 12181 13192
rect 12069 13150 12181 13158
rect 12619 13192 12731 13200
rect 12619 13158 12658 13192
rect 12692 13158 12731 13192
rect 12619 13150 12731 13158
rect 13169 13192 13281 13200
rect 13169 13158 13208 13192
rect 13242 13158 13281 13192
rect 13169 13150 13281 13158
rect 13719 13192 13800 13200
rect 13719 13158 13758 13192
rect 13792 13158 13800 13192
rect 13719 13150 13800 13158
rect -550 12650 -500 13150
rect 0 13119 50 13150
rect 550 13119 600 13150
rect 1100 13119 1150 13150
rect 0 12650 50 12681
rect 1650 13119 1700 13150
rect 2200 13119 2250 13150
rect 550 12650 600 12681
rect 1100 12650 1150 12681
rect 2750 13119 2800 13150
rect 3300 13119 3350 13150
rect 1650 12650 1700 12681
rect 2200 12650 2250 12681
rect 3850 13119 3900 13150
rect 4400 13119 4450 13150
rect 2750 12650 2800 12681
rect 3300 12650 3350 12681
rect 4950 13119 5000 13150
rect 5500 13119 5550 13150
rect 3850 12650 3900 12681
rect 4400 12650 4450 12681
rect 6050 13119 6100 13150
rect 6600 13119 6650 13150
rect 4950 12650 5000 12681
rect 5500 12650 5550 12681
rect 7150 13119 7200 13150
rect 7700 13119 7750 13150
rect 6050 12650 6100 12681
rect 6600 12650 6650 12681
rect 8250 13119 8300 13150
rect 8800 13119 8850 13150
rect 7150 12650 7200 12681
rect 7700 12650 7750 12681
rect 9350 13119 9400 13150
rect 9900 13119 9950 13150
rect 8250 12650 8300 12681
rect 8800 12650 8850 12681
rect 10450 13119 10500 13150
rect 11000 13119 11050 13150
rect 9350 12650 9400 12681
rect 9900 12650 9950 12681
rect 11550 13119 11600 13150
rect 12100 13119 12150 13150
rect 10450 12650 10500 12681
rect 11000 12650 11050 12681
rect 12650 13119 12700 13150
rect 13200 13119 13250 13150
rect 11550 12650 11600 12681
rect 12100 12650 12150 12681
rect 12650 12650 12700 12681
rect 13200 12650 13250 12681
rect 13750 12650 13800 13150
rect -550 12642 -469 12650
rect -550 12608 -542 12642
rect -508 12608 -469 12642
rect -550 12600 -469 12608
rect -31 12642 81 12650
rect -31 12608 8 12642
rect 42 12608 81 12642
rect -31 12600 81 12608
rect 519 12642 631 12650
rect 519 12608 558 12642
rect 592 12608 631 12642
rect 519 12600 631 12608
rect 1069 12642 1181 12650
rect 1069 12608 1108 12642
rect 1142 12608 1181 12642
rect 1069 12600 1181 12608
rect 1619 12642 1731 12650
rect 1619 12608 1658 12642
rect 1692 12608 1731 12642
rect 1619 12600 1731 12608
rect 2169 12642 2281 12650
rect 2169 12608 2208 12642
rect 2242 12608 2281 12642
rect 2169 12600 2281 12608
rect 2719 12642 2831 12650
rect 2719 12608 2758 12642
rect 2792 12608 2831 12642
rect 2719 12600 2831 12608
rect 3269 12642 3381 12650
rect 3269 12608 3308 12642
rect 3342 12608 3381 12642
rect 3269 12600 3381 12608
rect 3819 12642 3931 12650
rect 3819 12608 3858 12642
rect 3892 12608 3931 12642
rect 3819 12600 3931 12608
rect 4369 12642 4481 12650
rect 4369 12608 4408 12642
rect 4442 12608 4481 12642
rect 4369 12600 4481 12608
rect 4919 12642 5031 12650
rect 4919 12608 4958 12642
rect 4992 12608 5031 12642
rect 4919 12600 5031 12608
rect 5469 12642 5581 12650
rect 5469 12608 5508 12642
rect 5542 12608 5581 12642
rect 5469 12600 5581 12608
rect 6019 12642 6131 12650
rect 6019 12608 6058 12642
rect 6092 12608 6131 12642
rect 6019 12600 6131 12608
rect 6569 12642 6681 12650
rect 6569 12608 6608 12642
rect 6642 12608 6681 12642
rect 6569 12600 6681 12608
rect 7119 12642 7231 12650
rect 7119 12608 7158 12642
rect 7192 12608 7231 12642
rect 7119 12600 7231 12608
rect 7669 12642 7781 12650
rect 7669 12608 7708 12642
rect 7742 12608 7781 12642
rect 7669 12600 7781 12608
rect 8219 12642 8331 12650
rect 8219 12608 8258 12642
rect 8292 12608 8331 12642
rect 8219 12600 8331 12608
rect 8769 12642 8881 12650
rect 8769 12608 8808 12642
rect 8842 12608 8881 12642
rect 8769 12600 8881 12608
rect 9319 12642 9431 12650
rect 9319 12608 9358 12642
rect 9392 12608 9431 12642
rect 9319 12600 9431 12608
rect 9869 12642 9981 12650
rect 9869 12608 9908 12642
rect 9942 12608 9981 12642
rect 9869 12600 9981 12608
rect 10419 12642 10531 12650
rect 10419 12608 10458 12642
rect 10492 12608 10531 12642
rect 10419 12600 10531 12608
rect 10969 12642 11081 12650
rect 10969 12608 11008 12642
rect 11042 12608 11081 12642
rect 10969 12600 11081 12608
rect 11519 12642 11631 12650
rect 11519 12608 11558 12642
rect 11592 12608 11631 12642
rect 11519 12600 11631 12608
rect 12069 12642 12181 12650
rect 12069 12608 12108 12642
rect 12142 12608 12181 12642
rect 12069 12600 12181 12608
rect 12619 12642 12731 12650
rect 12619 12608 12658 12642
rect 12692 12608 12731 12642
rect 12619 12600 12731 12608
rect 13169 12642 13281 12650
rect 13169 12608 13208 12642
rect 13242 12608 13281 12642
rect 13169 12600 13281 12608
rect 13719 12642 13800 12650
rect 13719 12608 13758 12642
rect 13792 12608 13800 12642
rect 13719 12600 13800 12608
rect -550 12100 -500 12600
rect 0 12569 50 12600
rect 550 12569 600 12600
rect 1100 12569 1150 12600
rect 1650 12569 1700 12600
rect 0 12100 50 12131
rect 550 12100 600 12131
rect 2200 12569 2250 12600
rect 2750 12569 2800 12600
rect 1100 12100 1150 12131
rect 1650 12100 1700 12131
rect 3300 12569 3350 12600
rect 3850 12569 3900 12600
rect 2200 12100 2250 12131
rect 2750 12100 2800 12131
rect 4400 12569 4450 12600
rect 4950 12569 5000 12600
rect 3300 12100 3350 12131
rect 3850 12100 3900 12131
rect 5500 12569 5550 12600
rect 6050 12569 6100 12600
rect 4400 12100 4450 12131
rect 4950 12100 5000 12131
rect 6600 12569 6650 12600
rect 7150 12569 7200 12600
rect 5500 12100 5550 12131
rect 6050 12100 6100 12131
rect 7700 12569 7750 12600
rect 8250 12569 8300 12600
rect 6600 12100 6650 12131
rect 7150 12100 7200 12131
rect 8800 12569 8850 12600
rect 9350 12569 9400 12600
rect 7700 12100 7750 12131
rect 8250 12100 8300 12131
rect 9900 12569 9950 12600
rect 10450 12569 10500 12600
rect 8800 12100 8850 12131
rect 9350 12100 9400 12131
rect 11000 12569 11050 12600
rect 11550 12569 11600 12600
rect 9900 12100 9950 12131
rect 10450 12100 10500 12131
rect 12100 12569 12150 12600
rect 12650 12569 12700 12600
rect 11000 12100 11050 12131
rect 11550 12100 11600 12131
rect 13200 12569 13250 12600
rect 12100 12100 12150 12131
rect 12650 12100 12700 12131
rect 13200 12100 13250 12131
rect 13750 12100 13800 12600
rect -550 12092 -469 12100
rect -550 12058 -542 12092
rect -508 12058 -469 12092
rect -550 12050 -469 12058
rect -31 12092 81 12100
rect -31 12058 8 12092
rect 42 12058 81 12092
rect -31 12050 81 12058
rect 519 12092 631 12100
rect 519 12058 558 12092
rect 592 12058 631 12092
rect 519 12050 631 12058
rect 1069 12092 1181 12100
rect 1069 12058 1108 12092
rect 1142 12058 1181 12092
rect 1069 12050 1181 12058
rect 1619 12092 1731 12100
rect 1619 12058 1658 12092
rect 1692 12058 1731 12092
rect 1619 12050 1731 12058
rect 2169 12092 2281 12100
rect 2169 12058 2208 12092
rect 2242 12058 2281 12092
rect 2169 12050 2281 12058
rect 2719 12092 2831 12100
rect 2719 12058 2758 12092
rect 2792 12058 2831 12092
rect 2719 12050 2831 12058
rect 3269 12092 3381 12100
rect 3269 12058 3308 12092
rect 3342 12058 3381 12092
rect 3269 12050 3381 12058
rect 3819 12092 3931 12100
rect 3819 12058 3858 12092
rect 3892 12058 3931 12092
rect 3819 12050 3931 12058
rect 4369 12092 4481 12100
rect 4369 12058 4408 12092
rect 4442 12058 4481 12092
rect 4369 12050 4481 12058
rect 4919 12092 5031 12100
rect 4919 12058 4958 12092
rect 4992 12058 5031 12092
rect 4919 12050 5031 12058
rect 5469 12092 5581 12100
rect 5469 12058 5508 12092
rect 5542 12058 5581 12092
rect 5469 12050 5581 12058
rect 6019 12092 6131 12100
rect 6019 12058 6058 12092
rect 6092 12058 6131 12092
rect 6019 12050 6131 12058
rect 6569 12092 6681 12100
rect 6569 12058 6608 12092
rect 6642 12058 6681 12092
rect 6569 12050 6681 12058
rect 7119 12092 7231 12100
rect 7119 12058 7158 12092
rect 7192 12058 7231 12092
rect 7119 12050 7231 12058
rect 7669 12092 7781 12100
rect 7669 12058 7708 12092
rect 7742 12058 7781 12092
rect 7669 12050 7781 12058
rect 8219 12092 8331 12100
rect 8219 12058 8258 12092
rect 8292 12058 8331 12092
rect 8219 12050 8331 12058
rect 8769 12092 8881 12100
rect 8769 12058 8808 12092
rect 8842 12058 8881 12092
rect 8769 12050 8881 12058
rect 9319 12092 9431 12100
rect 9319 12058 9358 12092
rect 9392 12058 9431 12092
rect 9319 12050 9431 12058
rect 9869 12092 9981 12100
rect 9869 12058 9908 12092
rect 9942 12058 9981 12092
rect 9869 12050 9981 12058
rect 10419 12092 10531 12100
rect 10419 12058 10458 12092
rect 10492 12058 10531 12092
rect 10419 12050 10531 12058
rect 10969 12092 11081 12100
rect 10969 12058 11008 12092
rect 11042 12058 11081 12092
rect 10969 12050 11081 12058
rect 11519 12092 11631 12100
rect 11519 12058 11558 12092
rect 11592 12058 11631 12092
rect 11519 12050 11631 12058
rect 12069 12092 12181 12100
rect 12069 12058 12108 12092
rect 12142 12058 12181 12092
rect 12069 12050 12181 12058
rect 12619 12092 12731 12100
rect 12619 12058 12658 12092
rect 12692 12058 12731 12092
rect 12619 12050 12731 12058
rect 13169 12092 13281 12100
rect 13169 12058 13208 12092
rect 13242 12058 13281 12092
rect 13169 12050 13281 12058
rect 13719 12092 13800 12100
rect 13719 12058 13758 12092
rect 13792 12058 13800 12092
rect 13719 12050 13800 12058
rect -550 11550 -500 12050
rect 0 12019 50 12050
rect 550 12019 600 12050
rect 1100 12019 1150 12050
rect 0 11550 50 11581
rect 1650 12019 1700 12050
rect 2200 12019 2250 12050
rect 550 11550 600 11581
rect 1100 11550 1150 11581
rect 2750 12019 2800 12050
rect 3300 12019 3350 12050
rect 1650 11550 1700 11581
rect 2200 11550 2250 11581
rect 3850 12019 3900 12050
rect 4400 12019 4450 12050
rect 2750 11550 2800 11581
rect 3300 11550 3350 11581
rect 4950 12019 5000 12050
rect 5500 12019 5550 12050
rect 3850 11550 3900 11581
rect 4400 11550 4450 11581
rect 6050 12019 6100 12050
rect 6600 12019 6650 12050
rect 4950 11550 5000 11581
rect 5500 11550 5550 11581
rect 7150 12019 7200 12050
rect 7700 12019 7750 12050
rect 6050 11550 6100 11581
rect 6600 11550 6650 11581
rect 8250 12019 8300 12050
rect 8800 12019 8850 12050
rect 7150 11550 7200 11581
rect 7700 11550 7750 11581
rect 9350 12019 9400 12050
rect 9900 12019 9950 12050
rect 8250 11550 8300 11581
rect 8800 11550 8850 11581
rect 10450 12019 10500 12050
rect 11000 12019 11050 12050
rect 9350 11550 9400 11581
rect 9900 11550 9950 11581
rect 11550 12019 11600 12050
rect 12100 12019 12150 12050
rect 10450 11550 10500 11581
rect 11000 11550 11050 11581
rect 12650 12019 12700 12050
rect 13200 12019 13250 12050
rect 11550 11550 11600 11581
rect 12100 11550 12150 11581
rect 12650 11550 12700 11581
rect 13200 11550 13250 11581
rect 13750 11550 13800 12050
rect -550 11542 -469 11550
rect -550 11508 -542 11542
rect -508 11508 -469 11542
rect -550 11500 -469 11508
rect -31 11542 81 11550
rect -31 11508 8 11542
rect 42 11508 81 11542
rect -31 11500 81 11508
rect 519 11542 631 11550
rect 519 11508 558 11542
rect 592 11508 631 11542
rect 519 11500 631 11508
rect 1069 11542 1181 11550
rect 1069 11508 1108 11542
rect 1142 11508 1181 11542
rect 1069 11500 1181 11508
rect 1619 11542 1731 11550
rect 1619 11508 1658 11542
rect 1692 11508 1731 11542
rect 1619 11500 1731 11508
rect 2169 11542 2281 11550
rect 2169 11508 2208 11542
rect 2242 11508 2281 11542
rect 2169 11500 2281 11508
rect 2719 11542 2831 11550
rect 2719 11508 2758 11542
rect 2792 11508 2831 11542
rect 2719 11500 2831 11508
rect 3269 11542 3381 11550
rect 3269 11508 3308 11542
rect 3342 11508 3381 11542
rect 3269 11500 3381 11508
rect 3819 11542 3931 11550
rect 3819 11508 3858 11542
rect 3892 11508 3931 11542
rect 3819 11500 3931 11508
rect 4369 11542 4481 11550
rect 4369 11508 4408 11542
rect 4442 11508 4481 11542
rect 4369 11500 4481 11508
rect 4919 11542 5031 11550
rect 4919 11508 4958 11542
rect 4992 11508 5031 11542
rect 4919 11500 5031 11508
rect 5469 11542 5581 11550
rect 5469 11508 5508 11542
rect 5542 11508 5581 11542
rect 5469 11500 5581 11508
rect 6019 11542 6131 11550
rect 6019 11508 6058 11542
rect 6092 11508 6131 11542
rect 6019 11500 6131 11508
rect 6569 11542 6681 11550
rect 6569 11508 6608 11542
rect 6642 11508 6681 11542
rect 6569 11500 6681 11508
rect 7119 11542 7231 11550
rect 7119 11508 7158 11542
rect 7192 11508 7231 11542
rect 7119 11500 7231 11508
rect 7669 11542 7781 11550
rect 7669 11508 7708 11542
rect 7742 11508 7781 11542
rect 7669 11500 7781 11508
rect 8219 11542 8331 11550
rect 8219 11508 8258 11542
rect 8292 11508 8331 11542
rect 8219 11500 8331 11508
rect 8769 11542 8881 11550
rect 8769 11508 8808 11542
rect 8842 11508 8881 11542
rect 8769 11500 8881 11508
rect 9319 11542 9431 11550
rect 9319 11508 9358 11542
rect 9392 11508 9431 11542
rect 9319 11500 9431 11508
rect 9869 11542 9981 11550
rect 9869 11508 9908 11542
rect 9942 11508 9981 11542
rect 9869 11500 9981 11508
rect 10419 11542 10531 11550
rect 10419 11508 10458 11542
rect 10492 11508 10531 11542
rect 10419 11500 10531 11508
rect 10969 11542 11081 11550
rect 10969 11508 11008 11542
rect 11042 11508 11081 11542
rect 10969 11500 11081 11508
rect 11519 11542 11631 11550
rect 11519 11508 11558 11542
rect 11592 11508 11631 11542
rect 11519 11500 11631 11508
rect 12069 11542 12181 11550
rect 12069 11508 12108 11542
rect 12142 11508 12181 11542
rect 12069 11500 12181 11508
rect 12619 11542 12731 11550
rect 12619 11508 12658 11542
rect 12692 11508 12731 11542
rect 12619 11500 12731 11508
rect 13169 11542 13281 11550
rect 13169 11508 13208 11542
rect 13242 11508 13281 11542
rect 13169 11500 13281 11508
rect 13719 11542 13800 11550
rect 13719 11508 13758 11542
rect 13792 11508 13800 11542
rect 13719 11500 13800 11508
rect -550 11000 -500 11500
rect 0 11469 50 11500
rect 550 11469 600 11500
rect 1100 11469 1150 11500
rect 1650 11469 1700 11500
rect 0 11000 50 11031
rect 550 11000 600 11031
rect 2200 11469 2250 11500
rect 2750 11469 2800 11500
rect 1100 11000 1150 11031
rect 1650 11000 1700 11031
rect 3300 11469 3350 11500
rect 3850 11469 3900 11500
rect 2200 11000 2250 11031
rect 2750 11000 2800 11031
rect 4400 11469 4450 11500
rect 4950 11469 5000 11500
rect 3300 11000 3350 11031
rect 3850 11000 3900 11031
rect 5500 11469 5550 11500
rect 6050 11469 6100 11500
rect 4400 11000 4450 11031
rect 4950 11000 5000 11031
rect 6600 11469 6650 11500
rect 7150 11469 7200 11500
rect 5500 11000 5550 11031
rect 6050 11000 6100 11031
rect 7700 11469 7750 11500
rect 8250 11469 8300 11500
rect 6600 11000 6650 11031
rect 7150 11000 7200 11031
rect 8800 11469 8850 11500
rect 9350 11469 9400 11500
rect 7700 11000 7750 11031
rect 8250 11000 8300 11031
rect 9900 11469 9950 11500
rect 10450 11469 10500 11500
rect 8800 11000 8850 11031
rect 9350 11000 9400 11031
rect 11000 11469 11050 11500
rect 11550 11469 11600 11500
rect 9900 11000 9950 11031
rect 10450 11000 10500 11031
rect 12100 11469 12150 11500
rect 12650 11469 12700 11500
rect 11000 11000 11050 11031
rect 11550 11000 11600 11031
rect 13200 11469 13250 11500
rect 12100 11000 12150 11031
rect 12650 11000 12700 11031
rect 13200 11000 13250 11031
rect 13750 11000 13800 11500
rect -550 10992 -469 11000
rect -550 10958 -542 10992
rect -508 10958 -469 10992
rect -550 10950 -469 10958
rect -31 10992 81 11000
rect -31 10958 8 10992
rect 42 10958 81 10992
rect -31 10950 81 10958
rect 519 10992 631 11000
rect 519 10958 558 10992
rect 592 10958 631 10992
rect 519 10950 631 10958
rect 1069 10992 1181 11000
rect 1069 10958 1108 10992
rect 1142 10958 1181 10992
rect 1069 10950 1181 10958
rect 1619 10992 1731 11000
rect 1619 10958 1658 10992
rect 1692 10958 1731 10992
rect 1619 10950 1731 10958
rect 2169 10992 2281 11000
rect 2169 10958 2208 10992
rect 2242 10958 2281 10992
rect 2169 10950 2281 10958
rect 2719 10992 2831 11000
rect 2719 10958 2758 10992
rect 2792 10958 2831 10992
rect 2719 10950 2831 10958
rect 3269 10992 3381 11000
rect 3269 10958 3308 10992
rect 3342 10958 3381 10992
rect 3269 10950 3381 10958
rect 3819 10992 3931 11000
rect 3819 10958 3858 10992
rect 3892 10958 3931 10992
rect 3819 10950 3931 10958
rect 4369 10992 4481 11000
rect 4369 10958 4408 10992
rect 4442 10958 4481 10992
rect 4369 10950 4481 10958
rect 4919 10992 5031 11000
rect 4919 10958 4958 10992
rect 4992 10958 5031 10992
rect 4919 10950 5031 10958
rect 5469 10992 5581 11000
rect 5469 10958 5508 10992
rect 5542 10958 5581 10992
rect 5469 10950 5581 10958
rect 6019 10992 6131 11000
rect 6019 10958 6058 10992
rect 6092 10958 6131 10992
rect 6019 10950 6131 10958
rect 6569 10992 6681 11000
rect 6569 10958 6608 10992
rect 6642 10958 6681 10992
rect 6569 10950 6681 10958
rect 7119 10992 7231 11000
rect 7119 10958 7158 10992
rect 7192 10958 7231 10992
rect 7119 10950 7231 10958
rect 7669 10992 7781 11000
rect 7669 10958 7708 10992
rect 7742 10958 7781 10992
rect 7669 10950 7781 10958
rect 8219 10992 8331 11000
rect 8219 10958 8258 10992
rect 8292 10958 8331 10992
rect 8219 10950 8331 10958
rect 8769 10992 8881 11000
rect 8769 10958 8808 10992
rect 8842 10958 8881 10992
rect 8769 10950 8881 10958
rect 9319 10992 9431 11000
rect 9319 10958 9358 10992
rect 9392 10958 9431 10992
rect 9319 10950 9431 10958
rect 9869 10992 9981 11000
rect 9869 10958 9908 10992
rect 9942 10958 9981 10992
rect 9869 10950 9981 10958
rect 10419 10992 10531 11000
rect 10419 10958 10458 10992
rect 10492 10958 10531 10992
rect 10419 10950 10531 10958
rect 10969 10992 11081 11000
rect 10969 10958 11008 10992
rect 11042 10958 11081 10992
rect 10969 10950 11081 10958
rect 11519 10992 11631 11000
rect 11519 10958 11558 10992
rect 11592 10958 11631 10992
rect 11519 10950 11631 10958
rect 12069 10992 12181 11000
rect 12069 10958 12108 10992
rect 12142 10958 12181 10992
rect 12069 10950 12181 10958
rect 12619 10992 12731 11000
rect 12619 10958 12658 10992
rect 12692 10958 12731 10992
rect 12619 10950 12731 10958
rect 13169 10992 13281 11000
rect 13169 10958 13208 10992
rect 13242 10958 13281 10992
rect 13169 10950 13281 10958
rect 13719 10992 13800 11000
rect 13719 10958 13758 10992
rect 13792 10958 13800 10992
rect 13719 10950 13800 10958
rect -550 10450 -500 10950
rect 0 10919 50 10950
rect 550 10919 600 10950
rect 1100 10919 1150 10950
rect 0 10450 50 10481
rect 1650 10919 1700 10950
rect 2200 10919 2250 10950
rect 550 10450 600 10481
rect 1100 10450 1150 10481
rect 2750 10919 2800 10950
rect 3300 10919 3350 10950
rect 1650 10450 1700 10481
rect 2200 10450 2250 10481
rect 3850 10919 3900 10950
rect 4400 10919 4450 10950
rect 2750 10450 2800 10481
rect 3300 10450 3350 10481
rect 4950 10919 5000 10950
rect 5500 10919 5550 10950
rect 3850 10450 3900 10481
rect 4400 10450 4450 10481
rect 6050 10919 6100 10950
rect 6600 10919 6650 10950
rect 4950 10450 5000 10481
rect 5500 10450 5550 10481
rect 7150 10919 7200 10950
rect 7700 10919 7750 10950
rect 6050 10450 6100 10481
rect 6600 10450 6650 10481
rect 8250 10919 8300 10950
rect 8800 10919 8850 10950
rect 7150 10450 7200 10481
rect 7700 10450 7750 10481
rect 9350 10919 9400 10950
rect 9900 10919 9950 10950
rect 8250 10450 8300 10481
rect 8800 10450 8850 10481
rect 10450 10919 10500 10950
rect 11000 10919 11050 10950
rect 9350 10450 9400 10481
rect 9900 10450 9950 10481
rect 11550 10919 11600 10950
rect 12100 10919 12150 10950
rect 10450 10450 10500 10481
rect 11000 10450 11050 10481
rect 12650 10919 12700 10950
rect 13200 10919 13250 10950
rect 11550 10450 11600 10481
rect 12100 10450 12150 10481
rect 12650 10450 12700 10481
rect 13200 10450 13250 10481
rect 13750 10450 13800 10950
rect -550 10442 -469 10450
rect -550 10408 -542 10442
rect -508 10408 -469 10442
rect -550 10400 -469 10408
rect -31 10442 81 10450
rect -31 10408 8 10442
rect 42 10408 81 10442
rect -31 10400 81 10408
rect 519 10442 631 10450
rect 519 10408 558 10442
rect 592 10408 631 10442
rect 519 10400 631 10408
rect 1069 10442 1181 10450
rect 1069 10408 1108 10442
rect 1142 10408 1181 10442
rect 1069 10400 1181 10408
rect 1619 10442 1731 10450
rect 1619 10408 1658 10442
rect 1692 10408 1731 10442
rect 1619 10400 1731 10408
rect 2169 10442 2281 10450
rect 2169 10408 2208 10442
rect 2242 10408 2281 10442
rect 2169 10400 2281 10408
rect 2719 10442 2831 10450
rect 2719 10408 2758 10442
rect 2792 10408 2831 10442
rect 2719 10400 2831 10408
rect 3269 10442 3381 10450
rect 3269 10408 3308 10442
rect 3342 10408 3381 10442
rect 3269 10400 3381 10408
rect 3819 10442 3931 10450
rect 3819 10408 3858 10442
rect 3892 10408 3931 10442
rect 3819 10400 3931 10408
rect 4369 10442 4481 10450
rect 4369 10408 4408 10442
rect 4442 10408 4481 10442
rect 4369 10400 4481 10408
rect 4919 10442 5031 10450
rect 4919 10408 4958 10442
rect 4992 10408 5031 10442
rect 4919 10400 5031 10408
rect 5469 10442 5581 10450
rect 5469 10408 5508 10442
rect 5542 10408 5581 10442
rect 5469 10400 5581 10408
rect 6019 10442 6131 10450
rect 6019 10408 6058 10442
rect 6092 10408 6131 10442
rect 6019 10400 6131 10408
rect 6569 10442 6681 10450
rect 6569 10408 6608 10442
rect 6642 10408 6681 10442
rect 6569 10400 6681 10408
rect 7119 10442 7231 10450
rect 7119 10408 7158 10442
rect 7192 10408 7231 10442
rect 7119 10400 7231 10408
rect 7669 10442 7781 10450
rect 7669 10408 7708 10442
rect 7742 10408 7781 10442
rect 7669 10400 7781 10408
rect 8219 10442 8331 10450
rect 8219 10408 8258 10442
rect 8292 10408 8331 10442
rect 8219 10400 8331 10408
rect 8769 10442 8881 10450
rect 8769 10408 8808 10442
rect 8842 10408 8881 10442
rect 8769 10400 8881 10408
rect 9319 10442 9431 10450
rect 9319 10408 9358 10442
rect 9392 10408 9431 10442
rect 9319 10400 9431 10408
rect 9869 10442 9981 10450
rect 9869 10408 9908 10442
rect 9942 10408 9981 10442
rect 9869 10400 9981 10408
rect 10419 10442 10531 10450
rect 10419 10408 10458 10442
rect 10492 10408 10531 10442
rect 10419 10400 10531 10408
rect 10969 10442 11081 10450
rect 10969 10408 11008 10442
rect 11042 10408 11081 10442
rect 10969 10400 11081 10408
rect 11519 10442 11631 10450
rect 11519 10408 11558 10442
rect 11592 10408 11631 10442
rect 11519 10400 11631 10408
rect 12069 10442 12181 10450
rect 12069 10408 12108 10442
rect 12142 10408 12181 10442
rect 12069 10400 12181 10408
rect 12619 10442 12731 10450
rect 12619 10408 12658 10442
rect 12692 10408 12731 10442
rect 12619 10400 12731 10408
rect 13169 10442 13281 10450
rect 13169 10408 13208 10442
rect 13242 10408 13281 10442
rect 13169 10400 13281 10408
rect 13719 10442 13800 10450
rect 13719 10408 13758 10442
rect 13792 10408 13800 10442
rect 13719 10400 13800 10408
rect -550 9900 -500 10400
rect 0 10369 50 10400
rect 550 10369 600 10400
rect 1100 10369 1150 10400
rect 1650 10369 1700 10400
rect 0 9900 50 9931
rect 550 9900 600 9931
rect 2200 10369 2250 10400
rect 2750 10369 2800 10400
rect 1100 9900 1150 9931
rect 1650 9900 1700 9931
rect 3300 10369 3350 10400
rect 3850 10369 3900 10400
rect 2200 9900 2250 9931
rect 2750 9900 2800 9931
rect 4400 10369 4450 10400
rect 4950 10369 5000 10400
rect 3300 9900 3350 9931
rect 3850 9900 3900 9931
rect 5500 10369 5550 10400
rect 6050 10369 6100 10400
rect 4400 9900 4450 9931
rect 4950 9900 5000 9931
rect 6600 10369 6650 10400
rect 7150 10369 7200 10400
rect 5500 9900 5550 9931
rect 6050 9900 6100 9931
rect 7700 10369 7750 10400
rect 8250 10369 8300 10400
rect 6600 9900 6650 9931
rect 7150 9900 7200 9931
rect 8800 10369 8850 10400
rect 9350 10369 9400 10400
rect 7700 9900 7750 9931
rect 8250 9900 8300 9931
rect 9900 10369 9950 10400
rect 10450 10369 10500 10400
rect 8800 9900 8850 9931
rect 9350 9900 9400 9931
rect 11000 10369 11050 10400
rect 11550 10369 11600 10400
rect 9900 9900 9950 9931
rect 10450 9900 10500 9931
rect 12100 10369 12150 10400
rect 12650 10369 12700 10400
rect 11000 9900 11050 9931
rect 11550 9900 11600 9931
rect 13200 10369 13250 10400
rect 12100 9900 12150 9931
rect 12650 9900 12700 9931
rect 13200 9900 13250 9931
rect 13750 9900 13800 10400
rect -550 9892 -469 9900
rect -550 9858 -542 9892
rect -508 9858 -469 9892
rect -550 9850 -469 9858
rect -31 9892 81 9900
rect -31 9858 8 9892
rect 42 9858 81 9892
rect -31 9850 81 9858
rect 519 9892 631 9900
rect 519 9858 558 9892
rect 592 9858 631 9892
rect 519 9850 631 9858
rect 1069 9892 1181 9900
rect 1069 9858 1108 9892
rect 1142 9858 1181 9892
rect 1069 9850 1181 9858
rect 1619 9892 1731 9900
rect 1619 9858 1658 9892
rect 1692 9858 1731 9892
rect 1619 9850 1731 9858
rect 2169 9892 2281 9900
rect 2169 9858 2208 9892
rect 2242 9858 2281 9892
rect 2169 9850 2281 9858
rect 2719 9892 2831 9900
rect 2719 9858 2758 9892
rect 2792 9858 2831 9892
rect 2719 9850 2831 9858
rect 3269 9892 3381 9900
rect 3269 9858 3308 9892
rect 3342 9858 3381 9892
rect 3269 9850 3381 9858
rect 3819 9892 3931 9900
rect 3819 9858 3858 9892
rect 3892 9858 3931 9892
rect 3819 9850 3931 9858
rect 4369 9892 4481 9900
rect 4369 9858 4408 9892
rect 4442 9858 4481 9892
rect 4369 9850 4481 9858
rect 4919 9892 5031 9900
rect 4919 9858 4958 9892
rect 4992 9858 5031 9892
rect 4919 9850 5031 9858
rect 5469 9892 5581 9900
rect 5469 9858 5508 9892
rect 5542 9858 5581 9892
rect 5469 9850 5581 9858
rect 6019 9892 6131 9900
rect 6019 9858 6058 9892
rect 6092 9858 6131 9892
rect 6019 9850 6131 9858
rect 6569 9892 6681 9900
rect 6569 9858 6608 9892
rect 6642 9858 6681 9892
rect 6569 9850 6681 9858
rect 7119 9892 7231 9900
rect 7119 9858 7158 9892
rect 7192 9858 7231 9892
rect 7119 9850 7231 9858
rect 7669 9892 7781 9900
rect 7669 9858 7708 9892
rect 7742 9858 7781 9892
rect 7669 9850 7781 9858
rect 8219 9892 8331 9900
rect 8219 9858 8258 9892
rect 8292 9858 8331 9892
rect 8219 9850 8331 9858
rect 8769 9892 8881 9900
rect 8769 9858 8808 9892
rect 8842 9858 8881 9892
rect 8769 9850 8881 9858
rect 9319 9892 9431 9900
rect 9319 9858 9358 9892
rect 9392 9858 9431 9892
rect 9319 9850 9431 9858
rect 9869 9892 9981 9900
rect 9869 9858 9908 9892
rect 9942 9858 9981 9892
rect 9869 9850 9981 9858
rect 10419 9892 10531 9900
rect 10419 9858 10458 9892
rect 10492 9858 10531 9892
rect 10419 9850 10531 9858
rect 10969 9892 11081 9900
rect 10969 9858 11008 9892
rect 11042 9858 11081 9892
rect 10969 9850 11081 9858
rect 11519 9892 11631 9900
rect 11519 9858 11558 9892
rect 11592 9858 11631 9892
rect 11519 9850 11631 9858
rect 12069 9892 12181 9900
rect 12069 9858 12108 9892
rect 12142 9858 12181 9892
rect 12069 9850 12181 9858
rect 12619 9892 12731 9900
rect 12619 9858 12658 9892
rect 12692 9858 12731 9892
rect 12619 9850 12731 9858
rect 13169 9892 13281 9900
rect 13169 9858 13208 9892
rect 13242 9858 13281 9892
rect 13169 9850 13281 9858
rect 13719 9892 13800 9900
rect 13719 9858 13758 9892
rect 13792 9858 13800 9892
rect 13719 9850 13800 9858
rect -550 9350 -500 9850
rect 0 9819 50 9850
rect 550 9819 600 9850
rect 1100 9819 1150 9850
rect 0 9350 50 9381
rect 1650 9819 1700 9850
rect 2200 9819 2250 9850
rect 550 9350 600 9381
rect 1100 9350 1150 9381
rect 2750 9819 2800 9850
rect 3300 9819 3350 9850
rect 1650 9350 1700 9381
rect 2200 9350 2250 9381
rect 3850 9819 3900 9850
rect 4400 9819 4450 9850
rect 2750 9350 2800 9381
rect 3300 9350 3350 9381
rect 4950 9819 5000 9850
rect 5500 9819 5550 9850
rect 3850 9350 3900 9381
rect 4400 9350 4450 9381
rect 6050 9819 6100 9850
rect 6600 9819 6650 9850
rect 4950 9350 5000 9381
rect 5500 9350 5550 9381
rect 7150 9819 7200 9850
rect 7700 9819 7750 9850
rect 6050 9350 6100 9381
rect 6600 9350 6650 9381
rect 8250 9819 8300 9850
rect 8800 9819 8850 9850
rect 7150 9350 7200 9381
rect 7700 9350 7750 9381
rect 9350 9819 9400 9850
rect 9900 9819 9950 9850
rect 8250 9350 8300 9381
rect 8800 9350 8850 9381
rect 10450 9819 10500 9850
rect 11000 9819 11050 9850
rect 9350 9350 9400 9381
rect 9900 9350 9950 9381
rect 11550 9819 11600 9850
rect 12100 9819 12150 9850
rect 10450 9350 10500 9381
rect 11000 9350 11050 9381
rect 12650 9819 12700 9850
rect 13200 9819 13250 9850
rect 11550 9350 11600 9381
rect 12100 9350 12150 9381
rect 12650 9350 12700 9381
rect 13200 9350 13250 9381
rect 13750 9350 13800 9850
rect -550 9342 -469 9350
rect -550 9308 -542 9342
rect -508 9308 -469 9342
rect -550 9300 -469 9308
rect -31 9342 81 9350
rect -31 9308 8 9342
rect 42 9308 81 9342
rect -31 9300 81 9308
rect 519 9342 631 9350
rect 519 9308 558 9342
rect 592 9308 631 9342
rect 519 9300 631 9308
rect 1069 9342 1181 9350
rect 1069 9308 1108 9342
rect 1142 9308 1181 9342
rect 1069 9300 1181 9308
rect 1619 9342 1731 9350
rect 1619 9308 1658 9342
rect 1692 9308 1731 9342
rect 1619 9300 1731 9308
rect 2169 9342 2281 9350
rect 2169 9308 2208 9342
rect 2242 9308 2281 9342
rect 2169 9300 2281 9308
rect 2719 9342 2831 9350
rect 2719 9308 2758 9342
rect 2792 9308 2831 9342
rect 2719 9300 2831 9308
rect 3269 9342 3381 9350
rect 3269 9308 3308 9342
rect 3342 9308 3381 9342
rect 3269 9300 3381 9308
rect 3819 9342 3931 9350
rect 3819 9308 3858 9342
rect 3892 9308 3931 9342
rect 3819 9300 3931 9308
rect 4369 9342 4481 9350
rect 4369 9308 4408 9342
rect 4442 9308 4481 9342
rect 4369 9300 4481 9308
rect 4919 9342 5031 9350
rect 4919 9308 4958 9342
rect 4992 9308 5031 9342
rect 4919 9300 5031 9308
rect 5469 9342 5581 9350
rect 5469 9308 5508 9342
rect 5542 9308 5581 9342
rect 5469 9300 5581 9308
rect 6019 9342 6131 9350
rect 6019 9308 6058 9342
rect 6092 9308 6131 9342
rect 6019 9300 6131 9308
rect 6569 9342 6681 9350
rect 6569 9308 6608 9342
rect 6642 9308 6681 9342
rect 6569 9300 6681 9308
rect 7119 9342 7231 9350
rect 7119 9308 7158 9342
rect 7192 9308 7231 9342
rect 7119 9300 7231 9308
rect 7669 9342 7781 9350
rect 7669 9308 7708 9342
rect 7742 9308 7781 9342
rect 7669 9300 7781 9308
rect 8219 9342 8331 9350
rect 8219 9308 8258 9342
rect 8292 9308 8331 9342
rect 8219 9300 8331 9308
rect 8769 9342 8881 9350
rect 8769 9308 8808 9342
rect 8842 9308 8881 9342
rect 8769 9300 8881 9308
rect 9319 9342 9431 9350
rect 9319 9308 9358 9342
rect 9392 9308 9431 9342
rect 9319 9300 9431 9308
rect 9869 9342 9981 9350
rect 9869 9308 9908 9342
rect 9942 9308 9981 9342
rect 9869 9300 9981 9308
rect 10419 9342 10531 9350
rect 10419 9308 10458 9342
rect 10492 9308 10531 9342
rect 10419 9300 10531 9308
rect 10969 9342 11081 9350
rect 10969 9308 11008 9342
rect 11042 9308 11081 9342
rect 10969 9300 11081 9308
rect 11519 9342 11631 9350
rect 11519 9308 11558 9342
rect 11592 9308 11631 9342
rect 11519 9300 11631 9308
rect 12069 9342 12181 9350
rect 12069 9308 12108 9342
rect 12142 9308 12181 9342
rect 12069 9300 12181 9308
rect 12619 9342 12731 9350
rect 12619 9308 12658 9342
rect 12692 9308 12731 9342
rect 12619 9300 12731 9308
rect 13169 9342 13281 9350
rect 13169 9308 13208 9342
rect 13242 9308 13281 9342
rect 13169 9300 13281 9308
rect 13719 9342 13800 9350
rect 13719 9308 13758 9342
rect 13792 9308 13800 9342
rect 13719 9300 13800 9308
rect -550 8800 -500 9300
rect 0 9269 50 9300
rect 550 9269 600 9300
rect 1100 9269 1150 9300
rect 1650 9269 1700 9300
rect 0 8800 50 8831
rect 550 8800 600 8831
rect 2200 9269 2250 9300
rect 2750 9269 2800 9300
rect 1100 8800 1150 8831
rect 1650 8800 1700 8831
rect 3300 9269 3350 9300
rect 3850 9269 3900 9300
rect 2200 8800 2250 8831
rect 2750 8800 2800 8831
rect 4400 9269 4450 9300
rect 4950 9269 5000 9300
rect 3300 8800 3350 8831
rect 3850 8800 3900 8831
rect 5500 9269 5550 9300
rect 6050 9269 6100 9300
rect 4400 8800 4450 8831
rect 4950 8800 5000 8831
rect 6600 9269 6650 9300
rect 7150 9269 7200 9300
rect 5500 8800 5550 8831
rect 6050 8800 6100 8831
rect 7700 9269 7750 9300
rect 8250 9269 8300 9300
rect 6600 8800 6650 8831
rect 7150 8800 7200 8831
rect 8800 9269 8850 9300
rect 9350 9269 9400 9300
rect 7700 8800 7750 8831
rect 8250 8800 8300 8831
rect 9900 9269 9950 9300
rect 10450 9269 10500 9300
rect 8800 8800 8850 8831
rect 9350 8800 9400 8831
rect 11000 9269 11050 9300
rect 11550 9269 11600 9300
rect 9900 8800 9950 8831
rect 10450 8800 10500 8831
rect 12100 9269 12150 9300
rect 12650 9269 12700 9300
rect 11000 8800 11050 8831
rect 11550 8800 11600 8831
rect 13200 9269 13250 9300
rect 12100 8800 12150 8831
rect 12650 8800 12700 8831
rect 13200 8800 13250 8831
rect 13750 8800 13800 9300
rect -550 8792 -469 8800
rect -550 8758 -542 8792
rect -508 8758 -469 8792
rect -550 8750 -469 8758
rect -31 8792 81 8800
rect -31 8758 8 8792
rect 42 8758 81 8792
rect -31 8750 81 8758
rect 519 8792 631 8800
rect 519 8758 558 8792
rect 592 8758 631 8792
rect 519 8750 631 8758
rect 1069 8792 1181 8800
rect 1069 8758 1108 8792
rect 1142 8758 1181 8792
rect 1069 8750 1181 8758
rect 1619 8792 1731 8800
rect 1619 8758 1658 8792
rect 1692 8758 1731 8792
rect 1619 8750 1731 8758
rect 2169 8792 2281 8800
rect 2169 8758 2208 8792
rect 2242 8758 2281 8792
rect 2169 8750 2281 8758
rect 2719 8792 2831 8800
rect 2719 8758 2758 8792
rect 2792 8758 2831 8792
rect 2719 8750 2831 8758
rect 3269 8792 3381 8800
rect 3269 8758 3308 8792
rect 3342 8758 3381 8792
rect 3269 8750 3381 8758
rect 3819 8792 3931 8800
rect 3819 8758 3858 8792
rect 3892 8758 3931 8792
rect 3819 8750 3931 8758
rect 4369 8792 4481 8800
rect 4369 8758 4408 8792
rect 4442 8758 4481 8792
rect 4369 8750 4481 8758
rect 4919 8792 5031 8800
rect 4919 8758 4958 8792
rect 4992 8758 5031 8792
rect 4919 8750 5031 8758
rect 5469 8792 5581 8800
rect 5469 8758 5508 8792
rect 5542 8758 5581 8792
rect 5469 8750 5581 8758
rect 6019 8792 6131 8800
rect 6019 8758 6058 8792
rect 6092 8758 6131 8792
rect 6019 8750 6131 8758
rect 6569 8792 6681 8800
rect 6569 8758 6608 8792
rect 6642 8758 6681 8792
rect 6569 8750 6681 8758
rect 7119 8792 7231 8800
rect 7119 8758 7158 8792
rect 7192 8758 7231 8792
rect 7119 8750 7231 8758
rect 7669 8792 7781 8800
rect 7669 8758 7708 8792
rect 7742 8758 7781 8792
rect 7669 8750 7781 8758
rect 8219 8792 8331 8800
rect 8219 8758 8258 8792
rect 8292 8758 8331 8792
rect 8219 8750 8331 8758
rect 8769 8792 8881 8800
rect 8769 8758 8808 8792
rect 8842 8758 8881 8792
rect 8769 8750 8881 8758
rect 9319 8792 9431 8800
rect 9319 8758 9358 8792
rect 9392 8758 9431 8792
rect 9319 8750 9431 8758
rect 9869 8792 9981 8800
rect 9869 8758 9908 8792
rect 9942 8758 9981 8792
rect 9869 8750 9981 8758
rect 10419 8792 10531 8800
rect 10419 8758 10458 8792
rect 10492 8758 10531 8792
rect 10419 8750 10531 8758
rect 10969 8792 11081 8800
rect 10969 8758 11008 8792
rect 11042 8758 11081 8792
rect 10969 8750 11081 8758
rect 11519 8792 11631 8800
rect 11519 8758 11558 8792
rect 11592 8758 11631 8792
rect 11519 8750 11631 8758
rect 12069 8792 12181 8800
rect 12069 8758 12108 8792
rect 12142 8758 12181 8792
rect 12069 8750 12181 8758
rect 12619 8792 12731 8800
rect 12619 8758 12658 8792
rect 12692 8758 12731 8792
rect 12619 8750 12731 8758
rect 13169 8792 13281 8800
rect 13169 8758 13208 8792
rect 13242 8758 13281 8792
rect 13169 8750 13281 8758
rect 13719 8792 13800 8800
rect 13719 8758 13758 8792
rect 13792 8758 13800 8792
rect 13719 8750 13800 8758
rect -550 8250 -500 8750
rect 0 8719 50 8750
rect 550 8719 600 8750
rect 1100 8719 1150 8750
rect 0 8250 50 8281
rect 1650 8719 1700 8750
rect 2200 8719 2250 8750
rect 550 8250 600 8281
rect 1100 8250 1150 8281
rect 2750 8719 2800 8750
rect 3300 8719 3350 8750
rect 1650 8250 1700 8281
rect 2200 8250 2250 8281
rect 3850 8719 3900 8750
rect 4400 8719 4450 8750
rect 2750 8250 2800 8281
rect 3300 8250 3350 8281
rect 4950 8719 5000 8750
rect 5500 8719 5550 8750
rect 3850 8250 3900 8281
rect 4400 8250 4450 8281
rect 6050 8719 6100 8750
rect 6600 8719 6650 8750
rect 4950 8250 5000 8281
rect 5500 8250 5550 8281
rect 7150 8719 7200 8750
rect 7700 8719 7750 8750
rect 6050 8250 6100 8281
rect 6600 8250 6650 8281
rect 8250 8719 8300 8750
rect 8800 8719 8850 8750
rect 7150 8250 7200 8281
rect 7700 8250 7750 8281
rect 9350 8719 9400 8750
rect 9900 8719 9950 8750
rect 8250 8250 8300 8281
rect 8800 8250 8850 8281
rect 10450 8719 10500 8750
rect 11000 8719 11050 8750
rect 9350 8250 9400 8281
rect 9900 8250 9950 8281
rect 11550 8719 11600 8750
rect 12100 8719 12150 8750
rect 10450 8250 10500 8281
rect 11000 8250 11050 8281
rect 12650 8719 12700 8750
rect 13200 8719 13250 8750
rect 11550 8250 11600 8281
rect 12100 8250 12150 8281
rect 12650 8250 12700 8281
rect 13200 8250 13250 8281
rect 13750 8250 13800 8750
rect -550 8242 -469 8250
rect -550 8208 -542 8242
rect -508 8208 -469 8242
rect -550 8200 -469 8208
rect -31 8242 81 8250
rect -31 8208 8 8242
rect 42 8208 81 8242
rect -31 8200 81 8208
rect 519 8242 631 8250
rect 519 8208 558 8242
rect 592 8208 631 8242
rect 519 8200 631 8208
rect 1069 8242 1181 8250
rect 1069 8208 1108 8242
rect 1142 8208 1181 8242
rect 1069 8200 1181 8208
rect 1619 8242 1731 8250
rect 1619 8208 1658 8242
rect 1692 8208 1731 8242
rect 1619 8200 1731 8208
rect 2169 8242 2281 8250
rect 2169 8208 2208 8242
rect 2242 8208 2281 8242
rect 2169 8200 2281 8208
rect 2719 8242 2831 8250
rect 2719 8208 2758 8242
rect 2792 8208 2831 8242
rect 2719 8200 2831 8208
rect 3269 8242 3381 8250
rect 3269 8208 3308 8242
rect 3342 8208 3381 8242
rect 3269 8200 3381 8208
rect 3819 8242 3931 8250
rect 3819 8208 3858 8242
rect 3892 8208 3931 8242
rect 3819 8200 3931 8208
rect 4369 8242 4481 8250
rect 4369 8208 4408 8242
rect 4442 8208 4481 8242
rect 4369 8200 4481 8208
rect 4919 8242 5031 8250
rect 4919 8208 4958 8242
rect 4992 8208 5031 8242
rect 4919 8200 5031 8208
rect 5469 8242 5581 8250
rect 5469 8208 5508 8242
rect 5542 8208 5581 8242
rect 5469 8200 5581 8208
rect 6019 8242 6131 8250
rect 6019 8208 6058 8242
rect 6092 8208 6131 8242
rect 6019 8200 6131 8208
rect 6569 8242 6681 8250
rect 6569 8208 6608 8242
rect 6642 8208 6681 8242
rect 6569 8200 6681 8208
rect 7119 8242 7231 8250
rect 7119 8208 7158 8242
rect 7192 8208 7231 8242
rect 7119 8200 7231 8208
rect 7669 8242 7781 8250
rect 7669 8208 7708 8242
rect 7742 8208 7781 8242
rect 7669 8200 7781 8208
rect 8219 8242 8331 8250
rect 8219 8208 8258 8242
rect 8292 8208 8331 8242
rect 8219 8200 8331 8208
rect 8769 8242 8881 8250
rect 8769 8208 8808 8242
rect 8842 8208 8881 8242
rect 8769 8200 8881 8208
rect 9319 8242 9431 8250
rect 9319 8208 9358 8242
rect 9392 8208 9431 8242
rect 9319 8200 9431 8208
rect 9869 8242 9981 8250
rect 9869 8208 9908 8242
rect 9942 8208 9981 8242
rect 9869 8200 9981 8208
rect 10419 8242 10531 8250
rect 10419 8208 10458 8242
rect 10492 8208 10531 8242
rect 10419 8200 10531 8208
rect 10969 8242 11081 8250
rect 10969 8208 11008 8242
rect 11042 8208 11081 8242
rect 10969 8200 11081 8208
rect 11519 8242 11631 8250
rect 11519 8208 11558 8242
rect 11592 8208 11631 8242
rect 11519 8200 11631 8208
rect 12069 8242 12181 8250
rect 12069 8208 12108 8242
rect 12142 8208 12181 8242
rect 12069 8200 12181 8208
rect 12619 8242 12731 8250
rect 12619 8208 12658 8242
rect 12692 8208 12731 8242
rect 12619 8200 12731 8208
rect 13169 8242 13281 8250
rect 13169 8208 13208 8242
rect 13242 8208 13281 8242
rect 13169 8200 13281 8208
rect 13719 8242 13800 8250
rect 13719 8208 13758 8242
rect 13792 8208 13800 8242
rect 13719 8200 13800 8208
rect -550 7700 -500 8200
rect 0 8169 50 8200
rect 550 8169 600 8200
rect 1100 8169 1150 8200
rect 1650 8169 1700 8200
rect 0 7700 50 7731
rect 550 7700 600 7731
rect 2200 8169 2250 8200
rect 2750 8169 2800 8200
rect 1100 7700 1150 7731
rect 1650 7700 1700 7731
rect 3300 8169 3350 8200
rect 3850 8169 3900 8200
rect 2200 7700 2250 7731
rect 2750 7700 2800 7731
rect 4400 8169 4450 8200
rect 4950 8169 5000 8200
rect 3300 7700 3350 7731
rect 3850 7700 3900 7731
rect 5500 8169 5550 8200
rect 6050 8169 6100 8200
rect 4400 7700 4450 7731
rect 4950 7700 5000 7731
rect 6600 8169 6650 8200
rect 7150 8169 7200 8200
rect 5500 7700 5550 7731
rect 6050 7700 6100 7731
rect 7700 8169 7750 8200
rect 8250 8169 8300 8200
rect 6600 7700 6650 7731
rect 7150 7700 7200 7731
rect 8800 8169 8850 8200
rect 9350 8169 9400 8200
rect 7700 7700 7750 7731
rect 8250 7700 8300 7731
rect 9900 8169 9950 8200
rect 10450 8169 10500 8200
rect 8800 7700 8850 7731
rect 9350 7700 9400 7731
rect 11000 8169 11050 8200
rect 11550 8169 11600 8200
rect 9900 7700 9950 7731
rect 10450 7700 10500 7731
rect 12100 8169 12150 8200
rect 12650 8169 12700 8200
rect 11000 7700 11050 7731
rect 11550 7700 11600 7731
rect 13200 8169 13250 8200
rect 12100 7700 12150 7731
rect 12650 7700 12700 7731
rect 13200 7700 13250 7731
rect 13750 7700 13800 8200
rect -550 7692 -469 7700
rect -550 7658 -542 7692
rect -508 7658 -469 7692
rect -550 7650 -469 7658
rect -31 7692 81 7700
rect -31 7658 8 7692
rect 42 7658 81 7692
rect -31 7650 81 7658
rect 519 7692 631 7700
rect 519 7658 558 7692
rect 592 7658 631 7692
rect 519 7650 631 7658
rect 1069 7692 1181 7700
rect 1069 7658 1108 7692
rect 1142 7658 1181 7692
rect 1069 7650 1181 7658
rect 1619 7692 1731 7700
rect 1619 7658 1658 7692
rect 1692 7658 1731 7692
rect 1619 7650 1731 7658
rect 2169 7692 2281 7700
rect 2169 7658 2208 7692
rect 2242 7658 2281 7692
rect 2169 7650 2281 7658
rect 2719 7692 2831 7700
rect 2719 7658 2758 7692
rect 2792 7658 2831 7692
rect 2719 7650 2831 7658
rect 3269 7692 3381 7700
rect 3269 7658 3308 7692
rect 3342 7658 3381 7692
rect 3269 7650 3381 7658
rect 3819 7692 3931 7700
rect 3819 7658 3858 7692
rect 3892 7658 3931 7692
rect 3819 7650 3931 7658
rect 4369 7692 4481 7700
rect 4369 7658 4408 7692
rect 4442 7658 4481 7692
rect 4369 7650 4481 7658
rect 4919 7692 5031 7700
rect 4919 7658 4958 7692
rect 4992 7658 5031 7692
rect 4919 7650 5031 7658
rect 5469 7692 5581 7700
rect 5469 7658 5508 7692
rect 5542 7658 5581 7692
rect 5469 7650 5581 7658
rect 6019 7692 6131 7700
rect 6019 7658 6058 7692
rect 6092 7658 6131 7692
rect 6019 7650 6131 7658
rect 6569 7692 6681 7700
rect 6569 7658 6608 7692
rect 6642 7658 6681 7692
rect 6569 7650 6681 7658
rect 7119 7692 7231 7700
rect 7119 7658 7158 7692
rect 7192 7658 7231 7692
rect 7119 7650 7231 7658
rect 7669 7692 7781 7700
rect 7669 7658 7708 7692
rect 7742 7658 7781 7692
rect 7669 7650 7781 7658
rect 8219 7692 8331 7700
rect 8219 7658 8258 7692
rect 8292 7658 8331 7692
rect 8219 7650 8331 7658
rect 8769 7692 8881 7700
rect 8769 7658 8808 7692
rect 8842 7658 8881 7692
rect 8769 7650 8881 7658
rect 9319 7692 9431 7700
rect 9319 7658 9358 7692
rect 9392 7658 9431 7692
rect 9319 7650 9431 7658
rect 9869 7692 9981 7700
rect 9869 7658 9908 7692
rect 9942 7658 9981 7692
rect 9869 7650 9981 7658
rect 10419 7692 10531 7700
rect 10419 7658 10458 7692
rect 10492 7658 10531 7692
rect 10419 7650 10531 7658
rect 10969 7692 11081 7700
rect 10969 7658 11008 7692
rect 11042 7658 11081 7692
rect 10969 7650 11081 7658
rect 11519 7692 11631 7700
rect 11519 7658 11558 7692
rect 11592 7658 11631 7692
rect 11519 7650 11631 7658
rect 12069 7692 12181 7700
rect 12069 7658 12108 7692
rect 12142 7658 12181 7692
rect 12069 7650 12181 7658
rect 12619 7692 12731 7700
rect 12619 7658 12658 7692
rect 12692 7658 12731 7692
rect 12619 7650 12731 7658
rect 13169 7692 13281 7700
rect 13169 7658 13208 7692
rect 13242 7658 13281 7692
rect 13169 7650 13281 7658
rect 13719 7692 13800 7700
rect 13719 7658 13758 7692
rect 13792 7658 13800 7692
rect 13719 7650 13800 7658
rect -550 7150 -500 7650
rect 0 7619 50 7650
rect 550 7619 600 7650
rect 1100 7619 1150 7650
rect 0 7150 50 7181
rect 1650 7619 1700 7650
rect 2200 7619 2250 7650
rect 550 7150 600 7181
rect 1100 7150 1150 7181
rect 2750 7619 2800 7650
rect 3300 7619 3350 7650
rect 1650 7150 1700 7181
rect 2200 7150 2250 7181
rect 3850 7619 3900 7650
rect 4400 7619 4450 7650
rect 2750 7150 2800 7181
rect 3300 7150 3350 7181
rect 4950 7619 5000 7650
rect 5500 7619 5550 7650
rect 3850 7150 3900 7181
rect 4400 7150 4450 7181
rect 6050 7619 6100 7650
rect 6600 7619 6650 7650
rect 4950 7150 5000 7181
rect 5500 7150 5550 7181
rect 7150 7619 7200 7650
rect 7700 7619 7750 7650
rect 6050 7150 6100 7181
rect 6600 7150 6650 7181
rect 8250 7619 8300 7650
rect 8800 7619 8850 7650
rect 7150 7150 7200 7181
rect 7700 7150 7750 7181
rect 9350 7619 9400 7650
rect 9900 7619 9950 7650
rect 8250 7150 8300 7181
rect 8800 7150 8850 7181
rect 10450 7619 10500 7650
rect 11000 7619 11050 7650
rect 9350 7150 9400 7181
rect 9900 7150 9950 7181
rect 11550 7619 11600 7650
rect 12100 7619 12150 7650
rect 10450 7150 10500 7181
rect 11000 7150 11050 7181
rect 12650 7619 12700 7650
rect 13200 7619 13250 7650
rect 11550 7150 11600 7181
rect 12100 7150 12150 7181
rect 12650 7150 12700 7181
rect 13200 7150 13250 7181
rect 13750 7150 13800 7650
rect -550 7142 -469 7150
rect -550 7108 -542 7142
rect -508 7108 -469 7142
rect -550 7100 -469 7108
rect -31 7142 81 7150
rect -31 7108 8 7142
rect 42 7108 81 7142
rect -31 7100 81 7108
rect 519 7142 631 7150
rect 519 7108 558 7142
rect 592 7108 631 7142
rect 519 7100 631 7108
rect 1069 7142 1181 7150
rect 1069 7108 1108 7142
rect 1142 7108 1181 7142
rect 1069 7100 1181 7108
rect 1619 7142 1731 7150
rect 1619 7108 1658 7142
rect 1692 7108 1731 7142
rect 1619 7100 1731 7108
rect 2169 7142 2281 7150
rect 2169 7108 2208 7142
rect 2242 7108 2281 7142
rect 2169 7100 2281 7108
rect 2719 7142 2831 7150
rect 2719 7108 2758 7142
rect 2792 7108 2831 7142
rect 2719 7100 2831 7108
rect 3269 7142 3381 7150
rect 3269 7108 3308 7142
rect 3342 7108 3381 7142
rect 3269 7100 3381 7108
rect 3819 7142 3931 7150
rect 3819 7108 3858 7142
rect 3892 7108 3931 7142
rect 3819 7100 3931 7108
rect 4369 7142 4481 7150
rect 4369 7108 4408 7142
rect 4442 7108 4481 7142
rect 4369 7100 4481 7108
rect 4919 7142 5031 7150
rect 4919 7108 4958 7142
rect 4992 7108 5031 7142
rect 4919 7100 5031 7108
rect 5469 7142 5581 7150
rect 5469 7108 5508 7142
rect 5542 7108 5581 7142
rect 5469 7100 5581 7108
rect 6019 7142 6131 7150
rect 6019 7108 6058 7142
rect 6092 7108 6131 7142
rect 6019 7100 6131 7108
rect 6569 7142 6681 7150
rect 6569 7108 6608 7142
rect 6642 7108 6681 7142
rect 6569 7100 6681 7108
rect 7119 7142 7231 7150
rect 7119 7108 7158 7142
rect 7192 7108 7231 7142
rect 7119 7100 7231 7108
rect 7669 7142 7781 7150
rect 7669 7108 7708 7142
rect 7742 7108 7781 7142
rect 7669 7100 7781 7108
rect 8219 7142 8331 7150
rect 8219 7108 8258 7142
rect 8292 7108 8331 7142
rect 8219 7100 8331 7108
rect 8769 7142 8881 7150
rect 8769 7108 8808 7142
rect 8842 7108 8881 7142
rect 8769 7100 8881 7108
rect 9319 7142 9431 7150
rect 9319 7108 9358 7142
rect 9392 7108 9431 7142
rect 9319 7100 9431 7108
rect 9869 7142 9981 7150
rect 9869 7108 9908 7142
rect 9942 7108 9981 7142
rect 9869 7100 9981 7108
rect 10419 7142 10531 7150
rect 10419 7108 10458 7142
rect 10492 7108 10531 7142
rect 10419 7100 10531 7108
rect 10969 7142 11081 7150
rect 10969 7108 11008 7142
rect 11042 7108 11081 7142
rect 10969 7100 11081 7108
rect 11519 7142 11631 7150
rect 11519 7108 11558 7142
rect 11592 7108 11631 7142
rect 11519 7100 11631 7108
rect 12069 7142 12181 7150
rect 12069 7108 12108 7142
rect 12142 7108 12181 7142
rect 12069 7100 12181 7108
rect 12619 7142 12731 7150
rect 12619 7108 12658 7142
rect 12692 7108 12731 7142
rect 12619 7100 12731 7108
rect 13169 7142 13281 7150
rect 13169 7108 13208 7142
rect 13242 7108 13281 7142
rect 13169 7100 13281 7108
rect 13719 7142 13800 7150
rect 13719 7108 13758 7142
rect 13792 7108 13800 7142
rect 13719 7100 13800 7108
rect -550 6600 -500 7100
rect 0 7069 50 7100
rect 550 7069 600 7100
rect 1100 7069 1150 7100
rect 1650 7069 1700 7100
rect 0 6600 50 6631
rect 550 6600 600 6631
rect 2200 7069 2250 7100
rect 2750 7069 2800 7100
rect 1100 6600 1150 6631
rect 1650 6600 1700 6631
rect 3300 7069 3350 7100
rect 3850 7069 3900 7100
rect 2200 6600 2250 6631
rect 2750 6600 2800 6631
rect 4400 7069 4450 7100
rect 4950 7069 5000 7100
rect 3300 6600 3350 6631
rect 3850 6600 3900 6631
rect 5500 7069 5550 7100
rect 6050 7069 6100 7100
rect 4400 6600 4450 6631
rect 4950 6600 5000 6631
rect 6600 7069 6650 7100
rect 7150 7069 7200 7100
rect 5500 6600 5550 6631
rect 6050 6600 6100 6631
rect 7700 7069 7750 7100
rect 8250 7069 8300 7100
rect 6600 6600 6650 6631
rect 7150 6600 7200 6631
rect 8800 7069 8850 7100
rect 9350 7069 9400 7100
rect 7700 6600 7750 6631
rect 8250 6600 8300 6631
rect 9900 7069 9950 7100
rect 10450 7069 10500 7100
rect 8800 6600 8850 6631
rect 9350 6600 9400 6631
rect 11000 7069 11050 7100
rect 11550 7069 11600 7100
rect 9900 6600 9950 6631
rect 10450 6600 10500 6631
rect 12100 7069 12150 7100
rect 12650 7069 12700 7100
rect 11000 6600 11050 6631
rect 11550 6600 11600 6631
rect 13200 7069 13250 7100
rect 12100 6600 12150 6631
rect 12650 6600 12700 6631
rect 13200 6600 13250 6631
rect 13750 6600 13800 7100
rect -550 6592 -469 6600
rect -550 6558 -542 6592
rect -508 6558 -469 6592
rect -550 6550 -469 6558
rect -31 6592 81 6600
rect -31 6558 8 6592
rect 42 6558 81 6592
rect -31 6550 81 6558
rect 519 6592 631 6600
rect 519 6558 558 6592
rect 592 6558 631 6592
rect 519 6550 631 6558
rect 1069 6592 1181 6600
rect 1069 6558 1108 6592
rect 1142 6558 1181 6592
rect 1069 6550 1181 6558
rect 1619 6592 1731 6600
rect 1619 6558 1658 6592
rect 1692 6558 1731 6592
rect 1619 6550 1731 6558
rect 2169 6592 2281 6600
rect 2169 6558 2208 6592
rect 2242 6558 2281 6592
rect 2169 6550 2281 6558
rect 2719 6592 2831 6600
rect 2719 6558 2758 6592
rect 2792 6558 2831 6592
rect 2719 6550 2831 6558
rect 3269 6592 3381 6600
rect 3269 6558 3308 6592
rect 3342 6558 3381 6592
rect 3269 6550 3381 6558
rect 3819 6592 3931 6600
rect 3819 6558 3858 6592
rect 3892 6558 3931 6592
rect 3819 6550 3931 6558
rect 4369 6592 4481 6600
rect 4369 6558 4408 6592
rect 4442 6558 4481 6592
rect 4369 6550 4481 6558
rect 4919 6592 5031 6600
rect 4919 6558 4958 6592
rect 4992 6558 5031 6592
rect 4919 6550 5031 6558
rect 5469 6592 5581 6600
rect 5469 6558 5508 6592
rect 5542 6558 5581 6592
rect 5469 6550 5581 6558
rect 6019 6592 6131 6600
rect 6019 6558 6058 6592
rect 6092 6558 6131 6592
rect 6019 6550 6131 6558
rect 6569 6592 6681 6600
rect 6569 6558 6608 6592
rect 6642 6558 6681 6592
rect 6569 6550 6681 6558
rect 7119 6592 7231 6600
rect 7119 6558 7158 6592
rect 7192 6558 7231 6592
rect 7119 6550 7231 6558
rect 7669 6592 7781 6600
rect 7669 6558 7708 6592
rect 7742 6558 7781 6592
rect 7669 6550 7781 6558
rect 8219 6592 8331 6600
rect 8219 6558 8258 6592
rect 8292 6558 8331 6592
rect 8219 6550 8331 6558
rect 8769 6592 8881 6600
rect 8769 6558 8808 6592
rect 8842 6558 8881 6592
rect 8769 6550 8881 6558
rect 9319 6592 9431 6600
rect 9319 6558 9358 6592
rect 9392 6558 9431 6592
rect 9319 6550 9431 6558
rect 9869 6592 9981 6600
rect 9869 6558 9908 6592
rect 9942 6558 9981 6592
rect 9869 6550 9981 6558
rect 10419 6592 10531 6600
rect 10419 6558 10458 6592
rect 10492 6558 10531 6592
rect 10419 6550 10531 6558
rect 10969 6592 11081 6600
rect 10969 6558 11008 6592
rect 11042 6558 11081 6592
rect 10969 6550 11081 6558
rect 11519 6592 11631 6600
rect 11519 6558 11558 6592
rect 11592 6558 11631 6592
rect 11519 6550 11631 6558
rect 12069 6592 12181 6600
rect 12069 6558 12108 6592
rect 12142 6558 12181 6592
rect 12069 6550 12181 6558
rect 12619 6592 12731 6600
rect 12619 6558 12658 6592
rect 12692 6558 12731 6592
rect 12619 6550 12731 6558
rect 13169 6592 13281 6600
rect 13169 6558 13208 6592
rect 13242 6558 13281 6592
rect 13169 6550 13281 6558
rect 13719 6592 13800 6600
rect 13719 6558 13758 6592
rect 13792 6558 13800 6592
rect 13719 6550 13800 6558
rect -550 6050 -500 6550
rect 0 6519 50 6550
rect 550 6519 600 6550
rect 1100 6519 1150 6550
rect 0 6050 50 6081
rect 1650 6519 1700 6550
rect 2200 6519 2250 6550
rect 550 6050 600 6081
rect 1100 6050 1150 6081
rect 2750 6519 2800 6550
rect 3300 6519 3350 6550
rect 1650 6050 1700 6081
rect 2200 6050 2250 6081
rect 3850 6519 3900 6550
rect 4400 6519 4450 6550
rect 2750 6050 2800 6081
rect 3300 6050 3350 6081
rect 4950 6519 5000 6550
rect 5500 6519 5550 6550
rect 3850 6050 3900 6081
rect 4400 6050 4450 6081
rect 6050 6519 6100 6550
rect 6600 6519 6650 6550
rect 4950 6050 5000 6081
rect 5500 6050 5550 6081
rect 7150 6519 7200 6550
rect 7700 6519 7750 6550
rect 6050 6050 6100 6081
rect 6600 6050 6650 6081
rect 8250 6519 8300 6550
rect 8800 6519 8850 6550
rect 7150 6050 7200 6081
rect 7700 6050 7750 6081
rect 9350 6519 9400 6550
rect 9900 6519 9950 6550
rect 8250 6050 8300 6081
rect 8800 6050 8850 6081
rect 10450 6519 10500 6550
rect 11000 6519 11050 6550
rect 9350 6050 9400 6081
rect 9900 6050 9950 6081
rect 11550 6519 11600 6550
rect 12100 6519 12150 6550
rect 10450 6050 10500 6081
rect 11000 6050 11050 6081
rect 12650 6519 12700 6550
rect 13200 6519 13250 6550
rect 11550 6050 11600 6081
rect 12100 6050 12150 6081
rect 12650 6050 12700 6081
rect 13200 6050 13250 6081
rect 13750 6050 13800 6550
rect -550 6042 -469 6050
rect -550 6008 -542 6042
rect -508 6008 -469 6042
rect -550 6000 -469 6008
rect -31 6042 81 6050
rect -31 6008 8 6042
rect 42 6008 81 6042
rect -31 6000 81 6008
rect 519 6042 631 6050
rect 519 6008 558 6042
rect 592 6008 631 6042
rect 519 6000 631 6008
rect 1069 6042 1181 6050
rect 1069 6008 1108 6042
rect 1142 6008 1181 6042
rect 1069 6000 1181 6008
rect 1619 6042 1731 6050
rect 1619 6008 1658 6042
rect 1692 6008 1731 6042
rect 1619 6000 1731 6008
rect 2169 6042 2281 6050
rect 2169 6008 2208 6042
rect 2242 6008 2281 6042
rect 2169 6000 2281 6008
rect 2719 6042 2831 6050
rect 2719 6008 2758 6042
rect 2792 6008 2831 6042
rect 2719 6000 2831 6008
rect 3269 6042 3381 6050
rect 3269 6008 3308 6042
rect 3342 6008 3381 6042
rect 3269 6000 3381 6008
rect 3819 6042 3931 6050
rect 3819 6008 3858 6042
rect 3892 6008 3931 6042
rect 3819 6000 3931 6008
rect 4369 6042 4481 6050
rect 4369 6008 4408 6042
rect 4442 6008 4481 6042
rect 4369 6000 4481 6008
rect 4919 6042 5031 6050
rect 4919 6008 4958 6042
rect 4992 6008 5031 6042
rect 4919 6000 5031 6008
rect 5469 6042 5581 6050
rect 5469 6008 5508 6042
rect 5542 6008 5581 6042
rect 5469 6000 5581 6008
rect 6019 6042 6131 6050
rect 6019 6008 6058 6042
rect 6092 6008 6131 6042
rect 6019 6000 6131 6008
rect 6569 6042 6681 6050
rect 6569 6008 6608 6042
rect 6642 6008 6681 6042
rect 6569 6000 6681 6008
rect 7119 6042 7231 6050
rect 7119 6008 7158 6042
rect 7192 6008 7231 6042
rect 7119 6000 7231 6008
rect 7669 6042 7781 6050
rect 7669 6008 7708 6042
rect 7742 6008 7781 6042
rect 7669 6000 7781 6008
rect 8219 6042 8331 6050
rect 8219 6008 8258 6042
rect 8292 6008 8331 6042
rect 8219 6000 8331 6008
rect 8769 6042 8881 6050
rect 8769 6008 8808 6042
rect 8842 6008 8881 6042
rect 8769 6000 8881 6008
rect 9319 6042 9431 6050
rect 9319 6008 9358 6042
rect 9392 6008 9431 6042
rect 9319 6000 9431 6008
rect 9869 6042 9981 6050
rect 9869 6008 9908 6042
rect 9942 6008 9981 6042
rect 9869 6000 9981 6008
rect 10419 6042 10531 6050
rect 10419 6008 10458 6042
rect 10492 6008 10531 6042
rect 10419 6000 10531 6008
rect 10969 6042 11081 6050
rect 10969 6008 11008 6042
rect 11042 6008 11081 6042
rect 10969 6000 11081 6008
rect 11519 6042 11631 6050
rect 11519 6008 11558 6042
rect 11592 6008 11631 6042
rect 11519 6000 11631 6008
rect 12069 6042 12181 6050
rect 12069 6008 12108 6042
rect 12142 6008 12181 6042
rect 12069 6000 12181 6008
rect 12619 6042 12731 6050
rect 12619 6008 12658 6042
rect 12692 6008 12731 6042
rect 12619 6000 12731 6008
rect 13169 6042 13281 6050
rect 13169 6008 13208 6042
rect 13242 6008 13281 6042
rect 13169 6000 13281 6008
rect 13719 6042 13800 6050
rect 13719 6008 13758 6042
rect 13792 6008 13800 6042
rect 13719 6000 13800 6008
rect -550 5500 -500 6000
rect 0 5969 50 6000
rect 550 5969 600 6000
rect 1100 5969 1150 6000
rect 1650 5969 1700 6000
rect 0 5500 50 5531
rect 550 5500 600 5531
rect 2200 5969 2250 6000
rect 2750 5969 2800 6000
rect 1100 5500 1150 5531
rect 1650 5500 1700 5531
rect 3300 5969 3350 6000
rect 3850 5969 3900 6000
rect 2200 5500 2250 5531
rect 2750 5500 2800 5531
rect 4400 5969 4450 6000
rect 4950 5969 5000 6000
rect 3300 5500 3350 5531
rect 3850 5500 3900 5531
rect 5500 5969 5550 6000
rect 6050 5969 6100 6000
rect 4400 5500 4450 5531
rect 4950 5500 5000 5531
rect 6600 5969 6650 6000
rect 7150 5969 7200 6000
rect 5500 5500 5550 5531
rect 6050 5500 6100 5531
rect 7700 5969 7750 6000
rect 8250 5969 8300 6000
rect 6600 5500 6650 5531
rect 7150 5500 7200 5531
rect 8800 5969 8850 6000
rect 9350 5969 9400 6000
rect 7700 5500 7750 5531
rect 8250 5500 8300 5531
rect 9900 5969 9950 6000
rect 10450 5969 10500 6000
rect 8800 5500 8850 5531
rect 9350 5500 9400 5531
rect 11000 5969 11050 6000
rect 11550 5969 11600 6000
rect 9900 5500 9950 5531
rect 10450 5500 10500 5531
rect 12100 5969 12150 6000
rect 12650 5969 12700 6000
rect 11000 5500 11050 5531
rect 11550 5500 11600 5531
rect 13200 5969 13250 6000
rect 12100 5500 12150 5531
rect 12650 5500 12700 5531
rect 13200 5500 13250 5531
rect 13750 5500 13800 6000
rect -550 5492 -469 5500
rect -550 5458 -542 5492
rect -508 5458 -469 5492
rect -550 5450 -469 5458
rect -31 5492 81 5500
rect -31 5458 8 5492
rect 42 5458 81 5492
rect -31 5450 81 5458
rect 519 5492 631 5500
rect 519 5458 558 5492
rect 592 5458 631 5492
rect 519 5450 631 5458
rect 1069 5492 1181 5500
rect 1069 5458 1108 5492
rect 1142 5458 1181 5492
rect 1069 5450 1181 5458
rect 1619 5492 1731 5500
rect 1619 5458 1658 5492
rect 1692 5458 1731 5492
rect 1619 5450 1731 5458
rect 2169 5492 2281 5500
rect 2169 5458 2208 5492
rect 2242 5458 2281 5492
rect 2169 5450 2281 5458
rect 2719 5492 2831 5500
rect 2719 5458 2758 5492
rect 2792 5458 2831 5492
rect 2719 5450 2831 5458
rect 3269 5492 3381 5500
rect 3269 5458 3308 5492
rect 3342 5458 3381 5492
rect 3269 5450 3381 5458
rect 3819 5492 3931 5500
rect 3819 5458 3858 5492
rect 3892 5458 3931 5492
rect 3819 5450 3931 5458
rect 4369 5492 4481 5500
rect 4369 5458 4408 5492
rect 4442 5458 4481 5492
rect 4369 5450 4481 5458
rect 4919 5492 5031 5500
rect 4919 5458 4958 5492
rect 4992 5458 5031 5492
rect 4919 5450 5031 5458
rect 5469 5492 5581 5500
rect 5469 5458 5508 5492
rect 5542 5458 5581 5492
rect 5469 5450 5581 5458
rect 6019 5492 6131 5500
rect 6019 5458 6058 5492
rect 6092 5458 6131 5492
rect 6019 5450 6131 5458
rect 6569 5492 6681 5500
rect 6569 5458 6608 5492
rect 6642 5458 6681 5492
rect 6569 5450 6681 5458
rect 7119 5492 7231 5500
rect 7119 5458 7158 5492
rect 7192 5458 7231 5492
rect 7119 5450 7231 5458
rect 7669 5492 7781 5500
rect 7669 5458 7708 5492
rect 7742 5458 7781 5492
rect 7669 5450 7781 5458
rect 8219 5492 8331 5500
rect 8219 5458 8258 5492
rect 8292 5458 8331 5492
rect 8219 5450 8331 5458
rect 8769 5492 8881 5500
rect 8769 5458 8808 5492
rect 8842 5458 8881 5492
rect 8769 5450 8881 5458
rect 9319 5492 9431 5500
rect 9319 5458 9358 5492
rect 9392 5458 9431 5492
rect 9319 5450 9431 5458
rect 9869 5492 9981 5500
rect 9869 5458 9908 5492
rect 9942 5458 9981 5492
rect 9869 5450 9981 5458
rect 10419 5492 10531 5500
rect 10419 5458 10458 5492
rect 10492 5458 10531 5492
rect 10419 5450 10531 5458
rect 10969 5492 11081 5500
rect 10969 5458 11008 5492
rect 11042 5458 11081 5492
rect 10969 5450 11081 5458
rect 11519 5492 11631 5500
rect 11519 5458 11558 5492
rect 11592 5458 11631 5492
rect 11519 5450 11631 5458
rect 12069 5492 12181 5500
rect 12069 5458 12108 5492
rect 12142 5458 12181 5492
rect 12069 5450 12181 5458
rect 12619 5492 12731 5500
rect 12619 5458 12658 5492
rect 12692 5458 12731 5492
rect 12619 5450 12731 5458
rect 13169 5492 13281 5500
rect 13169 5458 13208 5492
rect 13242 5458 13281 5492
rect 13169 5450 13281 5458
rect 13719 5492 13800 5500
rect 13719 5458 13758 5492
rect 13792 5458 13800 5492
rect 13719 5450 13800 5458
rect -550 4950 -500 5450
rect 0 5419 50 5450
rect 550 5419 600 5450
rect 1100 5419 1150 5450
rect 0 4950 50 4981
rect 1650 5419 1700 5450
rect 2200 5419 2250 5450
rect 550 4950 600 4981
rect 1100 4950 1150 4981
rect 2750 5419 2800 5450
rect 3300 5419 3350 5450
rect 1650 4950 1700 4981
rect 2200 4950 2250 4981
rect 3850 5419 3900 5450
rect 4400 5419 4450 5450
rect 2750 4950 2800 4981
rect 3300 4950 3350 4981
rect 4950 5419 5000 5450
rect 5500 5419 5550 5450
rect 3850 4950 3900 4981
rect 4400 4950 4450 4981
rect 6050 5419 6100 5450
rect 6600 5419 6650 5450
rect 4950 4950 5000 4981
rect 5500 4950 5550 4981
rect 7150 5419 7200 5450
rect 7700 5419 7750 5450
rect 6050 4950 6100 4981
rect 6600 4950 6650 4981
rect 8250 5419 8300 5450
rect 8800 5419 8850 5450
rect 7150 4950 7200 4981
rect 7700 4950 7750 4981
rect 9350 5419 9400 5450
rect 9900 5419 9950 5450
rect 8250 4950 8300 4981
rect 8800 4950 8850 4981
rect 10450 5419 10500 5450
rect 11000 5419 11050 5450
rect 9350 4950 9400 4981
rect 9900 4950 9950 4981
rect 11550 5419 11600 5450
rect 12100 5419 12150 5450
rect 10450 4950 10500 4981
rect 11000 4950 11050 4981
rect 12650 5419 12700 5450
rect 13200 5419 13250 5450
rect 11550 4950 11600 4981
rect 12100 4950 12150 4981
rect 12650 4950 12700 4981
rect 13200 4950 13250 4981
rect 13750 4950 13800 5450
rect -550 4942 -469 4950
rect -550 4908 -542 4942
rect -508 4908 -469 4942
rect -550 4900 -469 4908
rect -31 4942 81 4950
rect -31 4908 8 4942
rect 42 4908 81 4942
rect -31 4900 81 4908
rect 519 4942 631 4950
rect 519 4908 558 4942
rect 592 4908 631 4942
rect 519 4900 631 4908
rect 1069 4942 1181 4950
rect 1069 4908 1108 4942
rect 1142 4908 1181 4942
rect 1069 4900 1181 4908
rect 1619 4942 1731 4950
rect 1619 4908 1658 4942
rect 1692 4908 1731 4942
rect 1619 4900 1731 4908
rect 2169 4942 2281 4950
rect 2169 4908 2208 4942
rect 2242 4908 2281 4942
rect 2169 4900 2281 4908
rect 2719 4942 2831 4950
rect 2719 4908 2758 4942
rect 2792 4908 2831 4942
rect 2719 4900 2831 4908
rect 3269 4942 3381 4950
rect 3269 4908 3308 4942
rect 3342 4908 3381 4942
rect 3269 4900 3381 4908
rect 3819 4942 3931 4950
rect 3819 4908 3858 4942
rect 3892 4908 3931 4942
rect 3819 4900 3931 4908
rect 4369 4942 4481 4950
rect 4369 4908 4408 4942
rect 4442 4908 4481 4942
rect 4369 4900 4481 4908
rect 4919 4942 5031 4950
rect 4919 4908 4958 4942
rect 4992 4908 5031 4942
rect 4919 4900 5031 4908
rect 5469 4942 5581 4950
rect 5469 4908 5508 4942
rect 5542 4908 5581 4942
rect 5469 4900 5581 4908
rect 6019 4942 6131 4950
rect 6019 4908 6058 4942
rect 6092 4908 6131 4942
rect 6019 4900 6131 4908
rect 6569 4942 6681 4950
rect 6569 4908 6608 4942
rect 6642 4908 6681 4942
rect 6569 4900 6681 4908
rect 7119 4942 7231 4950
rect 7119 4908 7158 4942
rect 7192 4908 7231 4942
rect 7119 4900 7231 4908
rect 7669 4942 7781 4950
rect 7669 4908 7708 4942
rect 7742 4908 7781 4942
rect 7669 4900 7781 4908
rect 8219 4942 8331 4950
rect 8219 4908 8258 4942
rect 8292 4908 8331 4942
rect 8219 4900 8331 4908
rect 8769 4942 8881 4950
rect 8769 4908 8808 4942
rect 8842 4908 8881 4942
rect 8769 4900 8881 4908
rect 9319 4942 9431 4950
rect 9319 4908 9358 4942
rect 9392 4908 9431 4942
rect 9319 4900 9431 4908
rect 9869 4942 9981 4950
rect 9869 4908 9908 4942
rect 9942 4908 9981 4942
rect 9869 4900 9981 4908
rect 10419 4942 10531 4950
rect 10419 4908 10458 4942
rect 10492 4908 10531 4942
rect 10419 4900 10531 4908
rect 10969 4942 11081 4950
rect 10969 4908 11008 4942
rect 11042 4908 11081 4942
rect 10969 4900 11081 4908
rect 11519 4942 11631 4950
rect 11519 4908 11558 4942
rect 11592 4908 11631 4942
rect 11519 4900 11631 4908
rect 12069 4942 12181 4950
rect 12069 4908 12108 4942
rect 12142 4908 12181 4942
rect 12069 4900 12181 4908
rect 12619 4942 12731 4950
rect 12619 4908 12658 4942
rect 12692 4908 12731 4942
rect 12619 4900 12731 4908
rect 13169 4942 13281 4950
rect 13169 4908 13208 4942
rect 13242 4908 13281 4942
rect 13169 4900 13281 4908
rect 13719 4942 13800 4950
rect 13719 4908 13758 4942
rect 13792 4908 13800 4942
rect 13719 4900 13800 4908
rect -550 4400 -500 4900
rect 0 4869 50 4900
rect 550 4869 600 4900
rect 1100 4869 1150 4900
rect 1650 4869 1700 4900
rect 0 4400 50 4431
rect 550 4400 600 4431
rect 2200 4869 2250 4900
rect 2750 4869 2800 4900
rect 1100 4400 1150 4431
rect 1650 4400 1700 4431
rect 3300 4869 3350 4900
rect 3850 4869 3900 4900
rect 2200 4400 2250 4431
rect 2750 4400 2800 4431
rect 4400 4869 4450 4900
rect 4950 4869 5000 4900
rect 3300 4400 3350 4431
rect 3850 4400 3900 4431
rect 5500 4869 5550 4900
rect 6050 4869 6100 4900
rect 4400 4400 4450 4431
rect 4950 4400 5000 4431
rect 6600 4869 6650 4900
rect 7150 4869 7200 4900
rect 5500 4400 5550 4431
rect 6050 4400 6100 4431
rect 7700 4869 7750 4900
rect 8250 4869 8300 4900
rect 6600 4400 6650 4431
rect 7150 4400 7200 4431
rect 8800 4869 8850 4900
rect 9350 4869 9400 4900
rect 7700 4400 7750 4431
rect 8250 4400 8300 4431
rect 9900 4869 9950 4900
rect 10450 4869 10500 4900
rect 8800 4400 8850 4431
rect 9350 4400 9400 4431
rect 11000 4869 11050 4900
rect 11550 4869 11600 4900
rect 9900 4400 9950 4431
rect 10450 4400 10500 4431
rect 12100 4869 12150 4900
rect 12650 4869 12700 4900
rect 11000 4400 11050 4431
rect 11550 4400 11600 4431
rect 13200 4869 13250 4900
rect 12100 4400 12150 4431
rect 12650 4400 12700 4431
rect 13200 4400 13250 4431
rect 13750 4400 13800 4900
rect -550 4392 -469 4400
rect -550 4358 -542 4392
rect -508 4358 -469 4392
rect -550 4350 -469 4358
rect -31 4392 81 4400
rect -31 4358 8 4392
rect 42 4358 81 4392
rect -31 4350 81 4358
rect 519 4392 631 4400
rect 519 4358 558 4392
rect 592 4358 631 4392
rect 519 4350 631 4358
rect 1069 4392 1181 4400
rect 1069 4358 1108 4392
rect 1142 4358 1181 4392
rect 1069 4350 1181 4358
rect 1619 4392 1731 4400
rect 1619 4358 1658 4392
rect 1692 4358 1731 4392
rect 1619 4350 1731 4358
rect 2169 4392 2281 4400
rect 2169 4358 2208 4392
rect 2242 4358 2281 4392
rect 2169 4350 2281 4358
rect 2719 4392 2831 4400
rect 2719 4358 2758 4392
rect 2792 4358 2831 4392
rect 2719 4350 2831 4358
rect 3269 4392 3381 4400
rect 3269 4358 3308 4392
rect 3342 4358 3381 4392
rect 3269 4350 3381 4358
rect 3819 4392 3931 4400
rect 3819 4358 3858 4392
rect 3892 4358 3931 4392
rect 3819 4350 3931 4358
rect 4369 4392 4481 4400
rect 4369 4358 4408 4392
rect 4442 4358 4481 4392
rect 4369 4350 4481 4358
rect 4919 4392 5031 4400
rect 4919 4358 4958 4392
rect 4992 4358 5031 4392
rect 4919 4350 5031 4358
rect 5469 4392 5581 4400
rect 5469 4358 5508 4392
rect 5542 4358 5581 4392
rect 5469 4350 5581 4358
rect 6019 4392 6131 4400
rect 6019 4358 6058 4392
rect 6092 4358 6131 4392
rect 6019 4350 6131 4358
rect 6569 4392 6681 4400
rect 6569 4358 6608 4392
rect 6642 4358 6681 4392
rect 6569 4350 6681 4358
rect 7119 4392 7231 4400
rect 7119 4358 7158 4392
rect 7192 4358 7231 4392
rect 7119 4350 7231 4358
rect 7669 4392 7781 4400
rect 7669 4358 7708 4392
rect 7742 4358 7781 4392
rect 7669 4350 7781 4358
rect 8219 4392 8331 4400
rect 8219 4358 8258 4392
rect 8292 4358 8331 4392
rect 8219 4350 8331 4358
rect 8769 4392 8881 4400
rect 8769 4358 8808 4392
rect 8842 4358 8881 4392
rect 8769 4350 8881 4358
rect 9319 4392 9431 4400
rect 9319 4358 9358 4392
rect 9392 4358 9431 4392
rect 9319 4350 9431 4358
rect 9869 4392 9981 4400
rect 9869 4358 9908 4392
rect 9942 4358 9981 4392
rect 9869 4350 9981 4358
rect 10419 4392 10531 4400
rect 10419 4358 10458 4392
rect 10492 4358 10531 4392
rect 10419 4350 10531 4358
rect 10969 4392 11081 4400
rect 10969 4358 11008 4392
rect 11042 4358 11081 4392
rect 10969 4350 11081 4358
rect 11519 4392 11631 4400
rect 11519 4358 11558 4392
rect 11592 4358 11631 4392
rect 11519 4350 11631 4358
rect 12069 4392 12181 4400
rect 12069 4358 12108 4392
rect 12142 4358 12181 4392
rect 12069 4350 12181 4358
rect 12619 4392 12731 4400
rect 12619 4358 12658 4392
rect 12692 4358 12731 4392
rect 12619 4350 12731 4358
rect 13169 4392 13281 4400
rect 13169 4358 13208 4392
rect 13242 4358 13281 4392
rect 13169 4350 13281 4358
rect 13719 4392 13800 4400
rect 13719 4358 13758 4392
rect 13792 4358 13800 4392
rect 13719 4350 13800 4358
rect -550 3850 -500 4350
rect 0 4319 50 4350
rect 550 4319 600 4350
rect 1100 4319 1150 4350
rect 0 3850 50 3881
rect 1650 4319 1700 4350
rect 2200 4319 2250 4350
rect 550 3850 600 3881
rect 1100 3850 1150 3881
rect 2750 4319 2800 4350
rect 3300 4319 3350 4350
rect 1650 3850 1700 3881
rect 2200 3850 2250 3881
rect 3850 4319 3900 4350
rect 4400 4319 4450 4350
rect 2750 3850 2800 3881
rect 3300 3850 3350 3881
rect 4950 4319 5000 4350
rect 5500 4319 5550 4350
rect 3850 3850 3900 3881
rect 4400 3850 4450 3881
rect 6050 4319 6100 4350
rect 6600 4319 6650 4350
rect 4950 3850 5000 3881
rect 5500 3850 5550 3881
rect 7150 4319 7200 4350
rect 7700 4319 7750 4350
rect 6050 3850 6100 3881
rect 6600 3850 6650 3881
rect 8250 4319 8300 4350
rect 8800 4319 8850 4350
rect 7150 3850 7200 3881
rect 7700 3850 7750 3881
rect 9350 4319 9400 4350
rect 9900 4319 9950 4350
rect 8250 3850 8300 3881
rect 8800 3850 8850 3881
rect 10450 4319 10500 4350
rect 11000 4319 11050 4350
rect 9350 3850 9400 3881
rect 9900 3850 9950 3881
rect 11550 4319 11600 4350
rect 12100 4319 12150 4350
rect 10450 3850 10500 3881
rect 11000 3850 11050 3881
rect 12650 4319 12700 4350
rect 13200 4319 13250 4350
rect 11550 3850 11600 3881
rect 12100 3850 12150 3881
rect 12650 3850 12700 3881
rect 13200 3850 13250 3881
rect 13750 3850 13800 4350
rect -550 3842 -469 3850
rect -550 3808 -542 3842
rect -508 3808 -469 3842
rect -550 3800 -469 3808
rect -31 3842 81 3850
rect -31 3808 8 3842
rect 42 3808 81 3842
rect -31 3800 81 3808
rect 519 3842 631 3850
rect 519 3808 558 3842
rect 592 3808 631 3842
rect 519 3800 631 3808
rect 1069 3842 1181 3850
rect 1069 3808 1108 3842
rect 1142 3808 1181 3842
rect 1069 3800 1181 3808
rect 1619 3842 1731 3850
rect 1619 3808 1658 3842
rect 1692 3808 1731 3842
rect 1619 3800 1731 3808
rect 2169 3842 2281 3850
rect 2169 3808 2208 3842
rect 2242 3808 2281 3842
rect 2169 3800 2281 3808
rect 2719 3842 2831 3850
rect 2719 3808 2758 3842
rect 2792 3808 2831 3842
rect 2719 3800 2831 3808
rect 3269 3842 3381 3850
rect 3269 3808 3308 3842
rect 3342 3808 3381 3842
rect 3269 3800 3381 3808
rect 3819 3842 3931 3850
rect 3819 3808 3858 3842
rect 3892 3808 3931 3842
rect 3819 3800 3931 3808
rect 4369 3842 4481 3850
rect 4369 3808 4408 3842
rect 4442 3808 4481 3842
rect 4369 3800 4481 3808
rect 4919 3842 5031 3850
rect 4919 3808 4958 3842
rect 4992 3808 5031 3842
rect 4919 3800 5031 3808
rect 5469 3842 5581 3850
rect 5469 3808 5508 3842
rect 5542 3808 5581 3842
rect 5469 3800 5581 3808
rect 6019 3842 6131 3850
rect 6019 3808 6058 3842
rect 6092 3808 6131 3842
rect 6019 3800 6131 3808
rect 6569 3842 6681 3850
rect 6569 3808 6608 3842
rect 6642 3808 6681 3842
rect 6569 3800 6681 3808
rect 7119 3842 7231 3850
rect 7119 3808 7158 3842
rect 7192 3808 7231 3842
rect 7119 3800 7231 3808
rect 7669 3842 7781 3850
rect 7669 3808 7708 3842
rect 7742 3808 7781 3842
rect 7669 3800 7781 3808
rect 8219 3842 8331 3850
rect 8219 3808 8258 3842
rect 8292 3808 8331 3842
rect 8219 3800 8331 3808
rect 8769 3842 8881 3850
rect 8769 3808 8808 3842
rect 8842 3808 8881 3842
rect 8769 3800 8881 3808
rect 9319 3842 9431 3850
rect 9319 3808 9358 3842
rect 9392 3808 9431 3842
rect 9319 3800 9431 3808
rect 9869 3842 9981 3850
rect 9869 3808 9908 3842
rect 9942 3808 9981 3842
rect 9869 3800 9981 3808
rect 10419 3842 10531 3850
rect 10419 3808 10458 3842
rect 10492 3808 10531 3842
rect 10419 3800 10531 3808
rect 10969 3842 11081 3850
rect 10969 3808 11008 3842
rect 11042 3808 11081 3842
rect 10969 3800 11081 3808
rect 11519 3842 11631 3850
rect 11519 3808 11558 3842
rect 11592 3808 11631 3842
rect 11519 3800 11631 3808
rect 12069 3842 12181 3850
rect 12069 3808 12108 3842
rect 12142 3808 12181 3842
rect 12069 3800 12181 3808
rect 12619 3842 12731 3850
rect 12619 3808 12658 3842
rect 12692 3808 12731 3842
rect 12619 3800 12731 3808
rect 13169 3842 13281 3850
rect 13169 3808 13208 3842
rect 13242 3808 13281 3842
rect 13169 3800 13281 3808
rect 13719 3842 13800 3850
rect 13719 3808 13758 3842
rect 13792 3808 13800 3842
rect 13719 3800 13800 3808
rect -550 3300 -500 3800
rect 0 3769 50 3800
rect 550 3769 600 3800
rect 1100 3769 1150 3800
rect 1650 3769 1700 3800
rect 0 3300 50 3331
rect 550 3300 600 3331
rect 2200 3769 2250 3800
rect 2750 3769 2800 3800
rect 1100 3300 1150 3331
rect 1650 3300 1700 3331
rect 3300 3769 3350 3800
rect 3850 3769 3900 3800
rect 2200 3300 2250 3331
rect 2750 3300 2800 3331
rect 4400 3769 4450 3800
rect 4950 3769 5000 3800
rect 3300 3300 3350 3331
rect 3850 3300 3900 3331
rect 5500 3769 5550 3800
rect 6050 3769 6100 3800
rect 4400 3300 4450 3331
rect 4950 3300 5000 3331
rect 6600 3769 6650 3800
rect 7150 3769 7200 3800
rect 5500 3300 5550 3331
rect 6050 3300 6100 3331
rect 7700 3769 7750 3800
rect 8250 3769 8300 3800
rect 6600 3300 6650 3331
rect 7150 3300 7200 3331
rect 8800 3769 8850 3800
rect 9350 3769 9400 3800
rect 7700 3300 7750 3331
rect 8250 3300 8300 3331
rect 9900 3769 9950 3800
rect 10450 3769 10500 3800
rect 8800 3300 8850 3331
rect 9350 3300 9400 3331
rect 11000 3769 11050 3800
rect 11550 3769 11600 3800
rect 9900 3300 9950 3331
rect 10450 3300 10500 3331
rect 12100 3769 12150 3800
rect 12650 3769 12700 3800
rect 11000 3300 11050 3331
rect 11550 3300 11600 3331
rect 13200 3769 13250 3800
rect 12100 3300 12150 3331
rect 12650 3300 12700 3331
rect 13200 3300 13250 3331
rect 13750 3300 13800 3800
rect -550 3292 -469 3300
rect -550 3258 -542 3292
rect -508 3258 -469 3292
rect -550 3250 -469 3258
rect -31 3292 81 3300
rect -31 3258 8 3292
rect 42 3258 81 3292
rect -31 3250 81 3258
rect 519 3292 631 3300
rect 519 3258 558 3292
rect 592 3258 631 3292
rect 519 3250 631 3258
rect 1069 3292 1181 3300
rect 1069 3258 1108 3292
rect 1142 3258 1181 3292
rect 1069 3250 1181 3258
rect 1619 3292 1731 3300
rect 1619 3258 1658 3292
rect 1692 3258 1731 3292
rect 1619 3250 1731 3258
rect 2169 3292 2281 3300
rect 2169 3258 2208 3292
rect 2242 3258 2281 3292
rect 2169 3250 2281 3258
rect 2719 3292 2831 3300
rect 2719 3258 2758 3292
rect 2792 3258 2831 3292
rect 2719 3250 2831 3258
rect 3269 3292 3381 3300
rect 3269 3258 3308 3292
rect 3342 3258 3381 3292
rect 3269 3250 3381 3258
rect 3819 3292 3931 3300
rect 3819 3258 3858 3292
rect 3892 3258 3931 3292
rect 3819 3250 3931 3258
rect 4369 3292 4481 3300
rect 4369 3258 4408 3292
rect 4442 3258 4481 3292
rect 4369 3250 4481 3258
rect 4919 3292 5031 3300
rect 4919 3258 4958 3292
rect 4992 3258 5031 3292
rect 4919 3250 5031 3258
rect 5469 3292 5581 3300
rect 5469 3258 5508 3292
rect 5542 3258 5581 3292
rect 5469 3250 5581 3258
rect 6019 3292 6131 3300
rect 6019 3258 6058 3292
rect 6092 3258 6131 3292
rect 6019 3250 6131 3258
rect 6569 3292 6681 3300
rect 6569 3258 6608 3292
rect 6642 3258 6681 3292
rect 6569 3250 6681 3258
rect 7119 3292 7231 3300
rect 7119 3258 7158 3292
rect 7192 3258 7231 3292
rect 7119 3250 7231 3258
rect 7669 3292 7781 3300
rect 7669 3258 7708 3292
rect 7742 3258 7781 3292
rect 7669 3250 7781 3258
rect 8219 3292 8331 3300
rect 8219 3258 8258 3292
rect 8292 3258 8331 3292
rect 8219 3250 8331 3258
rect 8769 3292 8881 3300
rect 8769 3258 8808 3292
rect 8842 3258 8881 3292
rect 8769 3250 8881 3258
rect 9319 3292 9431 3300
rect 9319 3258 9358 3292
rect 9392 3258 9431 3292
rect 9319 3250 9431 3258
rect 9869 3292 9981 3300
rect 9869 3258 9908 3292
rect 9942 3258 9981 3292
rect 9869 3250 9981 3258
rect 10419 3292 10531 3300
rect 10419 3258 10458 3292
rect 10492 3258 10531 3292
rect 10419 3250 10531 3258
rect 10969 3292 11081 3300
rect 10969 3258 11008 3292
rect 11042 3258 11081 3292
rect 10969 3250 11081 3258
rect 11519 3292 11631 3300
rect 11519 3258 11558 3292
rect 11592 3258 11631 3292
rect 11519 3250 11631 3258
rect 12069 3292 12181 3300
rect 12069 3258 12108 3292
rect 12142 3258 12181 3292
rect 12069 3250 12181 3258
rect 12619 3292 12731 3300
rect 12619 3258 12658 3292
rect 12692 3258 12731 3292
rect 12619 3250 12731 3258
rect 13169 3292 13281 3300
rect 13169 3258 13208 3292
rect 13242 3258 13281 3292
rect 13169 3250 13281 3258
rect 13719 3292 13800 3300
rect 13719 3258 13758 3292
rect 13792 3258 13800 3292
rect 13719 3250 13800 3258
rect -550 2750 -500 3250
rect 0 3219 50 3250
rect 550 3219 600 3250
rect 1100 3219 1150 3250
rect 0 2750 50 2781
rect 1650 3219 1700 3250
rect 2200 3219 2250 3250
rect 550 2750 600 2781
rect 1100 2750 1150 2781
rect 2750 3219 2800 3250
rect 3300 3219 3350 3250
rect 1650 2750 1700 2781
rect 2200 2750 2250 2781
rect 3850 3219 3900 3250
rect 4400 3219 4450 3250
rect 2750 2750 2800 2781
rect 3300 2750 3350 2781
rect 4950 3219 5000 3250
rect 5500 3219 5550 3250
rect 3850 2750 3900 2781
rect 4400 2750 4450 2781
rect 6050 3219 6100 3250
rect 6600 3219 6650 3250
rect 4950 2750 5000 2781
rect 5500 2750 5550 2781
rect 7150 3219 7200 3250
rect 7700 3219 7750 3250
rect 6050 2750 6100 2781
rect 6600 2750 6650 2781
rect 8250 3219 8300 3250
rect 8800 3219 8850 3250
rect 7150 2750 7200 2781
rect 7700 2750 7750 2781
rect 9350 3219 9400 3250
rect 9900 3219 9950 3250
rect 8250 2750 8300 2781
rect 8800 2750 8850 2781
rect 10450 3219 10500 3250
rect 11000 3219 11050 3250
rect 9350 2750 9400 2781
rect 9900 2750 9950 2781
rect 11550 3219 11600 3250
rect 12100 3219 12150 3250
rect 10450 2750 10500 2781
rect 11000 2750 11050 2781
rect 12650 3219 12700 3250
rect 13200 3219 13250 3250
rect 11550 2750 11600 2781
rect 12100 2750 12150 2781
rect 12650 2750 12700 2781
rect 13200 2750 13250 2781
rect 13750 2750 13800 3250
rect -550 2742 -469 2750
rect -550 2708 -542 2742
rect -508 2708 -469 2742
rect -550 2700 -469 2708
rect -31 2742 81 2750
rect -31 2708 8 2742
rect 42 2708 81 2742
rect -31 2700 81 2708
rect 519 2742 631 2750
rect 519 2708 558 2742
rect 592 2708 631 2742
rect 519 2700 631 2708
rect 1069 2742 1181 2750
rect 1069 2708 1108 2742
rect 1142 2708 1181 2742
rect 1069 2700 1181 2708
rect 1619 2742 1731 2750
rect 1619 2708 1658 2742
rect 1692 2708 1731 2742
rect 1619 2700 1731 2708
rect 2169 2742 2281 2750
rect 2169 2708 2208 2742
rect 2242 2708 2281 2742
rect 2169 2700 2281 2708
rect 2719 2742 2831 2750
rect 2719 2708 2758 2742
rect 2792 2708 2831 2742
rect 2719 2700 2831 2708
rect 3269 2742 3381 2750
rect 3269 2708 3308 2742
rect 3342 2708 3381 2742
rect 3269 2700 3381 2708
rect 3819 2742 3931 2750
rect 3819 2708 3858 2742
rect 3892 2708 3931 2742
rect 3819 2700 3931 2708
rect 4369 2742 4481 2750
rect 4369 2708 4408 2742
rect 4442 2708 4481 2742
rect 4369 2700 4481 2708
rect 4919 2742 5031 2750
rect 4919 2708 4958 2742
rect 4992 2708 5031 2742
rect 4919 2700 5031 2708
rect 5469 2742 5581 2750
rect 5469 2708 5508 2742
rect 5542 2708 5581 2742
rect 5469 2700 5581 2708
rect 6019 2742 6131 2750
rect 6019 2708 6058 2742
rect 6092 2708 6131 2742
rect 6019 2700 6131 2708
rect 6569 2742 6681 2750
rect 6569 2708 6608 2742
rect 6642 2708 6681 2742
rect 6569 2700 6681 2708
rect 7119 2742 7231 2750
rect 7119 2708 7158 2742
rect 7192 2708 7231 2742
rect 7119 2700 7231 2708
rect 7669 2742 7781 2750
rect 7669 2708 7708 2742
rect 7742 2708 7781 2742
rect 7669 2700 7781 2708
rect 8219 2742 8331 2750
rect 8219 2708 8258 2742
rect 8292 2708 8331 2742
rect 8219 2700 8331 2708
rect 8769 2742 8881 2750
rect 8769 2708 8808 2742
rect 8842 2708 8881 2742
rect 8769 2700 8881 2708
rect 9319 2742 9431 2750
rect 9319 2708 9358 2742
rect 9392 2708 9431 2742
rect 9319 2700 9431 2708
rect 9869 2742 9981 2750
rect 9869 2708 9908 2742
rect 9942 2708 9981 2742
rect 9869 2700 9981 2708
rect 10419 2742 10531 2750
rect 10419 2708 10458 2742
rect 10492 2708 10531 2742
rect 10419 2700 10531 2708
rect 10969 2742 11081 2750
rect 10969 2708 11008 2742
rect 11042 2708 11081 2742
rect 10969 2700 11081 2708
rect 11519 2742 11631 2750
rect 11519 2708 11558 2742
rect 11592 2708 11631 2742
rect 11519 2700 11631 2708
rect 12069 2742 12181 2750
rect 12069 2708 12108 2742
rect 12142 2708 12181 2742
rect 12069 2700 12181 2708
rect 12619 2742 12731 2750
rect 12619 2708 12658 2742
rect 12692 2708 12731 2742
rect 12619 2700 12731 2708
rect 13169 2742 13281 2750
rect 13169 2708 13208 2742
rect 13242 2708 13281 2742
rect 13169 2700 13281 2708
rect 13719 2742 13800 2750
rect 13719 2708 13758 2742
rect 13792 2708 13800 2742
rect 13719 2700 13800 2708
rect -550 2200 -500 2700
rect 0 2669 50 2700
rect 550 2669 600 2700
rect 1100 2669 1150 2700
rect 1650 2669 1700 2700
rect 0 2200 50 2231
rect 550 2200 600 2231
rect 2200 2669 2250 2700
rect 2750 2669 2800 2700
rect 1100 2200 1150 2231
rect 1650 2200 1700 2231
rect 3300 2669 3350 2700
rect 3850 2669 3900 2700
rect 2200 2200 2250 2231
rect 2750 2200 2800 2231
rect 4400 2669 4450 2700
rect 4950 2669 5000 2700
rect 3300 2200 3350 2231
rect 3850 2200 3900 2231
rect 5500 2669 5550 2700
rect 6050 2669 6100 2700
rect 4400 2200 4450 2231
rect 4950 2200 5000 2231
rect 6600 2669 6650 2700
rect 7150 2669 7200 2700
rect 5500 2200 5550 2231
rect 6050 2200 6100 2231
rect 7700 2669 7750 2700
rect 8250 2669 8300 2700
rect 6600 2200 6650 2231
rect 7150 2200 7200 2231
rect 8800 2669 8850 2700
rect 9350 2669 9400 2700
rect 7700 2200 7750 2231
rect 8250 2200 8300 2231
rect 9900 2669 9950 2700
rect 10450 2669 10500 2700
rect 8800 2200 8850 2231
rect 9350 2200 9400 2231
rect 11000 2669 11050 2700
rect 11550 2669 11600 2700
rect 9900 2200 9950 2231
rect 10450 2200 10500 2231
rect 12100 2669 12150 2700
rect 12650 2669 12700 2700
rect 11000 2200 11050 2231
rect 11550 2200 11600 2231
rect 13200 2669 13250 2700
rect 12100 2200 12150 2231
rect 12650 2200 12700 2231
rect 13200 2200 13250 2231
rect 13750 2200 13800 2700
rect -550 2192 -469 2200
rect -550 2158 -542 2192
rect -508 2158 -469 2192
rect -550 2150 -469 2158
rect -31 2192 81 2200
rect -31 2158 8 2192
rect 42 2158 81 2192
rect -31 2150 81 2158
rect 519 2192 631 2200
rect 519 2158 558 2192
rect 592 2158 631 2192
rect 519 2150 631 2158
rect 1069 2192 1181 2200
rect 1069 2158 1108 2192
rect 1142 2158 1181 2192
rect 1069 2150 1181 2158
rect 1619 2192 1731 2200
rect 1619 2158 1658 2192
rect 1692 2158 1731 2192
rect 1619 2150 1731 2158
rect 2169 2192 2281 2200
rect 2169 2158 2208 2192
rect 2242 2158 2281 2192
rect 2169 2150 2281 2158
rect 2719 2192 2831 2200
rect 2719 2158 2758 2192
rect 2792 2158 2831 2192
rect 2719 2150 2831 2158
rect 3269 2192 3381 2200
rect 3269 2158 3308 2192
rect 3342 2158 3381 2192
rect 3269 2150 3381 2158
rect 3819 2192 3931 2200
rect 3819 2158 3858 2192
rect 3892 2158 3931 2192
rect 3819 2150 3931 2158
rect 4369 2192 4481 2200
rect 4369 2158 4408 2192
rect 4442 2158 4481 2192
rect 4369 2150 4481 2158
rect 4919 2192 5031 2200
rect 4919 2158 4958 2192
rect 4992 2158 5031 2192
rect 4919 2150 5031 2158
rect 5469 2192 5581 2200
rect 5469 2158 5508 2192
rect 5542 2158 5581 2192
rect 5469 2150 5581 2158
rect 6019 2192 6131 2200
rect 6019 2158 6058 2192
rect 6092 2158 6131 2192
rect 6019 2150 6131 2158
rect 6569 2192 6681 2200
rect 6569 2158 6608 2192
rect 6642 2158 6681 2192
rect 6569 2150 6681 2158
rect 7119 2192 7231 2200
rect 7119 2158 7158 2192
rect 7192 2158 7231 2192
rect 7119 2150 7231 2158
rect 7669 2192 7781 2200
rect 7669 2158 7708 2192
rect 7742 2158 7781 2192
rect 7669 2150 7781 2158
rect 8219 2192 8331 2200
rect 8219 2158 8258 2192
rect 8292 2158 8331 2192
rect 8219 2150 8331 2158
rect 8769 2192 8881 2200
rect 8769 2158 8808 2192
rect 8842 2158 8881 2192
rect 8769 2150 8881 2158
rect 9319 2192 9431 2200
rect 9319 2158 9358 2192
rect 9392 2158 9431 2192
rect 9319 2150 9431 2158
rect 9869 2192 9981 2200
rect 9869 2158 9908 2192
rect 9942 2158 9981 2192
rect 9869 2150 9981 2158
rect 10419 2192 10531 2200
rect 10419 2158 10458 2192
rect 10492 2158 10531 2192
rect 10419 2150 10531 2158
rect 10969 2192 11081 2200
rect 10969 2158 11008 2192
rect 11042 2158 11081 2192
rect 10969 2150 11081 2158
rect 11519 2192 11631 2200
rect 11519 2158 11558 2192
rect 11592 2158 11631 2192
rect 11519 2150 11631 2158
rect 12069 2192 12181 2200
rect 12069 2158 12108 2192
rect 12142 2158 12181 2192
rect 12069 2150 12181 2158
rect 12619 2192 12731 2200
rect 12619 2158 12658 2192
rect 12692 2158 12731 2192
rect 12619 2150 12731 2158
rect 13169 2192 13281 2200
rect 13169 2158 13208 2192
rect 13242 2158 13281 2192
rect 13169 2150 13281 2158
rect 13719 2192 13800 2200
rect 13719 2158 13758 2192
rect 13792 2158 13800 2192
rect 13719 2150 13800 2158
rect -550 1650 -500 2150
rect 0 2119 50 2150
rect 550 2119 600 2150
rect 1100 2119 1150 2150
rect 0 1650 50 1681
rect 1650 2119 1700 2150
rect 2200 2119 2250 2150
rect 550 1650 600 1681
rect 1100 1650 1150 1681
rect 2750 2119 2800 2150
rect 3300 2119 3350 2150
rect 1650 1650 1700 1681
rect 2200 1650 2250 1681
rect 3850 2119 3900 2150
rect 4400 2119 4450 2150
rect 2750 1650 2800 1681
rect 3300 1650 3350 1681
rect 4950 2119 5000 2150
rect 5500 2119 5550 2150
rect 3850 1650 3900 1681
rect 4400 1650 4450 1681
rect 6050 2119 6100 2150
rect 6600 2119 6650 2150
rect 4950 1650 5000 1681
rect 5500 1650 5550 1681
rect 7150 2119 7200 2150
rect 7700 2119 7750 2150
rect 6050 1650 6100 1681
rect 6600 1650 6650 1681
rect 8250 2119 8300 2150
rect 8800 2119 8850 2150
rect 7150 1650 7200 1681
rect 7700 1650 7750 1681
rect 9350 2119 9400 2150
rect 9900 2119 9950 2150
rect 8250 1650 8300 1681
rect 8800 1650 8850 1681
rect 10450 2119 10500 2150
rect 11000 2119 11050 2150
rect 9350 1650 9400 1681
rect 9900 1650 9950 1681
rect 11550 2119 11600 2150
rect 12100 2119 12150 2150
rect 10450 1650 10500 1681
rect 11000 1650 11050 1681
rect 12650 2119 12700 2150
rect 13200 2119 13250 2150
rect 11550 1650 11600 1681
rect 12100 1650 12150 1681
rect 12650 1650 12700 1681
rect 13200 1650 13250 1681
rect 13750 1650 13800 2150
rect -550 1642 -469 1650
rect -550 1608 -542 1642
rect -508 1608 -469 1642
rect -550 1600 -469 1608
rect -31 1642 81 1650
rect -31 1608 8 1642
rect 42 1608 81 1642
rect -31 1600 81 1608
rect 519 1642 631 1650
rect 519 1608 558 1642
rect 592 1608 631 1642
rect 519 1600 631 1608
rect 1069 1642 1181 1650
rect 1069 1608 1108 1642
rect 1142 1608 1181 1642
rect 1069 1600 1181 1608
rect 1619 1642 1731 1650
rect 1619 1608 1658 1642
rect 1692 1608 1731 1642
rect 1619 1600 1731 1608
rect 2169 1642 2281 1650
rect 2169 1608 2208 1642
rect 2242 1608 2281 1642
rect 2169 1600 2281 1608
rect 2719 1642 2831 1650
rect 2719 1608 2758 1642
rect 2792 1608 2831 1642
rect 2719 1600 2831 1608
rect 3269 1642 3381 1650
rect 3269 1608 3308 1642
rect 3342 1608 3381 1642
rect 3269 1600 3381 1608
rect 3819 1642 3931 1650
rect 3819 1608 3858 1642
rect 3892 1608 3931 1642
rect 3819 1600 3931 1608
rect 4369 1642 4481 1650
rect 4369 1608 4408 1642
rect 4442 1608 4481 1642
rect 4369 1600 4481 1608
rect 4919 1642 5031 1650
rect 4919 1608 4958 1642
rect 4992 1608 5031 1642
rect 4919 1600 5031 1608
rect 5469 1642 5581 1650
rect 5469 1608 5508 1642
rect 5542 1608 5581 1642
rect 5469 1600 5581 1608
rect 6019 1642 6131 1650
rect 6019 1608 6058 1642
rect 6092 1608 6131 1642
rect 6019 1600 6131 1608
rect 6569 1642 6681 1650
rect 6569 1608 6608 1642
rect 6642 1608 6681 1642
rect 6569 1600 6681 1608
rect 7119 1642 7231 1650
rect 7119 1608 7158 1642
rect 7192 1608 7231 1642
rect 7119 1600 7231 1608
rect 7669 1642 7781 1650
rect 7669 1608 7708 1642
rect 7742 1608 7781 1642
rect 7669 1600 7781 1608
rect 8219 1642 8331 1650
rect 8219 1608 8258 1642
rect 8292 1608 8331 1642
rect 8219 1600 8331 1608
rect 8769 1642 8881 1650
rect 8769 1608 8808 1642
rect 8842 1608 8881 1642
rect 8769 1600 8881 1608
rect 9319 1642 9431 1650
rect 9319 1608 9358 1642
rect 9392 1608 9431 1642
rect 9319 1600 9431 1608
rect 9869 1642 9981 1650
rect 9869 1608 9908 1642
rect 9942 1608 9981 1642
rect 9869 1600 9981 1608
rect 10419 1642 10531 1650
rect 10419 1608 10458 1642
rect 10492 1608 10531 1642
rect 10419 1600 10531 1608
rect 10969 1642 11081 1650
rect 10969 1608 11008 1642
rect 11042 1608 11081 1642
rect 10969 1600 11081 1608
rect 11519 1642 11631 1650
rect 11519 1608 11558 1642
rect 11592 1608 11631 1642
rect 11519 1600 11631 1608
rect 12069 1642 12181 1650
rect 12069 1608 12108 1642
rect 12142 1608 12181 1642
rect 12069 1600 12181 1608
rect 12619 1642 12731 1650
rect 12619 1608 12658 1642
rect 12692 1608 12731 1642
rect 12619 1600 12731 1608
rect 13169 1642 13281 1650
rect 13169 1608 13208 1642
rect 13242 1608 13281 1642
rect 13169 1600 13281 1608
rect 13719 1642 13800 1650
rect 13719 1608 13758 1642
rect 13792 1608 13800 1642
rect 13719 1600 13800 1608
rect -550 1100 -500 1600
rect 0 1569 50 1600
rect 550 1569 600 1600
rect 1100 1569 1150 1600
rect 1650 1569 1700 1600
rect 0 1100 50 1131
rect 550 1100 600 1131
rect 2200 1569 2250 1600
rect 2750 1569 2800 1600
rect 1100 1100 1150 1131
rect 1650 1100 1700 1131
rect 3300 1569 3350 1600
rect 3850 1569 3900 1600
rect 2200 1100 2250 1131
rect 2750 1100 2800 1131
rect 4400 1569 4450 1600
rect 4950 1569 5000 1600
rect 3300 1100 3350 1131
rect 3850 1100 3900 1131
rect 5500 1569 5550 1600
rect 6050 1569 6100 1600
rect 4400 1100 4450 1131
rect 4950 1100 5000 1131
rect 6600 1569 6650 1600
rect 7150 1569 7200 1600
rect 5500 1100 5550 1131
rect 6050 1100 6100 1131
rect 7700 1569 7750 1600
rect 8250 1569 8300 1600
rect 6600 1100 6650 1131
rect 7150 1100 7200 1131
rect 8800 1569 8850 1600
rect 9350 1569 9400 1600
rect 7700 1100 7750 1131
rect 8250 1100 8300 1131
rect 9900 1569 9950 1600
rect 10450 1569 10500 1600
rect 8800 1100 8850 1131
rect 9350 1100 9400 1131
rect 11000 1569 11050 1600
rect 11550 1569 11600 1600
rect 9900 1100 9950 1131
rect 10450 1100 10500 1131
rect 12100 1569 12150 1600
rect 12650 1569 12700 1600
rect 11000 1100 11050 1131
rect 11550 1100 11600 1131
rect 13200 1569 13250 1600
rect 12100 1100 12150 1131
rect 12650 1100 12700 1131
rect 13200 1100 13250 1131
rect 13750 1100 13800 1600
rect -550 1092 -469 1100
rect -550 1058 -542 1092
rect -508 1058 -469 1092
rect -550 1050 -469 1058
rect -31 1092 81 1100
rect -31 1058 8 1092
rect 42 1058 81 1092
rect -31 1050 81 1058
rect 519 1092 631 1100
rect 519 1058 558 1092
rect 592 1058 631 1092
rect 519 1050 631 1058
rect 1069 1092 1181 1100
rect 1069 1058 1108 1092
rect 1142 1058 1181 1092
rect 1069 1050 1181 1058
rect 1619 1092 1731 1100
rect 1619 1058 1658 1092
rect 1692 1058 1731 1092
rect 1619 1050 1731 1058
rect 2169 1092 2281 1100
rect 2169 1058 2208 1092
rect 2242 1058 2281 1092
rect 2169 1050 2281 1058
rect 2719 1092 2831 1100
rect 2719 1058 2758 1092
rect 2792 1058 2831 1092
rect 2719 1050 2831 1058
rect 3269 1092 3381 1100
rect 3269 1058 3308 1092
rect 3342 1058 3381 1092
rect 3269 1050 3381 1058
rect 3819 1092 3931 1100
rect 3819 1058 3858 1092
rect 3892 1058 3931 1092
rect 3819 1050 3931 1058
rect 4369 1092 4481 1100
rect 4369 1058 4408 1092
rect 4442 1058 4481 1092
rect 4369 1050 4481 1058
rect 4919 1092 5031 1100
rect 4919 1058 4958 1092
rect 4992 1058 5031 1092
rect 4919 1050 5031 1058
rect 5469 1092 5581 1100
rect 5469 1058 5508 1092
rect 5542 1058 5581 1092
rect 5469 1050 5581 1058
rect 6019 1092 6131 1100
rect 6019 1058 6058 1092
rect 6092 1058 6131 1092
rect 6019 1050 6131 1058
rect 6569 1092 6681 1100
rect 6569 1058 6608 1092
rect 6642 1058 6681 1092
rect 6569 1050 6681 1058
rect 7119 1092 7231 1100
rect 7119 1058 7158 1092
rect 7192 1058 7231 1092
rect 7119 1050 7231 1058
rect 7669 1092 7781 1100
rect 7669 1058 7708 1092
rect 7742 1058 7781 1092
rect 7669 1050 7781 1058
rect 8219 1092 8331 1100
rect 8219 1058 8258 1092
rect 8292 1058 8331 1092
rect 8219 1050 8331 1058
rect 8769 1092 8881 1100
rect 8769 1058 8808 1092
rect 8842 1058 8881 1092
rect 8769 1050 8881 1058
rect 9319 1092 9431 1100
rect 9319 1058 9358 1092
rect 9392 1058 9431 1092
rect 9319 1050 9431 1058
rect 9869 1092 9981 1100
rect 9869 1058 9908 1092
rect 9942 1058 9981 1092
rect 9869 1050 9981 1058
rect 10419 1092 10531 1100
rect 10419 1058 10458 1092
rect 10492 1058 10531 1092
rect 10419 1050 10531 1058
rect 10969 1092 11081 1100
rect 10969 1058 11008 1092
rect 11042 1058 11081 1092
rect 10969 1050 11081 1058
rect 11519 1092 11631 1100
rect 11519 1058 11558 1092
rect 11592 1058 11631 1092
rect 11519 1050 11631 1058
rect 12069 1092 12181 1100
rect 12069 1058 12108 1092
rect 12142 1058 12181 1092
rect 12069 1050 12181 1058
rect 12619 1092 12731 1100
rect 12619 1058 12658 1092
rect 12692 1058 12731 1092
rect 12619 1050 12731 1058
rect 13169 1092 13281 1100
rect 13169 1058 13208 1092
rect 13242 1058 13281 1092
rect 13169 1050 13281 1058
rect 13719 1092 13800 1100
rect 13719 1058 13758 1092
rect 13792 1058 13800 1092
rect 13719 1050 13800 1058
rect -550 550 -500 1050
rect 0 1019 50 1050
rect 550 1019 600 1050
rect 1100 1019 1150 1050
rect 0 550 50 581
rect 1650 1019 1700 1050
rect 2200 1019 2250 1050
rect 550 550 600 581
rect 1100 550 1150 581
rect 2750 1019 2800 1050
rect 3300 1019 3350 1050
rect 1650 550 1700 581
rect 2200 550 2250 581
rect 3850 1019 3900 1050
rect 4400 1019 4450 1050
rect 2750 550 2800 581
rect 3300 550 3350 581
rect 4950 1019 5000 1050
rect 5500 1019 5550 1050
rect 3850 550 3900 581
rect 4400 550 4450 581
rect 6050 1019 6100 1050
rect 6600 1019 6650 1050
rect 4950 550 5000 581
rect 5500 550 5550 581
rect 7150 1019 7200 1050
rect 7700 1019 7750 1050
rect 6050 550 6100 581
rect 6600 550 6650 581
rect 8250 1019 8300 1050
rect 8800 1019 8850 1050
rect 7150 550 7200 581
rect 7700 550 7750 581
rect 9350 1019 9400 1050
rect 9900 1019 9950 1050
rect 8250 550 8300 581
rect 8800 550 8850 581
rect 10450 1019 10500 1050
rect 11000 1019 11050 1050
rect 9350 550 9400 581
rect 9900 550 9950 581
rect 11550 1019 11600 1050
rect 12100 1019 12150 1050
rect 10450 550 10500 581
rect 11000 550 11050 581
rect 12650 1019 12700 1050
rect 13200 1019 13250 1050
rect 11550 550 11600 581
rect 12100 550 12150 581
rect 12650 550 12700 581
rect 13200 550 13250 581
rect 13750 550 13800 1050
rect -550 542 -469 550
rect -550 508 -542 542
rect -508 508 -469 542
rect -550 500 -469 508
rect -31 542 81 550
rect -31 508 8 542
rect 42 508 81 542
rect -31 500 81 508
rect 519 542 631 550
rect 519 508 558 542
rect 592 508 631 542
rect 519 500 631 508
rect 1069 542 1181 550
rect 1069 508 1108 542
rect 1142 508 1181 542
rect 1069 500 1181 508
rect 1619 542 1731 550
rect 1619 508 1658 542
rect 1692 508 1731 542
rect 1619 500 1731 508
rect 2169 542 2281 550
rect 2169 508 2208 542
rect 2242 508 2281 542
rect 2169 500 2281 508
rect 2719 542 2831 550
rect 2719 508 2758 542
rect 2792 508 2831 542
rect 2719 500 2831 508
rect 3269 542 3381 550
rect 3269 508 3308 542
rect 3342 508 3381 542
rect 3269 500 3381 508
rect 3819 542 3931 550
rect 3819 508 3858 542
rect 3892 508 3931 542
rect 3819 500 3931 508
rect 4369 542 4481 550
rect 4369 508 4408 542
rect 4442 508 4481 542
rect 4369 500 4481 508
rect 4919 542 5031 550
rect 4919 508 4958 542
rect 4992 508 5031 542
rect 4919 500 5031 508
rect 5469 542 5581 550
rect 5469 508 5508 542
rect 5542 508 5581 542
rect 5469 500 5581 508
rect 6019 542 6131 550
rect 6019 508 6058 542
rect 6092 508 6131 542
rect 6019 500 6131 508
rect 6569 542 6681 550
rect 6569 508 6608 542
rect 6642 508 6681 542
rect 6569 500 6681 508
rect 7119 542 7231 550
rect 7119 508 7158 542
rect 7192 508 7231 542
rect 7119 500 7231 508
rect 7669 542 7781 550
rect 7669 508 7708 542
rect 7742 508 7781 542
rect 7669 500 7781 508
rect 8219 542 8331 550
rect 8219 508 8258 542
rect 8292 508 8331 542
rect 8219 500 8331 508
rect 8769 542 8881 550
rect 8769 508 8808 542
rect 8842 508 8881 542
rect 8769 500 8881 508
rect 9319 542 9431 550
rect 9319 508 9358 542
rect 9392 508 9431 542
rect 9319 500 9431 508
rect 9869 542 9981 550
rect 9869 508 9908 542
rect 9942 508 9981 542
rect 9869 500 9981 508
rect 10419 542 10531 550
rect 10419 508 10458 542
rect 10492 508 10531 542
rect 10419 500 10531 508
rect 10969 542 11081 550
rect 10969 508 11008 542
rect 11042 508 11081 542
rect 10969 500 11081 508
rect 11519 542 11631 550
rect 11519 508 11558 542
rect 11592 508 11631 542
rect 11519 500 11631 508
rect 12069 542 12181 550
rect 12069 508 12108 542
rect 12142 508 12181 542
rect 12069 500 12181 508
rect 12619 542 12731 550
rect 12619 508 12658 542
rect 12692 508 12731 542
rect 12619 500 12731 508
rect 13169 542 13281 550
rect 13169 508 13208 542
rect 13242 508 13281 542
rect 13169 500 13281 508
rect 13719 542 13800 550
rect 13719 508 13758 542
rect 13792 508 13800 542
rect 13719 500 13800 508
rect -550 0 -500 500
rect 0 469 50 500
rect 550 469 600 500
rect 1100 469 1150 500
rect 1650 469 1700 500
rect 0 0 50 31
rect 550 0 600 31
rect 2200 469 2250 500
rect 2750 469 2800 500
rect 1100 0 1150 31
rect 1650 0 1700 31
rect 3300 469 3350 500
rect 3850 469 3900 500
rect 2200 0 2250 31
rect 2750 0 2800 31
rect 4400 469 4450 500
rect 4950 469 5000 500
rect 3300 0 3350 31
rect 3850 0 3900 31
rect 5500 469 5550 500
rect 6050 469 6100 500
rect 4400 0 4450 31
rect 4950 0 5000 31
rect 6600 469 6650 500
rect 7150 469 7200 500
rect 5500 0 5550 31
rect 6050 0 6100 31
rect 7700 469 7750 500
rect 8250 469 8300 500
rect 6600 0 6650 31
rect 7150 0 7200 31
rect 8800 469 8850 500
rect 9350 469 9400 500
rect 7700 0 7750 31
rect 8250 0 8300 31
rect 9900 469 9950 500
rect 10450 469 10500 500
rect 8800 0 8850 31
rect 9350 0 9400 31
rect 11000 469 11050 500
rect 11550 469 11600 500
rect 9900 0 9950 31
rect 10450 0 10500 31
rect 12100 469 12150 500
rect 12650 469 12700 500
rect 11000 0 11050 31
rect 11550 0 11600 31
rect 13200 469 13250 500
rect 12100 0 12150 31
rect 12650 0 12700 31
rect 13200 0 13250 31
rect 13750 0 13800 500
rect -550 -8 -469 0
rect -550 -42 -542 -8
rect -508 -42 -469 -8
rect -550 -50 -469 -42
rect -31 -8 81 0
rect -31 -42 8 -8
rect 42 -42 81 -8
rect -31 -50 81 -42
rect 519 -8 631 0
rect 519 -42 558 -8
rect 592 -42 631 -8
rect 519 -50 631 -42
rect 1069 -8 1181 0
rect 1069 -42 1108 -8
rect 1142 -42 1181 -8
rect 1069 -50 1181 -42
rect 1619 -8 1731 0
rect 1619 -42 1658 -8
rect 1692 -42 1731 -8
rect 1619 -50 1731 -42
rect 2169 -8 2281 0
rect 2169 -42 2208 -8
rect 2242 -42 2281 -8
rect 2169 -50 2281 -42
rect 2719 -8 2831 0
rect 2719 -42 2758 -8
rect 2792 -42 2831 -8
rect 2719 -50 2831 -42
rect 3269 -8 3381 0
rect 3269 -42 3308 -8
rect 3342 -42 3381 -8
rect 3269 -50 3381 -42
rect 3819 -8 3931 0
rect 3819 -42 3858 -8
rect 3892 -42 3931 -8
rect 3819 -50 3931 -42
rect 4369 -8 4481 0
rect 4369 -42 4408 -8
rect 4442 -42 4481 -8
rect 4369 -50 4481 -42
rect 4919 -8 5031 0
rect 4919 -42 4958 -8
rect 4992 -42 5031 -8
rect 4919 -50 5031 -42
rect 5469 -8 5581 0
rect 5469 -42 5508 -8
rect 5542 -42 5581 -8
rect 5469 -50 5581 -42
rect 6019 -8 6131 0
rect 6019 -42 6058 -8
rect 6092 -42 6131 -8
rect 6019 -50 6131 -42
rect 6569 -8 6681 0
rect 6569 -42 6608 -8
rect 6642 -42 6681 -8
rect 6569 -50 6681 -42
rect 7119 -8 7231 0
rect 7119 -42 7158 -8
rect 7192 -42 7231 -8
rect 7119 -50 7231 -42
rect 7669 -8 7781 0
rect 7669 -42 7708 -8
rect 7742 -42 7781 -8
rect 7669 -50 7781 -42
rect 8219 -8 8331 0
rect 8219 -42 8258 -8
rect 8292 -42 8331 -8
rect 8219 -50 8331 -42
rect 8769 -8 8881 0
rect 8769 -42 8808 -8
rect 8842 -42 8881 -8
rect 8769 -50 8881 -42
rect 9319 -8 9431 0
rect 9319 -42 9358 -8
rect 9392 -42 9431 -8
rect 9319 -50 9431 -42
rect 9869 -8 9981 0
rect 9869 -42 9908 -8
rect 9942 -42 9981 -8
rect 9869 -50 9981 -42
rect 10419 -8 10531 0
rect 10419 -42 10458 -8
rect 10492 -42 10531 -8
rect 10419 -50 10531 -42
rect 10969 -8 11081 0
rect 10969 -42 11008 -8
rect 11042 -42 11081 -8
rect 10969 -50 11081 -42
rect 11519 -8 11631 0
rect 11519 -42 11558 -8
rect 11592 -42 11631 -8
rect 11519 -50 11631 -42
rect 12069 -8 12181 0
rect 12069 -42 12108 -8
rect 12142 -42 12181 -8
rect 12069 -50 12181 -42
rect 12619 -8 12731 0
rect 12619 -42 12658 -8
rect 12692 -42 12731 -8
rect 12619 -50 12731 -42
rect 13169 -8 13281 0
rect 13169 -42 13208 -8
rect 13242 -42 13281 -8
rect 13169 -50 13281 -42
rect 13719 -8 13800 0
rect 13719 -42 13758 -8
rect 13792 -42 13800 -8
rect 13719 -50 13800 -42
rect -550 -550 -500 -50
rect 0 -81 50 -50
rect 550 -81 600 -50
rect 1100 -81 1150 -50
rect 1650 -81 1700 -50
rect 2200 -81 2250 -50
rect 2750 -81 2800 -50
rect 3300 -81 3350 -50
rect 3850 -81 3900 -50
rect 4400 -81 4450 -50
rect 4950 -81 5000 -50
rect 5500 -81 5550 -50
rect 6050 -81 6100 -50
rect 6600 -81 6650 -50
rect 7150 -81 7200 -50
rect 7700 -81 7750 -50
rect 8250 -81 8300 -50
rect 8800 -81 8850 -50
rect 9350 -81 9400 -50
rect 9900 -81 9950 -50
rect 10450 -81 10500 -50
rect 11000 -81 11050 -50
rect 11550 -81 11600 -50
rect 12100 -81 12150 -50
rect 12650 -81 12700 -50
rect 13200 -81 13250 -50
rect 0 -550 50 -519
rect 550 -550 600 -519
rect 1100 -550 1150 -519
rect 1650 -550 1700 -519
rect 2200 -550 2250 -519
rect 2750 -550 2800 -519
rect 3300 -550 3350 -519
rect 3850 -550 3900 -519
rect 4400 -550 4450 -519
rect 4950 -550 5000 -519
rect 5500 -550 5550 -519
rect 6050 -550 6100 -519
rect 6600 -550 6650 -519
rect 7150 -550 7200 -519
rect 7700 -550 7750 -519
rect 8250 -550 8300 -519
rect 8800 -550 8850 -519
rect 9350 -550 9400 -519
rect 9900 -550 9950 -519
rect 10450 -550 10500 -519
rect 11000 -550 11050 -519
rect 11550 -550 11600 -519
rect 12100 -550 12150 -519
rect 12650 -550 12700 -519
rect 13200 -550 13250 -519
rect 13750 -550 13800 -50
rect -550 -558 13800 -550
rect -550 -592 -542 -558
rect -508 -592 8 -558
rect 42 -592 558 -558
rect 592 -592 1108 -558
rect 1142 -592 1658 -558
rect 1692 -592 2208 -558
rect 2242 -592 2758 -558
rect 2792 -592 3308 -558
rect 3342 -592 3858 -558
rect 3892 -592 4408 -558
rect 4442 -592 4958 -558
rect 4992 -592 5508 -558
rect 5542 -592 6058 -558
rect 6092 -592 6608 -558
rect 6642 -592 7158 -558
rect 7192 -592 7708 -558
rect 7742 -592 8258 -558
rect 8292 -592 8808 -558
rect 8842 -592 9358 -558
rect 9392 -592 9908 -558
rect 9942 -592 10458 -558
rect 10492 -592 11008 -558
rect 11042 -592 11558 -558
rect 11592 -592 12108 -558
rect 12142 -592 12658 -558
rect 12692 -592 13208 -558
rect 13242 -592 13758 -558
rect 13792 -592 13800 -558
rect -550 -600 13800 -592
<< polycont >>
rect -542 13708 -508 13742
rect 8 13708 42 13742
rect 558 13708 592 13742
rect 1108 13708 1142 13742
rect 1658 13708 1692 13742
rect 2208 13708 2242 13742
rect 2758 13708 2792 13742
rect 3308 13708 3342 13742
rect 3858 13708 3892 13742
rect 4408 13708 4442 13742
rect 4958 13708 4992 13742
rect 5508 13708 5542 13742
rect 6058 13708 6092 13742
rect 6608 13708 6642 13742
rect 7158 13708 7192 13742
rect 7708 13708 7742 13742
rect 8258 13708 8292 13742
rect 8808 13708 8842 13742
rect 9358 13708 9392 13742
rect 9908 13708 9942 13742
rect 10458 13708 10492 13742
rect 11008 13708 11042 13742
rect 11558 13708 11592 13742
rect 12108 13708 12142 13742
rect 12658 13708 12692 13742
rect 13208 13708 13242 13742
rect 13758 13708 13792 13742
rect -542 13158 -508 13192
rect 8 13158 42 13192
rect 558 13158 592 13192
rect 1108 13158 1142 13192
rect 1658 13158 1692 13192
rect 2208 13158 2242 13192
rect 2758 13158 2792 13192
rect 3308 13158 3342 13192
rect 3858 13158 3892 13192
rect 4408 13158 4442 13192
rect 4958 13158 4992 13192
rect 5508 13158 5542 13192
rect 6058 13158 6092 13192
rect 6608 13158 6642 13192
rect 7158 13158 7192 13192
rect 7708 13158 7742 13192
rect 8258 13158 8292 13192
rect 8808 13158 8842 13192
rect 9358 13158 9392 13192
rect 9908 13158 9942 13192
rect 10458 13158 10492 13192
rect 11008 13158 11042 13192
rect 11558 13158 11592 13192
rect 12108 13158 12142 13192
rect 12658 13158 12692 13192
rect 13208 13158 13242 13192
rect 13758 13158 13792 13192
rect -542 12608 -508 12642
rect 8 12608 42 12642
rect 558 12608 592 12642
rect 1108 12608 1142 12642
rect 1658 12608 1692 12642
rect 2208 12608 2242 12642
rect 2758 12608 2792 12642
rect 3308 12608 3342 12642
rect 3858 12608 3892 12642
rect 4408 12608 4442 12642
rect 4958 12608 4992 12642
rect 5508 12608 5542 12642
rect 6058 12608 6092 12642
rect 6608 12608 6642 12642
rect 7158 12608 7192 12642
rect 7708 12608 7742 12642
rect 8258 12608 8292 12642
rect 8808 12608 8842 12642
rect 9358 12608 9392 12642
rect 9908 12608 9942 12642
rect 10458 12608 10492 12642
rect 11008 12608 11042 12642
rect 11558 12608 11592 12642
rect 12108 12608 12142 12642
rect 12658 12608 12692 12642
rect 13208 12608 13242 12642
rect 13758 12608 13792 12642
rect -542 12058 -508 12092
rect 8 12058 42 12092
rect 558 12058 592 12092
rect 1108 12058 1142 12092
rect 1658 12058 1692 12092
rect 2208 12058 2242 12092
rect 2758 12058 2792 12092
rect 3308 12058 3342 12092
rect 3858 12058 3892 12092
rect 4408 12058 4442 12092
rect 4958 12058 4992 12092
rect 5508 12058 5542 12092
rect 6058 12058 6092 12092
rect 6608 12058 6642 12092
rect 7158 12058 7192 12092
rect 7708 12058 7742 12092
rect 8258 12058 8292 12092
rect 8808 12058 8842 12092
rect 9358 12058 9392 12092
rect 9908 12058 9942 12092
rect 10458 12058 10492 12092
rect 11008 12058 11042 12092
rect 11558 12058 11592 12092
rect 12108 12058 12142 12092
rect 12658 12058 12692 12092
rect 13208 12058 13242 12092
rect 13758 12058 13792 12092
rect -542 11508 -508 11542
rect 8 11508 42 11542
rect 558 11508 592 11542
rect 1108 11508 1142 11542
rect 1658 11508 1692 11542
rect 2208 11508 2242 11542
rect 2758 11508 2792 11542
rect 3308 11508 3342 11542
rect 3858 11508 3892 11542
rect 4408 11508 4442 11542
rect 4958 11508 4992 11542
rect 5508 11508 5542 11542
rect 6058 11508 6092 11542
rect 6608 11508 6642 11542
rect 7158 11508 7192 11542
rect 7708 11508 7742 11542
rect 8258 11508 8292 11542
rect 8808 11508 8842 11542
rect 9358 11508 9392 11542
rect 9908 11508 9942 11542
rect 10458 11508 10492 11542
rect 11008 11508 11042 11542
rect 11558 11508 11592 11542
rect 12108 11508 12142 11542
rect 12658 11508 12692 11542
rect 13208 11508 13242 11542
rect 13758 11508 13792 11542
rect -542 10958 -508 10992
rect 8 10958 42 10992
rect 558 10958 592 10992
rect 1108 10958 1142 10992
rect 1658 10958 1692 10992
rect 2208 10958 2242 10992
rect 2758 10958 2792 10992
rect 3308 10958 3342 10992
rect 3858 10958 3892 10992
rect 4408 10958 4442 10992
rect 4958 10958 4992 10992
rect 5508 10958 5542 10992
rect 6058 10958 6092 10992
rect 6608 10958 6642 10992
rect 7158 10958 7192 10992
rect 7708 10958 7742 10992
rect 8258 10958 8292 10992
rect 8808 10958 8842 10992
rect 9358 10958 9392 10992
rect 9908 10958 9942 10992
rect 10458 10958 10492 10992
rect 11008 10958 11042 10992
rect 11558 10958 11592 10992
rect 12108 10958 12142 10992
rect 12658 10958 12692 10992
rect 13208 10958 13242 10992
rect 13758 10958 13792 10992
rect -542 10408 -508 10442
rect 8 10408 42 10442
rect 558 10408 592 10442
rect 1108 10408 1142 10442
rect 1658 10408 1692 10442
rect 2208 10408 2242 10442
rect 2758 10408 2792 10442
rect 3308 10408 3342 10442
rect 3858 10408 3892 10442
rect 4408 10408 4442 10442
rect 4958 10408 4992 10442
rect 5508 10408 5542 10442
rect 6058 10408 6092 10442
rect 6608 10408 6642 10442
rect 7158 10408 7192 10442
rect 7708 10408 7742 10442
rect 8258 10408 8292 10442
rect 8808 10408 8842 10442
rect 9358 10408 9392 10442
rect 9908 10408 9942 10442
rect 10458 10408 10492 10442
rect 11008 10408 11042 10442
rect 11558 10408 11592 10442
rect 12108 10408 12142 10442
rect 12658 10408 12692 10442
rect 13208 10408 13242 10442
rect 13758 10408 13792 10442
rect -542 9858 -508 9892
rect 8 9858 42 9892
rect 558 9858 592 9892
rect 1108 9858 1142 9892
rect 1658 9858 1692 9892
rect 2208 9858 2242 9892
rect 2758 9858 2792 9892
rect 3308 9858 3342 9892
rect 3858 9858 3892 9892
rect 4408 9858 4442 9892
rect 4958 9858 4992 9892
rect 5508 9858 5542 9892
rect 6058 9858 6092 9892
rect 6608 9858 6642 9892
rect 7158 9858 7192 9892
rect 7708 9858 7742 9892
rect 8258 9858 8292 9892
rect 8808 9858 8842 9892
rect 9358 9858 9392 9892
rect 9908 9858 9942 9892
rect 10458 9858 10492 9892
rect 11008 9858 11042 9892
rect 11558 9858 11592 9892
rect 12108 9858 12142 9892
rect 12658 9858 12692 9892
rect 13208 9858 13242 9892
rect 13758 9858 13792 9892
rect -542 9308 -508 9342
rect 8 9308 42 9342
rect 558 9308 592 9342
rect 1108 9308 1142 9342
rect 1658 9308 1692 9342
rect 2208 9308 2242 9342
rect 2758 9308 2792 9342
rect 3308 9308 3342 9342
rect 3858 9308 3892 9342
rect 4408 9308 4442 9342
rect 4958 9308 4992 9342
rect 5508 9308 5542 9342
rect 6058 9308 6092 9342
rect 6608 9308 6642 9342
rect 7158 9308 7192 9342
rect 7708 9308 7742 9342
rect 8258 9308 8292 9342
rect 8808 9308 8842 9342
rect 9358 9308 9392 9342
rect 9908 9308 9942 9342
rect 10458 9308 10492 9342
rect 11008 9308 11042 9342
rect 11558 9308 11592 9342
rect 12108 9308 12142 9342
rect 12658 9308 12692 9342
rect 13208 9308 13242 9342
rect 13758 9308 13792 9342
rect -542 8758 -508 8792
rect 8 8758 42 8792
rect 558 8758 592 8792
rect 1108 8758 1142 8792
rect 1658 8758 1692 8792
rect 2208 8758 2242 8792
rect 2758 8758 2792 8792
rect 3308 8758 3342 8792
rect 3858 8758 3892 8792
rect 4408 8758 4442 8792
rect 4958 8758 4992 8792
rect 5508 8758 5542 8792
rect 6058 8758 6092 8792
rect 6608 8758 6642 8792
rect 7158 8758 7192 8792
rect 7708 8758 7742 8792
rect 8258 8758 8292 8792
rect 8808 8758 8842 8792
rect 9358 8758 9392 8792
rect 9908 8758 9942 8792
rect 10458 8758 10492 8792
rect 11008 8758 11042 8792
rect 11558 8758 11592 8792
rect 12108 8758 12142 8792
rect 12658 8758 12692 8792
rect 13208 8758 13242 8792
rect 13758 8758 13792 8792
rect -542 8208 -508 8242
rect 8 8208 42 8242
rect 558 8208 592 8242
rect 1108 8208 1142 8242
rect 1658 8208 1692 8242
rect 2208 8208 2242 8242
rect 2758 8208 2792 8242
rect 3308 8208 3342 8242
rect 3858 8208 3892 8242
rect 4408 8208 4442 8242
rect 4958 8208 4992 8242
rect 5508 8208 5542 8242
rect 6058 8208 6092 8242
rect 6608 8208 6642 8242
rect 7158 8208 7192 8242
rect 7708 8208 7742 8242
rect 8258 8208 8292 8242
rect 8808 8208 8842 8242
rect 9358 8208 9392 8242
rect 9908 8208 9942 8242
rect 10458 8208 10492 8242
rect 11008 8208 11042 8242
rect 11558 8208 11592 8242
rect 12108 8208 12142 8242
rect 12658 8208 12692 8242
rect 13208 8208 13242 8242
rect 13758 8208 13792 8242
rect -542 7658 -508 7692
rect 8 7658 42 7692
rect 558 7658 592 7692
rect 1108 7658 1142 7692
rect 1658 7658 1692 7692
rect 2208 7658 2242 7692
rect 2758 7658 2792 7692
rect 3308 7658 3342 7692
rect 3858 7658 3892 7692
rect 4408 7658 4442 7692
rect 4958 7658 4992 7692
rect 5508 7658 5542 7692
rect 6058 7658 6092 7692
rect 6608 7658 6642 7692
rect 7158 7658 7192 7692
rect 7708 7658 7742 7692
rect 8258 7658 8292 7692
rect 8808 7658 8842 7692
rect 9358 7658 9392 7692
rect 9908 7658 9942 7692
rect 10458 7658 10492 7692
rect 11008 7658 11042 7692
rect 11558 7658 11592 7692
rect 12108 7658 12142 7692
rect 12658 7658 12692 7692
rect 13208 7658 13242 7692
rect 13758 7658 13792 7692
rect -542 7108 -508 7142
rect 8 7108 42 7142
rect 558 7108 592 7142
rect 1108 7108 1142 7142
rect 1658 7108 1692 7142
rect 2208 7108 2242 7142
rect 2758 7108 2792 7142
rect 3308 7108 3342 7142
rect 3858 7108 3892 7142
rect 4408 7108 4442 7142
rect 4958 7108 4992 7142
rect 5508 7108 5542 7142
rect 6058 7108 6092 7142
rect 6608 7108 6642 7142
rect 7158 7108 7192 7142
rect 7708 7108 7742 7142
rect 8258 7108 8292 7142
rect 8808 7108 8842 7142
rect 9358 7108 9392 7142
rect 9908 7108 9942 7142
rect 10458 7108 10492 7142
rect 11008 7108 11042 7142
rect 11558 7108 11592 7142
rect 12108 7108 12142 7142
rect 12658 7108 12692 7142
rect 13208 7108 13242 7142
rect 13758 7108 13792 7142
rect -542 6558 -508 6592
rect 8 6558 42 6592
rect 558 6558 592 6592
rect 1108 6558 1142 6592
rect 1658 6558 1692 6592
rect 2208 6558 2242 6592
rect 2758 6558 2792 6592
rect 3308 6558 3342 6592
rect 3858 6558 3892 6592
rect 4408 6558 4442 6592
rect 4958 6558 4992 6592
rect 5508 6558 5542 6592
rect 6058 6558 6092 6592
rect 6608 6558 6642 6592
rect 7158 6558 7192 6592
rect 7708 6558 7742 6592
rect 8258 6558 8292 6592
rect 8808 6558 8842 6592
rect 9358 6558 9392 6592
rect 9908 6558 9942 6592
rect 10458 6558 10492 6592
rect 11008 6558 11042 6592
rect 11558 6558 11592 6592
rect 12108 6558 12142 6592
rect 12658 6558 12692 6592
rect 13208 6558 13242 6592
rect 13758 6558 13792 6592
rect -542 6008 -508 6042
rect 8 6008 42 6042
rect 558 6008 592 6042
rect 1108 6008 1142 6042
rect 1658 6008 1692 6042
rect 2208 6008 2242 6042
rect 2758 6008 2792 6042
rect 3308 6008 3342 6042
rect 3858 6008 3892 6042
rect 4408 6008 4442 6042
rect 4958 6008 4992 6042
rect 5508 6008 5542 6042
rect 6058 6008 6092 6042
rect 6608 6008 6642 6042
rect 7158 6008 7192 6042
rect 7708 6008 7742 6042
rect 8258 6008 8292 6042
rect 8808 6008 8842 6042
rect 9358 6008 9392 6042
rect 9908 6008 9942 6042
rect 10458 6008 10492 6042
rect 11008 6008 11042 6042
rect 11558 6008 11592 6042
rect 12108 6008 12142 6042
rect 12658 6008 12692 6042
rect 13208 6008 13242 6042
rect 13758 6008 13792 6042
rect -542 5458 -508 5492
rect 8 5458 42 5492
rect 558 5458 592 5492
rect 1108 5458 1142 5492
rect 1658 5458 1692 5492
rect 2208 5458 2242 5492
rect 2758 5458 2792 5492
rect 3308 5458 3342 5492
rect 3858 5458 3892 5492
rect 4408 5458 4442 5492
rect 4958 5458 4992 5492
rect 5508 5458 5542 5492
rect 6058 5458 6092 5492
rect 6608 5458 6642 5492
rect 7158 5458 7192 5492
rect 7708 5458 7742 5492
rect 8258 5458 8292 5492
rect 8808 5458 8842 5492
rect 9358 5458 9392 5492
rect 9908 5458 9942 5492
rect 10458 5458 10492 5492
rect 11008 5458 11042 5492
rect 11558 5458 11592 5492
rect 12108 5458 12142 5492
rect 12658 5458 12692 5492
rect 13208 5458 13242 5492
rect 13758 5458 13792 5492
rect -542 4908 -508 4942
rect 8 4908 42 4942
rect 558 4908 592 4942
rect 1108 4908 1142 4942
rect 1658 4908 1692 4942
rect 2208 4908 2242 4942
rect 2758 4908 2792 4942
rect 3308 4908 3342 4942
rect 3858 4908 3892 4942
rect 4408 4908 4442 4942
rect 4958 4908 4992 4942
rect 5508 4908 5542 4942
rect 6058 4908 6092 4942
rect 6608 4908 6642 4942
rect 7158 4908 7192 4942
rect 7708 4908 7742 4942
rect 8258 4908 8292 4942
rect 8808 4908 8842 4942
rect 9358 4908 9392 4942
rect 9908 4908 9942 4942
rect 10458 4908 10492 4942
rect 11008 4908 11042 4942
rect 11558 4908 11592 4942
rect 12108 4908 12142 4942
rect 12658 4908 12692 4942
rect 13208 4908 13242 4942
rect 13758 4908 13792 4942
rect -542 4358 -508 4392
rect 8 4358 42 4392
rect 558 4358 592 4392
rect 1108 4358 1142 4392
rect 1658 4358 1692 4392
rect 2208 4358 2242 4392
rect 2758 4358 2792 4392
rect 3308 4358 3342 4392
rect 3858 4358 3892 4392
rect 4408 4358 4442 4392
rect 4958 4358 4992 4392
rect 5508 4358 5542 4392
rect 6058 4358 6092 4392
rect 6608 4358 6642 4392
rect 7158 4358 7192 4392
rect 7708 4358 7742 4392
rect 8258 4358 8292 4392
rect 8808 4358 8842 4392
rect 9358 4358 9392 4392
rect 9908 4358 9942 4392
rect 10458 4358 10492 4392
rect 11008 4358 11042 4392
rect 11558 4358 11592 4392
rect 12108 4358 12142 4392
rect 12658 4358 12692 4392
rect 13208 4358 13242 4392
rect 13758 4358 13792 4392
rect -542 3808 -508 3842
rect 8 3808 42 3842
rect 558 3808 592 3842
rect 1108 3808 1142 3842
rect 1658 3808 1692 3842
rect 2208 3808 2242 3842
rect 2758 3808 2792 3842
rect 3308 3808 3342 3842
rect 3858 3808 3892 3842
rect 4408 3808 4442 3842
rect 4958 3808 4992 3842
rect 5508 3808 5542 3842
rect 6058 3808 6092 3842
rect 6608 3808 6642 3842
rect 7158 3808 7192 3842
rect 7708 3808 7742 3842
rect 8258 3808 8292 3842
rect 8808 3808 8842 3842
rect 9358 3808 9392 3842
rect 9908 3808 9942 3842
rect 10458 3808 10492 3842
rect 11008 3808 11042 3842
rect 11558 3808 11592 3842
rect 12108 3808 12142 3842
rect 12658 3808 12692 3842
rect 13208 3808 13242 3842
rect 13758 3808 13792 3842
rect -542 3258 -508 3292
rect 8 3258 42 3292
rect 558 3258 592 3292
rect 1108 3258 1142 3292
rect 1658 3258 1692 3292
rect 2208 3258 2242 3292
rect 2758 3258 2792 3292
rect 3308 3258 3342 3292
rect 3858 3258 3892 3292
rect 4408 3258 4442 3292
rect 4958 3258 4992 3292
rect 5508 3258 5542 3292
rect 6058 3258 6092 3292
rect 6608 3258 6642 3292
rect 7158 3258 7192 3292
rect 7708 3258 7742 3292
rect 8258 3258 8292 3292
rect 8808 3258 8842 3292
rect 9358 3258 9392 3292
rect 9908 3258 9942 3292
rect 10458 3258 10492 3292
rect 11008 3258 11042 3292
rect 11558 3258 11592 3292
rect 12108 3258 12142 3292
rect 12658 3258 12692 3292
rect 13208 3258 13242 3292
rect 13758 3258 13792 3292
rect -542 2708 -508 2742
rect 8 2708 42 2742
rect 558 2708 592 2742
rect 1108 2708 1142 2742
rect 1658 2708 1692 2742
rect 2208 2708 2242 2742
rect 2758 2708 2792 2742
rect 3308 2708 3342 2742
rect 3858 2708 3892 2742
rect 4408 2708 4442 2742
rect 4958 2708 4992 2742
rect 5508 2708 5542 2742
rect 6058 2708 6092 2742
rect 6608 2708 6642 2742
rect 7158 2708 7192 2742
rect 7708 2708 7742 2742
rect 8258 2708 8292 2742
rect 8808 2708 8842 2742
rect 9358 2708 9392 2742
rect 9908 2708 9942 2742
rect 10458 2708 10492 2742
rect 11008 2708 11042 2742
rect 11558 2708 11592 2742
rect 12108 2708 12142 2742
rect 12658 2708 12692 2742
rect 13208 2708 13242 2742
rect 13758 2708 13792 2742
rect -542 2158 -508 2192
rect 8 2158 42 2192
rect 558 2158 592 2192
rect 1108 2158 1142 2192
rect 1658 2158 1692 2192
rect 2208 2158 2242 2192
rect 2758 2158 2792 2192
rect 3308 2158 3342 2192
rect 3858 2158 3892 2192
rect 4408 2158 4442 2192
rect 4958 2158 4992 2192
rect 5508 2158 5542 2192
rect 6058 2158 6092 2192
rect 6608 2158 6642 2192
rect 7158 2158 7192 2192
rect 7708 2158 7742 2192
rect 8258 2158 8292 2192
rect 8808 2158 8842 2192
rect 9358 2158 9392 2192
rect 9908 2158 9942 2192
rect 10458 2158 10492 2192
rect 11008 2158 11042 2192
rect 11558 2158 11592 2192
rect 12108 2158 12142 2192
rect 12658 2158 12692 2192
rect 13208 2158 13242 2192
rect 13758 2158 13792 2192
rect -542 1608 -508 1642
rect 8 1608 42 1642
rect 558 1608 592 1642
rect 1108 1608 1142 1642
rect 1658 1608 1692 1642
rect 2208 1608 2242 1642
rect 2758 1608 2792 1642
rect 3308 1608 3342 1642
rect 3858 1608 3892 1642
rect 4408 1608 4442 1642
rect 4958 1608 4992 1642
rect 5508 1608 5542 1642
rect 6058 1608 6092 1642
rect 6608 1608 6642 1642
rect 7158 1608 7192 1642
rect 7708 1608 7742 1642
rect 8258 1608 8292 1642
rect 8808 1608 8842 1642
rect 9358 1608 9392 1642
rect 9908 1608 9942 1642
rect 10458 1608 10492 1642
rect 11008 1608 11042 1642
rect 11558 1608 11592 1642
rect 12108 1608 12142 1642
rect 12658 1608 12692 1642
rect 13208 1608 13242 1642
rect 13758 1608 13792 1642
rect -542 1058 -508 1092
rect 8 1058 42 1092
rect 558 1058 592 1092
rect 1108 1058 1142 1092
rect 1658 1058 1692 1092
rect 2208 1058 2242 1092
rect 2758 1058 2792 1092
rect 3308 1058 3342 1092
rect 3858 1058 3892 1092
rect 4408 1058 4442 1092
rect 4958 1058 4992 1092
rect 5508 1058 5542 1092
rect 6058 1058 6092 1092
rect 6608 1058 6642 1092
rect 7158 1058 7192 1092
rect 7708 1058 7742 1092
rect 8258 1058 8292 1092
rect 8808 1058 8842 1092
rect 9358 1058 9392 1092
rect 9908 1058 9942 1092
rect 10458 1058 10492 1092
rect 11008 1058 11042 1092
rect 11558 1058 11592 1092
rect 12108 1058 12142 1092
rect 12658 1058 12692 1092
rect 13208 1058 13242 1092
rect 13758 1058 13792 1092
rect -542 508 -508 542
rect 8 508 42 542
rect 558 508 592 542
rect 1108 508 1142 542
rect 1658 508 1692 542
rect 2208 508 2242 542
rect 2758 508 2792 542
rect 3308 508 3342 542
rect 3858 508 3892 542
rect 4408 508 4442 542
rect 4958 508 4992 542
rect 5508 508 5542 542
rect 6058 508 6092 542
rect 6608 508 6642 542
rect 7158 508 7192 542
rect 7708 508 7742 542
rect 8258 508 8292 542
rect 8808 508 8842 542
rect 9358 508 9392 542
rect 9908 508 9942 542
rect 10458 508 10492 542
rect 11008 508 11042 542
rect 11558 508 11592 542
rect 12108 508 12142 542
rect 12658 508 12692 542
rect 13208 508 13242 542
rect 13758 508 13792 542
rect -542 -42 -508 -8
rect 8 -42 42 -8
rect 558 -42 592 -8
rect 1108 -42 1142 -8
rect 1658 -42 1692 -8
rect 2208 -42 2242 -8
rect 2758 -42 2792 -8
rect 3308 -42 3342 -8
rect 3858 -42 3892 -8
rect 4408 -42 4442 -8
rect 4958 -42 4992 -8
rect 5508 -42 5542 -8
rect 6058 -42 6092 -8
rect 6608 -42 6642 -8
rect 7158 -42 7192 -8
rect 7708 -42 7742 -8
rect 8258 -42 8292 -8
rect 8808 -42 8842 -8
rect 9358 -42 9392 -8
rect 9908 -42 9942 -8
rect 10458 -42 10492 -8
rect 11008 -42 11042 -8
rect 11558 -42 11592 -8
rect 12108 -42 12142 -8
rect 12658 -42 12692 -8
rect 13208 -42 13242 -8
rect 13758 -42 13792 -8
rect -542 -592 -508 -558
rect 8 -592 42 -558
rect 558 -592 592 -558
rect 1108 -592 1142 -558
rect 1658 -592 1692 -558
rect 2208 -592 2242 -558
rect 2758 -592 2792 -558
rect 3308 -592 3342 -558
rect 3858 -592 3892 -558
rect 4408 -592 4442 -558
rect 4958 -592 4992 -558
rect 5508 -592 5542 -558
rect 6058 -592 6092 -558
rect 6608 -592 6642 -558
rect 7158 -592 7192 -558
rect 7708 -592 7742 -558
rect 8258 -592 8292 -558
rect 8808 -592 8842 -558
rect 9358 -592 9392 -558
rect 9908 -592 9942 -558
rect 10458 -592 10492 -558
rect 11008 -592 11042 -558
rect 11558 -592 11592 -558
rect 12108 -592 12142 -558
rect 12658 -592 12692 -558
rect 13208 -592 13242 -558
rect 13758 -592 13792 -558
<< locali >>
rect -5525 18713 18775 18725
rect -5525 -5563 -5513 18713
rect -1537 14725 14787 14737
rect -1537 -1575 -1525 14725
rect -1025 14213 14275 14225
rect -1025 13217 -1013 14213
rect -17 13937 0 14213
rect 533 13937 550 14213
rect 1083 13937 1100 14213
rect 1633 13937 1650 14213
rect 2183 13937 2200 14213
rect 2733 13937 2750 14213
rect 3283 13937 3300 14213
rect 3833 13937 3850 14213
rect 4383 13937 4400 14213
rect 4933 13937 4950 14213
rect 5483 13937 5500 14213
rect 6033 13937 6050 14213
rect 6583 13937 6600 14213
rect 7133 13937 7150 14213
rect 7683 13937 7700 14213
rect 8233 13937 8250 14213
rect 8783 13937 8800 14213
rect 9333 13937 9350 14213
rect 9883 13937 9900 14213
rect 10433 13937 10450 14213
rect 10983 13937 11000 14213
rect 11533 13937 11550 14213
rect 12083 13937 12100 14213
rect 12633 13937 12650 14213
rect 13183 13937 13200 14213
rect -737 13925 13987 13937
rect -737 13217 -725 13925
rect -550 13742 -500 13750
rect -550 13708 -542 13742
rect -508 13708 -500 13742
rect -550 13700 -500 13708
rect 0 13742 50 13750
rect 0 13708 8 13742
rect 42 13708 50 13742
rect 0 13700 50 13708
rect 550 13742 600 13750
rect 550 13708 558 13742
rect 592 13708 600 13742
rect 550 13700 600 13708
rect 1100 13742 1150 13750
rect 1100 13708 1108 13742
rect 1142 13708 1150 13742
rect 1100 13700 1150 13708
rect 1650 13742 1700 13750
rect 1650 13708 1658 13742
rect 1692 13708 1700 13742
rect 1650 13700 1700 13708
rect 2200 13742 2250 13750
rect 2200 13708 2208 13742
rect 2242 13708 2250 13742
rect 2200 13700 2250 13708
rect 2750 13742 2800 13750
rect 2750 13708 2758 13742
rect 2792 13708 2800 13742
rect 2750 13700 2800 13708
rect 3300 13742 3350 13750
rect 3300 13708 3308 13742
rect 3342 13708 3350 13742
rect 3300 13700 3350 13708
rect 3850 13742 3900 13750
rect 3850 13708 3858 13742
rect 3892 13708 3900 13742
rect 3850 13700 3900 13708
rect 4400 13742 4450 13750
rect 4400 13708 4408 13742
rect 4442 13708 4450 13742
rect 4400 13700 4450 13708
rect 4950 13742 5000 13750
rect 4950 13708 4958 13742
rect 4992 13708 5000 13742
rect 4950 13700 5000 13708
rect 5500 13742 5550 13750
rect 5500 13708 5508 13742
rect 5542 13708 5550 13742
rect 5500 13700 5550 13708
rect 6050 13742 6100 13750
rect 6050 13708 6058 13742
rect 6092 13708 6100 13742
rect 6050 13700 6100 13708
rect 6600 13742 6650 13750
rect 6600 13708 6608 13742
rect 6642 13708 6650 13742
rect 6600 13700 6650 13708
rect 7150 13742 7200 13750
rect 7150 13708 7158 13742
rect 7192 13708 7200 13742
rect 7150 13700 7200 13708
rect 7700 13742 7750 13750
rect 7700 13708 7708 13742
rect 7742 13708 7750 13742
rect 7700 13700 7750 13708
rect 8250 13742 8300 13750
rect 8250 13708 8258 13742
rect 8292 13708 8300 13742
rect 8250 13700 8300 13708
rect 8800 13742 8850 13750
rect 8800 13708 8808 13742
rect 8842 13708 8850 13742
rect 8800 13700 8850 13708
rect 9350 13742 9400 13750
rect 9350 13708 9358 13742
rect 9392 13708 9400 13742
rect 9350 13700 9400 13708
rect 9900 13742 9950 13750
rect 9900 13708 9908 13742
rect 9942 13708 9950 13742
rect 9900 13700 9950 13708
rect 10450 13742 10500 13750
rect 10450 13708 10458 13742
rect 10492 13708 10500 13742
rect 10450 13700 10500 13708
rect 11000 13742 11050 13750
rect 11000 13708 11008 13742
rect 11042 13708 11050 13742
rect 11000 13700 11050 13708
rect 11550 13742 11600 13750
rect 11550 13708 11558 13742
rect 11592 13708 11600 13742
rect 11550 13700 11600 13708
rect 12100 13742 12150 13750
rect 12100 13708 12108 13742
rect 12142 13708 12150 13742
rect 12100 13700 12150 13708
rect 12650 13742 12700 13750
rect 12650 13708 12658 13742
rect 12692 13708 12700 13742
rect 12650 13700 12700 13708
rect 13200 13742 13250 13750
rect 13200 13708 13208 13742
rect 13242 13708 13250 13742
rect 13200 13700 13250 13708
rect 13750 13742 13800 13750
rect 13750 13708 13758 13742
rect 13792 13708 13800 13742
rect 13750 13700 13800 13708
rect 73 13671 527 13677
rect 1173 13671 1627 13677
rect 2273 13671 2727 13677
rect 3373 13671 3827 13677
rect 4473 13671 4927 13677
rect 5573 13671 6027 13677
rect 6673 13671 7127 13677
rect 7773 13671 8227 13677
rect 8873 13671 9327 13677
rect 9973 13671 10427 13677
rect 11073 13671 11527 13677
rect 12173 13671 12627 13677
rect 13273 13671 13727 13677
rect -23 13663 -6 13671
rect -64 13237 -23 13264
rect -64 13229 -6 13237
rect 56 13663 544 13671
rect 73 13615 527 13663
rect 73 13285 135 13615
rect 465 13285 527 13615
rect 73 13237 527 13285
rect 56 13229 544 13237
rect 606 13663 623 13671
rect 1077 13663 1094 13671
rect 623 13237 664 13264
rect 606 13229 664 13237
rect -64 13223 -29 13229
rect 73 13223 527 13229
rect 629 13223 664 13229
rect 1036 13237 1077 13264
rect 1036 13229 1094 13237
rect 1156 13663 1644 13671
rect 1173 13615 1627 13663
rect 1173 13285 1235 13615
rect 1565 13285 1627 13615
rect 1173 13237 1627 13285
rect 1156 13229 1644 13237
rect 1706 13663 1723 13671
rect 2177 13663 2194 13671
rect 1723 13237 1764 13264
rect 1706 13229 1764 13237
rect 1036 13223 1071 13229
rect 1173 13223 1627 13229
rect 1729 13223 1764 13229
rect 2136 13237 2177 13264
rect 2136 13229 2194 13237
rect 2256 13663 2744 13671
rect 2273 13615 2727 13663
rect 2273 13285 2335 13615
rect 2665 13285 2727 13615
rect 2273 13237 2727 13285
rect 2256 13229 2744 13237
rect 2806 13663 2823 13671
rect 3277 13663 3294 13671
rect 2823 13237 2864 13264
rect 2806 13229 2864 13237
rect 2136 13223 2171 13229
rect 2273 13223 2727 13229
rect 2829 13223 2864 13229
rect 3236 13237 3277 13264
rect 3236 13229 3294 13237
rect 3356 13663 3844 13671
rect 3373 13615 3827 13663
rect 3373 13285 3435 13615
rect 3765 13285 3827 13615
rect 3373 13237 3827 13285
rect 3356 13229 3844 13237
rect 3906 13663 3923 13671
rect 4377 13663 4394 13671
rect 3923 13237 3964 13264
rect 3906 13229 3964 13237
rect 3236 13223 3271 13229
rect 3373 13223 3827 13229
rect 3929 13223 3964 13229
rect 4336 13237 4377 13264
rect 4336 13229 4394 13237
rect 4456 13663 4944 13671
rect 4473 13615 4927 13663
rect 4473 13285 4535 13615
rect 4865 13285 4927 13615
rect 4473 13237 4927 13285
rect 4456 13229 4944 13237
rect 5006 13663 5023 13671
rect 5477 13663 5494 13671
rect 5023 13237 5064 13264
rect 5006 13229 5064 13237
rect 4336 13223 4371 13229
rect 4473 13223 4927 13229
rect 5029 13223 5064 13229
rect 5436 13237 5477 13264
rect 5436 13229 5494 13237
rect 5556 13663 6044 13671
rect 5573 13615 6027 13663
rect 5573 13285 5635 13615
rect 5965 13285 6027 13615
rect 5573 13237 6027 13285
rect 5556 13229 6044 13237
rect 6106 13663 6123 13671
rect 6577 13663 6594 13671
rect 6123 13237 6164 13264
rect 6106 13229 6164 13237
rect 5436 13223 5471 13229
rect 5573 13223 6027 13229
rect 6129 13223 6164 13229
rect 6536 13237 6577 13264
rect 6536 13229 6594 13237
rect 6656 13663 7144 13671
rect 6673 13615 7127 13663
rect 6673 13285 6735 13615
rect 7065 13285 7127 13615
rect 6673 13237 7127 13285
rect 6656 13229 7144 13237
rect 7206 13663 7223 13671
rect 7677 13663 7694 13671
rect 7223 13237 7264 13264
rect 7206 13229 7264 13237
rect 6536 13223 6571 13229
rect 6673 13223 7127 13229
rect 7229 13223 7264 13229
rect 7636 13237 7677 13264
rect 7636 13229 7694 13237
rect 7756 13663 8244 13671
rect 7773 13615 8227 13663
rect 7773 13285 7835 13615
rect 8165 13285 8227 13615
rect 7773 13237 8227 13285
rect 7756 13229 8244 13237
rect 8306 13663 8323 13671
rect 8777 13663 8794 13671
rect 8323 13237 8364 13264
rect 8306 13229 8364 13237
rect 7636 13223 7671 13229
rect 7773 13223 8227 13229
rect 8329 13223 8364 13229
rect 8736 13237 8777 13264
rect 8736 13229 8794 13237
rect 8856 13663 9344 13671
rect 8873 13615 9327 13663
rect 8873 13285 8935 13615
rect 9265 13285 9327 13615
rect 8873 13237 9327 13285
rect 8856 13229 9344 13237
rect 9406 13663 9423 13671
rect 9877 13663 9894 13671
rect 9423 13237 9464 13264
rect 9406 13229 9464 13237
rect 8736 13223 8771 13229
rect 8873 13223 9327 13229
rect 9429 13223 9464 13229
rect 9836 13237 9877 13264
rect 9836 13229 9894 13237
rect 9956 13663 10444 13671
rect 9973 13615 10427 13663
rect 9973 13285 10035 13615
rect 10365 13285 10427 13615
rect 9973 13237 10427 13285
rect 9956 13229 10444 13237
rect 10506 13663 10523 13671
rect 10977 13663 10994 13671
rect 10523 13237 10564 13264
rect 10506 13229 10564 13237
rect 9836 13223 9871 13229
rect 9973 13223 10427 13229
rect 10529 13223 10564 13229
rect 10936 13237 10977 13264
rect 10936 13229 10994 13237
rect 11056 13663 11544 13671
rect 11073 13615 11527 13663
rect 11073 13285 11135 13615
rect 11465 13285 11527 13615
rect 11073 13237 11527 13285
rect 11056 13229 11544 13237
rect 11606 13663 11623 13671
rect 12077 13663 12094 13671
rect 11623 13237 11664 13264
rect 11606 13229 11664 13237
rect 10936 13223 10971 13229
rect 11073 13223 11527 13229
rect 11629 13223 11664 13229
rect 12036 13237 12077 13264
rect 12036 13229 12094 13237
rect 12156 13663 12644 13671
rect 12173 13615 12627 13663
rect 12173 13285 12235 13615
rect 12565 13285 12627 13615
rect 12173 13237 12627 13285
rect 12156 13229 12644 13237
rect 12706 13663 12723 13671
rect 13177 13663 13194 13671
rect 12723 13237 12764 13264
rect 12706 13229 12764 13237
rect 12036 13223 12071 13229
rect 12173 13223 12627 13229
rect 12729 13223 12764 13229
rect 13136 13237 13177 13264
rect 13136 13229 13194 13237
rect 13256 13663 13727 13671
rect 13273 13615 13727 13663
rect 13273 13285 13335 13615
rect 13665 13285 13727 13615
rect 13273 13237 13727 13285
rect 13256 13229 13727 13237
rect 13136 13223 13171 13229
rect 13273 13223 13727 13229
rect -1025 13200 -725 13217
rect -471 13206 -463 13223
rect -37 13206 -29 13223
rect 79 13206 87 13223
rect 513 13206 521 13223
rect 629 13206 637 13223
rect 1063 13206 1071 13223
rect 1179 13206 1187 13223
rect 1613 13206 1621 13223
rect 1729 13206 1737 13223
rect 2163 13206 2171 13223
rect 2279 13206 2287 13223
rect 2713 13206 2721 13223
rect 2829 13206 2837 13223
rect 3263 13206 3271 13223
rect 3379 13206 3387 13223
rect 3813 13206 3821 13223
rect 3929 13206 3937 13223
rect 4363 13206 4371 13223
rect 4479 13206 4487 13223
rect 4913 13206 4921 13223
rect 5029 13206 5037 13223
rect 5463 13206 5471 13223
rect 5579 13206 5587 13223
rect 6013 13206 6021 13223
rect 6129 13206 6137 13223
rect 6563 13206 6571 13223
rect 6679 13206 6687 13223
rect 7113 13206 7121 13223
rect 7229 13206 7237 13223
rect 7663 13206 7671 13223
rect 7779 13206 7787 13223
rect 8213 13206 8221 13223
rect 8329 13206 8337 13223
rect 8763 13206 8771 13223
rect 8879 13206 8887 13223
rect 9313 13206 9321 13223
rect 9429 13206 9437 13223
rect 9863 13206 9871 13223
rect 9979 13206 9987 13223
rect 10413 13206 10421 13223
rect 10529 13206 10537 13223
rect 10963 13206 10971 13223
rect 11079 13206 11087 13223
rect 11513 13206 11521 13223
rect 11629 13206 11637 13223
rect 12063 13206 12071 13223
rect 12179 13206 12187 13223
rect 12613 13206 12621 13223
rect 12729 13206 12737 13223
rect 13163 13206 13171 13223
rect 13279 13206 13287 13223
rect 13713 13206 13721 13223
rect 13975 13217 13987 13925
rect 14263 13217 14275 14213
rect 13975 13200 14275 13217
rect -1025 12667 -1013 13200
rect -737 12667 -725 13200
rect -550 13192 -500 13200
rect -550 13158 -542 13192
rect -508 13158 -500 13192
rect -550 13150 -500 13158
rect 0 13192 50 13200
rect 0 13158 8 13192
rect 42 13158 50 13192
rect 0 13150 50 13158
rect 550 13192 600 13200
rect 550 13158 558 13192
rect 592 13158 600 13192
rect 550 13150 600 13158
rect 1100 13192 1150 13200
rect 1100 13158 1108 13192
rect 1142 13158 1150 13192
rect 1100 13150 1150 13158
rect 1650 13192 1700 13200
rect 1650 13158 1658 13192
rect 1692 13158 1700 13192
rect 1650 13150 1700 13158
rect 2200 13192 2250 13200
rect 2200 13158 2208 13192
rect 2242 13158 2250 13192
rect 2200 13150 2250 13158
rect 2750 13192 2800 13200
rect 2750 13158 2758 13192
rect 2792 13158 2800 13192
rect 2750 13150 2800 13158
rect 3300 13192 3350 13200
rect 3300 13158 3308 13192
rect 3342 13158 3350 13192
rect 3300 13150 3350 13158
rect 3850 13192 3900 13200
rect 3850 13158 3858 13192
rect 3892 13158 3900 13192
rect 3850 13150 3900 13158
rect 4400 13192 4450 13200
rect 4400 13158 4408 13192
rect 4442 13158 4450 13192
rect 4400 13150 4450 13158
rect 4950 13192 5000 13200
rect 4950 13158 4958 13192
rect 4992 13158 5000 13192
rect 4950 13150 5000 13158
rect 5500 13192 5550 13200
rect 5500 13158 5508 13192
rect 5542 13158 5550 13192
rect 5500 13150 5550 13158
rect 6050 13192 6100 13200
rect 6050 13158 6058 13192
rect 6092 13158 6100 13192
rect 6050 13150 6100 13158
rect 6600 13192 6650 13200
rect 6600 13158 6608 13192
rect 6642 13158 6650 13192
rect 6600 13150 6650 13158
rect 7150 13192 7200 13200
rect 7150 13158 7158 13192
rect 7192 13158 7200 13192
rect 7150 13150 7200 13158
rect 7700 13192 7750 13200
rect 7700 13158 7708 13192
rect 7742 13158 7750 13192
rect 7700 13150 7750 13158
rect 8250 13192 8300 13200
rect 8250 13158 8258 13192
rect 8292 13158 8300 13192
rect 8250 13150 8300 13158
rect 8800 13192 8850 13200
rect 8800 13158 8808 13192
rect 8842 13158 8850 13192
rect 8800 13150 8850 13158
rect 9350 13192 9400 13200
rect 9350 13158 9358 13192
rect 9392 13158 9400 13192
rect 9350 13150 9400 13158
rect 9900 13192 9950 13200
rect 9900 13158 9908 13192
rect 9942 13158 9950 13192
rect 9900 13150 9950 13158
rect 10450 13192 10500 13200
rect 10450 13158 10458 13192
rect 10492 13158 10500 13192
rect 10450 13150 10500 13158
rect 11000 13192 11050 13200
rect 11000 13158 11008 13192
rect 11042 13158 11050 13192
rect 11000 13150 11050 13158
rect 11550 13192 11600 13200
rect 11550 13158 11558 13192
rect 11592 13158 11600 13192
rect 11550 13150 11600 13158
rect 12100 13192 12150 13200
rect 12100 13158 12108 13192
rect 12142 13158 12150 13192
rect 12100 13150 12150 13158
rect 12650 13192 12700 13200
rect 12650 13158 12658 13192
rect 12692 13158 12700 13192
rect 12650 13150 12700 13158
rect 13200 13192 13250 13200
rect 13200 13158 13208 13192
rect 13242 13158 13250 13192
rect 13200 13150 13250 13158
rect 13750 13192 13800 13200
rect 13750 13158 13758 13192
rect 13792 13158 13800 13192
rect 13750 13150 13800 13158
rect -471 13127 -463 13144
rect -37 13127 -29 13144
rect 79 13127 87 13144
rect 513 13127 521 13144
rect 629 13127 637 13144
rect 1063 13127 1071 13144
rect 1179 13127 1187 13144
rect 1613 13127 1621 13144
rect 1729 13127 1737 13144
rect 2163 13127 2171 13144
rect 2279 13127 2287 13144
rect 2713 13127 2721 13144
rect 2829 13127 2837 13144
rect 3263 13127 3271 13144
rect 3379 13127 3387 13144
rect 3813 13127 3821 13144
rect 3929 13127 3937 13144
rect 4363 13127 4371 13144
rect 4479 13127 4487 13144
rect 4913 13127 4921 13144
rect 5029 13127 5037 13144
rect 5463 13127 5471 13144
rect 5579 13127 5587 13144
rect 6013 13127 6021 13144
rect 6129 13127 6137 13144
rect 6563 13127 6571 13144
rect 6679 13127 6687 13144
rect 7113 13127 7121 13144
rect 7229 13127 7237 13144
rect 7663 13127 7671 13144
rect 7779 13127 7787 13144
rect 8213 13127 8221 13144
rect 8329 13127 8337 13144
rect 8763 13127 8771 13144
rect 8879 13127 8887 13144
rect 9313 13127 9321 13144
rect 9429 13127 9437 13144
rect 9863 13127 9871 13144
rect 9979 13127 9987 13144
rect 10413 13127 10421 13144
rect 10529 13127 10537 13144
rect 10963 13127 10971 13144
rect 11079 13127 11087 13144
rect 11513 13127 11521 13144
rect 11629 13127 11637 13144
rect 12063 13127 12071 13144
rect 12179 13127 12187 13144
rect 12613 13127 12621 13144
rect 12729 13127 12737 13144
rect 13163 13127 13171 13144
rect 13279 13127 13287 13144
rect 13713 13127 13721 13144
rect -477 13121 -23 13127
rect 79 13121 114 13127
rect -477 13113 -6 13121
rect -477 13065 -23 13113
rect -477 12735 -415 13065
rect -85 12735 -23 13065
rect -477 12687 -23 12735
rect -477 12679 -6 12687
rect 56 13113 114 13121
rect 73 13086 114 13113
rect 486 13121 521 13127
rect 623 13121 1077 13127
rect 1179 13121 1214 13127
rect 486 13113 544 13121
rect 486 13086 527 13113
rect 73 12687 114 12714
rect 56 12679 114 12687
rect -477 12673 -23 12679
rect 79 12673 114 12679
rect 486 12687 527 12714
rect 486 12679 544 12687
rect 606 13113 1094 13121
rect 623 13065 1077 13113
rect 623 12735 685 13065
rect 1015 12735 1077 13065
rect 623 12687 1077 12735
rect 606 12679 1094 12687
rect 1156 13113 1214 13121
rect 1173 13086 1214 13113
rect 1586 13121 1621 13127
rect 1723 13121 2177 13127
rect 2279 13121 2314 13127
rect 1586 13113 1644 13121
rect 1586 13086 1627 13113
rect 1173 12687 1214 12714
rect 1156 12679 1214 12687
rect 486 12673 521 12679
rect 623 12673 1077 12679
rect 1179 12673 1214 12679
rect 1586 12687 1627 12714
rect 1586 12679 1644 12687
rect 1706 13113 2194 13121
rect 1723 13065 2177 13113
rect 1723 12735 1785 13065
rect 2115 12735 2177 13065
rect 1723 12687 2177 12735
rect 1706 12679 2194 12687
rect 2256 13113 2314 13121
rect 2273 13086 2314 13113
rect 2686 13121 2721 13127
rect 2823 13121 3277 13127
rect 3379 13121 3414 13127
rect 2686 13113 2744 13121
rect 2686 13086 2727 13113
rect 2273 12687 2314 12714
rect 2256 12679 2314 12687
rect 1586 12673 1621 12679
rect 1723 12673 2177 12679
rect 2279 12673 2314 12679
rect 2686 12687 2727 12714
rect 2686 12679 2744 12687
rect 2806 13113 3294 13121
rect 2823 13065 3277 13113
rect 2823 12735 2885 13065
rect 3215 12735 3277 13065
rect 2823 12687 3277 12735
rect 2806 12679 3294 12687
rect 3356 13113 3414 13121
rect 3373 13086 3414 13113
rect 3786 13121 3821 13127
rect 3923 13121 4377 13127
rect 4479 13121 4514 13127
rect 3786 13113 3844 13121
rect 3786 13086 3827 13113
rect 3373 12687 3414 12714
rect 3356 12679 3414 12687
rect 2686 12673 2721 12679
rect 2823 12673 3277 12679
rect 3379 12673 3414 12679
rect 3786 12687 3827 12714
rect 3786 12679 3844 12687
rect 3906 13113 4394 13121
rect 3923 13065 4377 13113
rect 3923 12735 3985 13065
rect 4315 12735 4377 13065
rect 3923 12687 4377 12735
rect 3906 12679 4394 12687
rect 4456 13113 4514 13121
rect 4473 13086 4514 13113
rect 4886 13121 4921 13127
rect 5023 13121 5477 13127
rect 5579 13121 5614 13127
rect 4886 13113 4944 13121
rect 4886 13086 4927 13113
rect 4473 12687 4514 12714
rect 4456 12679 4514 12687
rect 3786 12673 3821 12679
rect 3923 12673 4377 12679
rect 4479 12673 4514 12679
rect 4886 12687 4927 12714
rect 4886 12679 4944 12687
rect 5006 13113 5494 13121
rect 5023 13065 5477 13113
rect 5023 12735 5085 13065
rect 5415 12735 5477 13065
rect 5023 12687 5477 12735
rect 5006 12679 5494 12687
rect 5556 13113 5614 13121
rect 5573 13086 5614 13113
rect 5986 13121 6021 13127
rect 6123 13121 6577 13127
rect 6679 13121 6714 13127
rect 5986 13113 6044 13121
rect 5986 13086 6027 13113
rect 5573 12687 5614 12714
rect 5556 12679 5614 12687
rect 4886 12673 4921 12679
rect 5023 12673 5477 12679
rect 5579 12673 5614 12679
rect 5986 12687 6027 12714
rect 5986 12679 6044 12687
rect 6106 13113 6594 13121
rect 6123 13065 6577 13113
rect 6123 12735 6185 13065
rect 6515 12735 6577 13065
rect 6123 12687 6577 12735
rect 6106 12679 6594 12687
rect 6656 13113 6714 13121
rect 6673 13086 6714 13113
rect 7086 13121 7121 13127
rect 7223 13121 7677 13127
rect 7779 13121 7814 13127
rect 7086 13113 7144 13121
rect 7086 13086 7127 13113
rect 6673 12687 6714 12714
rect 6656 12679 6714 12687
rect 5986 12673 6021 12679
rect 6123 12673 6577 12679
rect 6679 12673 6714 12679
rect 7086 12687 7127 12714
rect 7086 12679 7144 12687
rect 7206 13113 7694 13121
rect 7223 13065 7677 13113
rect 7223 12735 7285 13065
rect 7615 12735 7677 13065
rect 7223 12687 7677 12735
rect 7206 12679 7694 12687
rect 7756 13113 7814 13121
rect 7773 13086 7814 13113
rect 8186 13121 8221 13127
rect 8323 13121 8777 13127
rect 8879 13121 8914 13127
rect 8186 13113 8244 13121
rect 8186 13086 8227 13113
rect 7773 12687 7814 12714
rect 7756 12679 7814 12687
rect 7086 12673 7121 12679
rect 7223 12673 7677 12679
rect 7779 12673 7814 12679
rect 8186 12687 8227 12714
rect 8186 12679 8244 12687
rect 8306 13113 8794 13121
rect 8323 13065 8777 13113
rect 8323 12735 8385 13065
rect 8715 12735 8777 13065
rect 8323 12687 8777 12735
rect 8306 12679 8794 12687
rect 8856 13113 8914 13121
rect 8873 13086 8914 13113
rect 9286 13121 9321 13127
rect 9423 13121 9877 13127
rect 9979 13121 10014 13127
rect 9286 13113 9344 13121
rect 9286 13086 9327 13113
rect 8873 12687 8914 12714
rect 8856 12679 8914 12687
rect 8186 12673 8221 12679
rect 8323 12673 8777 12679
rect 8879 12673 8914 12679
rect 9286 12687 9327 12714
rect 9286 12679 9344 12687
rect 9406 13113 9894 13121
rect 9423 13065 9877 13113
rect 9423 12735 9485 13065
rect 9815 12735 9877 13065
rect 9423 12687 9877 12735
rect 9406 12679 9894 12687
rect 9956 13113 10014 13121
rect 9973 13086 10014 13113
rect 10386 13121 10421 13127
rect 10523 13121 10977 13127
rect 11079 13121 11114 13127
rect 10386 13113 10444 13121
rect 10386 13086 10427 13113
rect 9973 12687 10014 12714
rect 9956 12679 10014 12687
rect 9286 12673 9321 12679
rect 9423 12673 9877 12679
rect 9979 12673 10014 12679
rect 10386 12687 10427 12714
rect 10386 12679 10444 12687
rect 10506 13113 10994 13121
rect 10523 13065 10977 13113
rect 10523 12735 10585 13065
rect 10915 12735 10977 13065
rect 10523 12687 10977 12735
rect 10506 12679 10994 12687
rect 11056 13113 11114 13121
rect 11073 13086 11114 13113
rect 11486 13121 11521 13127
rect 11623 13121 12077 13127
rect 12179 13121 12214 13127
rect 11486 13113 11544 13121
rect 11486 13086 11527 13113
rect 11073 12687 11114 12714
rect 11056 12679 11114 12687
rect 10386 12673 10421 12679
rect 10523 12673 10977 12679
rect 11079 12673 11114 12679
rect 11486 12687 11527 12714
rect 11486 12679 11544 12687
rect 11606 13113 12094 13121
rect 11623 13065 12077 13113
rect 11623 12735 11685 13065
rect 12015 12735 12077 13065
rect 11623 12687 12077 12735
rect 11606 12679 12094 12687
rect 12156 13113 12214 13121
rect 12173 13086 12214 13113
rect 12586 13121 12621 13127
rect 12723 13121 13177 13127
rect 13279 13121 13314 13127
rect 12586 13113 12644 13121
rect 12586 13086 12627 13113
rect 12173 12687 12214 12714
rect 12156 12679 12214 12687
rect 11486 12673 11521 12679
rect 11623 12673 12077 12679
rect 12179 12673 12214 12679
rect 12586 12687 12627 12714
rect 12586 12679 12644 12687
rect 12706 13113 13194 13121
rect 12723 13065 13177 13113
rect 12723 12735 12785 13065
rect 13115 12735 13177 13065
rect 12723 12687 13177 12735
rect 12706 12679 13194 12687
rect 13256 13113 13314 13121
rect 13273 13086 13314 13113
rect 13273 12687 13314 12714
rect 13256 12679 13314 12687
rect 12586 12673 12621 12679
rect 12723 12673 13177 12679
rect 13279 12673 13314 12679
rect -1025 12650 -725 12667
rect -471 12656 -463 12673
rect -37 12656 -29 12673
rect 79 12656 87 12673
rect 513 12656 521 12673
rect 629 12656 637 12673
rect 1063 12656 1071 12673
rect 1179 12656 1187 12673
rect 1613 12656 1621 12673
rect 1729 12656 1737 12673
rect 2163 12656 2171 12673
rect 2279 12656 2287 12673
rect 2713 12656 2721 12673
rect 2829 12656 2837 12673
rect 3263 12656 3271 12673
rect 3379 12656 3387 12673
rect 3813 12656 3821 12673
rect 3929 12656 3937 12673
rect 4363 12656 4371 12673
rect 4479 12656 4487 12673
rect 4913 12656 4921 12673
rect 5029 12656 5037 12673
rect 5463 12656 5471 12673
rect 5579 12656 5587 12673
rect 6013 12656 6021 12673
rect 6129 12656 6137 12673
rect 6563 12656 6571 12673
rect 6679 12656 6687 12673
rect 7113 12656 7121 12673
rect 7229 12656 7237 12673
rect 7663 12656 7671 12673
rect 7779 12656 7787 12673
rect 8213 12656 8221 12673
rect 8329 12656 8337 12673
rect 8763 12656 8771 12673
rect 8879 12656 8887 12673
rect 9313 12656 9321 12673
rect 9429 12656 9437 12673
rect 9863 12656 9871 12673
rect 9979 12656 9987 12673
rect 10413 12656 10421 12673
rect 10529 12656 10537 12673
rect 10963 12656 10971 12673
rect 11079 12656 11087 12673
rect 11513 12656 11521 12673
rect 11629 12656 11637 12673
rect 12063 12656 12071 12673
rect 12179 12656 12187 12673
rect 12613 12656 12621 12673
rect 12729 12656 12737 12673
rect 13163 12656 13171 12673
rect 13279 12656 13287 12673
rect 13713 12656 13721 12673
rect 13975 12669 13987 13200
rect 14263 12669 14275 13200
rect 13975 12650 14275 12669
rect -1025 12117 -1013 12650
rect -737 12117 -725 12650
rect -550 12642 -500 12650
rect -550 12608 -542 12642
rect -508 12608 -500 12642
rect -550 12600 -500 12608
rect 0 12642 50 12650
rect 0 12608 8 12642
rect 42 12608 50 12642
rect 0 12600 50 12608
rect 550 12642 600 12650
rect 550 12608 558 12642
rect 592 12608 600 12642
rect 550 12600 600 12608
rect 1100 12642 1150 12650
rect 1100 12608 1108 12642
rect 1142 12608 1150 12642
rect 1100 12600 1150 12608
rect 1650 12642 1700 12650
rect 1650 12608 1658 12642
rect 1692 12608 1700 12642
rect 1650 12600 1700 12608
rect 2200 12642 2250 12650
rect 2200 12608 2208 12642
rect 2242 12608 2250 12642
rect 2200 12600 2250 12608
rect 2750 12642 2800 12650
rect 2750 12608 2758 12642
rect 2792 12608 2800 12642
rect 2750 12600 2800 12608
rect 3300 12642 3350 12650
rect 3300 12608 3308 12642
rect 3342 12608 3350 12642
rect 3300 12600 3350 12608
rect 3850 12642 3900 12650
rect 3850 12608 3858 12642
rect 3892 12608 3900 12642
rect 3850 12600 3900 12608
rect 4400 12642 4450 12650
rect 4400 12608 4408 12642
rect 4442 12608 4450 12642
rect 4400 12600 4450 12608
rect 4950 12642 5000 12650
rect 4950 12608 4958 12642
rect 4992 12608 5000 12642
rect 4950 12600 5000 12608
rect 5500 12642 5550 12650
rect 5500 12608 5508 12642
rect 5542 12608 5550 12642
rect 5500 12600 5550 12608
rect 6050 12642 6100 12650
rect 6050 12608 6058 12642
rect 6092 12608 6100 12642
rect 6050 12600 6100 12608
rect 6600 12642 6650 12650
rect 6600 12608 6608 12642
rect 6642 12608 6650 12642
rect 6600 12600 6650 12608
rect 7150 12642 7200 12650
rect 7150 12608 7158 12642
rect 7192 12608 7200 12642
rect 7150 12600 7200 12608
rect 7700 12642 7750 12650
rect 7700 12608 7708 12642
rect 7742 12608 7750 12642
rect 7700 12600 7750 12608
rect 8250 12642 8300 12650
rect 8250 12608 8258 12642
rect 8292 12608 8300 12642
rect 8250 12600 8300 12608
rect 8800 12642 8850 12650
rect 8800 12608 8808 12642
rect 8842 12608 8850 12642
rect 8800 12600 8850 12608
rect 9350 12642 9400 12650
rect 9350 12608 9358 12642
rect 9392 12608 9400 12642
rect 9350 12600 9400 12608
rect 9900 12642 9950 12650
rect 9900 12608 9908 12642
rect 9942 12608 9950 12642
rect 9900 12600 9950 12608
rect 10450 12642 10500 12650
rect 10450 12608 10458 12642
rect 10492 12608 10500 12642
rect 10450 12600 10500 12608
rect 11000 12642 11050 12650
rect 11000 12608 11008 12642
rect 11042 12608 11050 12642
rect 11000 12600 11050 12608
rect 11550 12642 11600 12650
rect 11550 12608 11558 12642
rect 11592 12608 11600 12642
rect 11550 12600 11600 12608
rect 12100 12642 12150 12650
rect 12100 12608 12108 12642
rect 12142 12608 12150 12642
rect 12100 12600 12150 12608
rect 12650 12642 12700 12650
rect 12650 12608 12658 12642
rect 12692 12608 12700 12642
rect 12650 12600 12700 12608
rect 13200 12642 13250 12650
rect 13200 12608 13208 12642
rect 13242 12608 13250 12642
rect 13200 12600 13250 12608
rect 13750 12642 13800 12650
rect 13750 12608 13758 12642
rect 13792 12608 13800 12642
rect 13750 12600 13800 12608
rect -471 12577 -463 12594
rect -37 12577 -29 12594
rect 79 12577 87 12594
rect 513 12577 521 12594
rect 629 12577 637 12594
rect 1063 12577 1071 12594
rect 1179 12577 1187 12594
rect 1613 12577 1621 12594
rect 1729 12577 1737 12594
rect 2163 12577 2171 12594
rect 2279 12577 2287 12594
rect 2713 12577 2721 12594
rect 2829 12577 2837 12594
rect 3263 12577 3271 12594
rect 3379 12577 3387 12594
rect 3813 12577 3821 12594
rect 3929 12577 3937 12594
rect 4363 12577 4371 12594
rect 4479 12577 4487 12594
rect 4913 12577 4921 12594
rect 5029 12577 5037 12594
rect 5463 12577 5471 12594
rect 5579 12577 5587 12594
rect 6013 12577 6021 12594
rect 6129 12577 6137 12594
rect 6563 12577 6571 12594
rect 6679 12577 6687 12594
rect 7113 12577 7121 12594
rect 7229 12577 7237 12594
rect 7663 12577 7671 12594
rect 7779 12577 7787 12594
rect 8213 12577 8221 12594
rect 8329 12577 8337 12594
rect 8763 12577 8771 12594
rect 8879 12577 8887 12594
rect 9313 12577 9321 12594
rect 9429 12577 9437 12594
rect 9863 12577 9871 12594
rect 9979 12577 9987 12594
rect 10413 12577 10421 12594
rect 10529 12577 10537 12594
rect 10963 12577 10971 12594
rect 11079 12577 11087 12594
rect 11513 12577 11521 12594
rect 11629 12577 11637 12594
rect 12063 12577 12071 12594
rect 12179 12577 12187 12594
rect 12613 12577 12621 12594
rect 12729 12577 12737 12594
rect 13163 12577 13171 12594
rect 13279 12577 13287 12594
rect 13713 12577 13721 12594
rect -64 12571 -29 12577
rect 73 12571 527 12577
rect 629 12571 664 12577
rect -64 12563 -6 12571
rect -64 12536 -23 12563
rect -64 12137 -23 12164
rect -64 12129 -6 12137
rect 56 12563 544 12571
rect 73 12515 527 12563
rect 73 12185 135 12515
rect 465 12185 527 12515
rect 73 12137 527 12185
rect 56 12129 544 12137
rect 606 12563 664 12571
rect 623 12536 664 12563
rect 1036 12571 1071 12577
rect 1173 12571 1627 12577
rect 1729 12571 1764 12577
rect 1036 12563 1094 12571
rect 1036 12536 1077 12563
rect 623 12137 664 12164
rect 606 12129 664 12137
rect -64 12123 -29 12129
rect 73 12123 527 12129
rect 629 12123 664 12129
rect 1036 12137 1077 12164
rect 1036 12129 1094 12137
rect 1156 12563 1644 12571
rect 1173 12515 1627 12563
rect 1173 12185 1235 12515
rect 1565 12185 1627 12515
rect 1173 12137 1627 12185
rect 1156 12129 1644 12137
rect 1706 12563 1764 12571
rect 1723 12536 1764 12563
rect 2136 12571 2171 12577
rect 2273 12571 2727 12577
rect 2829 12571 2864 12577
rect 2136 12563 2194 12571
rect 2136 12536 2177 12563
rect 1723 12137 1764 12164
rect 1706 12129 1764 12137
rect 1036 12123 1071 12129
rect 1173 12123 1627 12129
rect 1729 12123 1764 12129
rect 2136 12137 2177 12164
rect 2136 12129 2194 12137
rect 2256 12563 2744 12571
rect 2273 12515 2727 12563
rect 2273 12185 2335 12515
rect 2665 12185 2727 12515
rect 2273 12137 2727 12185
rect 2256 12129 2744 12137
rect 2806 12563 2864 12571
rect 2823 12536 2864 12563
rect 3236 12571 3271 12577
rect 3373 12571 3827 12577
rect 3929 12571 3964 12577
rect 3236 12563 3294 12571
rect 3236 12536 3277 12563
rect 2823 12137 2864 12164
rect 2806 12129 2864 12137
rect 2136 12123 2171 12129
rect 2273 12123 2727 12129
rect 2829 12123 2864 12129
rect 3236 12137 3277 12164
rect 3236 12129 3294 12137
rect 3356 12563 3844 12571
rect 3373 12515 3827 12563
rect 3373 12185 3435 12515
rect 3765 12185 3827 12515
rect 3373 12137 3827 12185
rect 3356 12129 3844 12137
rect 3906 12563 3964 12571
rect 3923 12536 3964 12563
rect 4336 12571 4371 12577
rect 4473 12571 4927 12577
rect 5029 12571 5064 12577
rect 4336 12563 4394 12571
rect 4336 12536 4377 12563
rect 3923 12137 3964 12164
rect 3906 12129 3964 12137
rect 3236 12123 3271 12129
rect 3373 12123 3827 12129
rect 3929 12123 3964 12129
rect 4336 12137 4377 12164
rect 4336 12129 4394 12137
rect 4456 12563 4944 12571
rect 4473 12515 4927 12563
rect 4473 12185 4535 12515
rect 4865 12185 4927 12515
rect 4473 12137 4927 12185
rect 4456 12129 4944 12137
rect 5006 12563 5064 12571
rect 5023 12536 5064 12563
rect 5436 12571 5471 12577
rect 5573 12571 6027 12577
rect 6129 12571 6164 12577
rect 5436 12563 5494 12571
rect 5436 12536 5477 12563
rect 5023 12137 5064 12164
rect 5006 12129 5064 12137
rect 4336 12123 4371 12129
rect 4473 12123 4927 12129
rect 5029 12123 5064 12129
rect 5436 12137 5477 12164
rect 5436 12129 5494 12137
rect 5556 12563 6044 12571
rect 5573 12515 6027 12563
rect 5573 12185 5635 12515
rect 5965 12185 6027 12515
rect 5573 12137 6027 12185
rect 5556 12129 6044 12137
rect 6106 12563 6164 12571
rect 6123 12536 6164 12563
rect 6536 12571 6571 12577
rect 6673 12571 7127 12577
rect 7229 12571 7264 12577
rect 6536 12563 6594 12571
rect 6536 12536 6577 12563
rect 6123 12137 6164 12164
rect 6106 12129 6164 12137
rect 5436 12123 5471 12129
rect 5573 12123 6027 12129
rect 6129 12123 6164 12129
rect 6536 12137 6577 12164
rect 6536 12129 6594 12137
rect 6656 12563 7144 12571
rect 6673 12515 7127 12563
rect 6673 12185 6735 12515
rect 7065 12185 7127 12515
rect 6673 12137 7127 12185
rect 6656 12129 7144 12137
rect 7206 12563 7264 12571
rect 7223 12536 7264 12563
rect 7636 12571 7671 12577
rect 7773 12571 8227 12577
rect 8329 12571 8364 12577
rect 7636 12563 7694 12571
rect 7636 12536 7677 12563
rect 7223 12137 7264 12164
rect 7206 12129 7264 12137
rect 6536 12123 6571 12129
rect 6673 12123 7127 12129
rect 7229 12123 7264 12129
rect 7636 12137 7677 12164
rect 7636 12129 7694 12137
rect 7756 12563 8244 12571
rect 7773 12515 8227 12563
rect 7773 12185 7835 12515
rect 8165 12185 8227 12515
rect 7773 12137 8227 12185
rect 7756 12129 8244 12137
rect 8306 12563 8364 12571
rect 8323 12536 8364 12563
rect 8736 12571 8771 12577
rect 8873 12571 9327 12577
rect 9429 12571 9464 12577
rect 8736 12563 8794 12571
rect 8736 12536 8777 12563
rect 8323 12137 8364 12164
rect 8306 12129 8364 12137
rect 7636 12123 7671 12129
rect 7773 12123 8227 12129
rect 8329 12123 8364 12129
rect 8736 12137 8777 12164
rect 8736 12129 8794 12137
rect 8856 12563 9344 12571
rect 8873 12515 9327 12563
rect 8873 12185 8935 12515
rect 9265 12185 9327 12515
rect 8873 12137 9327 12185
rect 8856 12129 9344 12137
rect 9406 12563 9464 12571
rect 9423 12536 9464 12563
rect 9836 12571 9871 12577
rect 9973 12571 10427 12577
rect 10529 12571 10564 12577
rect 9836 12563 9894 12571
rect 9836 12536 9877 12563
rect 9423 12137 9464 12164
rect 9406 12129 9464 12137
rect 8736 12123 8771 12129
rect 8873 12123 9327 12129
rect 9429 12123 9464 12129
rect 9836 12137 9877 12164
rect 9836 12129 9894 12137
rect 9956 12563 10444 12571
rect 9973 12515 10427 12563
rect 9973 12185 10035 12515
rect 10365 12185 10427 12515
rect 9973 12137 10427 12185
rect 9956 12129 10444 12137
rect 10506 12563 10564 12571
rect 10523 12536 10564 12563
rect 10936 12571 10971 12577
rect 11073 12571 11527 12577
rect 11629 12571 11664 12577
rect 10936 12563 10994 12571
rect 10936 12536 10977 12563
rect 10523 12137 10564 12164
rect 10506 12129 10564 12137
rect 9836 12123 9871 12129
rect 9973 12123 10427 12129
rect 10529 12123 10564 12129
rect 10936 12137 10977 12164
rect 10936 12129 10994 12137
rect 11056 12563 11544 12571
rect 11073 12515 11527 12563
rect 11073 12185 11135 12515
rect 11465 12185 11527 12515
rect 11073 12137 11527 12185
rect 11056 12129 11544 12137
rect 11606 12563 11664 12571
rect 11623 12536 11664 12563
rect 12036 12571 12071 12577
rect 12173 12571 12627 12577
rect 12729 12571 12764 12577
rect 12036 12563 12094 12571
rect 12036 12536 12077 12563
rect 11623 12137 11664 12164
rect 11606 12129 11664 12137
rect 10936 12123 10971 12129
rect 11073 12123 11527 12129
rect 11629 12123 11664 12129
rect 12036 12137 12077 12164
rect 12036 12129 12094 12137
rect 12156 12563 12644 12571
rect 12173 12515 12627 12563
rect 12173 12185 12235 12515
rect 12565 12185 12627 12515
rect 12173 12137 12627 12185
rect 12156 12129 12644 12137
rect 12706 12563 12764 12571
rect 12723 12536 12764 12563
rect 13136 12571 13171 12577
rect 13273 12571 13727 12577
rect 13136 12563 13194 12571
rect 13136 12536 13177 12563
rect 12723 12137 12764 12164
rect 12706 12129 12764 12137
rect 12036 12123 12071 12129
rect 12173 12123 12627 12129
rect 12729 12123 12764 12129
rect 13136 12137 13177 12164
rect 13136 12129 13194 12137
rect 13256 12563 13727 12571
rect 13273 12515 13727 12563
rect 13273 12185 13335 12515
rect 13665 12185 13727 12515
rect 13273 12137 13727 12185
rect 13256 12129 13727 12137
rect 13136 12123 13171 12129
rect 13273 12123 13727 12129
rect -1025 12100 -725 12117
rect -471 12106 -463 12123
rect -37 12106 -29 12123
rect 79 12106 87 12123
rect 513 12106 521 12123
rect 629 12106 637 12123
rect 1063 12106 1071 12123
rect 1179 12106 1187 12123
rect 1613 12106 1621 12123
rect 1729 12106 1737 12123
rect 2163 12106 2171 12123
rect 2279 12106 2287 12123
rect 2713 12106 2721 12123
rect 2829 12106 2837 12123
rect 3263 12106 3271 12123
rect 3379 12106 3387 12123
rect 3813 12106 3821 12123
rect 3929 12106 3937 12123
rect 4363 12106 4371 12123
rect 4479 12106 4487 12123
rect 4913 12106 4921 12123
rect 5029 12106 5037 12123
rect 5463 12106 5471 12123
rect 5579 12106 5587 12123
rect 6013 12106 6021 12123
rect 6129 12106 6137 12123
rect 6563 12106 6571 12123
rect 6679 12106 6687 12123
rect 7113 12106 7121 12123
rect 7229 12106 7237 12123
rect 7663 12106 7671 12123
rect 7779 12106 7787 12123
rect 8213 12106 8221 12123
rect 8329 12106 8337 12123
rect 8763 12106 8771 12123
rect 8879 12106 8887 12123
rect 9313 12106 9321 12123
rect 9429 12106 9437 12123
rect 9863 12106 9871 12123
rect 9979 12106 9987 12123
rect 10413 12106 10421 12123
rect 10529 12106 10537 12123
rect 10963 12106 10971 12123
rect 11079 12106 11087 12123
rect 11513 12106 11521 12123
rect 11629 12106 11637 12123
rect 12063 12106 12071 12123
rect 12179 12106 12187 12123
rect 12613 12106 12621 12123
rect 12729 12106 12737 12123
rect 13163 12106 13171 12123
rect 13279 12106 13287 12123
rect 13713 12106 13721 12123
rect 13975 12117 13987 12650
rect 14263 12117 14275 12650
rect 13975 12100 14275 12117
rect -1025 11567 -1013 12100
rect -737 11567 -725 12100
rect -550 12092 -500 12100
rect -550 12058 -542 12092
rect -508 12058 -500 12092
rect -550 12050 -500 12058
rect 0 12092 50 12100
rect 0 12058 8 12092
rect 42 12058 50 12092
rect 0 12050 50 12058
rect 550 12092 600 12100
rect 550 12058 558 12092
rect 592 12058 600 12092
rect 550 12050 600 12058
rect 1100 12092 1150 12100
rect 1100 12058 1108 12092
rect 1142 12058 1150 12092
rect 1100 12050 1150 12058
rect 1650 12092 1700 12100
rect 1650 12058 1658 12092
rect 1692 12058 1700 12092
rect 1650 12050 1700 12058
rect 2200 12092 2250 12100
rect 2200 12058 2208 12092
rect 2242 12058 2250 12092
rect 2200 12050 2250 12058
rect 2750 12092 2800 12100
rect 2750 12058 2758 12092
rect 2792 12058 2800 12092
rect 2750 12050 2800 12058
rect 3300 12092 3350 12100
rect 3300 12058 3308 12092
rect 3342 12058 3350 12092
rect 3300 12050 3350 12058
rect 3850 12092 3900 12100
rect 3850 12058 3858 12092
rect 3892 12058 3900 12092
rect 3850 12050 3900 12058
rect 4400 12092 4450 12100
rect 4400 12058 4408 12092
rect 4442 12058 4450 12092
rect 4400 12050 4450 12058
rect 4950 12092 5000 12100
rect 4950 12058 4958 12092
rect 4992 12058 5000 12092
rect 4950 12050 5000 12058
rect 5500 12092 5550 12100
rect 5500 12058 5508 12092
rect 5542 12058 5550 12092
rect 5500 12050 5550 12058
rect 6050 12092 6100 12100
rect 6050 12058 6058 12092
rect 6092 12058 6100 12092
rect 6050 12050 6100 12058
rect 6600 12092 6650 12100
rect 6600 12058 6608 12092
rect 6642 12058 6650 12092
rect 6600 12050 6650 12058
rect 7150 12092 7200 12100
rect 7150 12058 7158 12092
rect 7192 12058 7200 12092
rect 7150 12050 7200 12058
rect 7700 12092 7750 12100
rect 7700 12058 7708 12092
rect 7742 12058 7750 12092
rect 7700 12050 7750 12058
rect 8250 12092 8300 12100
rect 8250 12058 8258 12092
rect 8292 12058 8300 12092
rect 8250 12050 8300 12058
rect 8800 12092 8850 12100
rect 8800 12058 8808 12092
rect 8842 12058 8850 12092
rect 8800 12050 8850 12058
rect 9350 12092 9400 12100
rect 9350 12058 9358 12092
rect 9392 12058 9400 12092
rect 9350 12050 9400 12058
rect 9900 12092 9950 12100
rect 9900 12058 9908 12092
rect 9942 12058 9950 12092
rect 9900 12050 9950 12058
rect 10450 12092 10500 12100
rect 10450 12058 10458 12092
rect 10492 12058 10500 12092
rect 10450 12050 10500 12058
rect 11000 12092 11050 12100
rect 11000 12058 11008 12092
rect 11042 12058 11050 12092
rect 11000 12050 11050 12058
rect 11550 12092 11600 12100
rect 11550 12058 11558 12092
rect 11592 12058 11600 12092
rect 11550 12050 11600 12058
rect 12100 12092 12150 12100
rect 12100 12058 12108 12092
rect 12142 12058 12150 12092
rect 12100 12050 12150 12058
rect 12650 12092 12700 12100
rect 12650 12058 12658 12092
rect 12692 12058 12700 12092
rect 12650 12050 12700 12058
rect 13200 12092 13250 12100
rect 13200 12058 13208 12092
rect 13242 12058 13250 12092
rect 13200 12050 13250 12058
rect 13750 12092 13800 12100
rect 13750 12058 13758 12092
rect 13792 12058 13800 12092
rect 13750 12050 13800 12058
rect -471 12027 -463 12044
rect -37 12027 -29 12044
rect 79 12027 87 12044
rect 513 12027 521 12044
rect 629 12027 637 12044
rect 1063 12027 1071 12044
rect 1179 12027 1187 12044
rect 1613 12027 1621 12044
rect 1729 12027 1737 12044
rect 2163 12027 2171 12044
rect 2279 12027 2287 12044
rect 2713 12027 2721 12044
rect 2829 12027 2837 12044
rect 3263 12027 3271 12044
rect 3379 12027 3387 12044
rect 3813 12027 3821 12044
rect 3929 12027 3937 12044
rect 4363 12027 4371 12044
rect 4479 12027 4487 12044
rect 4913 12027 4921 12044
rect 5029 12027 5037 12044
rect 5463 12027 5471 12044
rect 5579 12027 5587 12044
rect 6013 12027 6021 12044
rect 6129 12027 6137 12044
rect 6563 12027 6571 12044
rect 6679 12027 6687 12044
rect 7113 12027 7121 12044
rect 7229 12027 7237 12044
rect 7663 12027 7671 12044
rect 7779 12027 7787 12044
rect 8213 12027 8221 12044
rect 8329 12027 8337 12044
rect 8763 12027 8771 12044
rect 8879 12027 8887 12044
rect 9313 12027 9321 12044
rect 9429 12027 9437 12044
rect 9863 12027 9871 12044
rect 9979 12027 9987 12044
rect 10413 12027 10421 12044
rect 10529 12027 10537 12044
rect 10963 12027 10971 12044
rect 11079 12027 11087 12044
rect 11513 12027 11521 12044
rect 11629 12027 11637 12044
rect 12063 12027 12071 12044
rect 12179 12027 12187 12044
rect 12613 12027 12621 12044
rect 12729 12027 12737 12044
rect 13163 12027 13171 12044
rect 13279 12027 13287 12044
rect 13713 12027 13721 12044
rect -477 12021 -23 12027
rect 79 12021 114 12027
rect -477 12013 -6 12021
rect -477 11965 -23 12013
rect -477 11635 -415 11965
rect -85 11635 -23 11965
rect -477 11587 -23 11635
rect -477 11579 -6 11587
rect 56 12013 114 12021
rect 73 11986 114 12013
rect 486 12021 521 12027
rect 623 12021 1077 12027
rect 1179 12021 1214 12027
rect 486 12013 544 12021
rect 486 11986 527 12013
rect 73 11587 114 11614
rect 56 11579 114 11587
rect -477 11573 -23 11579
rect 79 11573 114 11579
rect 486 11587 527 11614
rect 486 11579 544 11587
rect 606 12013 1094 12021
rect 623 11965 1077 12013
rect 623 11635 685 11965
rect 1015 11635 1077 11965
rect 623 11587 1077 11635
rect 606 11579 1094 11587
rect 1156 12013 1214 12021
rect 1173 11986 1214 12013
rect 1586 12021 1621 12027
rect 1723 12021 2177 12027
rect 2279 12021 2314 12027
rect 1586 12013 1644 12021
rect 1586 11986 1627 12013
rect 1173 11587 1214 11614
rect 1156 11579 1214 11587
rect 486 11573 521 11579
rect 623 11573 1077 11579
rect 1179 11573 1214 11579
rect 1586 11587 1627 11614
rect 1586 11579 1644 11587
rect 1706 12013 2194 12021
rect 1723 11965 2177 12013
rect 1723 11635 1785 11965
rect 2115 11635 2177 11965
rect 1723 11587 2177 11635
rect 1706 11579 2194 11587
rect 2256 12013 2314 12021
rect 2273 11986 2314 12013
rect 2686 12021 2721 12027
rect 2823 12021 3277 12027
rect 3379 12021 3414 12027
rect 2686 12013 2744 12021
rect 2686 11986 2727 12013
rect 2273 11587 2314 11614
rect 2256 11579 2314 11587
rect 1586 11573 1621 11579
rect 1723 11573 2177 11579
rect 2279 11573 2314 11579
rect 2686 11587 2727 11614
rect 2686 11579 2744 11587
rect 2806 12013 3294 12021
rect 2823 11965 3277 12013
rect 2823 11635 2885 11965
rect 3215 11635 3277 11965
rect 2823 11587 3277 11635
rect 2806 11579 3294 11587
rect 3356 12013 3414 12021
rect 3373 11986 3414 12013
rect 3786 12021 3821 12027
rect 3923 12021 4377 12027
rect 4479 12021 4514 12027
rect 3786 12013 3844 12021
rect 3786 11986 3827 12013
rect 3373 11587 3414 11614
rect 3356 11579 3414 11587
rect 2686 11573 2721 11579
rect 2823 11573 3277 11579
rect 3379 11573 3414 11579
rect 3786 11587 3827 11614
rect 3786 11579 3844 11587
rect 3906 12013 4394 12021
rect 3923 11965 4377 12013
rect 3923 11635 3985 11965
rect 4315 11635 4377 11965
rect 3923 11587 4377 11635
rect 3906 11579 4394 11587
rect 4456 12013 4514 12021
rect 4473 11986 4514 12013
rect 4886 12021 4921 12027
rect 5023 12021 5477 12027
rect 5579 12021 5614 12027
rect 4886 12013 4944 12021
rect 4886 11986 4927 12013
rect 4473 11587 4514 11614
rect 4456 11579 4514 11587
rect 3786 11573 3821 11579
rect 3923 11573 4377 11579
rect 4479 11573 4514 11579
rect 4886 11587 4927 11614
rect 4886 11579 4944 11587
rect 5006 12013 5494 12021
rect 5023 11965 5477 12013
rect 5023 11635 5085 11965
rect 5415 11635 5477 11965
rect 5023 11587 5477 11635
rect 5006 11579 5494 11587
rect 5556 12013 5614 12021
rect 5573 11986 5614 12013
rect 5986 12021 6021 12027
rect 6123 12021 6577 12027
rect 6679 12021 6714 12027
rect 5986 12013 6044 12021
rect 5986 11986 6027 12013
rect 5573 11587 5614 11614
rect 5556 11579 5614 11587
rect 4886 11573 4921 11579
rect 5023 11573 5477 11579
rect 5579 11573 5614 11579
rect 5986 11587 6027 11614
rect 5986 11579 6044 11587
rect 6106 12013 6594 12021
rect 6123 11965 6577 12013
rect 6123 11635 6185 11965
rect 6515 11635 6577 11965
rect 6123 11587 6577 11635
rect 6106 11579 6594 11587
rect 6656 12013 6714 12021
rect 6673 11986 6714 12013
rect 7086 12021 7121 12027
rect 7223 12021 7677 12027
rect 7779 12021 7814 12027
rect 7086 12013 7144 12021
rect 7086 11986 7127 12013
rect 6673 11587 6714 11614
rect 6656 11579 6714 11587
rect 5986 11573 6021 11579
rect 6123 11573 6577 11579
rect 6679 11573 6714 11579
rect 7086 11587 7127 11614
rect 7086 11579 7144 11587
rect 7206 12013 7694 12021
rect 7223 11965 7677 12013
rect 7223 11635 7285 11965
rect 7615 11635 7677 11965
rect 7223 11587 7677 11635
rect 7206 11579 7694 11587
rect 7756 12013 7814 12021
rect 7773 11986 7814 12013
rect 8186 12021 8221 12027
rect 8323 12021 8777 12027
rect 8879 12021 8914 12027
rect 8186 12013 8244 12021
rect 8186 11986 8227 12013
rect 7773 11587 7814 11614
rect 7756 11579 7814 11587
rect 7086 11573 7121 11579
rect 7223 11573 7677 11579
rect 7779 11573 7814 11579
rect 8186 11587 8227 11614
rect 8186 11579 8244 11587
rect 8306 12013 8794 12021
rect 8323 11965 8777 12013
rect 8323 11635 8385 11965
rect 8715 11635 8777 11965
rect 8323 11587 8777 11635
rect 8306 11579 8794 11587
rect 8856 12013 8914 12021
rect 8873 11986 8914 12013
rect 9286 12021 9321 12027
rect 9423 12021 9877 12027
rect 9979 12021 10014 12027
rect 9286 12013 9344 12021
rect 9286 11986 9327 12013
rect 8873 11587 8914 11614
rect 8856 11579 8914 11587
rect 8186 11573 8221 11579
rect 8323 11573 8777 11579
rect 8879 11573 8914 11579
rect 9286 11587 9327 11614
rect 9286 11579 9344 11587
rect 9406 12013 9894 12021
rect 9423 11965 9877 12013
rect 9423 11635 9485 11965
rect 9815 11635 9877 11965
rect 9423 11587 9877 11635
rect 9406 11579 9894 11587
rect 9956 12013 10014 12021
rect 9973 11986 10014 12013
rect 10386 12021 10421 12027
rect 10523 12021 10977 12027
rect 11079 12021 11114 12027
rect 10386 12013 10444 12021
rect 10386 11986 10427 12013
rect 9973 11587 10014 11614
rect 9956 11579 10014 11587
rect 9286 11573 9321 11579
rect 9423 11573 9877 11579
rect 9979 11573 10014 11579
rect 10386 11587 10427 11614
rect 10386 11579 10444 11587
rect 10506 12013 10994 12021
rect 10523 11965 10977 12013
rect 10523 11635 10585 11965
rect 10915 11635 10977 11965
rect 10523 11587 10977 11635
rect 10506 11579 10994 11587
rect 11056 12013 11114 12021
rect 11073 11986 11114 12013
rect 11486 12021 11521 12027
rect 11623 12021 12077 12027
rect 12179 12021 12214 12027
rect 11486 12013 11544 12021
rect 11486 11986 11527 12013
rect 11073 11587 11114 11614
rect 11056 11579 11114 11587
rect 10386 11573 10421 11579
rect 10523 11573 10977 11579
rect 11079 11573 11114 11579
rect 11486 11587 11527 11614
rect 11486 11579 11544 11587
rect 11606 12013 12094 12021
rect 11623 11965 12077 12013
rect 11623 11635 11685 11965
rect 12015 11635 12077 11965
rect 11623 11587 12077 11635
rect 11606 11579 12094 11587
rect 12156 12013 12214 12021
rect 12173 11986 12214 12013
rect 12586 12021 12621 12027
rect 12723 12021 13177 12027
rect 13279 12021 13314 12027
rect 12586 12013 12644 12021
rect 12586 11986 12627 12013
rect 12173 11587 12214 11614
rect 12156 11579 12214 11587
rect 11486 11573 11521 11579
rect 11623 11573 12077 11579
rect 12179 11573 12214 11579
rect 12586 11587 12627 11614
rect 12586 11579 12644 11587
rect 12706 12013 13194 12021
rect 12723 11965 13177 12013
rect 12723 11635 12785 11965
rect 13115 11635 13177 11965
rect 12723 11587 13177 11635
rect 12706 11579 13194 11587
rect 13256 12013 13314 12021
rect 13273 11986 13314 12013
rect 13273 11587 13314 11614
rect 13256 11579 13314 11587
rect 12586 11573 12621 11579
rect 12723 11573 13177 11579
rect 13279 11573 13314 11579
rect -1025 11550 -725 11567
rect -471 11556 -463 11573
rect -37 11556 -29 11573
rect 79 11556 87 11573
rect 513 11556 521 11573
rect 629 11556 637 11573
rect 1063 11556 1071 11573
rect 1179 11556 1187 11573
rect 1613 11556 1621 11573
rect 1729 11556 1737 11573
rect 2163 11556 2171 11573
rect 2279 11556 2287 11573
rect 2713 11556 2721 11573
rect 2829 11556 2837 11573
rect 3263 11556 3271 11573
rect 3379 11556 3387 11573
rect 3813 11556 3821 11573
rect 3929 11556 3937 11573
rect 4363 11556 4371 11573
rect 4479 11556 4487 11573
rect 4913 11556 4921 11573
rect 5029 11556 5037 11573
rect 5463 11556 5471 11573
rect 5579 11556 5587 11573
rect 6013 11556 6021 11573
rect 6129 11556 6137 11573
rect 6563 11556 6571 11573
rect 6679 11556 6687 11573
rect 7113 11556 7121 11573
rect 7229 11556 7237 11573
rect 7663 11556 7671 11573
rect 7779 11556 7787 11573
rect 8213 11556 8221 11573
rect 8329 11556 8337 11573
rect 8763 11556 8771 11573
rect 8879 11556 8887 11573
rect 9313 11556 9321 11573
rect 9429 11556 9437 11573
rect 9863 11556 9871 11573
rect 9979 11556 9987 11573
rect 10413 11556 10421 11573
rect 10529 11556 10537 11573
rect 10963 11556 10971 11573
rect 11079 11556 11087 11573
rect 11513 11556 11521 11573
rect 11629 11556 11637 11573
rect 12063 11556 12071 11573
rect 12179 11556 12187 11573
rect 12613 11556 12621 11573
rect 12729 11556 12737 11573
rect 13163 11556 13171 11573
rect 13279 11556 13287 11573
rect 13713 11556 13721 11573
rect 13975 11569 13987 12100
rect 14263 11569 14275 12100
rect 13975 11550 14275 11569
rect -1025 11017 -1013 11550
rect -737 11017 -725 11550
rect -550 11542 -500 11550
rect -550 11508 -542 11542
rect -508 11508 -500 11542
rect -550 11500 -500 11508
rect 0 11542 50 11550
rect 0 11508 8 11542
rect 42 11508 50 11542
rect 0 11500 50 11508
rect 550 11542 600 11550
rect 550 11508 558 11542
rect 592 11508 600 11542
rect 550 11500 600 11508
rect 1100 11542 1150 11550
rect 1100 11508 1108 11542
rect 1142 11508 1150 11542
rect 1100 11500 1150 11508
rect 1650 11542 1700 11550
rect 1650 11508 1658 11542
rect 1692 11508 1700 11542
rect 1650 11500 1700 11508
rect 2200 11542 2250 11550
rect 2200 11508 2208 11542
rect 2242 11508 2250 11542
rect 2200 11500 2250 11508
rect 2750 11542 2800 11550
rect 2750 11508 2758 11542
rect 2792 11508 2800 11542
rect 2750 11500 2800 11508
rect 3300 11542 3350 11550
rect 3300 11508 3308 11542
rect 3342 11508 3350 11542
rect 3300 11500 3350 11508
rect 3850 11542 3900 11550
rect 3850 11508 3858 11542
rect 3892 11508 3900 11542
rect 3850 11500 3900 11508
rect 4400 11542 4450 11550
rect 4400 11508 4408 11542
rect 4442 11508 4450 11542
rect 4400 11500 4450 11508
rect 4950 11542 5000 11550
rect 4950 11508 4958 11542
rect 4992 11508 5000 11542
rect 4950 11500 5000 11508
rect 5500 11542 5550 11550
rect 5500 11508 5508 11542
rect 5542 11508 5550 11542
rect 5500 11500 5550 11508
rect 6050 11542 6100 11550
rect 6050 11508 6058 11542
rect 6092 11508 6100 11542
rect 6050 11500 6100 11508
rect 6600 11542 6650 11550
rect 6600 11508 6608 11542
rect 6642 11508 6650 11542
rect 6600 11500 6650 11508
rect 7150 11542 7200 11550
rect 7150 11508 7158 11542
rect 7192 11508 7200 11542
rect 7150 11500 7200 11508
rect 7700 11542 7750 11550
rect 7700 11508 7708 11542
rect 7742 11508 7750 11542
rect 7700 11500 7750 11508
rect 8250 11542 8300 11550
rect 8250 11508 8258 11542
rect 8292 11508 8300 11542
rect 8250 11500 8300 11508
rect 8800 11542 8850 11550
rect 8800 11508 8808 11542
rect 8842 11508 8850 11542
rect 8800 11500 8850 11508
rect 9350 11542 9400 11550
rect 9350 11508 9358 11542
rect 9392 11508 9400 11542
rect 9350 11500 9400 11508
rect 9900 11542 9950 11550
rect 9900 11508 9908 11542
rect 9942 11508 9950 11542
rect 9900 11500 9950 11508
rect 10450 11542 10500 11550
rect 10450 11508 10458 11542
rect 10492 11508 10500 11542
rect 10450 11500 10500 11508
rect 11000 11542 11050 11550
rect 11000 11508 11008 11542
rect 11042 11508 11050 11542
rect 11000 11500 11050 11508
rect 11550 11542 11600 11550
rect 11550 11508 11558 11542
rect 11592 11508 11600 11542
rect 11550 11500 11600 11508
rect 12100 11542 12150 11550
rect 12100 11508 12108 11542
rect 12142 11508 12150 11542
rect 12100 11500 12150 11508
rect 12650 11542 12700 11550
rect 12650 11508 12658 11542
rect 12692 11508 12700 11542
rect 12650 11500 12700 11508
rect 13200 11542 13250 11550
rect 13200 11508 13208 11542
rect 13242 11508 13250 11542
rect 13200 11500 13250 11508
rect 13750 11542 13800 11550
rect 13750 11508 13758 11542
rect 13792 11508 13800 11542
rect 13750 11500 13800 11508
rect -471 11477 -463 11494
rect -37 11477 -29 11494
rect 79 11477 87 11494
rect 513 11477 521 11494
rect 629 11477 637 11494
rect 1063 11477 1071 11494
rect 1179 11477 1187 11494
rect 1613 11477 1621 11494
rect 1729 11477 1737 11494
rect 2163 11477 2171 11494
rect 2279 11477 2287 11494
rect 2713 11477 2721 11494
rect 2829 11477 2837 11494
rect 3263 11477 3271 11494
rect 3379 11477 3387 11494
rect 3813 11477 3821 11494
rect 3929 11477 3937 11494
rect 4363 11477 4371 11494
rect 4479 11477 4487 11494
rect 4913 11477 4921 11494
rect 5029 11477 5037 11494
rect 5463 11477 5471 11494
rect 5579 11477 5587 11494
rect 6013 11477 6021 11494
rect 6129 11477 6137 11494
rect 6563 11477 6571 11494
rect 6679 11477 6687 11494
rect 7113 11477 7121 11494
rect 7229 11477 7237 11494
rect 7663 11477 7671 11494
rect 7779 11477 7787 11494
rect 8213 11477 8221 11494
rect 8329 11477 8337 11494
rect 8763 11477 8771 11494
rect 8879 11477 8887 11494
rect 9313 11477 9321 11494
rect 9429 11477 9437 11494
rect 9863 11477 9871 11494
rect 9979 11477 9987 11494
rect 10413 11477 10421 11494
rect 10529 11477 10537 11494
rect 10963 11477 10971 11494
rect 11079 11477 11087 11494
rect 11513 11477 11521 11494
rect 11629 11477 11637 11494
rect 12063 11477 12071 11494
rect 12179 11477 12187 11494
rect 12613 11477 12621 11494
rect 12729 11477 12737 11494
rect 13163 11477 13171 11494
rect 13279 11477 13287 11494
rect 13713 11477 13721 11494
rect -64 11471 -29 11477
rect 73 11471 527 11477
rect 629 11471 664 11477
rect -64 11463 -6 11471
rect -64 11436 -23 11463
rect -64 11037 -23 11064
rect -64 11029 -6 11037
rect 56 11463 544 11471
rect 73 11415 527 11463
rect 73 11085 135 11415
rect 465 11085 527 11415
rect 73 11037 527 11085
rect 56 11029 544 11037
rect 606 11463 664 11471
rect 623 11436 664 11463
rect 1036 11471 1071 11477
rect 1173 11471 1627 11477
rect 1729 11471 1764 11477
rect 1036 11463 1094 11471
rect 1036 11436 1077 11463
rect 623 11037 664 11064
rect 606 11029 664 11037
rect -64 11023 -29 11029
rect 73 11023 527 11029
rect 629 11023 664 11029
rect 1036 11037 1077 11064
rect 1036 11029 1094 11037
rect 1156 11463 1644 11471
rect 1173 11415 1627 11463
rect 1173 11085 1235 11415
rect 1565 11085 1627 11415
rect 1173 11037 1627 11085
rect 1156 11029 1644 11037
rect 1706 11463 1764 11471
rect 1723 11436 1764 11463
rect 2136 11471 2171 11477
rect 2273 11471 2727 11477
rect 2829 11471 2864 11477
rect 2136 11463 2194 11471
rect 2136 11436 2177 11463
rect 1723 11037 1764 11064
rect 1706 11029 1764 11037
rect 1036 11023 1071 11029
rect 1173 11023 1627 11029
rect 1729 11023 1764 11029
rect 2136 11037 2177 11064
rect 2136 11029 2194 11037
rect 2256 11463 2744 11471
rect 2273 11415 2727 11463
rect 2273 11085 2335 11415
rect 2665 11085 2727 11415
rect 2273 11037 2727 11085
rect 2256 11029 2744 11037
rect 2806 11463 2864 11471
rect 2823 11436 2864 11463
rect 3236 11471 3271 11477
rect 3373 11471 3827 11477
rect 3929 11471 3964 11477
rect 3236 11463 3294 11471
rect 3236 11436 3277 11463
rect 2823 11037 2864 11064
rect 2806 11029 2864 11037
rect 2136 11023 2171 11029
rect 2273 11023 2727 11029
rect 2829 11023 2864 11029
rect 3236 11037 3277 11064
rect 3236 11029 3294 11037
rect 3356 11463 3844 11471
rect 3373 11415 3827 11463
rect 3373 11085 3435 11415
rect 3765 11085 3827 11415
rect 3373 11037 3827 11085
rect 3356 11029 3844 11037
rect 3906 11463 3964 11471
rect 3923 11436 3964 11463
rect 4336 11471 4371 11477
rect 4473 11471 4927 11477
rect 5029 11471 5064 11477
rect 4336 11463 4394 11471
rect 4336 11436 4377 11463
rect 3923 11037 3964 11064
rect 3906 11029 3964 11037
rect 3236 11023 3271 11029
rect 3373 11023 3827 11029
rect 3929 11023 3964 11029
rect 4336 11037 4377 11064
rect 4336 11029 4394 11037
rect 4456 11463 4944 11471
rect 4473 11415 4927 11463
rect 4473 11085 4535 11415
rect 4865 11085 4927 11415
rect 4473 11037 4927 11085
rect 4456 11029 4944 11037
rect 5006 11463 5064 11471
rect 5023 11436 5064 11463
rect 5436 11471 5471 11477
rect 5573 11471 6027 11477
rect 6129 11471 6164 11477
rect 5436 11463 5494 11471
rect 5436 11436 5477 11463
rect 5023 11037 5064 11064
rect 5006 11029 5064 11037
rect 4336 11023 4371 11029
rect 4473 11023 4927 11029
rect 5029 11023 5064 11029
rect 5436 11037 5477 11064
rect 5436 11029 5494 11037
rect 5556 11463 6044 11471
rect 5573 11415 6027 11463
rect 5573 11085 5635 11415
rect 5965 11085 6027 11415
rect 5573 11037 6027 11085
rect 5556 11029 6044 11037
rect 6106 11463 6164 11471
rect 6123 11436 6164 11463
rect 6536 11471 6571 11477
rect 6673 11471 7127 11477
rect 7229 11471 7264 11477
rect 6536 11463 6594 11471
rect 6536 11436 6577 11463
rect 6123 11037 6164 11064
rect 6106 11029 6164 11037
rect 5436 11023 5471 11029
rect 5573 11023 6027 11029
rect 6129 11023 6164 11029
rect 6536 11037 6577 11064
rect 6536 11029 6594 11037
rect 6656 11463 7144 11471
rect 6673 11415 7127 11463
rect 6673 11085 6735 11415
rect 7065 11085 7127 11415
rect 6673 11037 7127 11085
rect 6656 11029 7144 11037
rect 7206 11463 7264 11471
rect 7223 11436 7264 11463
rect 7636 11471 7671 11477
rect 7773 11471 8227 11477
rect 8329 11471 8364 11477
rect 7636 11463 7694 11471
rect 7636 11436 7677 11463
rect 7223 11037 7264 11064
rect 7206 11029 7264 11037
rect 6536 11023 6571 11029
rect 6673 11023 7127 11029
rect 7229 11023 7264 11029
rect 7636 11037 7677 11064
rect 7636 11029 7694 11037
rect 7756 11463 8244 11471
rect 7773 11415 8227 11463
rect 7773 11085 7835 11415
rect 8165 11085 8227 11415
rect 7773 11037 8227 11085
rect 7756 11029 8244 11037
rect 8306 11463 8364 11471
rect 8323 11436 8364 11463
rect 8736 11471 8771 11477
rect 8873 11471 9327 11477
rect 9429 11471 9464 11477
rect 8736 11463 8794 11471
rect 8736 11436 8777 11463
rect 8323 11037 8364 11064
rect 8306 11029 8364 11037
rect 7636 11023 7671 11029
rect 7773 11023 8227 11029
rect 8329 11023 8364 11029
rect 8736 11037 8777 11064
rect 8736 11029 8794 11037
rect 8856 11463 9344 11471
rect 8873 11415 9327 11463
rect 8873 11085 8935 11415
rect 9265 11085 9327 11415
rect 8873 11037 9327 11085
rect 8856 11029 9344 11037
rect 9406 11463 9464 11471
rect 9423 11436 9464 11463
rect 9836 11471 9871 11477
rect 9973 11471 10427 11477
rect 10529 11471 10564 11477
rect 9836 11463 9894 11471
rect 9836 11436 9877 11463
rect 9423 11037 9464 11064
rect 9406 11029 9464 11037
rect 8736 11023 8771 11029
rect 8873 11023 9327 11029
rect 9429 11023 9464 11029
rect 9836 11037 9877 11064
rect 9836 11029 9894 11037
rect 9956 11463 10444 11471
rect 9973 11415 10427 11463
rect 9973 11085 10035 11415
rect 10365 11085 10427 11415
rect 9973 11037 10427 11085
rect 9956 11029 10444 11037
rect 10506 11463 10564 11471
rect 10523 11436 10564 11463
rect 10936 11471 10971 11477
rect 11073 11471 11527 11477
rect 11629 11471 11664 11477
rect 10936 11463 10994 11471
rect 10936 11436 10977 11463
rect 10523 11037 10564 11064
rect 10506 11029 10564 11037
rect 9836 11023 9871 11029
rect 9973 11023 10427 11029
rect 10529 11023 10564 11029
rect 10936 11037 10977 11064
rect 10936 11029 10994 11037
rect 11056 11463 11544 11471
rect 11073 11415 11527 11463
rect 11073 11085 11135 11415
rect 11465 11085 11527 11415
rect 11073 11037 11527 11085
rect 11056 11029 11544 11037
rect 11606 11463 11664 11471
rect 11623 11436 11664 11463
rect 12036 11471 12071 11477
rect 12173 11471 12627 11477
rect 12729 11471 12764 11477
rect 12036 11463 12094 11471
rect 12036 11436 12077 11463
rect 11623 11037 11664 11064
rect 11606 11029 11664 11037
rect 10936 11023 10971 11029
rect 11073 11023 11527 11029
rect 11629 11023 11664 11029
rect 12036 11037 12077 11064
rect 12036 11029 12094 11037
rect 12156 11463 12644 11471
rect 12173 11415 12627 11463
rect 12173 11085 12235 11415
rect 12565 11085 12627 11415
rect 12173 11037 12627 11085
rect 12156 11029 12644 11037
rect 12706 11463 12764 11471
rect 12723 11436 12764 11463
rect 13136 11471 13171 11477
rect 13273 11471 13727 11477
rect 13136 11463 13194 11471
rect 13136 11436 13177 11463
rect 12723 11037 12764 11064
rect 12706 11029 12764 11037
rect 12036 11023 12071 11029
rect 12173 11023 12627 11029
rect 12729 11023 12764 11029
rect 13136 11037 13177 11064
rect 13136 11029 13194 11037
rect 13256 11463 13727 11471
rect 13273 11415 13727 11463
rect 13273 11085 13335 11415
rect 13665 11085 13727 11415
rect 13273 11037 13727 11085
rect 13256 11029 13727 11037
rect 13136 11023 13171 11029
rect 13273 11023 13727 11029
rect -1025 11000 -725 11017
rect -471 11006 -463 11023
rect -37 11006 -29 11023
rect 79 11006 87 11023
rect 513 11006 521 11023
rect 629 11006 637 11023
rect 1063 11006 1071 11023
rect 1179 11006 1187 11023
rect 1613 11006 1621 11023
rect 1729 11006 1737 11023
rect 2163 11006 2171 11023
rect 2279 11006 2287 11023
rect 2713 11006 2721 11023
rect 2829 11006 2837 11023
rect 3263 11006 3271 11023
rect 3379 11006 3387 11023
rect 3813 11006 3821 11023
rect 3929 11006 3937 11023
rect 4363 11006 4371 11023
rect 4479 11006 4487 11023
rect 4913 11006 4921 11023
rect 5029 11006 5037 11023
rect 5463 11006 5471 11023
rect 5579 11006 5587 11023
rect 6013 11006 6021 11023
rect 6129 11006 6137 11023
rect 6563 11006 6571 11023
rect 6679 11006 6687 11023
rect 7113 11006 7121 11023
rect 7229 11006 7237 11023
rect 7663 11006 7671 11023
rect 7779 11006 7787 11023
rect 8213 11006 8221 11023
rect 8329 11006 8337 11023
rect 8763 11006 8771 11023
rect 8879 11006 8887 11023
rect 9313 11006 9321 11023
rect 9429 11006 9437 11023
rect 9863 11006 9871 11023
rect 9979 11006 9987 11023
rect 10413 11006 10421 11023
rect 10529 11006 10537 11023
rect 10963 11006 10971 11023
rect 11079 11006 11087 11023
rect 11513 11006 11521 11023
rect 11629 11006 11637 11023
rect 12063 11006 12071 11023
rect 12179 11006 12187 11023
rect 12613 11006 12621 11023
rect 12729 11006 12737 11023
rect 13163 11006 13171 11023
rect 13279 11006 13287 11023
rect 13713 11006 13721 11023
rect 13975 11017 13987 11550
rect 14263 11017 14275 11550
rect 13975 11000 14275 11017
rect -1025 10467 -1013 11000
rect -737 10467 -725 11000
rect -550 10992 -500 11000
rect -550 10958 -542 10992
rect -508 10958 -500 10992
rect -550 10950 -500 10958
rect 0 10992 50 11000
rect 0 10958 8 10992
rect 42 10958 50 10992
rect 0 10950 50 10958
rect 550 10992 600 11000
rect 550 10958 558 10992
rect 592 10958 600 10992
rect 550 10950 600 10958
rect 1100 10992 1150 11000
rect 1100 10958 1108 10992
rect 1142 10958 1150 10992
rect 1100 10950 1150 10958
rect 1650 10992 1700 11000
rect 1650 10958 1658 10992
rect 1692 10958 1700 10992
rect 1650 10950 1700 10958
rect 2200 10992 2250 11000
rect 2200 10958 2208 10992
rect 2242 10958 2250 10992
rect 2200 10950 2250 10958
rect 2750 10992 2800 11000
rect 2750 10958 2758 10992
rect 2792 10958 2800 10992
rect 2750 10950 2800 10958
rect 3300 10992 3350 11000
rect 3300 10958 3308 10992
rect 3342 10958 3350 10992
rect 3300 10950 3350 10958
rect 3850 10992 3900 11000
rect 3850 10958 3858 10992
rect 3892 10958 3900 10992
rect 3850 10950 3900 10958
rect 4400 10992 4450 11000
rect 4400 10958 4408 10992
rect 4442 10958 4450 10992
rect 4400 10950 4450 10958
rect 4950 10992 5000 11000
rect 4950 10958 4958 10992
rect 4992 10958 5000 10992
rect 4950 10950 5000 10958
rect 5500 10992 5550 11000
rect 5500 10958 5508 10992
rect 5542 10958 5550 10992
rect 5500 10950 5550 10958
rect 6050 10992 6100 11000
rect 6050 10958 6058 10992
rect 6092 10958 6100 10992
rect 6050 10950 6100 10958
rect 6600 10992 6650 11000
rect 6600 10958 6608 10992
rect 6642 10958 6650 10992
rect 6600 10950 6650 10958
rect 7150 10992 7200 11000
rect 7150 10958 7158 10992
rect 7192 10958 7200 10992
rect 7150 10950 7200 10958
rect 7700 10992 7750 11000
rect 7700 10958 7708 10992
rect 7742 10958 7750 10992
rect 7700 10950 7750 10958
rect 8250 10992 8300 11000
rect 8250 10958 8258 10992
rect 8292 10958 8300 10992
rect 8250 10950 8300 10958
rect 8800 10992 8850 11000
rect 8800 10958 8808 10992
rect 8842 10958 8850 10992
rect 8800 10950 8850 10958
rect 9350 10992 9400 11000
rect 9350 10958 9358 10992
rect 9392 10958 9400 10992
rect 9350 10950 9400 10958
rect 9900 10992 9950 11000
rect 9900 10958 9908 10992
rect 9942 10958 9950 10992
rect 9900 10950 9950 10958
rect 10450 10992 10500 11000
rect 10450 10958 10458 10992
rect 10492 10958 10500 10992
rect 10450 10950 10500 10958
rect 11000 10992 11050 11000
rect 11000 10958 11008 10992
rect 11042 10958 11050 10992
rect 11000 10950 11050 10958
rect 11550 10992 11600 11000
rect 11550 10958 11558 10992
rect 11592 10958 11600 10992
rect 11550 10950 11600 10958
rect 12100 10992 12150 11000
rect 12100 10958 12108 10992
rect 12142 10958 12150 10992
rect 12100 10950 12150 10958
rect 12650 10992 12700 11000
rect 12650 10958 12658 10992
rect 12692 10958 12700 10992
rect 12650 10950 12700 10958
rect 13200 10992 13250 11000
rect 13200 10958 13208 10992
rect 13242 10958 13250 10992
rect 13200 10950 13250 10958
rect 13750 10992 13800 11000
rect 13750 10958 13758 10992
rect 13792 10958 13800 10992
rect 13750 10950 13800 10958
rect -471 10927 -463 10944
rect -37 10927 -29 10944
rect 79 10927 87 10944
rect 513 10927 521 10944
rect 629 10927 637 10944
rect 1063 10927 1071 10944
rect 1179 10927 1187 10944
rect 1613 10927 1621 10944
rect 1729 10927 1737 10944
rect 2163 10927 2171 10944
rect 2279 10927 2287 10944
rect 2713 10927 2721 10944
rect 2829 10927 2837 10944
rect 3263 10927 3271 10944
rect 3379 10927 3387 10944
rect 3813 10927 3821 10944
rect 3929 10927 3937 10944
rect 4363 10927 4371 10944
rect 4479 10927 4487 10944
rect 4913 10927 4921 10944
rect 5029 10927 5037 10944
rect 5463 10927 5471 10944
rect 5579 10927 5587 10944
rect 6013 10927 6021 10944
rect 6129 10927 6137 10944
rect 6563 10927 6571 10944
rect 6679 10927 6687 10944
rect 7113 10927 7121 10944
rect 7229 10927 7237 10944
rect 7663 10927 7671 10944
rect 7779 10927 7787 10944
rect 8213 10927 8221 10944
rect 8329 10927 8337 10944
rect 8763 10927 8771 10944
rect 8879 10927 8887 10944
rect 9313 10927 9321 10944
rect 9429 10927 9437 10944
rect 9863 10927 9871 10944
rect 9979 10927 9987 10944
rect 10413 10927 10421 10944
rect 10529 10927 10537 10944
rect 10963 10927 10971 10944
rect 11079 10927 11087 10944
rect 11513 10927 11521 10944
rect 11629 10927 11637 10944
rect 12063 10927 12071 10944
rect 12179 10927 12187 10944
rect 12613 10927 12621 10944
rect 12729 10927 12737 10944
rect 13163 10927 13171 10944
rect 13279 10927 13287 10944
rect 13713 10927 13721 10944
rect -477 10921 -23 10927
rect 79 10921 114 10927
rect -477 10913 -6 10921
rect -477 10865 -23 10913
rect -477 10535 -415 10865
rect -85 10535 -23 10865
rect -477 10487 -23 10535
rect -477 10479 -6 10487
rect 56 10913 114 10921
rect 73 10886 114 10913
rect 486 10921 521 10927
rect 623 10921 1077 10927
rect 1179 10921 1214 10927
rect 486 10913 544 10921
rect 486 10886 527 10913
rect 73 10487 114 10514
rect 56 10479 114 10487
rect -477 10473 -23 10479
rect 79 10473 114 10479
rect 486 10487 527 10514
rect 486 10479 544 10487
rect 606 10913 1094 10921
rect 623 10865 1077 10913
rect 623 10535 685 10865
rect 1015 10535 1077 10865
rect 623 10487 1077 10535
rect 606 10479 1094 10487
rect 1156 10913 1214 10921
rect 1173 10886 1214 10913
rect 1586 10921 1621 10927
rect 1723 10921 2177 10927
rect 2279 10921 2314 10927
rect 1586 10913 1644 10921
rect 1586 10886 1627 10913
rect 1173 10487 1214 10514
rect 1156 10479 1214 10487
rect 486 10473 521 10479
rect 623 10473 1077 10479
rect 1179 10473 1214 10479
rect 1586 10487 1627 10514
rect 1586 10479 1644 10487
rect 1706 10913 2194 10921
rect 1723 10865 2177 10913
rect 1723 10535 1785 10865
rect 2115 10535 2177 10865
rect 1723 10487 2177 10535
rect 1706 10479 2194 10487
rect 2256 10913 2314 10921
rect 2273 10886 2314 10913
rect 2686 10921 2721 10927
rect 2823 10921 3277 10927
rect 3379 10921 3414 10927
rect 2686 10913 2744 10921
rect 2686 10886 2727 10913
rect 2273 10487 2314 10514
rect 2256 10479 2314 10487
rect 1586 10473 1621 10479
rect 1723 10473 2177 10479
rect 2279 10473 2314 10479
rect 2686 10487 2727 10514
rect 2686 10479 2744 10487
rect 2806 10913 3294 10921
rect 2823 10865 3277 10913
rect 2823 10535 2885 10865
rect 3215 10535 3277 10865
rect 2823 10487 3277 10535
rect 2806 10479 3294 10487
rect 3356 10913 3414 10921
rect 3373 10886 3414 10913
rect 3786 10921 3821 10927
rect 3923 10921 4377 10927
rect 4479 10921 4514 10927
rect 3786 10913 3844 10921
rect 3786 10886 3827 10913
rect 3373 10487 3414 10514
rect 3356 10479 3414 10487
rect 2686 10473 2721 10479
rect 2823 10473 3277 10479
rect 3379 10473 3414 10479
rect 3786 10487 3827 10514
rect 3786 10479 3844 10487
rect 3906 10913 4394 10921
rect 3923 10865 4377 10913
rect 3923 10535 3985 10865
rect 4315 10535 4377 10865
rect 3923 10487 4377 10535
rect 3906 10479 4394 10487
rect 4456 10913 4514 10921
rect 4473 10886 4514 10913
rect 4886 10921 4921 10927
rect 5023 10921 5477 10927
rect 5579 10921 5614 10927
rect 4886 10913 4944 10921
rect 4886 10886 4927 10913
rect 4473 10487 4514 10514
rect 4456 10479 4514 10487
rect 3786 10473 3821 10479
rect 3923 10473 4377 10479
rect 4479 10473 4514 10479
rect 4886 10487 4927 10514
rect 4886 10479 4944 10487
rect 5006 10913 5494 10921
rect 5023 10865 5477 10913
rect 5023 10535 5085 10865
rect 5415 10535 5477 10865
rect 5023 10487 5477 10535
rect 5006 10479 5494 10487
rect 5556 10913 5614 10921
rect 5573 10886 5614 10913
rect 5986 10921 6021 10927
rect 6123 10921 6577 10927
rect 6679 10921 6714 10927
rect 5986 10913 6044 10921
rect 5986 10886 6027 10913
rect 5573 10487 5614 10514
rect 5556 10479 5614 10487
rect 4886 10473 4921 10479
rect 5023 10473 5477 10479
rect 5579 10473 5614 10479
rect 5986 10487 6027 10514
rect 5986 10479 6044 10487
rect 6106 10913 6594 10921
rect 6123 10865 6577 10913
rect 6123 10535 6185 10865
rect 6515 10535 6577 10865
rect 6123 10487 6577 10535
rect 6106 10479 6594 10487
rect 6656 10913 6714 10921
rect 6673 10886 6714 10913
rect 7086 10921 7121 10927
rect 7223 10921 7677 10927
rect 7779 10921 7814 10927
rect 7086 10913 7144 10921
rect 7086 10886 7127 10913
rect 6673 10487 6714 10514
rect 6656 10479 6714 10487
rect 5986 10473 6021 10479
rect 6123 10473 6577 10479
rect 6679 10473 6714 10479
rect 7086 10487 7127 10514
rect 7086 10479 7144 10487
rect 7206 10913 7694 10921
rect 7223 10865 7677 10913
rect 7223 10535 7285 10865
rect 7615 10535 7677 10865
rect 7223 10487 7677 10535
rect 7206 10479 7694 10487
rect 7756 10913 7814 10921
rect 7773 10886 7814 10913
rect 8186 10921 8221 10927
rect 8323 10921 8777 10927
rect 8879 10921 8914 10927
rect 8186 10913 8244 10921
rect 8186 10886 8227 10913
rect 7773 10487 7814 10514
rect 7756 10479 7814 10487
rect 7086 10473 7121 10479
rect 7223 10473 7677 10479
rect 7779 10473 7814 10479
rect 8186 10487 8227 10514
rect 8186 10479 8244 10487
rect 8306 10913 8794 10921
rect 8323 10865 8777 10913
rect 8323 10535 8385 10865
rect 8715 10535 8777 10865
rect 8323 10487 8777 10535
rect 8306 10479 8794 10487
rect 8856 10913 8914 10921
rect 8873 10886 8914 10913
rect 9286 10921 9321 10927
rect 9423 10921 9877 10927
rect 9979 10921 10014 10927
rect 9286 10913 9344 10921
rect 9286 10886 9327 10913
rect 8873 10487 8914 10514
rect 8856 10479 8914 10487
rect 8186 10473 8221 10479
rect 8323 10473 8777 10479
rect 8879 10473 8914 10479
rect 9286 10487 9327 10514
rect 9286 10479 9344 10487
rect 9406 10913 9894 10921
rect 9423 10865 9877 10913
rect 9423 10535 9485 10865
rect 9815 10535 9877 10865
rect 9423 10487 9877 10535
rect 9406 10479 9894 10487
rect 9956 10913 10014 10921
rect 9973 10886 10014 10913
rect 10386 10921 10421 10927
rect 10523 10921 10977 10927
rect 11079 10921 11114 10927
rect 10386 10913 10444 10921
rect 10386 10886 10427 10913
rect 9973 10487 10014 10514
rect 9956 10479 10014 10487
rect 9286 10473 9321 10479
rect 9423 10473 9877 10479
rect 9979 10473 10014 10479
rect 10386 10487 10427 10514
rect 10386 10479 10444 10487
rect 10506 10913 10994 10921
rect 10523 10865 10977 10913
rect 10523 10535 10585 10865
rect 10915 10535 10977 10865
rect 10523 10487 10977 10535
rect 10506 10479 10994 10487
rect 11056 10913 11114 10921
rect 11073 10886 11114 10913
rect 11486 10921 11521 10927
rect 11623 10921 12077 10927
rect 12179 10921 12214 10927
rect 11486 10913 11544 10921
rect 11486 10886 11527 10913
rect 11073 10487 11114 10514
rect 11056 10479 11114 10487
rect 10386 10473 10421 10479
rect 10523 10473 10977 10479
rect 11079 10473 11114 10479
rect 11486 10487 11527 10514
rect 11486 10479 11544 10487
rect 11606 10913 12094 10921
rect 11623 10865 12077 10913
rect 11623 10535 11685 10865
rect 12015 10535 12077 10865
rect 11623 10487 12077 10535
rect 11606 10479 12094 10487
rect 12156 10913 12214 10921
rect 12173 10886 12214 10913
rect 12586 10921 12621 10927
rect 12723 10921 13177 10927
rect 13279 10921 13314 10927
rect 12586 10913 12644 10921
rect 12586 10886 12627 10913
rect 12173 10487 12214 10514
rect 12156 10479 12214 10487
rect 11486 10473 11521 10479
rect 11623 10473 12077 10479
rect 12179 10473 12214 10479
rect 12586 10487 12627 10514
rect 12586 10479 12644 10487
rect 12706 10913 13194 10921
rect 12723 10865 13177 10913
rect 12723 10535 12785 10865
rect 13115 10535 13177 10865
rect 12723 10487 13177 10535
rect 12706 10479 13194 10487
rect 13256 10913 13314 10921
rect 13273 10886 13314 10913
rect 13273 10487 13314 10514
rect 13256 10479 13314 10487
rect 12586 10473 12621 10479
rect 12723 10473 13177 10479
rect 13279 10473 13314 10479
rect -1025 10450 -725 10467
rect -471 10456 -463 10473
rect -37 10456 -29 10473
rect 79 10456 87 10473
rect 513 10456 521 10473
rect 629 10456 637 10473
rect 1063 10456 1071 10473
rect 1179 10456 1187 10473
rect 1613 10456 1621 10473
rect 1729 10456 1737 10473
rect 2163 10456 2171 10473
rect 2279 10456 2287 10473
rect 2713 10456 2721 10473
rect 2829 10456 2837 10473
rect 3263 10456 3271 10473
rect 3379 10456 3387 10473
rect 3813 10456 3821 10473
rect 3929 10456 3937 10473
rect 4363 10456 4371 10473
rect 4479 10456 4487 10473
rect 4913 10456 4921 10473
rect 5029 10456 5037 10473
rect 5463 10456 5471 10473
rect 5579 10456 5587 10473
rect 6013 10456 6021 10473
rect 6129 10456 6137 10473
rect 6563 10456 6571 10473
rect 6679 10456 6687 10473
rect 7113 10456 7121 10473
rect 7229 10456 7237 10473
rect 7663 10456 7671 10473
rect 7779 10456 7787 10473
rect 8213 10456 8221 10473
rect 8329 10456 8337 10473
rect 8763 10456 8771 10473
rect 8879 10456 8887 10473
rect 9313 10456 9321 10473
rect 9429 10456 9437 10473
rect 9863 10456 9871 10473
rect 9979 10456 9987 10473
rect 10413 10456 10421 10473
rect 10529 10456 10537 10473
rect 10963 10456 10971 10473
rect 11079 10456 11087 10473
rect 11513 10456 11521 10473
rect 11629 10456 11637 10473
rect 12063 10456 12071 10473
rect 12179 10456 12187 10473
rect 12613 10456 12621 10473
rect 12729 10456 12737 10473
rect 13163 10456 13171 10473
rect 13279 10456 13287 10473
rect 13713 10456 13721 10473
rect 13975 10469 13987 11000
rect 14263 10469 14275 11000
rect 13975 10450 14275 10469
rect -1025 9917 -1013 10450
rect -737 9917 -725 10450
rect -550 10442 -500 10450
rect -550 10408 -542 10442
rect -508 10408 -500 10442
rect -550 10400 -500 10408
rect 0 10442 50 10450
rect 0 10408 8 10442
rect 42 10408 50 10442
rect 0 10400 50 10408
rect 550 10442 600 10450
rect 550 10408 558 10442
rect 592 10408 600 10442
rect 550 10400 600 10408
rect 1100 10442 1150 10450
rect 1100 10408 1108 10442
rect 1142 10408 1150 10442
rect 1100 10400 1150 10408
rect 1650 10442 1700 10450
rect 1650 10408 1658 10442
rect 1692 10408 1700 10442
rect 1650 10400 1700 10408
rect 2200 10442 2250 10450
rect 2200 10408 2208 10442
rect 2242 10408 2250 10442
rect 2200 10400 2250 10408
rect 2750 10442 2800 10450
rect 2750 10408 2758 10442
rect 2792 10408 2800 10442
rect 2750 10400 2800 10408
rect 3300 10442 3350 10450
rect 3300 10408 3308 10442
rect 3342 10408 3350 10442
rect 3300 10400 3350 10408
rect 3850 10442 3900 10450
rect 3850 10408 3858 10442
rect 3892 10408 3900 10442
rect 3850 10400 3900 10408
rect 4400 10442 4450 10450
rect 4400 10408 4408 10442
rect 4442 10408 4450 10442
rect 4400 10400 4450 10408
rect 4950 10442 5000 10450
rect 4950 10408 4958 10442
rect 4992 10408 5000 10442
rect 4950 10400 5000 10408
rect 5500 10442 5550 10450
rect 5500 10408 5508 10442
rect 5542 10408 5550 10442
rect 5500 10400 5550 10408
rect 6050 10442 6100 10450
rect 6050 10408 6058 10442
rect 6092 10408 6100 10442
rect 6050 10400 6100 10408
rect 6600 10442 6650 10450
rect 6600 10408 6608 10442
rect 6642 10408 6650 10442
rect 6600 10400 6650 10408
rect 7150 10442 7200 10450
rect 7150 10408 7158 10442
rect 7192 10408 7200 10442
rect 7150 10400 7200 10408
rect 7700 10442 7750 10450
rect 7700 10408 7708 10442
rect 7742 10408 7750 10442
rect 7700 10400 7750 10408
rect 8250 10442 8300 10450
rect 8250 10408 8258 10442
rect 8292 10408 8300 10442
rect 8250 10400 8300 10408
rect 8800 10442 8850 10450
rect 8800 10408 8808 10442
rect 8842 10408 8850 10442
rect 8800 10400 8850 10408
rect 9350 10442 9400 10450
rect 9350 10408 9358 10442
rect 9392 10408 9400 10442
rect 9350 10400 9400 10408
rect 9900 10442 9950 10450
rect 9900 10408 9908 10442
rect 9942 10408 9950 10442
rect 9900 10400 9950 10408
rect 10450 10442 10500 10450
rect 10450 10408 10458 10442
rect 10492 10408 10500 10442
rect 10450 10400 10500 10408
rect 11000 10442 11050 10450
rect 11000 10408 11008 10442
rect 11042 10408 11050 10442
rect 11000 10400 11050 10408
rect 11550 10442 11600 10450
rect 11550 10408 11558 10442
rect 11592 10408 11600 10442
rect 11550 10400 11600 10408
rect 12100 10442 12150 10450
rect 12100 10408 12108 10442
rect 12142 10408 12150 10442
rect 12100 10400 12150 10408
rect 12650 10442 12700 10450
rect 12650 10408 12658 10442
rect 12692 10408 12700 10442
rect 12650 10400 12700 10408
rect 13200 10442 13250 10450
rect 13200 10408 13208 10442
rect 13242 10408 13250 10442
rect 13200 10400 13250 10408
rect 13750 10442 13800 10450
rect 13750 10408 13758 10442
rect 13792 10408 13800 10442
rect 13750 10400 13800 10408
rect -471 10377 -463 10394
rect -37 10377 -29 10394
rect 79 10377 87 10394
rect 513 10377 521 10394
rect 629 10377 637 10394
rect 1063 10377 1071 10394
rect 1179 10377 1187 10394
rect 1613 10377 1621 10394
rect 1729 10377 1737 10394
rect 2163 10377 2171 10394
rect 2279 10377 2287 10394
rect 2713 10377 2721 10394
rect 2829 10377 2837 10394
rect 3263 10377 3271 10394
rect 3379 10377 3387 10394
rect 3813 10377 3821 10394
rect 3929 10377 3937 10394
rect 4363 10377 4371 10394
rect 4479 10377 4487 10394
rect 4913 10377 4921 10394
rect 5029 10377 5037 10394
rect 5463 10377 5471 10394
rect 5579 10377 5587 10394
rect 6013 10377 6021 10394
rect 6129 10377 6137 10394
rect 6563 10377 6571 10394
rect 6679 10377 6687 10394
rect 7113 10377 7121 10394
rect 7229 10377 7237 10394
rect 7663 10377 7671 10394
rect 7779 10377 7787 10394
rect 8213 10377 8221 10394
rect 8329 10377 8337 10394
rect 8763 10377 8771 10394
rect 8879 10377 8887 10394
rect 9313 10377 9321 10394
rect 9429 10377 9437 10394
rect 9863 10377 9871 10394
rect 9979 10377 9987 10394
rect 10413 10377 10421 10394
rect 10529 10377 10537 10394
rect 10963 10377 10971 10394
rect 11079 10377 11087 10394
rect 11513 10377 11521 10394
rect 11629 10377 11637 10394
rect 12063 10377 12071 10394
rect 12179 10377 12187 10394
rect 12613 10377 12621 10394
rect 12729 10377 12737 10394
rect 13163 10377 13171 10394
rect 13279 10377 13287 10394
rect 13713 10377 13721 10394
rect -64 10371 -29 10377
rect 73 10371 527 10377
rect 629 10371 664 10377
rect -64 10363 -6 10371
rect -64 10336 -23 10363
rect -64 9937 -23 9964
rect -64 9929 -6 9937
rect 56 10363 544 10371
rect 73 10315 527 10363
rect 73 9985 135 10315
rect 465 9985 527 10315
rect 73 9937 527 9985
rect 56 9929 544 9937
rect 606 10363 664 10371
rect 623 10336 664 10363
rect 1036 10371 1071 10377
rect 1173 10371 1627 10377
rect 1729 10371 1764 10377
rect 1036 10363 1094 10371
rect 1036 10336 1077 10363
rect 623 9937 664 9964
rect 606 9929 664 9937
rect -64 9923 -29 9929
rect 73 9923 527 9929
rect 629 9923 664 9929
rect 1036 9937 1077 9964
rect 1036 9929 1094 9937
rect 1156 10363 1644 10371
rect 1173 10315 1627 10363
rect 1173 9985 1235 10315
rect 1565 9985 1627 10315
rect 1173 9937 1627 9985
rect 1156 9929 1644 9937
rect 1706 10363 1764 10371
rect 1723 10336 1764 10363
rect 2136 10371 2171 10377
rect 2273 10371 2727 10377
rect 2829 10371 2864 10377
rect 2136 10363 2194 10371
rect 2136 10336 2177 10363
rect 1723 9937 1764 9964
rect 1706 9929 1764 9937
rect 1036 9923 1071 9929
rect 1173 9923 1627 9929
rect 1729 9923 1764 9929
rect 2136 9937 2177 9964
rect 2136 9929 2194 9937
rect 2256 10363 2744 10371
rect 2273 10315 2727 10363
rect 2273 9985 2335 10315
rect 2665 9985 2727 10315
rect 2273 9937 2727 9985
rect 2256 9929 2744 9937
rect 2806 10363 2864 10371
rect 2823 10336 2864 10363
rect 3236 10371 3271 10377
rect 3373 10371 3827 10377
rect 3929 10371 3964 10377
rect 3236 10363 3294 10371
rect 3236 10336 3277 10363
rect 2823 9937 2864 9964
rect 2806 9929 2864 9937
rect 2136 9923 2171 9929
rect 2273 9923 2727 9929
rect 2829 9923 2864 9929
rect 3236 9937 3277 9964
rect 3236 9929 3294 9937
rect 3356 10363 3844 10371
rect 3373 10315 3827 10363
rect 3373 9985 3435 10315
rect 3765 9985 3827 10315
rect 3373 9937 3827 9985
rect 3356 9929 3844 9937
rect 3906 10363 3964 10371
rect 3923 10336 3964 10363
rect 4336 10371 4371 10377
rect 4473 10371 4927 10377
rect 5029 10371 5064 10377
rect 4336 10363 4394 10371
rect 4336 10336 4377 10363
rect 3923 9937 3964 9964
rect 3906 9929 3964 9937
rect 3236 9923 3271 9929
rect 3373 9923 3827 9929
rect 3929 9923 3964 9929
rect 4336 9937 4377 9964
rect 4336 9929 4394 9937
rect 4456 10363 4944 10371
rect 4473 10315 4927 10363
rect 4473 9985 4535 10315
rect 4865 9985 4927 10315
rect 4473 9937 4927 9985
rect 4456 9929 4944 9937
rect 5006 10363 5064 10371
rect 5023 10336 5064 10363
rect 5436 10371 5471 10377
rect 5573 10371 6027 10377
rect 6129 10371 6164 10377
rect 5436 10363 5494 10371
rect 5436 10336 5477 10363
rect 5023 9937 5064 9964
rect 5006 9929 5064 9937
rect 4336 9923 4371 9929
rect 4473 9923 4927 9929
rect 5029 9923 5064 9929
rect 5436 9937 5477 9964
rect 5436 9929 5494 9937
rect 5556 10363 6044 10371
rect 5573 10315 6027 10363
rect 5573 9985 5635 10315
rect 5965 9985 6027 10315
rect 5573 9937 6027 9985
rect 5556 9929 6044 9937
rect 6106 10363 6164 10371
rect 6123 10336 6164 10363
rect 6536 10371 6571 10377
rect 6673 10371 7127 10377
rect 7229 10371 7264 10377
rect 6536 10363 6594 10371
rect 6536 10336 6577 10363
rect 6123 9937 6164 9964
rect 6106 9929 6164 9937
rect 5436 9923 5471 9929
rect 5573 9923 6027 9929
rect 6129 9923 6164 9929
rect 6536 9937 6577 9964
rect 6536 9929 6594 9937
rect 6656 10363 7144 10371
rect 6673 10315 7127 10363
rect 6673 9985 6735 10315
rect 7065 9985 7127 10315
rect 6673 9937 7127 9985
rect 6656 9929 7144 9937
rect 7206 10363 7264 10371
rect 7223 10336 7264 10363
rect 7636 10371 7671 10377
rect 7773 10371 8227 10377
rect 8329 10371 8364 10377
rect 7636 10363 7694 10371
rect 7636 10336 7677 10363
rect 7223 9937 7264 9964
rect 7206 9929 7264 9937
rect 6536 9923 6571 9929
rect 6673 9923 7127 9929
rect 7229 9923 7264 9929
rect 7636 9937 7677 9964
rect 7636 9929 7694 9937
rect 7756 10363 8244 10371
rect 7773 10315 8227 10363
rect 7773 9985 7835 10315
rect 8165 9985 8227 10315
rect 7773 9937 8227 9985
rect 7756 9929 8244 9937
rect 8306 10363 8364 10371
rect 8323 10336 8364 10363
rect 8736 10371 8771 10377
rect 8873 10371 9327 10377
rect 9429 10371 9464 10377
rect 8736 10363 8794 10371
rect 8736 10336 8777 10363
rect 8323 9937 8364 9964
rect 8306 9929 8364 9937
rect 7636 9923 7671 9929
rect 7773 9923 8227 9929
rect 8329 9923 8364 9929
rect 8736 9937 8777 9964
rect 8736 9929 8794 9937
rect 8856 10363 9344 10371
rect 8873 10315 9327 10363
rect 8873 9985 8935 10315
rect 9265 9985 9327 10315
rect 8873 9937 9327 9985
rect 8856 9929 9344 9937
rect 9406 10363 9464 10371
rect 9423 10336 9464 10363
rect 9836 10371 9871 10377
rect 9973 10371 10427 10377
rect 10529 10371 10564 10377
rect 9836 10363 9894 10371
rect 9836 10336 9877 10363
rect 9423 9937 9464 9964
rect 9406 9929 9464 9937
rect 8736 9923 8771 9929
rect 8873 9923 9327 9929
rect 9429 9923 9464 9929
rect 9836 9937 9877 9964
rect 9836 9929 9894 9937
rect 9956 10363 10444 10371
rect 9973 10315 10427 10363
rect 9973 9985 10035 10315
rect 10365 9985 10427 10315
rect 9973 9937 10427 9985
rect 9956 9929 10444 9937
rect 10506 10363 10564 10371
rect 10523 10336 10564 10363
rect 10936 10371 10971 10377
rect 11073 10371 11527 10377
rect 11629 10371 11664 10377
rect 10936 10363 10994 10371
rect 10936 10336 10977 10363
rect 10523 9937 10564 9964
rect 10506 9929 10564 9937
rect 9836 9923 9871 9929
rect 9973 9923 10427 9929
rect 10529 9923 10564 9929
rect 10936 9937 10977 9964
rect 10936 9929 10994 9937
rect 11056 10363 11544 10371
rect 11073 10315 11527 10363
rect 11073 9985 11135 10315
rect 11465 9985 11527 10315
rect 11073 9937 11527 9985
rect 11056 9929 11544 9937
rect 11606 10363 11664 10371
rect 11623 10336 11664 10363
rect 12036 10371 12071 10377
rect 12173 10371 12627 10377
rect 12729 10371 12764 10377
rect 12036 10363 12094 10371
rect 12036 10336 12077 10363
rect 11623 9937 11664 9964
rect 11606 9929 11664 9937
rect 10936 9923 10971 9929
rect 11073 9923 11527 9929
rect 11629 9923 11664 9929
rect 12036 9937 12077 9964
rect 12036 9929 12094 9937
rect 12156 10363 12644 10371
rect 12173 10315 12627 10363
rect 12173 9985 12235 10315
rect 12565 9985 12627 10315
rect 12173 9937 12627 9985
rect 12156 9929 12644 9937
rect 12706 10363 12764 10371
rect 12723 10336 12764 10363
rect 13136 10371 13171 10377
rect 13273 10371 13727 10377
rect 13136 10363 13194 10371
rect 13136 10336 13177 10363
rect 12723 9937 12764 9964
rect 12706 9929 12764 9937
rect 12036 9923 12071 9929
rect 12173 9923 12627 9929
rect 12729 9923 12764 9929
rect 13136 9937 13177 9964
rect 13136 9929 13194 9937
rect 13256 10363 13727 10371
rect 13273 10315 13727 10363
rect 13273 9985 13335 10315
rect 13665 9985 13727 10315
rect 13273 9937 13727 9985
rect 13256 9929 13727 9937
rect 13136 9923 13171 9929
rect 13273 9923 13727 9929
rect -1025 9900 -725 9917
rect -471 9906 -463 9923
rect -37 9906 -29 9923
rect 79 9906 87 9923
rect 513 9906 521 9923
rect 629 9906 637 9923
rect 1063 9906 1071 9923
rect 1179 9906 1187 9923
rect 1613 9906 1621 9923
rect 1729 9906 1737 9923
rect 2163 9906 2171 9923
rect 2279 9906 2287 9923
rect 2713 9906 2721 9923
rect 2829 9906 2837 9923
rect 3263 9906 3271 9923
rect 3379 9906 3387 9923
rect 3813 9906 3821 9923
rect 3929 9906 3937 9923
rect 4363 9906 4371 9923
rect 4479 9906 4487 9923
rect 4913 9906 4921 9923
rect 5029 9906 5037 9923
rect 5463 9906 5471 9923
rect 5579 9906 5587 9923
rect 6013 9906 6021 9923
rect 6129 9906 6137 9923
rect 6563 9906 6571 9923
rect 6679 9906 6687 9923
rect 7113 9906 7121 9923
rect 7229 9906 7237 9923
rect 7663 9906 7671 9923
rect 7779 9906 7787 9923
rect 8213 9906 8221 9923
rect 8329 9906 8337 9923
rect 8763 9906 8771 9923
rect 8879 9906 8887 9923
rect 9313 9906 9321 9923
rect 9429 9906 9437 9923
rect 9863 9906 9871 9923
rect 9979 9906 9987 9923
rect 10413 9906 10421 9923
rect 10529 9906 10537 9923
rect 10963 9906 10971 9923
rect 11079 9906 11087 9923
rect 11513 9906 11521 9923
rect 11629 9906 11637 9923
rect 12063 9906 12071 9923
rect 12179 9906 12187 9923
rect 12613 9906 12621 9923
rect 12729 9906 12737 9923
rect 13163 9906 13171 9923
rect 13279 9906 13287 9923
rect 13713 9906 13721 9923
rect 13975 9917 13987 10450
rect 14263 9917 14275 10450
rect 13975 9900 14275 9917
rect -1025 9367 -1013 9900
rect -737 9367 -725 9900
rect -550 9892 -500 9900
rect -550 9858 -542 9892
rect -508 9858 -500 9892
rect -550 9850 -500 9858
rect 0 9892 50 9900
rect 0 9858 8 9892
rect 42 9858 50 9892
rect 0 9850 50 9858
rect 550 9892 600 9900
rect 550 9858 558 9892
rect 592 9858 600 9892
rect 550 9850 600 9858
rect 1100 9892 1150 9900
rect 1100 9858 1108 9892
rect 1142 9858 1150 9892
rect 1100 9850 1150 9858
rect 1650 9892 1700 9900
rect 1650 9858 1658 9892
rect 1692 9858 1700 9892
rect 1650 9850 1700 9858
rect 2200 9892 2250 9900
rect 2200 9858 2208 9892
rect 2242 9858 2250 9892
rect 2200 9850 2250 9858
rect 2750 9892 2800 9900
rect 2750 9858 2758 9892
rect 2792 9858 2800 9892
rect 2750 9850 2800 9858
rect 3300 9892 3350 9900
rect 3300 9858 3308 9892
rect 3342 9858 3350 9892
rect 3300 9850 3350 9858
rect 3850 9892 3900 9900
rect 3850 9858 3858 9892
rect 3892 9858 3900 9892
rect 3850 9850 3900 9858
rect 4400 9892 4450 9900
rect 4400 9858 4408 9892
rect 4442 9858 4450 9892
rect 4400 9850 4450 9858
rect 4950 9892 5000 9900
rect 4950 9858 4958 9892
rect 4992 9858 5000 9892
rect 4950 9850 5000 9858
rect 5500 9892 5550 9900
rect 5500 9858 5508 9892
rect 5542 9858 5550 9892
rect 5500 9850 5550 9858
rect 6050 9892 6100 9900
rect 6050 9858 6058 9892
rect 6092 9858 6100 9892
rect 6050 9850 6100 9858
rect 6600 9892 6650 9900
rect 6600 9858 6608 9892
rect 6642 9858 6650 9892
rect 6600 9850 6650 9858
rect 7150 9892 7200 9900
rect 7150 9858 7158 9892
rect 7192 9858 7200 9892
rect 7150 9850 7200 9858
rect 7700 9892 7750 9900
rect 7700 9858 7708 9892
rect 7742 9858 7750 9892
rect 7700 9850 7750 9858
rect 8250 9892 8300 9900
rect 8250 9858 8258 9892
rect 8292 9858 8300 9892
rect 8250 9850 8300 9858
rect 8800 9892 8850 9900
rect 8800 9858 8808 9892
rect 8842 9858 8850 9892
rect 8800 9850 8850 9858
rect 9350 9892 9400 9900
rect 9350 9858 9358 9892
rect 9392 9858 9400 9892
rect 9350 9850 9400 9858
rect 9900 9892 9950 9900
rect 9900 9858 9908 9892
rect 9942 9858 9950 9892
rect 9900 9850 9950 9858
rect 10450 9892 10500 9900
rect 10450 9858 10458 9892
rect 10492 9858 10500 9892
rect 10450 9850 10500 9858
rect 11000 9892 11050 9900
rect 11000 9858 11008 9892
rect 11042 9858 11050 9892
rect 11000 9850 11050 9858
rect 11550 9892 11600 9900
rect 11550 9858 11558 9892
rect 11592 9858 11600 9892
rect 11550 9850 11600 9858
rect 12100 9892 12150 9900
rect 12100 9858 12108 9892
rect 12142 9858 12150 9892
rect 12100 9850 12150 9858
rect 12650 9892 12700 9900
rect 12650 9858 12658 9892
rect 12692 9858 12700 9892
rect 12650 9850 12700 9858
rect 13200 9892 13250 9900
rect 13200 9858 13208 9892
rect 13242 9858 13250 9892
rect 13200 9850 13250 9858
rect 13750 9892 13800 9900
rect 13750 9858 13758 9892
rect 13792 9858 13800 9892
rect 13750 9850 13800 9858
rect -471 9827 -463 9844
rect -37 9827 -29 9844
rect 79 9827 87 9844
rect 513 9827 521 9844
rect 629 9827 637 9844
rect 1063 9827 1071 9844
rect 1179 9827 1187 9844
rect 1613 9827 1621 9844
rect 1729 9827 1737 9844
rect 2163 9827 2171 9844
rect 2279 9827 2287 9844
rect 2713 9827 2721 9844
rect 2829 9827 2837 9844
rect 3263 9827 3271 9844
rect 3379 9827 3387 9844
rect 3813 9827 3821 9844
rect 3929 9827 3937 9844
rect 4363 9827 4371 9844
rect 4479 9827 4487 9844
rect 4913 9827 4921 9844
rect 5029 9827 5037 9844
rect 5463 9827 5471 9844
rect 5579 9827 5587 9844
rect 6013 9827 6021 9844
rect 6129 9827 6137 9844
rect 6563 9827 6571 9844
rect 6679 9827 6687 9844
rect 7113 9827 7121 9844
rect 7229 9827 7237 9844
rect 7663 9827 7671 9844
rect 7779 9827 7787 9844
rect 8213 9827 8221 9844
rect 8329 9827 8337 9844
rect 8763 9827 8771 9844
rect 8879 9827 8887 9844
rect 9313 9827 9321 9844
rect 9429 9827 9437 9844
rect 9863 9827 9871 9844
rect 9979 9827 9987 9844
rect 10413 9827 10421 9844
rect 10529 9827 10537 9844
rect 10963 9827 10971 9844
rect 11079 9827 11087 9844
rect 11513 9827 11521 9844
rect 11629 9827 11637 9844
rect 12063 9827 12071 9844
rect 12179 9827 12187 9844
rect 12613 9827 12621 9844
rect 12729 9827 12737 9844
rect 13163 9827 13171 9844
rect 13279 9827 13287 9844
rect 13713 9827 13721 9844
rect -477 9821 -23 9827
rect 79 9821 114 9827
rect -477 9813 -6 9821
rect -477 9765 -23 9813
rect -477 9435 -415 9765
rect -85 9435 -23 9765
rect -477 9387 -23 9435
rect -477 9379 -6 9387
rect 56 9813 114 9821
rect 73 9786 114 9813
rect 486 9821 521 9827
rect 623 9821 1077 9827
rect 1179 9821 1214 9827
rect 486 9813 544 9821
rect 486 9786 527 9813
rect 73 9387 114 9414
rect 56 9379 114 9387
rect -477 9373 -23 9379
rect 79 9373 114 9379
rect 486 9387 527 9414
rect 486 9379 544 9387
rect 606 9813 1094 9821
rect 623 9765 1077 9813
rect 623 9435 685 9765
rect 1015 9435 1077 9765
rect 623 9387 1077 9435
rect 606 9379 1094 9387
rect 1156 9813 1214 9821
rect 1173 9786 1214 9813
rect 1586 9821 1621 9827
rect 1723 9821 2177 9827
rect 2279 9821 2314 9827
rect 1586 9813 1644 9821
rect 1586 9786 1627 9813
rect 1173 9387 1214 9414
rect 1156 9379 1214 9387
rect 486 9373 521 9379
rect 623 9373 1077 9379
rect 1179 9373 1214 9379
rect 1586 9387 1627 9414
rect 1586 9379 1644 9387
rect 1706 9813 2194 9821
rect 1723 9765 2177 9813
rect 1723 9435 1785 9765
rect 2115 9435 2177 9765
rect 1723 9387 2177 9435
rect 1706 9379 2194 9387
rect 2256 9813 2314 9821
rect 2273 9786 2314 9813
rect 2686 9821 2721 9827
rect 2823 9821 3277 9827
rect 3379 9821 3414 9827
rect 2686 9813 2744 9821
rect 2686 9786 2727 9813
rect 2273 9387 2314 9414
rect 2256 9379 2314 9387
rect 1586 9373 1621 9379
rect 1723 9373 2177 9379
rect 2279 9373 2314 9379
rect 2686 9387 2727 9414
rect 2686 9379 2744 9387
rect 2806 9813 3294 9821
rect 2823 9765 3277 9813
rect 2823 9435 2885 9765
rect 3215 9435 3277 9765
rect 2823 9387 3277 9435
rect 2806 9379 3294 9387
rect 3356 9813 3414 9821
rect 3373 9786 3414 9813
rect 3786 9821 3821 9827
rect 3923 9821 4377 9827
rect 4479 9821 4514 9827
rect 3786 9813 3844 9821
rect 3786 9786 3827 9813
rect 3373 9387 3414 9414
rect 3356 9379 3414 9387
rect 2686 9373 2721 9379
rect 2823 9373 3277 9379
rect 3379 9373 3414 9379
rect 3786 9387 3827 9414
rect 3786 9379 3844 9387
rect 3906 9813 4394 9821
rect 3923 9765 4377 9813
rect 3923 9435 3985 9765
rect 4315 9435 4377 9765
rect 3923 9387 4377 9435
rect 3906 9379 4394 9387
rect 4456 9813 4514 9821
rect 4473 9786 4514 9813
rect 4886 9821 4921 9827
rect 5023 9821 5477 9827
rect 5579 9821 5614 9827
rect 4886 9813 4944 9821
rect 4886 9786 4927 9813
rect 4473 9387 4514 9414
rect 4456 9379 4514 9387
rect 3786 9373 3821 9379
rect 3923 9373 4377 9379
rect 4479 9373 4514 9379
rect 4886 9387 4927 9414
rect 4886 9379 4944 9387
rect 5006 9813 5494 9821
rect 5023 9765 5477 9813
rect 5023 9435 5085 9765
rect 5415 9435 5477 9765
rect 5023 9387 5477 9435
rect 5006 9379 5494 9387
rect 5556 9813 5614 9821
rect 5573 9786 5614 9813
rect 5986 9821 6021 9827
rect 6123 9821 6577 9827
rect 6679 9821 6714 9827
rect 5986 9813 6044 9821
rect 5986 9786 6027 9813
rect 5573 9387 5614 9414
rect 5556 9379 5614 9387
rect 4886 9373 4921 9379
rect 5023 9373 5477 9379
rect 5579 9373 5614 9379
rect 5986 9387 6027 9414
rect 5986 9379 6044 9387
rect 6106 9813 6594 9821
rect 6123 9765 6577 9813
rect 6123 9435 6185 9765
rect 6515 9435 6577 9765
rect 6123 9387 6577 9435
rect 6106 9379 6594 9387
rect 6656 9813 6714 9821
rect 6673 9786 6714 9813
rect 7086 9821 7121 9827
rect 7223 9821 7677 9827
rect 7779 9821 7814 9827
rect 7086 9813 7144 9821
rect 7086 9786 7127 9813
rect 6673 9387 6714 9414
rect 6656 9379 6714 9387
rect 5986 9373 6021 9379
rect 6123 9373 6577 9379
rect 6679 9373 6714 9379
rect 7086 9387 7127 9414
rect 7086 9379 7144 9387
rect 7206 9813 7694 9821
rect 7223 9765 7677 9813
rect 7223 9435 7285 9765
rect 7615 9435 7677 9765
rect 7223 9387 7677 9435
rect 7206 9379 7694 9387
rect 7756 9813 7814 9821
rect 7773 9786 7814 9813
rect 8186 9821 8221 9827
rect 8323 9821 8777 9827
rect 8879 9821 8914 9827
rect 8186 9813 8244 9821
rect 8186 9786 8227 9813
rect 7773 9387 7814 9414
rect 7756 9379 7814 9387
rect 7086 9373 7121 9379
rect 7223 9373 7677 9379
rect 7779 9373 7814 9379
rect 8186 9387 8227 9414
rect 8186 9379 8244 9387
rect 8306 9813 8794 9821
rect 8323 9765 8777 9813
rect 8323 9435 8385 9765
rect 8715 9435 8777 9765
rect 8323 9387 8777 9435
rect 8306 9379 8794 9387
rect 8856 9813 8914 9821
rect 8873 9786 8914 9813
rect 9286 9821 9321 9827
rect 9423 9821 9877 9827
rect 9979 9821 10014 9827
rect 9286 9813 9344 9821
rect 9286 9786 9327 9813
rect 8873 9387 8914 9414
rect 8856 9379 8914 9387
rect 8186 9373 8221 9379
rect 8323 9373 8777 9379
rect 8879 9373 8914 9379
rect 9286 9387 9327 9414
rect 9286 9379 9344 9387
rect 9406 9813 9894 9821
rect 9423 9765 9877 9813
rect 9423 9435 9485 9765
rect 9815 9435 9877 9765
rect 9423 9387 9877 9435
rect 9406 9379 9894 9387
rect 9956 9813 10014 9821
rect 9973 9786 10014 9813
rect 10386 9821 10421 9827
rect 10523 9821 10977 9827
rect 11079 9821 11114 9827
rect 10386 9813 10444 9821
rect 10386 9786 10427 9813
rect 9973 9387 10014 9414
rect 9956 9379 10014 9387
rect 9286 9373 9321 9379
rect 9423 9373 9877 9379
rect 9979 9373 10014 9379
rect 10386 9387 10427 9414
rect 10386 9379 10444 9387
rect 10506 9813 10994 9821
rect 10523 9765 10977 9813
rect 10523 9435 10585 9765
rect 10915 9435 10977 9765
rect 10523 9387 10977 9435
rect 10506 9379 10994 9387
rect 11056 9813 11114 9821
rect 11073 9786 11114 9813
rect 11486 9821 11521 9827
rect 11623 9821 12077 9827
rect 12179 9821 12214 9827
rect 11486 9813 11544 9821
rect 11486 9786 11527 9813
rect 11073 9387 11114 9414
rect 11056 9379 11114 9387
rect 10386 9373 10421 9379
rect 10523 9373 10977 9379
rect 11079 9373 11114 9379
rect 11486 9387 11527 9414
rect 11486 9379 11544 9387
rect 11606 9813 12094 9821
rect 11623 9765 12077 9813
rect 11623 9435 11685 9765
rect 12015 9435 12077 9765
rect 11623 9387 12077 9435
rect 11606 9379 12094 9387
rect 12156 9813 12214 9821
rect 12173 9786 12214 9813
rect 12586 9821 12621 9827
rect 12723 9821 13177 9827
rect 13279 9821 13314 9827
rect 12586 9813 12644 9821
rect 12586 9786 12627 9813
rect 12173 9387 12214 9414
rect 12156 9379 12214 9387
rect 11486 9373 11521 9379
rect 11623 9373 12077 9379
rect 12179 9373 12214 9379
rect 12586 9387 12627 9414
rect 12586 9379 12644 9387
rect 12706 9813 13194 9821
rect 12723 9765 13177 9813
rect 12723 9435 12785 9765
rect 13115 9435 13177 9765
rect 12723 9387 13177 9435
rect 12706 9379 13194 9387
rect 13256 9813 13314 9821
rect 13273 9786 13314 9813
rect 13273 9387 13314 9414
rect 13256 9379 13314 9387
rect 12586 9373 12621 9379
rect 12723 9373 13177 9379
rect 13279 9373 13314 9379
rect -1025 9350 -725 9367
rect -471 9356 -463 9373
rect -37 9356 -29 9373
rect 79 9356 87 9373
rect 513 9356 521 9373
rect 629 9356 637 9373
rect 1063 9356 1071 9373
rect 1179 9356 1187 9373
rect 1613 9356 1621 9373
rect 1729 9356 1737 9373
rect 2163 9356 2171 9373
rect 2279 9356 2287 9373
rect 2713 9356 2721 9373
rect 2829 9356 2837 9373
rect 3263 9356 3271 9373
rect 3379 9356 3387 9373
rect 3813 9356 3821 9373
rect 3929 9356 3937 9373
rect 4363 9356 4371 9373
rect 4479 9356 4487 9373
rect 4913 9356 4921 9373
rect 5029 9356 5037 9373
rect 5463 9356 5471 9373
rect 5579 9356 5587 9373
rect 6013 9356 6021 9373
rect 6129 9356 6137 9373
rect 6563 9356 6571 9373
rect 6679 9356 6687 9373
rect 7113 9356 7121 9373
rect 7229 9356 7237 9373
rect 7663 9356 7671 9373
rect 7779 9356 7787 9373
rect 8213 9356 8221 9373
rect 8329 9356 8337 9373
rect 8763 9356 8771 9373
rect 8879 9356 8887 9373
rect 9313 9356 9321 9373
rect 9429 9356 9437 9373
rect 9863 9356 9871 9373
rect 9979 9356 9987 9373
rect 10413 9356 10421 9373
rect 10529 9356 10537 9373
rect 10963 9356 10971 9373
rect 11079 9356 11087 9373
rect 11513 9356 11521 9373
rect 11629 9356 11637 9373
rect 12063 9356 12071 9373
rect 12179 9356 12187 9373
rect 12613 9356 12621 9373
rect 12729 9356 12737 9373
rect 13163 9356 13171 9373
rect 13279 9356 13287 9373
rect 13713 9356 13721 9373
rect 13975 9369 13987 9900
rect 14263 9369 14275 9900
rect 13975 9350 14275 9369
rect -1025 8817 -1013 9350
rect -737 8817 -725 9350
rect -550 9342 -500 9350
rect -550 9308 -542 9342
rect -508 9308 -500 9342
rect -550 9300 -500 9308
rect 0 9342 50 9350
rect 0 9308 8 9342
rect 42 9308 50 9342
rect 0 9300 50 9308
rect 550 9342 600 9350
rect 550 9308 558 9342
rect 592 9308 600 9342
rect 550 9300 600 9308
rect 1100 9342 1150 9350
rect 1100 9308 1108 9342
rect 1142 9308 1150 9342
rect 1100 9300 1150 9308
rect 1650 9342 1700 9350
rect 1650 9308 1658 9342
rect 1692 9308 1700 9342
rect 1650 9300 1700 9308
rect 2200 9342 2250 9350
rect 2200 9308 2208 9342
rect 2242 9308 2250 9342
rect 2200 9300 2250 9308
rect 2750 9342 2800 9350
rect 2750 9308 2758 9342
rect 2792 9308 2800 9342
rect 2750 9300 2800 9308
rect 3300 9342 3350 9350
rect 3300 9308 3308 9342
rect 3342 9308 3350 9342
rect 3300 9300 3350 9308
rect 3850 9342 3900 9350
rect 3850 9308 3858 9342
rect 3892 9308 3900 9342
rect 3850 9300 3900 9308
rect 4400 9342 4450 9350
rect 4400 9308 4408 9342
rect 4442 9308 4450 9342
rect 4400 9300 4450 9308
rect 4950 9342 5000 9350
rect 4950 9308 4958 9342
rect 4992 9308 5000 9342
rect 4950 9300 5000 9308
rect 5500 9342 5550 9350
rect 5500 9308 5508 9342
rect 5542 9308 5550 9342
rect 5500 9300 5550 9308
rect 6050 9342 6100 9350
rect 6050 9308 6058 9342
rect 6092 9308 6100 9342
rect 6050 9300 6100 9308
rect 6600 9342 6650 9350
rect 6600 9308 6608 9342
rect 6642 9308 6650 9342
rect 6600 9300 6650 9308
rect 7150 9342 7200 9350
rect 7150 9308 7158 9342
rect 7192 9308 7200 9342
rect 7150 9300 7200 9308
rect 7700 9342 7750 9350
rect 7700 9308 7708 9342
rect 7742 9308 7750 9342
rect 7700 9300 7750 9308
rect 8250 9342 8300 9350
rect 8250 9308 8258 9342
rect 8292 9308 8300 9342
rect 8250 9300 8300 9308
rect 8800 9342 8850 9350
rect 8800 9308 8808 9342
rect 8842 9308 8850 9342
rect 8800 9300 8850 9308
rect 9350 9342 9400 9350
rect 9350 9308 9358 9342
rect 9392 9308 9400 9342
rect 9350 9300 9400 9308
rect 9900 9342 9950 9350
rect 9900 9308 9908 9342
rect 9942 9308 9950 9342
rect 9900 9300 9950 9308
rect 10450 9342 10500 9350
rect 10450 9308 10458 9342
rect 10492 9308 10500 9342
rect 10450 9300 10500 9308
rect 11000 9342 11050 9350
rect 11000 9308 11008 9342
rect 11042 9308 11050 9342
rect 11000 9300 11050 9308
rect 11550 9342 11600 9350
rect 11550 9308 11558 9342
rect 11592 9308 11600 9342
rect 11550 9300 11600 9308
rect 12100 9342 12150 9350
rect 12100 9308 12108 9342
rect 12142 9308 12150 9342
rect 12100 9300 12150 9308
rect 12650 9342 12700 9350
rect 12650 9308 12658 9342
rect 12692 9308 12700 9342
rect 12650 9300 12700 9308
rect 13200 9342 13250 9350
rect 13200 9308 13208 9342
rect 13242 9308 13250 9342
rect 13200 9300 13250 9308
rect 13750 9342 13800 9350
rect 13750 9308 13758 9342
rect 13792 9308 13800 9342
rect 13750 9300 13800 9308
rect -471 9277 -463 9294
rect -37 9277 -29 9294
rect 79 9277 87 9294
rect 513 9277 521 9294
rect 629 9277 637 9294
rect 1063 9277 1071 9294
rect 1179 9277 1187 9294
rect 1613 9277 1621 9294
rect 1729 9277 1737 9294
rect 2163 9277 2171 9294
rect 2279 9277 2287 9294
rect 2713 9277 2721 9294
rect 2829 9277 2837 9294
rect 3263 9277 3271 9294
rect 3379 9277 3387 9294
rect 3813 9277 3821 9294
rect 3929 9277 3937 9294
rect 4363 9277 4371 9294
rect 4479 9277 4487 9294
rect 4913 9277 4921 9294
rect 5029 9277 5037 9294
rect 5463 9277 5471 9294
rect 5579 9277 5587 9294
rect 6013 9277 6021 9294
rect 6129 9277 6137 9294
rect 6563 9277 6571 9294
rect 6679 9277 6687 9294
rect 7113 9277 7121 9294
rect 7229 9277 7237 9294
rect 7663 9277 7671 9294
rect 7779 9277 7787 9294
rect 8213 9277 8221 9294
rect 8329 9277 8337 9294
rect 8763 9277 8771 9294
rect 8879 9277 8887 9294
rect 9313 9277 9321 9294
rect 9429 9277 9437 9294
rect 9863 9277 9871 9294
rect 9979 9277 9987 9294
rect 10413 9277 10421 9294
rect 10529 9277 10537 9294
rect 10963 9277 10971 9294
rect 11079 9277 11087 9294
rect 11513 9277 11521 9294
rect 11629 9277 11637 9294
rect 12063 9277 12071 9294
rect 12179 9277 12187 9294
rect 12613 9277 12621 9294
rect 12729 9277 12737 9294
rect 13163 9277 13171 9294
rect 13279 9277 13287 9294
rect 13713 9277 13721 9294
rect -64 9271 -29 9277
rect 73 9271 527 9277
rect 629 9271 664 9277
rect -64 9263 -6 9271
rect -64 9236 -23 9263
rect -64 8837 -23 8864
rect -64 8829 -6 8837
rect 56 9263 544 9271
rect 73 9215 527 9263
rect 73 8885 135 9215
rect 465 8885 527 9215
rect 73 8837 527 8885
rect 56 8829 544 8837
rect 606 9263 664 9271
rect 623 9236 664 9263
rect 1036 9271 1071 9277
rect 1173 9271 1627 9277
rect 1729 9271 1764 9277
rect 1036 9263 1094 9271
rect 1036 9236 1077 9263
rect 623 8837 664 8864
rect 606 8829 664 8837
rect -64 8823 -29 8829
rect 73 8823 527 8829
rect 629 8823 664 8829
rect 1036 8837 1077 8864
rect 1036 8829 1094 8837
rect 1156 9263 1644 9271
rect 1173 9215 1627 9263
rect 1173 8885 1235 9215
rect 1565 8885 1627 9215
rect 1173 8837 1627 8885
rect 1156 8829 1644 8837
rect 1706 9263 1764 9271
rect 1723 9236 1764 9263
rect 2136 9271 2171 9277
rect 2273 9271 2727 9277
rect 2829 9271 2864 9277
rect 2136 9263 2194 9271
rect 2136 9236 2177 9263
rect 1723 8837 1764 8864
rect 1706 8829 1764 8837
rect 1036 8823 1071 8829
rect 1173 8823 1627 8829
rect 1729 8823 1764 8829
rect 2136 8837 2177 8864
rect 2136 8829 2194 8837
rect 2256 9263 2744 9271
rect 2273 9215 2727 9263
rect 2273 8885 2335 9215
rect 2665 8885 2727 9215
rect 2273 8837 2727 8885
rect 2256 8829 2744 8837
rect 2806 9263 2864 9271
rect 2823 9236 2864 9263
rect 3236 9271 3271 9277
rect 3373 9271 3827 9277
rect 3929 9271 3964 9277
rect 3236 9263 3294 9271
rect 3236 9236 3277 9263
rect 2823 8837 2864 8864
rect 2806 8829 2864 8837
rect 2136 8823 2171 8829
rect 2273 8823 2727 8829
rect 2829 8823 2864 8829
rect 3236 8837 3277 8864
rect 3236 8829 3294 8837
rect 3356 9263 3844 9271
rect 3373 9215 3827 9263
rect 3373 8885 3435 9215
rect 3765 8885 3827 9215
rect 3373 8837 3827 8885
rect 3356 8829 3844 8837
rect 3906 9263 3964 9271
rect 3923 9236 3964 9263
rect 4336 9271 4371 9277
rect 4473 9271 4927 9277
rect 5029 9271 5064 9277
rect 4336 9263 4394 9271
rect 4336 9236 4377 9263
rect 3923 8837 3964 8864
rect 3906 8829 3964 8837
rect 3236 8823 3271 8829
rect 3373 8823 3827 8829
rect 3929 8823 3964 8829
rect 4336 8837 4377 8864
rect 4336 8829 4394 8837
rect 4456 9263 4944 9271
rect 4473 9215 4927 9263
rect 4473 8885 4535 9215
rect 4865 8885 4927 9215
rect 4473 8837 4927 8885
rect 4456 8829 4944 8837
rect 5006 9263 5064 9271
rect 5023 9236 5064 9263
rect 5436 9271 5471 9277
rect 5573 9271 6027 9277
rect 6129 9271 6164 9277
rect 5436 9263 5494 9271
rect 5436 9236 5477 9263
rect 5023 8837 5064 8864
rect 5006 8829 5064 8837
rect 4336 8823 4371 8829
rect 4473 8823 4927 8829
rect 5029 8823 5064 8829
rect 5436 8837 5477 8864
rect 5436 8829 5494 8837
rect 5556 9263 6044 9271
rect 5573 9215 6027 9263
rect 5573 8885 5635 9215
rect 5965 8885 6027 9215
rect 5573 8837 6027 8885
rect 5556 8829 6044 8837
rect 6106 9263 6164 9271
rect 6123 9236 6164 9263
rect 6536 9271 6571 9277
rect 6673 9271 7127 9277
rect 7229 9271 7264 9277
rect 6536 9263 6594 9271
rect 6536 9236 6577 9263
rect 6123 8837 6164 8864
rect 6106 8829 6164 8837
rect 5436 8823 5471 8829
rect 5573 8823 6027 8829
rect 6129 8823 6164 8829
rect 6536 8837 6577 8864
rect 6536 8829 6594 8837
rect 6656 9263 7144 9271
rect 6673 9215 7127 9263
rect 6673 8885 6735 9215
rect 7065 8885 7127 9215
rect 6673 8837 7127 8885
rect 6656 8829 7144 8837
rect 7206 9263 7264 9271
rect 7223 9236 7264 9263
rect 7636 9271 7671 9277
rect 7773 9271 8227 9277
rect 8329 9271 8364 9277
rect 7636 9263 7694 9271
rect 7636 9236 7677 9263
rect 7223 8837 7264 8864
rect 7206 8829 7264 8837
rect 6536 8823 6571 8829
rect 6673 8823 7127 8829
rect 7229 8823 7264 8829
rect 7636 8837 7677 8864
rect 7636 8829 7694 8837
rect 7756 9263 8244 9271
rect 7773 9215 8227 9263
rect 7773 8885 7835 9215
rect 8165 8885 8227 9215
rect 7773 8837 8227 8885
rect 7756 8829 8244 8837
rect 8306 9263 8364 9271
rect 8323 9236 8364 9263
rect 8736 9271 8771 9277
rect 8873 9271 9327 9277
rect 9429 9271 9464 9277
rect 8736 9263 8794 9271
rect 8736 9236 8777 9263
rect 8323 8837 8364 8864
rect 8306 8829 8364 8837
rect 7636 8823 7671 8829
rect 7773 8823 8227 8829
rect 8329 8823 8364 8829
rect 8736 8837 8777 8864
rect 8736 8829 8794 8837
rect 8856 9263 9344 9271
rect 8873 9215 9327 9263
rect 8873 8885 8935 9215
rect 9265 8885 9327 9215
rect 8873 8837 9327 8885
rect 8856 8829 9344 8837
rect 9406 9263 9464 9271
rect 9423 9236 9464 9263
rect 9836 9271 9871 9277
rect 9973 9271 10427 9277
rect 10529 9271 10564 9277
rect 9836 9263 9894 9271
rect 9836 9236 9877 9263
rect 9423 8837 9464 8864
rect 9406 8829 9464 8837
rect 8736 8823 8771 8829
rect 8873 8823 9327 8829
rect 9429 8823 9464 8829
rect 9836 8837 9877 8864
rect 9836 8829 9894 8837
rect 9956 9263 10444 9271
rect 9973 9215 10427 9263
rect 9973 8885 10035 9215
rect 10365 8885 10427 9215
rect 9973 8837 10427 8885
rect 9956 8829 10444 8837
rect 10506 9263 10564 9271
rect 10523 9236 10564 9263
rect 10936 9271 10971 9277
rect 11073 9271 11527 9277
rect 11629 9271 11664 9277
rect 10936 9263 10994 9271
rect 10936 9236 10977 9263
rect 10523 8837 10564 8864
rect 10506 8829 10564 8837
rect 9836 8823 9871 8829
rect 9973 8823 10427 8829
rect 10529 8823 10564 8829
rect 10936 8837 10977 8864
rect 10936 8829 10994 8837
rect 11056 9263 11544 9271
rect 11073 9215 11527 9263
rect 11073 8885 11135 9215
rect 11465 8885 11527 9215
rect 11073 8837 11527 8885
rect 11056 8829 11544 8837
rect 11606 9263 11664 9271
rect 11623 9236 11664 9263
rect 12036 9271 12071 9277
rect 12173 9271 12627 9277
rect 12729 9271 12764 9277
rect 12036 9263 12094 9271
rect 12036 9236 12077 9263
rect 11623 8837 11664 8864
rect 11606 8829 11664 8837
rect 10936 8823 10971 8829
rect 11073 8823 11527 8829
rect 11629 8823 11664 8829
rect 12036 8837 12077 8864
rect 12036 8829 12094 8837
rect 12156 9263 12644 9271
rect 12173 9215 12627 9263
rect 12173 8885 12235 9215
rect 12565 8885 12627 9215
rect 12173 8837 12627 8885
rect 12156 8829 12644 8837
rect 12706 9263 12764 9271
rect 12723 9236 12764 9263
rect 13136 9271 13171 9277
rect 13273 9271 13727 9277
rect 13136 9263 13194 9271
rect 13136 9236 13177 9263
rect 12723 8837 12764 8864
rect 12706 8829 12764 8837
rect 12036 8823 12071 8829
rect 12173 8823 12627 8829
rect 12729 8823 12764 8829
rect 13136 8837 13177 8864
rect 13136 8829 13194 8837
rect 13256 9263 13727 9271
rect 13273 9215 13727 9263
rect 13273 8885 13335 9215
rect 13665 8885 13727 9215
rect 13273 8837 13727 8885
rect 13256 8829 13727 8837
rect 13136 8823 13171 8829
rect 13273 8823 13727 8829
rect -1025 8800 -725 8817
rect -471 8806 -463 8823
rect -37 8806 -29 8823
rect 79 8806 87 8823
rect 513 8806 521 8823
rect 629 8806 637 8823
rect 1063 8806 1071 8823
rect 1179 8806 1187 8823
rect 1613 8806 1621 8823
rect 1729 8806 1737 8823
rect 2163 8806 2171 8823
rect 2279 8806 2287 8823
rect 2713 8806 2721 8823
rect 2829 8806 2837 8823
rect 3263 8806 3271 8823
rect 3379 8806 3387 8823
rect 3813 8806 3821 8823
rect 3929 8806 3937 8823
rect 4363 8806 4371 8823
rect 4479 8806 4487 8823
rect 4913 8806 4921 8823
rect 5029 8806 5037 8823
rect 5463 8806 5471 8823
rect 5579 8806 5587 8823
rect 6013 8806 6021 8823
rect 6129 8806 6137 8823
rect 6563 8806 6571 8823
rect 6679 8806 6687 8823
rect 7113 8806 7121 8823
rect 7229 8806 7237 8823
rect 7663 8806 7671 8823
rect 7779 8806 7787 8823
rect 8213 8806 8221 8823
rect 8329 8806 8337 8823
rect 8763 8806 8771 8823
rect 8879 8806 8887 8823
rect 9313 8806 9321 8823
rect 9429 8806 9437 8823
rect 9863 8806 9871 8823
rect 9979 8806 9987 8823
rect 10413 8806 10421 8823
rect 10529 8806 10537 8823
rect 10963 8806 10971 8823
rect 11079 8806 11087 8823
rect 11513 8806 11521 8823
rect 11629 8806 11637 8823
rect 12063 8806 12071 8823
rect 12179 8806 12187 8823
rect 12613 8806 12621 8823
rect 12729 8806 12737 8823
rect 13163 8806 13171 8823
rect 13279 8806 13287 8823
rect 13713 8806 13721 8823
rect 13975 8817 13987 9350
rect 14263 8817 14275 9350
rect 13975 8800 14275 8817
rect -1025 8267 -1013 8800
rect -737 8267 -725 8800
rect -550 8792 -500 8800
rect -550 8758 -542 8792
rect -508 8758 -500 8792
rect -550 8750 -500 8758
rect 0 8792 50 8800
rect 0 8758 8 8792
rect 42 8758 50 8792
rect 0 8750 50 8758
rect 550 8792 600 8800
rect 550 8758 558 8792
rect 592 8758 600 8792
rect 550 8750 600 8758
rect 1100 8792 1150 8800
rect 1100 8758 1108 8792
rect 1142 8758 1150 8792
rect 1100 8750 1150 8758
rect 1650 8792 1700 8800
rect 1650 8758 1658 8792
rect 1692 8758 1700 8792
rect 1650 8750 1700 8758
rect 2200 8792 2250 8800
rect 2200 8758 2208 8792
rect 2242 8758 2250 8792
rect 2200 8750 2250 8758
rect 2750 8792 2800 8800
rect 2750 8758 2758 8792
rect 2792 8758 2800 8792
rect 2750 8750 2800 8758
rect 3300 8792 3350 8800
rect 3300 8758 3308 8792
rect 3342 8758 3350 8792
rect 3300 8750 3350 8758
rect 3850 8792 3900 8800
rect 3850 8758 3858 8792
rect 3892 8758 3900 8792
rect 3850 8750 3900 8758
rect 4400 8792 4450 8800
rect 4400 8758 4408 8792
rect 4442 8758 4450 8792
rect 4400 8750 4450 8758
rect 4950 8792 5000 8800
rect 4950 8758 4958 8792
rect 4992 8758 5000 8792
rect 4950 8750 5000 8758
rect 5500 8792 5550 8800
rect 5500 8758 5508 8792
rect 5542 8758 5550 8792
rect 5500 8750 5550 8758
rect 6050 8792 6100 8800
rect 6050 8758 6058 8792
rect 6092 8758 6100 8792
rect 6050 8750 6100 8758
rect 6600 8792 6650 8800
rect 6600 8758 6608 8792
rect 6642 8758 6650 8792
rect 6600 8750 6650 8758
rect 7150 8792 7200 8800
rect 7150 8758 7158 8792
rect 7192 8758 7200 8792
rect 7150 8750 7200 8758
rect 7700 8792 7750 8800
rect 7700 8758 7708 8792
rect 7742 8758 7750 8792
rect 7700 8750 7750 8758
rect 8250 8792 8300 8800
rect 8250 8758 8258 8792
rect 8292 8758 8300 8792
rect 8250 8750 8300 8758
rect 8800 8792 8850 8800
rect 8800 8758 8808 8792
rect 8842 8758 8850 8792
rect 8800 8750 8850 8758
rect 9350 8792 9400 8800
rect 9350 8758 9358 8792
rect 9392 8758 9400 8792
rect 9350 8750 9400 8758
rect 9900 8792 9950 8800
rect 9900 8758 9908 8792
rect 9942 8758 9950 8792
rect 9900 8750 9950 8758
rect 10450 8792 10500 8800
rect 10450 8758 10458 8792
rect 10492 8758 10500 8792
rect 10450 8750 10500 8758
rect 11000 8792 11050 8800
rect 11000 8758 11008 8792
rect 11042 8758 11050 8792
rect 11000 8750 11050 8758
rect 11550 8792 11600 8800
rect 11550 8758 11558 8792
rect 11592 8758 11600 8792
rect 11550 8750 11600 8758
rect 12100 8792 12150 8800
rect 12100 8758 12108 8792
rect 12142 8758 12150 8792
rect 12100 8750 12150 8758
rect 12650 8792 12700 8800
rect 12650 8758 12658 8792
rect 12692 8758 12700 8792
rect 12650 8750 12700 8758
rect 13200 8792 13250 8800
rect 13200 8758 13208 8792
rect 13242 8758 13250 8792
rect 13200 8750 13250 8758
rect 13750 8792 13800 8800
rect 13750 8758 13758 8792
rect 13792 8758 13800 8792
rect 13750 8750 13800 8758
rect -471 8727 -463 8744
rect -37 8727 -29 8744
rect 79 8727 87 8744
rect 513 8727 521 8744
rect 629 8727 637 8744
rect 1063 8727 1071 8744
rect 1179 8727 1187 8744
rect 1613 8727 1621 8744
rect 1729 8727 1737 8744
rect 2163 8727 2171 8744
rect 2279 8727 2287 8744
rect 2713 8727 2721 8744
rect 2829 8727 2837 8744
rect 3263 8727 3271 8744
rect 3379 8727 3387 8744
rect 3813 8727 3821 8744
rect 3929 8727 3937 8744
rect 4363 8727 4371 8744
rect 4479 8727 4487 8744
rect 4913 8727 4921 8744
rect 5029 8727 5037 8744
rect 5463 8727 5471 8744
rect 5579 8727 5587 8744
rect 6013 8727 6021 8744
rect 6129 8727 6137 8744
rect 6563 8727 6571 8744
rect 6679 8727 6687 8744
rect 7113 8727 7121 8744
rect 7229 8727 7237 8744
rect 7663 8727 7671 8744
rect 7779 8727 7787 8744
rect 8213 8727 8221 8744
rect 8329 8727 8337 8744
rect 8763 8727 8771 8744
rect 8879 8727 8887 8744
rect 9313 8727 9321 8744
rect 9429 8727 9437 8744
rect 9863 8727 9871 8744
rect 9979 8727 9987 8744
rect 10413 8727 10421 8744
rect 10529 8727 10537 8744
rect 10963 8727 10971 8744
rect 11079 8727 11087 8744
rect 11513 8727 11521 8744
rect 11629 8727 11637 8744
rect 12063 8727 12071 8744
rect 12179 8727 12187 8744
rect 12613 8727 12621 8744
rect 12729 8727 12737 8744
rect 13163 8727 13171 8744
rect 13279 8727 13287 8744
rect 13713 8727 13721 8744
rect -477 8721 -23 8727
rect 79 8721 114 8727
rect -477 8713 -6 8721
rect -477 8665 -23 8713
rect -477 8335 -415 8665
rect -85 8335 -23 8665
rect -477 8287 -23 8335
rect -477 8279 -6 8287
rect 56 8713 114 8721
rect 73 8686 114 8713
rect 486 8721 521 8727
rect 623 8721 1077 8727
rect 1179 8721 1214 8727
rect 486 8713 544 8721
rect 486 8686 527 8713
rect 73 8287 114 8314
rect 56 8279 114 8287
rect -477 8273 -23 8279
rect 79 8273 114 8279
rect 486 8287 527 8314
rect 486 8279 544 8287
rect 606 8713 1094 8721
rect 623 8665 1077 8713
rect 623 8335 685 8665
rect 1015 8335 1077 8665
rect 623 8287 1077 8335
rect 606 8279 1094 8287
rect 1156 8713 1214 8721
rect 1173 8686 1214 8713
rect 1586 8721 1621 8727
rect 1723 8721 2177 8727
rect 2279 8721 2314 8727
rect 1586 8713 1644 8721
rect 1586 8686 1627 8713
rect 1173 8287 1214 8314
rect 1156 8279 1214 8287
rect 486 8273 521 8279
rect 623 8273 1077 8279
rect 1179 8273 1214 8279
rect 1586 8287 1627 8314
rect 1586 8279 1644 8287
rect 1706 8713 2194 8721
rect 1723 8665 2177 8713
rect 1723 8335 1785 8665
rect 2115 8335 2177 8665
rect 1723 8287 2177 8335
rect 1706 8279 2194 8287
rect 2256 8713 2314 8721
rect 2273 8686 2314 8713
rect 2686 8721 2721 8727
rect 2823 8721 3277 8727
rect 3379 8721 3414 8727
rect 2686 8713 2744 8721
rect 2686 8686 2727 8713
rect 2273 8287 2314 8314
rect 2256 8279 2314 8287
rect 1586 8273 1621 8279
rect 1723 8273 2177 8279
rect 2279 8273 2314 8279
rect 2686 8287 2727 8314
rect 2686 8279 2744 8287
rect 2806 8713 3294 8721
rect 2823 8665 3277 8713
rect 2823 8335 2885 8665
rect 3215 8335 3277 8665
rect 2823 8287 3277 8335
rect 2806 8279 3294 8287
rect 3356 8713 3414 8721
rect 3373 8686 3414 8713
rect 3786 8721 3821 8727
rect 3923 8721 4377 8727
rect 4479 8721 4514 8727
rect 3786 8713 3844 8721
rect 3786 8686 3827 8713
rect 3373 8287 3414 8314
rect 3356 8279 3414 8287
rect 2686 8273 2721 8279
rect 2823 8273 3277 8279
rect 3379 8273 3414 8279
rect 3786 8287 3827 8314
rect 3786 8279 3844 8287
rect 3906 8713 4394 8721
rect 3923 8665 4377 8713
rect 3923 8335 3985 8665
rect 4315 8335 4377 8665
rect 3923 8287 4377 8335
rect 3906 8279 4394 8287
rect 4456 8713 4514 8721
rect 4473 8686 4514 8713
rect 4886 8721 4921 8727
rect 5023 8721 5477 8727
rect 5579 8721 5614 8727
rect 4886 8713 4944 8721
rect 4886 8686 4927 8713
rect 4473 8287 4514 8314
rect 4456 8279 4514 8287
rect 3786 8273 3821 8279
rect 3923 8273 4377 8279
rect 4479 8273 4514 8279
rect 4886 8287 4927 8314
rect 4886 8279 4944 8287
rect 5006 8713 5494 8721
rect 5023 8665 5477 8713
rect 5023 8335 5085 8665
rect 5415 8335 5477 8665
rect 5023 8287 5477 8335
rect 5006 8279 5494 8287
rect 5556 8713 5614 8721
rect 5573 8686 5614 8713
rect 5986 8721 6021 8727
rect 6123 8721 6577 8727
rect 6679 8721 6714 8727
rect 5986 8713 6044 8721
rect 5986 8686 6027 8713
rect 5573 8287 5614 8314
rect 5556 8279 5614 8287
rect 4886 8273 4921 8279
rect 5023 8273 5477 8279
rect 5579 8273 5614 8279
rect 5986 8287 6027 8314
rect 5986 8279 6044 8287
rect 6106 8713 6594 8721
rect 6123 8665 6577 8713
rect 6123 8335 6185 8665
rect 6515 8335 6577 8665
rect 6123 8287 6577 8335
rect 6106 8279 6594 8287
rect 6656 8713 6714 8721
rect 6673 8686 6714 8713
rect 7086 8721 7121 8727
rect 7223 8721 7677 8727
rect 7779 8721 7814 8727
rect 7086 8713 7144 8721
rect 7086 8686 7127 8713
rect 6673 8287 6714 8314
rect 6656 8279 6714 8287
rect 5986 8273 6021 8279
rect 6123 8273 6577 8279
rect 6679 8273 6714 8279
rect 7086 8287 7127 8314
rect 7086 8279 7144 8287
rect 7206 8713 7694 8721
rect 7223 8665 7677 8713
rect 7223 8335 7285 8665
rect 7615 8335 7677 8665
rect 7223 8287 7677 8335
rect 7206 8279 7694 8287
rect 7756 8713 7814 8721
rect 7773 8686 7814 8713
rect 8186 8721 8221 8727
rect 8323 8721 8777 8727
rect 8879 8721 8914 8727
rect 8186 8713 8244 8721
rect 8186 8686 8227 8713
rect 7773 8287 7814 8314
rect 7756 8279 7814 8287
rect 7086 8273 7121 8279
rect 7223 8273 7677 8279
rect 7779 8273 7814 8279
rect 8186 8287 8227 8314
rect 8186 8279 8244 8287
rect 8306 8713 8794 8721
rect 8323 8665 8777 8713
rect 8323 8335 8385 8665
rect 8715 8335 8777 8665
rect 8323 8287 8777 8335
rect 8306 8279 8794 8287
rect 8856 8713 8914 8721
rect 8873 8686 8914 8713
rect 9286 8721 9321 8727
rect 9423 8721 9877 8727
rect 9979 8721 10014 8727
rect 9286 8713 9344 8721
rect 9286 8686 9327 8713
rect 8873 8287 8914 8314
rect 8856 8279 8914 8287
rect 8186 8273 8221 8279
rect 8323 8273 8777 8279
rect 8879 8273 8914 8279
rect 9286 8287 9327 8314
rect 9286 8279 9344 8287
rect 9406 8713 9894 8721
rect 9423 8665 9877 8713
rect 9423 8335 9485 8665
rect 9815 8335 9877 8665
rect 9423 8287 9877 8335
rect 9406 8279 9894 8287
rect 9956 8713 10014 8721
rect 9973 8686 10014 8713
rect 10386 8721 10421 8727
rect 10523 8721 10977 8727
rect 11079 8721 11114 8727
rect 10386 8713 10444 8721
rect 10386 8686 10427 8713
rect 9973 8287 10014 8314
rect 9956 8279 10014 8287
rect 9286 8273 9321 8279
rect 9423 8273 9877 8279
rect 9979 8273 10014 8279
rect 10386 8287 10427 8314
rect 10386 8279 10444 8287
rect 10506 8713 10994 8721
rect 10523 8665 10977 8713
rect 10523 8335 10585 8665
rect 10915 8335 10977 8665
rect 10523 8287 10977 8335
rect 10506 8279 10994 8287
rect 11056 8713 11114 8721
rect 11073 8686 11114 8713
rect 11486 8721 11521 8727
rect 11623 8721 12077 8727
rect 12179 8721 12214 8727
rect 11486 8713 11544 8721
rect 11486 8686 11527 8713
rect 11073 8287 11114 8314
rect 11056 8279 11114 8287
rect 10386 8273 10421 8279
rect 10523 8273 10977 8279
rect 11079 8273 11114 8279
rect 11486 8287 11527 8314
rect 11486 8279 11544 8287
rect 11606 8713 12094 8721
rect 11623 8665 12077 8713
rect 11623 8335 11685 8665
rect 12015 8335 12077 8665
rect 11623 8287 12077 8335
rect 11606 8279 12094 8287
rect 12156 8713 12214 8721
rect 12173 8686 12214 8713
rect 12586 8721 12621 8727
rect 12723 8721 13177 8727
rect 13279 8721 13314 8727
rect 12586 8713 12644 8721
rect 12586 8686 12627 8713
rect 12173 8287 12214 8314
rect 12156 8279 12214 8287
rect 11486 8273 11521 8279
rect 11623 8273 12077 8279
rect 12179 8273 12214 8279
rect 12586 8287 12627 8314
rect 12586 8279 12644 8287
rect 12706 8713 13194 8721
rect 12723 8665 13177 8713
rect 12723 8335 12785 8665
rect 13115 8335 13177 8665
rect 12723 8287 13177 8335
rect 12706 8279 13194 8287
rect 13256 8713 13314 8721
rect 13273 8686 13314 8713
rect 13273 8287 13314 8314
rect 13256 8279 13314 8287
rect 12586 8273 12621 8279
rect 12723 8273 13177 8279
rect 13279 8273 13314 8279
rect -1025 8250 -725 8267
rect -471 8256 -463 8273
rect -37 8256 -29 8273
rect 79 8256 87 8273
rect 513 8256 521 8273
rect 629 8256 637 8273
rect 1063 8256 1071 8273
rect 1179 8256 1187 8273
rect 1613 8256 1621 8273
rect 1729 8256 1737 8273
rect 2163 8256 2171 8273
rect 2279 8256 2287 8273
rect 2713 8256 2721 8273
rect 2829 8256 2837 8273
rect 3263 8256 3271 8273
rect 3379 8256 3387 8273
rect 3813 8256 3821 8273
rect 3929 8256 3937 8273
rect 4363 8256 4371 8273
rect 4479 8256 4487 8273
rect 4913 8256 4921 8273
rect 5029 8256 5037 8273
rect 5463 8256 5471 8273
rect 5579 8256 5587 8273
rect 6013 8256 6021 8273
rect 6129 8256 6137 8273
rect 6563 8256 6571 8273
rect 6679 8256 6687 8273
rect 7113 8256 7121 8273
rect 7229 8256 7237 8273
rect 7663 8256 7671 8273
rect 7779 8256 7787 8273
rect 8213 8256 8221 8273
rect 8329 8256 8337 8273
rect 8763 8256 8771 8273
rect 8879 8256 8887 8273
rect 9313 8256 9321 8273
rect 9429 8256 9437 8273
rect 9863 8256 9871 8273
rect 9979 8256 9987 8273
rect 10413 8256 10421 8273
rect 10529 8256 10537 8273
rect 10963 8256 10971 8273
rect 11079 8256 11087 8273
rect 11513 8256 11521 8273
rect 11629 8256 11637 8273
rect 12063 8256 12071 8273
rect 12179 8256 12187 8273
rect 12613 8256 12621 8273
rect 12729 8256 12737 8273
rect 13163 8256 13171 8273
rect 13279 8256 13287 8273
rect 13713 8256 13721 8273
rect 13975 8269 13987 8800
rect 14263 8269 14275 8800
rect 13975 8250 14275 8269
rect -1025 7717 -1013 8250
rect -737 7717 -725 8250
rect -550 8242 -500 8250
rect -550 8208 -542 8242
rect -508 8208 -500 8242
rect -550 8200 -500 8208
rect 0 8242 50 8250
rect 0 8208 8 8242
rect 42 8208 50 8242
rect 0 8200 50 8208
rect 550 8242 600 8250
rect 550 8208 558 8242
rect 592 8208 600 8242
rect 550 8200 600 8208
rect 1100 8242 1150 8250
rect 1100 8208 1108 8242
rect 1142 8208 1150 8242
rect 1100 8200 1150 8208
rect 1650 8242 1700 8250
rect 1650 8208 1658 8242
rect 1692 8208 1700 8242
rect 1650 8200 1700 8208
rect 2200 8242 2250 8250
rect 2200 8208 2208 8242
rect 2242 8208 2250 8242
rect 2200 8200 2250 8208
rect 2750 8242 2800 8250
rect 2750 8208 2758 8242
rect 2792 8208 2800 8242
rect 2750 8200 2800 8208
rect 3300 8242 3350 8250
rect 3300 8208 3308 8242
rect 3342 8208 3350 8242
rect 3300 8200 3350 8208
rect 3850 8242 3900 8250
rect 3850 8208 3858 8242
rect 3892 8208 3900 8242
rect 3850 8200 3900 8208
rect 4400 8242 4450 8250
rect 4400 8208 4408 8242
rect 4442 8208 4450 8242
rect 4400 8200 4450 8208
rect 4950 8242 5000 8250
rect 4950 8208 4958 8242
rect 4992 8208 5000 8242
rect 4950 8200 5000 8208
rect 5500 8242 5550 8250
rect 5500 8208 5508 8242
rect 5542 8208 5550 8242
rect 5500 8200 5550 8208
rect 6050 8242 6100 8250
rect 6050 8208 6058 8242
rect 6092 8208 6100 8242
rect 6050 8200 6100 8208
rect 6600 8242 6650 8250
rect 6600 8208 6608 8242
rect 6642 8208 6650 8242
rect 6600 8200 6650 8208
rect 7150 8242 7200 8250
rect 7150 8208 7158 8242
rect 7192 8208 7200 8242
rect 7150 8200 7200 8208
rect 7700 8242 7750 8250
rect 7700 8208 7708 8242
rect 7742 8208 7750 8242
rect 7700 8200 7750 8208
rect 8250 8242 8300 8250
rect 8250 8208 8258 8242
rect 8292 8208 8300 8242
rect 8250 8200 8300 8208
rect 8800 8242 8850 8250
rect 8800 8208 8808 8242
rect 8842 8208 8850 8242
rect 8800 8200 8850 8208
rect 9350 8242 9400 8250
rect 9350 8208 9358 8242
rect 9392 8208 9400 8242
rect 9350 8200 9400 8208
rect 9900 8242 9950 8250
rect 9900 8208 9908 8242
rect 9942 8208 9950 8242
rect 9900 8200 9950 8208
rect 10450 8242 10500 8250
rect 10450 8208 10458 8242
rect 10492 8208 10500 8242
rect 10450 8200 10500 8208
rect 11000 8242 11050 8250
rect 11000 8208 11008 8242
rect 11042 8208 11050 8242
rect 11000 8200 11050 8208
rect 11550 8242 11600 8250
rect 11550 8208 11558 8242
rect 11592 8208 11600 8242
rect 11550 8200 11600 8208
rect 12100 8242 12150 8250
rect 12100 8208 12108 8242
rect 12142 8208 12150 8242
rect 12100 8200 12150 8208
rect 12650 8242 12700 8250
rect 12650 8208 12658 8242
rect 12692 8208 12700 8242
rect 12650 8200 12700 8208
rect 13200 8242 13250 8250
rect 13200 8208 13208 8242
rect 13242 8208 13250 8242
rect 13200 8200 13250 8208
rect 13750 8242 13800 8250
rect 13750 8208 13758 8242
rect 13792 8208 13800 8242
rect 13750 8200 13800 8208
rect -471 8177 -463 8194
rect -37 8177 -29 8194
rect 79 8177 87 8194
rect 513 8177 521 8194
rect 629 8177 637 8194
rect 1063 8177 1071 8194
rect 1179 8177 1187 8194
rect 1613 8177 1621 8194
rect 1729 8177 1737 8194
rect 2163 8177 2171 8194
rect 2279 8177 2287 8194
rect 2713 8177 2721 8194
rect 2829 8177 2837 8194
rect 3263 8177 3271 8194
rect 3379 8177 3387 8194
rect 3813 8177 3821 8194
rect 3929 8177 3937 8194
rect 4363 8177 4371 8194
rect 4479 8177 4487 8194
rect 4913 8177 4921 8194
rect 5029 8177 5037 8194
rect 5463 8177 5471 8194
rect 5579 8177 5587 8194
rect 6013 8177 6021 8194
rect 6129 8177 6137 8194
rect 6563 8177 6571 8194
rect 6679 8177 6687 8194
rect 7113 8177 7121 8194
rect 7229 8177 7237 8194
rect 7663 8177 7671 8194
rect 7779 8177 7787 8194
rect 8213 8177 8221 8194
rect 8329 8177 8337 8194
rect 8763 8177 8771 8194
rect 8879 8177 8887 8194
rect 9313 8177 9321 8194
rect 9429 8177 9437 8194
rect 9863 8177 9871 8194
rect 9979 8177 9987 8194
rect 10413 8177 10421 8194
rect 10529 8177 10537 8194
rect 10963 8177 10971 8194
rect 11079 8177 11087 8194
rect 11513 8177 11521 8194
rect 11629 8177 11637 8194
rect 12063 8177 12071 8194
rect 12179 8177 12187 8194
rect 12613 8177 12621 8194
rect 12729 8177 12737 8194
rect 13163 8177 13171 8194
rect 13279 8177 13287 8194
rect 13713 8177 13721 8194
rect -64 8171 -29 8177
rect 73 8171 527 8177
rect 629 8171 664 8177
rect -64 8163 -6 8171
rect -64 8136 -23 8163
rect -64 7737 -23 7764
rect -64 7729 -6 7737
rect 56 8163 544 8171
rect 73 8115 527 8163
rect 73 7785 135 8115
rect 465 7785 527 8115
rect 73 7737 527 7785
rect 56 7729 544 7737
rect 606 8163 664 8171
rect 623 8136 664 8163
rect 1036 8171 1071 8177
rect 1173 8171 1627 8177
rect 1729 8171 1764 8177
rect 1036 8163 1094 8171
rect 1036 8136 1077 8163
rect 623 7737 664 7764
rect 606 7729 664 7737
rect -64 7723 -29 7729
rect 73 7723 527 7729
rect 629 7723 664 7729
rect 1036 7737 1077 7764
rect 1036 7729 1094 7737
rect 1156 8163 1644 8171
rect 1173 8115 1627 8163
rect 1173 7785 1235 8115
rect 1565 7785 1627 8115
rect 1173 7737 1627 7785
rect 1156 7729 1644 7737
rect 1706 8163 1764 8171
rect 1723 8136 1764 8163
rect 2136 8171 2171 8177
rect 2273 8171 2727 8177
rect 2829 8171 2864 8177
rect 2136 8163 2194 8171
rect 2136 8136 2177 8163
rect 1723 7737 1764 7764
rect 1706 7729 1764 7737
rect 1036 7723 1071 7729
rect 1173 7723 1627 7729
rect 1729 7723 1764 7729
rect 2136 7737 2177 7764
rect 2136 7729 2194 7737
rect 2256 8163 2744 8171
rect 2273 8115 2727 8163
rect 2273 7785 2335 8115
rect 2665 7785 2727 8115
rect 2273 7737 2727 7785
rect 2256 7729 2744 7737
rect 2806 8163 2864 8171
rect 2823 8136 2864 8163
rect 3236 8171 3271 8177
rect 3373 8171 3827 8177
rect 3929 8171 3964 8177
rect 3236 8163 3294 8171
rect 3236 8136 3277 8163
rect 2823 7737 2864 7764
rect 2806 7729 2864 7737
rect 2136 7723 2171 7729
rect 2273 7723 2727 7729
rect 2829 7723 2864 7729
rect 3236 7737 3277 7764
rect 3236 7729 3294 7737
rect 3356 8163 3844 8171
rect 3373 8115 3827 8163
rect 3373 7785 3435 8115
rect 3765 7785 3827 8115
rect 3373 7737 3827 7785
rect 3356 7729 3844 7737
rect 3906 8163 3964 8171
rect 3923 8136 3964 8163
rect 4336 8171 4371 8177
rect 4473 8171 4927 8177
rect 5029 8171 5064 8177
rect 4336 8163 4394 8171
rect 4336 8136 4377 8163
rect 3923 7737 3964 7764
rect 3906 7729 3964 7737
rect 3236 7723 3271 7729
rect 3373 7723 3827 7729
rect 3929 7723 3964 7729
rect 4336 7737 4377 7764
rect 4336 7729 4394 7737
rect 4456 8163 4944 8171
rect 4473 8115 4927 8163
rect 4473 7785 4535 8115
rect 4865 7785 4927 8115
rect 4473 7737 4927 7785
rect 4456 7729 4944 7737
rect 5006 8163 5064 8171
rect 5023 8136 5064 8163
rect 5436 8171 5471 8177
rect 5573 8171 6027 8177
rect 6129 8171 6164 8177
rect 5436 8163 5494 8171
rect 5436 8136 5477 8163
rect 5023 7737 5064 7764
rect 5006 7729 5064 7737
rect 4336 7723 4371 7729
rect 4473 7723 4927 7729
rect 5029 7723 5064 7729
rect 5436 7737 5477 7764
rect 5436 7729 5494 7737
rect 5556 8163 6044 8171
rect 5573 8115 6027 8163
rect 5573 7785 5635 8115
rect 5965 7785 6027 8115
rect 5573 7737 6027 7785
rect 5556 7729 6044 7737
rect 6106 8163 6164 8171
rect 6123 8136 6164 8163
rect 6536 8171 6571 8177
rect 6673 8171 7127 8177
rect 7229 8171 7264 8177
rect 6536 8163 6594 8171
rect 6536 8136 6577 8163
rect 6123 7737 6164 7764
rect 6106 7729 6164 7737
rect 5436 7723 5471 7729
rect 5573 7723 6027 7729
rect 6129 7723 6164 7729
rect 6536 7737 6577 7764
rect 6536 7729 6594 7737
rect 6656 8163 7144 8171
rect 6673 8115 7127 8163
rect 6673 7785 6735 8115
rect 7065 7785 7127 8115
rect 6673 7737 7127 7785
rect 6656 7729 7144 7737
rect 7206 8163 7264 8171
rect 7223 8136 7264 8163
rect 7636 8171 7671 8177
rect 7773 8171 8227 8177
rect 8329 8171 8364 8177
rect 7636 8163 7694 8171
rect 7636 8136 7677 8163
rect 7223 7737 7264 7764
rect 7206 7729 7264 7737
rect 6536 7723 6571 7729
rect 6673 7723 7127 7729
rect 7229 7723 7264 7729
rect 7636 7737 7677 7764
rect 7636 7729 7694 7737
rect 7756 8163 8244 8171
rect 7773 8115 8227 8163
rect 7773 7785 7835 8115
rect 8165 7785 8227 8115
rect 7773 7737 8227 7785
rect 7756 7729 8244 7737
rect 8306 8163 8364 8171
rect 8323 8136 8364 8163
rect 8736 8171 8771 8177
rect 8873 8171 9327 8177
rect 9429 8171 9464 8177
rect 8736 8163 8794 8171
rect 8736 8136 8777 8163
rect 8323 7737 8364 7764
rect 8306 7729 8364 7737
rect 7636 7723 7671 7729
rect 7773 7723 8227 7729
rect 8329 7723 8364 7729
rect 8736 7737 8777 7764
rect 8736 7729 8794 7737
rect 8856 8163 9344 8171
rect 8873 8115 9327 8163
rect 8873 7785 8935 8115
rect 9265 7785 9327 8115
rect 8873 7737 9327 7785
rect 8856 7729 9344 7737
rect 9406 8163 9464 8171
rect 9423 8136 9464 8163
rect 9836 8171 9871 8177
rect 9973 8171 10427 8177
rect 10529 8171 10564 8177
rect 9836 8163 9894 8171
rect 9836 8136 9877 8163
rect 9423 7737 9464 7764
rect 9406 7729 9464 7737
rect 8736 7723 8771 7729
rect 8873 7723 9327 7729
rect 9429 7723 9464 7729
rect 9836 7737 9877 7764
rect 9836 7729 9894 7737
rect 9956 8163 10444 8171
rect 9973 8115 10427 8163
rect 9973 7785 10035 8115
rect 10365 7785 10427 8115
rect 9973 7737 10427 7785
rect 9956 7729 10444 7737
rect 10506 8163 10564 8171
rect 10523 8136 10564 8163
rect 10936 8171 10971 8177
rect 11073 8171 11527 8177
rect 11629 8171 11664 8177
rect 10936 8163 10994 8171
rect 10936 8136 10977 8163
rect 10523 7737 10564 7764
rect 10506 7729 10564 7737
rect 9836 7723 9871 7729
rect 9973 7723 10427 7729
rect 10529 7723 10564 7729
rect 10936 7737 10977 7764
rect 10936 7729 10994 7737
rect 11056 8163 11544 8171
rect 11073 8115 11527 8163
rect 11073 7785 11135 8115
rect 11465 7785 11527 8115
rect 11073 7737 11527 7785
rect 11056 7729 11544 7737
rect 11606 8163 11664 8171
rect 11623 8136 11664 8163
rect 12036 8171 12071 8177
rect 12173 8171 12627 8177
rect 12729 8171 12764 8177
rect 12036 8163 12094 8171
rect 12036 8136 12077 8163
rect 11623 7737 11664 7764
rect 11606 7729 11664 7737
rect 10936 7723 10971 7729
rect 11073 7723 11527 7729
rect 11629 7723 11664 7729
rect 12036 7737 12077 7764
rect 12036 7729 12094 7737
rect 12156 8163 12644 8171
rect 12173 8115 12627 8163
rect 12173 7785 12235 8115
rect 12565 7785 12627 8115
rect 12173 7737 12627 7785
rect 12156 7729 12644 7737
rect 12706 8163 12764 8171
rect 12723 8136 12764 8163
rect 13136 8171 13171 8177
rect 13273 8171 13727 8177
rect 13136 8163 13194 8171
rect 13136 8136 13177 8163
rect 12723 7737 12764 7764
rect 12706 7729 12764 7737
rect 12036 7723 12071 7729
rect 12173 7723 12627 7729
rect 12729 7723 12764 7729
rect 13136 7737 13177 7764
rect 13136 7729 13194 7737
rect 13256 8163 13727 8171
rect 13273 8115 13727 8163
rect 13273 7785 13335 8115
rect 13665 7785 13727 8115
rect 13273 7737 13727 7785
rect 13256 7729 13727 7737
rect 13136 7723 13171 7729
rect 13273 7723 13727 7729
rect -1025 7700 -725 7717
rect -471 7706 -463 7723
rect -37 7706 -29 7723
rect 79 7706 87 7723
rect 513 7706 521 7723
rect 629 7706 637 7723
rect 1063 7706 1071 7723
rect 1179 7706 1187 7723
rect 1613 7706 1621 7723
rect 1729 7706 1737 7723
rect 2163 7706 2171 7723
rect 2279 7706 2287 7723
rect 2713 7706 2721 7723
rect 2829 7706 2837 7723
rect 3263 7706 3271 7723
rect 3379 7706 3387 7723
rect 3813 7706 3821 7723
rect 3929 7706 3937 7723
rect 4363 7706 4371 7723
rect 4479 7706 4487 7723
rect 4913 7706 4921 7723
rect 5029 7706 5037 7723
rect 5463 7706 5471 7723
rect 5579 7706 5587 7723
rect 6013 7706 6021 7723
rect 6129 7706 6137 7723
rect 6563 7706 6571 7723
rect 6679 7706 6687 7723
rect 7113 7706 7121 7723
rect 7229 7706 7237 7723
rect 7663 7706 7671 7723
rect 7779 7706 7787 7723
rect 8213 7706 8221 7723
rect 8329 7706 8337 7723
rect 8763 7706 8771 7723
rect 8879 7706 8887 7723
rect 9313 7706 9321 7723
rect 9429 7706 9437 7723
rect 9863 7706 9871 7723
rect 9979 7706 9987 7723
rect 10413 7706 10421 7723
rect 10529 7706 10537 7723
rect 10963 7706 10971 7723
rect 11079 7706 11087 7723
rect 11513 7706 11521 7723
rect 11629 7706 11637 7723
rect 12063 7706 12071 7723
rect 12179 7706 12187 7723
rect 12613 7706 12621 7723
rect 12729 7706 12737 7723
rect 13163 7706 13171 7723
rect 13279 7706 13287 7723
rect 13713 7706 13721 7723
rect 13975 7717 13987 8250
rect 14263 7717 14275 8250
rect 13975 7700 14275 7717
rect -1025 7167 -1013 7700
rect -737 7167 -725 7700
rect -550 7692 -500 7700
rect -550 7658 -542 7692
rect -508 7658 -500 7692
rect -550 7650 -500 7658
rect 0 7692 50 7700
rect 0 7658 8 7692
rect 42 7658 50 7692
rect 0 7650 50 7658
rect 550 7692 600 7700
rect 550 7658 558 7692
rect 592 7658 600 7692
rect 550 7650 600 7658
rect 1100 7692 1150 7700
rect 1100 7658 1108 7692
rect 1142 7658 1150 7692
rect 1100 7650 1150 7658
rect 1650 7692 1700 7700
rect 1650 7658 1658 7692
rect 1692 7658 1700 7692
rect 1650 7650 1700 7658
rect 2200 7692 2250 7700
rect 2200 7658 2208 7692
rect 2242 7658 2250 7692
rect 2200 7650 2250 7658
rect 2750 7692 2800 7700
rect 2750 7658 2758 7692
rect 2792 7658 2800 7692
rect 2750 7650 2800 7658
rect 3300 7692 3350 7700
rect 3300 7658 3308 7692
rect 3342 7658 3350 7692
rect 3300 7650 3350 7658
rect 3850 7692 3900 7700
rect 3850 7658 3858 7692
rect 3892 7658 3900 7692
rect 3850 7650 3900 7658
rect 4400 7692 4450 7700
rect 4400 7658 4408 7692
rect 4442 7658 4450 7692
rect 4400 7650 4450 7658
rect 4950 7692 5000 7700
rect 4950 7658 4958 7692
rect 4992 7658 5000 7692
rect 4950 7650 5000 7658
rect 5500 7692 5550 7700
rect 5500 7658 5508 7692
rect 5542 7658 5550 7692
rect 5500 7650 5550 7658
rect 6050 7692 6100 7700
rect 6050 7658 6058 7692
rect 6092 7658 6100 7692
rect 6050 7650 6100 7658
rect 6600 7692 6650 7700
rect 6600 7658 6608 7692
rect 6642 7658 6650 7692
rect 6600 7650 6650 7658
rect 7150 7692 7200 7700
rect 7150 7658 7158 7692
rect 7192 7658 7200 7692
rect 7150 7650 7200 7658
rect 7700 7692 7750 7700
rect 7700 7658 7708 7692
rect 7742 7658 7750 7692
rect 7700 7650 7750 7658
rect 8250 7692 8300 7700
rect 8250 7658 8258 7692
rect 8292 7658 8300 7692
rect 8250 7650 8300 7658
rect 8800 7692 8850 7700
rect 8800 7658 8808 7692
rect 8842 7658 8850 7692
rect 8800 7650 8850 7658
rect 9350 7692 9400 7700
rect 9350 7658 9358 7692
rect 9392 7658 9400 7692
rect 9350 7650 9400 7658
rect 9900 7692 9950 7700
rect 9900 7658 9908 7692
rect 9942 7658 9950 7692
rect 9900 7650 9950 7658
rect 10450 7692 10500 7700
rect 10450 7658 10458 7692
rect 10492 7658 10500 7692
rect 10450 7650 10500 7658
rect 11000 7692 11050 7700
rect 11000 7658 11008 7692
rect 11042 7658 11050 7692
rect 11000 7650 11050 7658
rect 11550 7692 11600 7700
rect 11550 7658 11558 7692
rect 11592 7658 11600 7692
rect 11550 7650 11600 7658
rect 12100 7692 12150 7700
rect 12100 7658 12108 7692
rect 12142 7658 12150 7692
rect 12100 7650 12150 7658
rect 12650 7692 12700 7700
rect 12650 7658 12658 7692
rect 12692 7658 12700 7692
rect 12650 7650 12700 7658
rect 13200 7692 13250 7700
rect 13200 7658 13208 7692
rect 13242 7658 13250 7692
rect 13200 7650 13250 7658
rect 13750 7692 13800 7700
rect 13750 7658 13758 7692
rect 13792 7658 13800 7692
rect 13750 7650 13800 7658
rect -471 7627 -463 7644
rect -37 7627 -29 7644
rect 79 7627 87 7644
rect 513 7627 521 7644
rect 629 7627 637 7644
rect 1063 7627 1071 7644
rect 1179 7627 1187 7644
rect 1613 7627 1621 7644
rect 1729 7627 1737 7644
rect 2163 7627 2171 7644
rect 2279 7627 2287 7644
rect 2713 7627 2721 7644
rect 2829 7627 2837 7644
rect 3263 7627 3271 7644
rect 3379 7627 3387 7644
rect 3813 7627 3821 7644
rect 3929 7627 3937 7644
rect 4363 7627 4371 7644
rect 4479 7627 4487 7644
rect 4913 7627 4921 7644
rect 5029 7627 5037 7644
rect 5463 7627 5471 7644
rect 5579 7627 5587 7644
rect 6013 7627 6021 7644
rect 6129 7627 6137 7644
rect 6563 7627 6571 7644
rect 6679 7627 6687 7644
rect 7113 7627 7121 7644
rect 7229 7627 7237 7644
rect 7663 7627 7671 7644
rect 7779 7627 7787 7644
rect 8213 7627 8221 7644
rect 8329 7627 8337 7644
rect 8763 7627 8771 7644
rect 8879 7627 8887 7644
rect 9313 7627 9321 7644
rect 9429 7627 9437 7644
rect 9863 7627 9871 7644
rect 9979 7627 9987 7644
rect 10413 7627 10421 7644
rect 10529 7627 10537 7644
rect 10963 7627 10971 7644
rect 11079 7627 11087 7644
rect 11513 7627 11521 7644
rect 11629 7627 11637 7644
rect 12063 7627 12071 7644
rect 12179 7627 12187 7644
rect 12613 7627 12621 7644
rect 12729 7627 12737 7644
rect 13163 7627 13171 7644
rect 13279 7627 13287 7644
rect 13713 7627 13721 7644
rect -477 7621 -23 7627
rect 79 7621 114 7627
rect -477 7613 -6 7621
rect -477 7565 -23 7613
rect -477 7235 -415 7565
rect -85 7235 -23 7565
rect -477 7187 -23 7235
rect -477 7179 -6 7187
rect 56 7613 114 7621
rect 73 7586 114 7613
rect 486 7621 521 7627
rect 623 7621 1077 7627
rect 1179 7621 1214 7627
rect 486 7613 544 7621
rect 486 7586 527 7613
rect 73 7187 114 7214
rect 56 7179 114 7187
rect -477 7173 -23 7179
rect 79 7173 114 7179
rect 486 7187 527 7214
rect 486 7179 544 7187
rect 606 7613 1094 7621
rect 623 7565 1077 7613
rect 623 7235 685 7565
rect 1015 7235 1077 7565
rect 623 7187 1077 7235
rect 606 7179 1094 7187
rect 1156 7613 1214 7621
rect 1173 7586 1214 7613
rect 1586 7621 1621 7627
rect 1723 7621 2177 7627
rect 2279 7621 2314 7627
rect 1586 7613 1644 7621
rect 1586 7586 1627 7613
rect 1173 7187 1214 7214
rect 1156 7179 1214 7187
rect 486 7173 521 7179
rect 623 7173 1077 7179
rect 1179 7173 1214 7179
rect 1586 7187 1627 7214
rect 1586 7179 1644 7187
rect 1706 7613 2194 7621
rect 1723 7565 2177 7613
rect 1723 7235 1785 7565
rect 2115 7235 2177 7565
rect 1723 7187 2177 7235
rect 1706 7179 2194 7187
rect 2256 7613 2314 7621
rect 2273 7586 2314 7613
rect 2686 7621 2721 7627
rect 2823 7621 3277 7627
rect 3379 7621 3414 7627
rect 2686 7613 2744 7621
rect 2686 7586 2727 7613
rect 2273 7187 2314 7214
rect 2256 7179 2314 7187
rect 1586 7173 1621 7179
rect 1723 7173 2177 7179
rect 2279 7173 2314 7179
rect 2686 7187 2727 7214
rect 2686 7179 2744 7187
rect 2806 7613 3294 7621
rect 2823 7565 3277 7613
rect 2823 7235 2885 7565
rect 3215 7235 3277 7565
rect 2823 7187 3277 7235
rect 2806 7179 3294 7187
rect 3356 7613 3414 7621
rect 3373 7586 3414 7613
rect 3786 7621 3821 7627
rect 3923 7621 4377 7627
rect 4479 7621 4514 7627
rect 3786 7613 3844 7621
rect 3786 7586 3827 7613
rect 3373 7187 3414 7214
rect 3356 7179 3414 7187
rect 2686 7173 2721 7179
rect 2823 7173 3277 7179
rect 3379 7173 3414 7179
rect 3786 7187 3827 7214
rect 3786 7179 3844 7187
rect 3906 7613 4394 7621
rect 3923 7565 4377 7613
rect 3923 7235 3985 7565
rect 4315 7235 4377 7565
rect 3923 7187 4377 7235
rect 3906 7179 4394 7187
rect 4456 7613 4514 7621
rect 4473 7586 4514 7613
rect 4886 7621 4921 7627
rect 5023 7621 5477 7627
rect 5579 7621 5614 7627
rect 4886 7613 4944 7621
rect 4886 7586 4927 7613
rect 4473 7187 4514 7214
rect 4456 7179 4514 7187
rect 3786 7173 3821 7179
rect 3923 7173 4377 7179
rect 4479 7173 4514 7179
rect 4886 7187 4927 7214
rect 4886 7179 4944 7187
rect 5006 7613 5494 7621
rect 5023 7565 5477 7613
rect 5023 7235 5085 7565
rect 5415 7235 5477 7565
rect 5023 7187 5477 7235
rect 5006 7179 5494 7187
rect 5556 7613 5614 7621
rect 5573 7586 5614 7613
rect 5986 7621 6021 7627
rect 6123 7621 6577 7627
rect 6679 7621 6714 7627
rect 5986 7613 6044 7621
rect 5986 7586 6027 7613
rect 5573 7187 5614 7214
rect 5556 7179 5614 7187
rect 4886 7173 4921 7179
rect 5023 7173 5477 7179
rect 5579 7173 5614 7179
rect 5986 7187 6027 7214
rect 5986 7179 6044 7187
rect 6106 7613 6594 7621
rect 6123 7565 6577 7613
rect 6123 7235 6185 7565
rect 6515 7235 6577 7565
rect 6123 7187 6577 7235
rect 6106 7179 6594 7187
rect 6656 7613 6714 7621
rect 6673 7586 6714 7613
rect 7086 7621 7121 7627
rect 7223 7621 7677 7627
rect 7779 7621 7814 7627
rect 7086 7613 7144 7621
rect 7086 7586 7127 7613
rect 6673 7187 6714 7214
rect 6656 7179 6714 7187
rect 5986 7173 6021 7179
rect 6123 7173 6577 7179
rect 6679 7173 6714 7179
rect 7086 7187 7127 7214
rect 7086 7179 7144 7187
rect 7206 7613 7694 7621
rect 7223 7565 7677 7613
rect 7223 7235 7285 7565
rect 7615 7235 7677 7565
rect 7223 7187 7677 7235
rect 7206 7179 7694 7187
rect 7756 7613 7814 7621
rect 7773 7586 7814 7613
rect 8186 7621 8221 7627
rect 8323 7621 8777 7627
rect 8879 7621 8914 7627
rect 8186 7613 8244 7621
rect 8186 7586 8227 7613
rect 7773 7187 7814 7214
rect 7756 7179 7814 7187
rect 7086 7173 7121 7179
rect 7223 7173 7677 7179
rect 7779 7173 7814 7179
rect 8186 7187 8227 7214
rect 8186 7179 8244 7187
rect 8306 7613 8794 7621
rect 8323 7565 8777 7613
rect 8323 7235 8385 7565
rect 8715 7235 8777 7565
rect 8323 7187 8777 7235
rect 8306 7179 8794 7187
rect 8856 7613 8914 7621
rect 8873 7586 8914 7613
rect 9286 7621 9321 7627
rect 9423 7621 9877 7627
rect 9979 7621 10014 7627
rect 9286 7613 9344 7621
rect 9286 7586 9327 7613
rect 8873 7187 8914 7214
rect 8856 7179 8914 7187
rect 8186 7173 8221 7179
rect 8323 7173 8777 7179
rect 8879 7173 8914 7179
rect 9286 7187 9327 7214
rect 9286 7179 9344 7187
rect 9406 7613 9894 7621
rect 9423 7565 9877 7613
rect 9423 7235 9485 7565
rect 9815 7235 9877 7565
rect 9423 7187 9877 7235
rect 9406 7179 9894 7187
rect 9956 7613 10014 7621
rect 9973 7586 10014 7613
rect 10386 7621 10421 7627
rect 10523 7621 10977 7627
rect 11079 7621 11114 7627
rect 10386 7613 10444 7621
rect 10386 7586 10427 7613
rect 9973 7187 10014 7214
rect 9956 7179 10014 7187
rect 9286 7173 9321 7179
rect 9423 7173 9877 7179
rect 9979 7173 10014 7179
rect 10386 7187 10427 7214
rect 10386 7179 10444 7187
rect 10506 7613 10994 7621
rect 10523 7565 10977 7613
rect 10523 7235 10585 7565
rect 10915 7235 10977 7565
rect 10523 7187 10977 7235
rect 10506 7179 10994 7187
rect 11056 7613 11114 7621
rect 11073 7586 11114 7613
rect 11486 7621 11521 7627
rect 11623 7621 12077 7627
rect 12179 7621 12214 7627
rect 11486 7613 11544 7621
rect 11486 7586 11527 7613
rect 11073 7187 11114 7214
rect 11056 7179 11114 7187
rect 10386 7173 10421 7179
rect 10523 7173 10977 7179
rect 11079 7173 11114 7179
rect 11486 7187 11527 7214
rect 11486 7179 11544 7187
rect 11606 7613 12094 7621
rect 11623 7565 12077 7613
rect 11623 7235 11685 7565
rect 12015 7235 12077 7565
rect 11623 7187 12077 7235
rect 11606 7179 12094 7187
rect 12156 7613 12214 7621
rect 12173 7586 12214 7613
rect 12586 7621 12621 7627
rect 12723 7621 13177 7627
rect 13279 7621 13314 7627
rect 12586 7613 12644 7621
rect 12586 7586 12627 7613
rect 12173 7187 12214 7214
rect 12156 7179 12214 7187
rect 11486 7173 11521 7179
rect 11623 7173 12077 7179
rect 12179 7173 12214 7179
rect 12586 7187 12627 7214
rect 12586 7179 12644 7187
rect 12706 7613 13194 7621
rect 12723 7565 13177 7613
rect 12723 7235 12785 7565
rect 13115 7235 13177 7565
rect 12723 7187 13177 7235
rect 12706 7179 13194 7187
rect 13256 7613 13314 7621
rect 13273 7586 13314 7613
rect 13273 7187 13314 7214
rect 13256 7179 13314 7187
rect 12586 7173 12621 7179
rect 12723 7173 13177 7179
rect 13279 7173 13314 7179
rect -1025 7150 -725 7167
rect -471 7156 -463 7173
rect -37 7156 -29 7173
rect 79 7156 87 7173
rect 513 7156 521 7173
rect 629 7156 637 7173
rect 1063 7156 1071 7173
rect 1179 7156 1187 7173
rect 1613 7156 1621 7173
rect 1729 7156 1737 7173
rect 2163 7156 2171 7173
rect 2279 7156 2287 7173
rect 2713 7156 2721 7173
rect 2829 7156 2837 7173
rect 3263 7156 3271 7173
rect 3379 7156 3387 7173
rect 3813 7156 3821 7173
rect 3929 7156 3937 7173
rect 4363 7156 4371 7173
rect 4479 7156 4487 7173
rect 4913 7156 4921 7173
rect 5029 7156 5037 7173
rect 5463 7156 5471 7173
rect 5579 7156 5587 7173
rect 6013 7156 6021 7173
rect 6129 7156 6137 7173
rect 6563 7156 6571 7173
rect 6679 7156 6687 7173
rect 7113 7156 7121 7173
rect 7229 7156 7237 7173
rect 7663 7156 7671 7173
rect 7779 7156 7787 7173
rect 8213 7156 8221 7173
rect 8329 7156 8337 7173
rect 8763 7156 8771 7173
rect 8879 7156 8887 7173
rect 9313 7156 9321 7173
rect 9429 7156 9437 7173
rect 9863 7156 9871 7173
rect 9979 7156 9987 7173
rect 10413 7156 10421 7173
rect 10529 7156 10537 7173
rect 10963 7156 10971 7173
rect 11079 7156 11087 7173
rect 11513 7156 11521 7173
rect 11629 7156 11637 7173
rect 12063 7156 12071 7173
rect 12179 7156 12187 7173
rect 12613 7156 12621 7173
rect 12729 7156 12737 7173
rect 13163 7156 13171 7173
rect 13279 7156 13287 7173
rect 13713 7156 13721 7173
rect 13975 7169 13987 7700
rect 14263 7169 14275 7700
rect 13975 7150 14275 7169
rect -1025 6617 -1013 7150
rect -737 6617 -725 7150
rect -550 7142 -500 7150
rect -550 7108 -542 7142
rect -508 7108 -500 7142
rect -550 7100 -500 7108
rect 0 7142 50 7150
rect 0 7108 8 7142
rect 42 7108 50 7142
rect 0 7100 50 7108
rect 550 7142 600 7150
rect 550 7108 558 7142
rect 592 7108 600 7142
rect 550 7100 600 7108
rect 1100 7142 1150 7150
rect 1100 7108 1108 7142
rect 1142 7108 1150 7142
rect 1100 7100 1150 7108
rect 1650 7142 1700 7150
rect 1650 7108 1658 7142
rect 1692 7108 1700 7142
rect 1650 7100 1700 7108
rect 2200 7142 2250 7150
rect 2200 7108 2208 7142
rect 2242 7108 2250 7142
rect 2200 7100 2250 7108
rect 2750 7142 2800 7150
rect 2750 7108 2758 7142
rect 2792 7108 2800 7142
rect 2750 7100 2800 7108
rect 3300 7142 3350 7150
rect 3300 7108 3308 7142
rect 3342 7108 3350 7142
rect 3300 7100 3350 7108
rect 3850 7142 3900 7150
rect 3850 7108 3858 7142
rect 3892 7108 3900 7142
rect 3850 7100 3900 7108
rect 4400 7142 4450 7150
rect 4400 7108 4408 7142
rect 4442 7108 4450 7142
rect 4400 7100 4450 7108
rect 4950 7142 5000 7150
rect 4950 7108 4958 7142
rect 4992 7108 5000 7142
rect 4950 7100 5000 7108
rect 5500 7142 5550 7150
rect 5500 7108 5508 7142
rect 5542 7108 5550 7142
rect 5500 7100 5550 7108
rect 6050 7142 6100 7150
rect 6050 7108 6058 7142
rect 6092 7108 6100 7142
rect 6050 7100 6100 7108
rect 6600 7142 6650 7150
rect 6600 7108 6608 7142
rect 6642 7108 6650 7142
rect 6600 7100 6650 7108
rect 7150 7142 7200 7150
rect 7150 7108 7158 7142
rect 7192 7108 7200 7142
rect 7150 7100 7200 7108
rect 7700 7142 7750 7150
rect 7700 7108 7708 7142
rect 7742 7108 7750 7142
rect 7700 7100 7750 7108
rect 8250 7142 8300 7150
rect 8250 7108 8258 7142
rect 8292 7108 8300 7142
rect 8250 7100 8300 7108
rect 8800 7142 8850 7150
rect 8800 7108 8808 7142
rect 8842 7108 8850 7142
rect 8800 7100 8850 7108
rect 9350 7142 9400 7150
rect 9350 7108 9358 7142
rect 9392 7108 9400 7142
rect 9350 7100 9400 7108
rect 9900 7142 9950 7150
rect 9900 7108 9908 7142
rect 9942 7108 9950 7142
rect 9900 7100 9950 7108
rect 10450 7142 10500 7150
rect 10450 7108 10458 7142
rect 10492 7108 10500 7142
rect 10450 7100 10500 7108
rect 11000 7142 11050 7150
rect 11000 7108 11008 7142
rect 11042 7108 11050 7142
rect 11000 7100 11050 7108
rect 11550 7142 11600 7150
rect 11550 7108 11558 7142
rect 11592 7108 11600 7142
rect 11550 7100 11600 7108
rect 12100 7142 12150 7150
rect 12100 7108 12108 7142
rect 12142 7108 12150 7142
rect 12100 7100 12150 7108
rect 12650 7142 12700 7150
rect 12650 7108 12658 7142
rect 12692 7108 12700 7142
rect 12650 7100 12700 7108
rect 13200 7142 13250 7150
rect 13200 7108 13208 7142
rect 13242 7108 13250 7142
rect 13200 7100 13250 7108
rect 13750 7142 13800 7150
rect 13750 7108 13758 7142
rect 13792 7108 13800 7142
rect 13750 7100 13800 7108
rect -471 7077 -463 7094
rect -37 7077 -29 7094
rect 79 7077 87 7094
rect 513 7077 521 7094
rect 629 7077 637 7094
rect 1063 7077 1071 7094
rect 1179 7077 1187 7094
rect 1613 7077 1621 7094
rect 1729 7077 1737 7094
rect 2163 7077 2171 7094
rect 2279 7077 2287 7094
rect 2713 7077 2721 7094
rect 2829 7077 2837 7094
rect 3263 7077 3271 7094
rect 3379 7077 3387 7094
rect 3813 7077 3821 7094
rect 3929 7077 3937 7094
rect 4363 7077 4371 7094
rect 4479 7077 4487 7094
rect 4913 7077 4921 7094
rect 5029 7077 5037 7094
rect 5463 7077 5471 7094
rect 5579 7077 5587 7094
rect 6013 7077 6021 7094
rect 6129 7077 6137 7094
rect 6563 7077 6571 7094
rect 6679 7077 6687 7094
rect 7113 7077 7121 7094
rect 7229 7077 7237 7094
rect 7663 7077 7671 7094
rect 7779 7077 7787 7094
rect 8213 7077 8221 7094
rect 8329 7077 8337 7094
rect 8763 7077 8771 7094
rect 8879 7077 8887 7094
rect 9313 7077 9321 7094
rect 9429 7077 9437 7094
rect 9863 7077 9871 7094
rect 9979 7077 9987 7094
rect 10413 7077 10421 7094
rect 10529 7077 10537 7094
rect 10963 7077 10971 7094
rect 11079 7077 11087 7094
rect 11513 7077 11521 7094
rect 11629 7077 11637 7094
rect 12063 7077 12071 7094
rect 12179 7077 12187 7094
rect 12613 7077 12621 7094
rect 12729 7077 12737 7094
rect 13163 7077 13171 7094
rect 13279 7077 13287 7094
rect 13713 7077 13721 7094
rect -64 7071 -29 7077
rect 73 7071 527 7077
rect 629 7071 664 7077
rect -64 7063 -6 7071
rect -64 7036 -23 7063
rect -64 6637 -23 6664
rect -64 6629 -6 6637
rect 56 7063 544 7071
rect 73 7015 527 7063
rect 73 6685 135 7015
rect 465 6685 527 7015
rect 73 6637 527 6685
rect 56 6629 544 6637
rect 606 7063 664 7071
rect 623 7036 664 7063
rect 1036 7071 1071 7077
rect 1173 7071 1627 7077
rect 1729 7071 1764 7077
rect 1036 7063 1094 7071
rect 1036 7036 1077 7063
rect 623 6637 664 6664
rect 606 6629 664 6637
rect -64 6623 -29 6629
rect 73 6623 527 6629
rect 629 6623 664 6629
rect 1036 6637 1077 6664
rect 1036 6629 1094 6637
rect 1156 7063 1644 7071
rect 1173 7015 1627 7063
rect 1173 6685 1235 7015
rect 1565 6685 1627 7015
rect 1173 6637 1627 6685
rect 1156 6629 1644 6637
rect 1706 7063 1764 7071
rect 1723 7036 1764 7063
rect 2136 7071 2171 7077
rect 2273 7071 2727 7077
rect 2829 7071 2864 7077
rect 2136 7063 2194 7071
rect 2136 7036 2177 7063
rect 1723 6637 1764 6664
rect 1706 6629 1764 6637
rect 1036 6623 1071 6629
rect 1173 6623 1627 6629
rect 1729 6623 1764 6629
rect 2136 6637 2177 6664
rect 2136 6629 2194 6637
rect 2256 7063 2744 7071
rect 2273 7015 2727 7063
rect 2273 6685 2335 7015
rect 2665 6685 2727 7015
rect 2273 6637 2727 6685
rect 2256 6629 2744 6637
rect 2806 7063 2864 7071
rect 2823 7036 2864 7063
rect 3236 7071 3271 7077
rect 3373 7071 3827 7077
rect 3929 7071 3964 7077
rect 3236 7063 3294 7071
rect 3236 7036 3277 7063
rect 2823 6637 2864 6664
rect 2806 6629 2864 6637
rect 2136 6623 2171 6629
rect 2273 6623 2727 6629
rect 2829 6623 2864 6629
rect 3236 6637 3277 6664
rect 3236 6629 3294 6637
rect 3356 7063 3844 7071
rect 3373 7015 3827 7063
rect 3373 6685 3435 7015
rect 3765 6685 3827 7015
rect 3373 6637 3827 6685
rect 3356 6629 3844 6637
rect 3906 7063 3964 7071
rect 3923 7036 3964 7063
rect 4336 7071 4371 7077
rect 4473 7071 4927 7077
rect 5029 7071 5064 7077
rect 4336 7063 4394 7071
rect 4336 7036 4377 7063
rect 3923 6637 3964 6664
rect 3906 6629 3964 6637
rect 3236 6623 3271 6629
rect 3373 6623 3827 6629
rect 3929 6623 3964 6629
rect 4336 6637 4377 6664
rect 4336 6629 4394 6637
rect 4456 7063 4944 7071
rect 4473 7015 4927 7063
rect 4473 6685 4535 7015
rect 4865 6685 4927 7015
rect 4473 6637 4927 6685
rect 4456 6629 4944 6637
rect 5006 7063 5064 7071
rect 5023 7036 5064 7063
rect 5436 7071 5471 7077
rect 5573 7071 6027 7077
rect 6129 7071 6164 7077
rect 5436 7063 5494 7071
rect 5436 7036 5477 7063
rect 5023 6637 5064 6664
rect 5006 6629 5064 6637
rect 4336 6623 4371 6629
rect 4473 6623 4927 6629
rect 5029 6623 5064 6629
rect 5436 6637 5477 6664
rect 5436 6629 5494 6637
rect 5556 7063 6044 7071
rect 5573 7015 6027 7063
rect 5573 6685 5635 7015
rect 5965 6685 6027 7015
rect 5573 6637 6027 6685
rect 5556 6629 6044 6637
rect 6106 7063 6164 7071
rect 6123 7036 6164 7063
rect 6536 7071 6571 7077
rect 6673 7071 7127 7077
rect 7229 7071 7264 7077
rect 6536 7063 6594 7071
rect 6536 7036 6577 7063
rect 6123 6637 6164 6664
rect 6106 6629 6164 6637
rect 5436 6623 5471 6629
rect 5573 6623 6027 6629
rect 6129 6623 6164 6629
rect 6536 6637 6577 6664
rect 6536 6629 6594 6637
rect 6656 7063 7144 7071
rect 6673 7015 7127 7063
rect 6673 6685 6735 7015
rect 7065 6685 7127 7015
rect 6673 6637 7127 6685
rect 6656 6629 7144 6637
rect 7206 7063 7264 7071
rect 7223 7036 7264 7063
rect 7636 7071 7671 7077
rect 7773 7071 8227 7077
rect 8329 7071 8364 7077
rect 7636 7063 7694 7071
rect 7636 7036 7677 7063
rect 7223 6637 7264 6664
rect 7206 6629 7264 6637
rect 6536 6623 6571 6629
rect 6673 6623 7127 6629
rect 7229 6623 7264 6629
rect 7636 6637 7677 6664
rect 7636 6629 7694 6637
rect 7756 7063 8244 7071
rect 7773 7015 8227 7063
rect 7773 6685 7835 7015
rect 8165 6685 8227 7015
rect 7773 6637 8227 6685
rect 7756 6629 8244 6637
rect 8306 7063 8364 7071
rect 8323 7036 8364 7063
rect 8736 7071 8771 7077
rect 8873 7071 9327 7077
rect 9429 7071 9464 7077
rect 8736 7063 8794 7071
rect 8736 7036 8777 7063
rect 8323 6637 8364 6664
rect 8306 6629 8364 6637
rect 7636 6623 7671 6629
rect 7773 6623 8227 6629
rect 8329 6623 8364 6629
rect 8736 6637 8777 6664
rect 8736 6629 8794 6637
rect 8856 7063 9344 7071
rect 8873 7015 9327 7063
rect 8873 6685 8935 7015
rect 9265 6685 9327 7015
rect 8873 6637 9327 6685
rect 8856 6629 9344 6637
rect 9406 7063 9464 7071
rect 9423 7036 9464 7063
rect 9836 7071 9871 7077
rect 9973 7071 10427 7077
rect 10529 7071 10564 7077
rect 9836 7063 9894 7071
rect 9836 7036 9877 7063
rect 9423 6637 9464 6664
rect 9406 6629 9464 6637
rect 8736 6623 8771 6629
rect 8873 6623 9327 6629
rect 9429 6623 9464 6629
rect 9836 6637 9877 6664
rect 9836 6629 9894 6637
rect 9956 7063 10444 7071
rect 9973 7015 10427 7063
rect 9973 6685 10035 7015
rect 10365 6685 10427 7015
rect 9973 6637 10427 6685
rect 9956 6629 10444 6637
rect 10506 7063 10564 7071
rect 10523 7036 10564 7063
rect 10936 7071 10971 7077
rect 11073 7071 11527 7077
rect 11629 7071 11664 7077
rect 10936 7063 10994 7071
rect 10936 7036 10977 7063
rect 10523 6637 10564 6664
rect 10506 6629 10564 6637
rect 9836 6623 9871 6629
rect 9973 6623 10427 6629
rect 10529 6623 10564 6629
rect 10936 6637 10977 6664
rect 10936 6629 10994 6637
rect 11056 7063 11544 7071
rect 11073 7015 11527 7063
rect 11073 6685 11135 7015
rect 11465 6685 11527 7015
rect 11073 6637 11527 6685
rect 11056 6629 11544 6637
rect 11606 7063 11664 7071
rect 11623 7036 11664 7063
rect 12036 7071 12071 7077
rect 12173 7071 12627 7077
rect 12729 7071 12764 7077
rect 12036 7063 12094 7071
rect 12036 7036 12077 7063
rect 11623 6637 11664 6664
rect 11606 6629 11664 6637
rect 10936 6623 10971 6629
rect 11073 6623 11527 6629
rect 11629 6623 11664 6629
rect 12036 6637 12077 6664
rect 12036 6629 12094 6637
rect 12156 7063 12644 7071
rect 12173 7015 12627 7063
rect 12173 6685 12235 7015
rect 12565 6685 12627 7015
rect 12173 6637 12627 6685
rect 12156 6629 12644 6637
rect 12706 7063 12764 7071
rect 12723 7036 12764 7063
rect 13136 7071 13171 7077
rect 13273 7071 13727 7077
rect 13136 7063 13194 7071
rect 13136 7036 13177 7063
rect 12723 6637 12764 6664
rect 12706 6629 12764 6637
rect 12036 6623 12071 6629
rect 12173 6623 12627 6629
rect 12729 6623 12764 6629
rect 13136 6637 13177 6664
rect 13136 6629 13194 6637
rect 13256 7063 13727 7071
rect 13273 7015 13727 7063
rect 13273 6685 13335 7015
rect 13665 6685 13727 7015
rect 13273 6637 13727 6685
rect 13256 6629 13727 6637
rect 13136 6623 13171 6629
rect 13273 6623 13727 6629
rect -1025 6600 -725 6617
rect -471 6606 -463 6623
rect -37 6606 -29 6623
rect 79 6606 87 6623
rect 513 6606 521 6623
rect 629 6606 637 6623
rect 1063 6606 1071 6623
rect 1179 6606 1187 6623
rect 1613 6606 1621 6623
rect 1729 6606 1737 6623
rect 2163 6606 2171 6623
rect 2279 6606 2287 6623
rect 2713 6606 2721 6623
rect 2829 6606 2837 6623
rect 3263 6606 3271 6623
rect 3379 6606 3387 6623
rect 3813 6606 3821 6623
rect 3929 6606 3937 6623
rect 4363 6606 4371 6623
rect 4479 6606 4487 6623
rect 4913 6606 4921 6623
rect 5029 6606 5037 6623
rect 5463 6606 5471 6623
rect 5579 6606 5587 6623
rect 6013 6606 6021 6623
rect 6129 6606 6137 6623
rect 6563 6606 6571 6623
rect 6679 6606 6687 6623
rect 7113 6606 7121 6623
rect 7229 6606 7237 6623
rect 7663 6606 7671 6623
rect 7779 6606 7787 6623
rect 8213 6606 8221 6623
rect 8329 6606 8337 6623
rect 8763 6606 8771 6623
rect 8879 6606 8887 6623
rect 9313 6606 9321 6623
rect 9429 6606 9437 6623
rect 9863 6606 9871 6623
rect 9979 6606 9987 6623
rect 10413 6606 10421 6623
rect 10529 6606 10537 6623
rect 10963 6606 10971 6623
rect 11079 6606 11087 6623
rect 11513 6606 11521 6623
rect 11629 6606 11637 6623
rect 12063 6606 12071 6623
rect 12179 6606 12187 6623
rect 12613 6606 12621 6623
rect 12729 6606 12737 6623
rect 13163 6606 13171 6623
rect 13279 6606 13287 6623
rect 13713 6606 13721 6623
rect 13975 6617 13987 7150
rect 14263 6617 14275 7150
rect 13975 6600 14275 6617
rect -1025 6067 -1013 6600
rect -737 6067 -725 6600
rect -550 6592 -500 6600
rect -550 6558 -542 6592
rect -508 6558 -500 6592
rect -550 6550 -500 6558
rect 0 6592 50 6600
rect 0 6558 8 6592
rect 42 6558 50 6592
rect 0 6550 50 6558
rect 550 6592 600 6600
rect 550 6558 558 6592
rect 592 6558 600 6592
rect 550 6550 600 6558
rect 1100 6592 1150 6600
rect 1100 6558 1108 6592
rect 1142 6558 1150 6592
rect 1100 6550 1150 6558
rect 1650 6592 1700 6600
rect 1650 6558 1658 6592
rect 1692 6558 1700 6592
rect 1650 6550 1700 6558
rect 2200 6592 2250 6600
rect 2200 6558 2208 6592
rect 2242 6558 2250 6592
rect 2200 6550 2250 6558
rect 2750 6592 2800 6600
rect 2750 6558 2758 6592
rect 2792 6558 2800 6592
rect 2750 6550 2800 6558
rect 3300 6592 3350 6600
rect 3300 6558 3308 6592
rect 3342 6558 3350 6592
rect 3300 6550 3350 6558
rect 3850 6592 3900 6600
rect 3850 6558 3858 6592
rect 3892 6558 3900 6592
rect 3850 6550 3900 6558
rect 4400 6592 4450 6600
rect 4400 6558 4408 6592
rect 4442 6558 4450 6592
rect 4400 6550 4450 6558
rect 4950 6592 5000 6600
rect 4950 6558 4958 6592
rect 4992 6558 5000 6592
rect 4950 6550 5000 6558
rect 5500 6592 5550 6600
rect 5500 6558 5508 6592
rect 5542 6558 5550 6592
rect 5500 6550 5550 6558
rect 6050 6592 6100 6600
rect 6050 6558 6058 6592
rect 6092 6558 6100 6592
rect 6050 6550 6100 6558
rect 6600 6592 6650 6600
rect 6600 6558 6608 6592
rect 6642 6558 6650 6592
rect 6600 6550 6650 6558
rect 7150 6592 7200 6600
rect 7150 6558 7158 6592
rect 7192 6558 7200 6592
rect 7150 6550 7200 6558
rect 7700 6592 7750 6600
rect 7700 6558 7708 6592
rect 7742 6558 7750 6592
rect 7700 6550 7750 6558
rect 8250 6592 8300 6600
rect 8250 6558 8258 6592
rect 8292 6558 8300 6592
rect 8250 6550 8300 6558
rect 8800 6592 8850 6600
rect 8800 6558 8808 6592
rect 8842 6558 8850 6592
rect 8800 6550 8850 6558
rect 9350 6592 9400 6600
rect 9350 6558 9358 6592
rect 9392 6558 9400 6592
rect 9350 6550 9400 6558
rect 9900 6592 9950 6600
rect 9900 6558 9908 6592
rect 9942 6558 9950 6592
rect 9900 6550 9950 6558
rect 10450 6592 10500 6600
rect 10450 6558 10458 6592
rect 10492 6558 10500 6592
rect 10450 6550 10500 6558
rect 11000 6592 11050 6600
rect 11000 6558 11008 6592
rect 11042 6558 11050 6592
rect 11000 6550 11050 6558
rect 11550 6592 11600 6600
rect 11550 6558 11558 6592
rect 11592 6558 11600 6592
rect 11550 6550 11600 6558
rect 12100 6592 12150 6600
rect 12100 6558 12108 6592
rect 12142 6558 12150 6592
rect 12100 6550 12150 6558
rect 12650 6592 12700 6600
rect 12650 6558 12658 6592
rect 12692 6558 12700 6592
rect 12650 6550 12700 6558
rect 13200 6592 13250 6600
rect 13200 6558 13208 6592
rect 13242 6558 13250 6592
rect 13200 6550 13250 6558
rect 13750 6592 13800 6600
rect 13750 6558 13758 6592
rect 13792 6558 13800 6592
rect 13750 6550 13800 6558
rect -471 6527 -463 6544
rect -37 6527 -29 6544
rect 79 6527 87 6544
rect 513 6527 521 6544
rect 629 6527 637 6544
rect 1063 6527 1071 6544
rect 1179 6527 1187 6544
rect 1613 6527 1621 6544
rect 1729 6527 1737 6544
rect 2163 6527 2171 6544
rect 2279 6527 2287 6544
rect 2713 6527 2721 6544
rect 2829 6527 2837 6544
rect 3263 6527 3271 6544
rect 3379 6527 3387 6544
rect 3813 6527 3821 6544
rect 3929 6527 3937 6544
rect 4363 6527 4371 6544
rect 4479 6527 4487 6544
rect 4913 6527 4921 6544
rect 5029 6527 5037 6544
rect 5463 6527 5471 6544
rect 5579 6527 5587 6544
rect 6013 6527 6021 6544
rect 6129 6527 6137 6544
rect 6563 6527 6571 6544
rect 6679 6527 6687 6544
rect 7113 6527 7121 6544
rect 7229 6527 7237 6544
rect 7663 6527 7671 6544
rect 7779 6527 7787 6544
rect 8213 6527 8221 6544
rect 8329 6527 8337 6544
rect 8763 6527 8771 6544
rect 8879 6527 8887 6544
rect 9313 6527 9321 6544
rect 9429 6527 9437 6544
rect 9863 6527 9871 6544
rect 9979 6527 9987 6544
rect 10413 6527 10421 6544
rect 10529 6527 10537 6544
rect 10963 6527 10971 6544
rect 11079 6527 11087 6544
rect 11513 6527 11521 6544
rect 11629 6527 11637 6544
rect 12063 6527 12071 6544
rect 12179 6527 12187 6544
rect 12613 6527 12621 6544
rect 12729 6527 12737 6544
rect 13163 6527 13171 6544
rect 13279 6527 13287 6544
rect 13713 6527 13721 6544
rect -477 6521 -23 6527
rect 79 6521 114 6527
rect -477 6513 -6 6521
rect -477 6465 -23 6513
rect -477 6135 -415 6465
rect -85 6135 -23 6465
rect -477 6087 -23 6135
rect -477 6079 -6 6087
rect 56 6513 114 6521
rect 73 6486 114 6513
rect 486 6521 521 6527
rect 623 6521 1077 6527
rect 1179 6521 1214 6527
rect 486 6513 544 6521
rect 486 6486 527 6513
rect 73 6087 114 6114
rect 56 6079 114 6087
rect -477 6073 -23 6079
rect 79 6073 114 6079
rect 486 6087 527 6114
rect 486 6079 544 6087
rect 606 6513 1094 6521
rect 623 6465 1077 6513
rect 623 6135 685 6465
rect 1015 6135 1077 6465
rect 623 6087 1077 6135
rect 606 6079 1094 6087
rect 1156 6513 1214 6521
rect 1173 6486 1214 6513
rect 1586 6521 1621 6527
rect 1723 6521 2177 6527
rect 2279 6521 2314 6527
rect 1586 6513 1644 6521
rect 1586 6486 1627 6513
rect 1173 6087 1214 6114
rect 1156 6079 1214 6087
rect 486 6073 521 6079
rect 623 6073 1077 6079
rect 1179 6073 1214 6079
rect 1586 6087 1627 6114
rect 1586 6079 1644 6087
rect 1706 6513 2194 6521
rect 1723 6465 2177 6513
rect 1723 6135 1785 6465
rect 2115 6135 2177 6465
rect 1723 6087 2177 6135
rect 1706 6079 2194 6087
rect 2256 6513 2314 6521
rect 2273 6486 2314 6513
rect 2686 6521 2721 6527
rect 2823 6521 3277 6527
rect 3379 6521 3414 6527
rect 2686 6513 2744 6521
rect 2686 6486 2727 6513
rect 2273 6087 2314 6114
rect 2256 6079 2314 6087
rect 1586 6073 1621 6079
rect 1723 6073 2177 6079
rect 2279 6073 2314 6079
rect 2686 6087 2727 6114
rect 2686 6079 2744 6087
rect 2806 6513 3294 6521
rect 2823 6465 3277 6513
rect 2823 6135 2885 6465
rect 3215 6135 3277 6465
rect 2823 6087 3277 6135
rect 2806 6079 3294 6087
rect 3356 6513 3414 6521
rect 3373 6486 3414 6513
rect 3786 6521 3821 6527
rect 3923 6521 4377 6527
rect 4479 6521 4514 6527
rect 3786 6513 3844 6521
rect 3786 6486 3827 6513
rect 3373 6087 3414 6114
rect 3356 6079 3414 6087
rect 2686 6073 2721 6079
rect 2823 6073 3277 6079
rect 3379 6073 3414 6079
rect 3786 6087 3827 6114
rect 3786 6079 3844 6087
rect 3906 6513 4394 6521
rect 3923 6465 4377 6513
rect 3923 6135 3985 6465
rect 4315 6135 4377 6465
rect 3923 6087 4377 6135
rect 3906 6079 4394 6087
rect 4456 6513 4514 6521
rect 4473 6486 4514 6513
rect 4886 6521 4921 6527
rect 5023 6521 5477 6527
rect 5579 6521 5614 6527
rect 4886 6513 4944 6521
rect 4886 6486 4927 6513
rect 4473 6087 4514 6114
rect 4456 6079 4514 6087
rect 3786 6073 3821 6079
rect 3923 6073 4377 6079
rect 4479 6073 4514 6079
rect 4886 6087 4927 6114
rect 4886 6079 4944 6087
rect 5006 6513 5494 6521
rect 5023 6465 5477 6513
rect 5023 6135 5085 6465
rect 5415 6135 5477 6465
rect 5023 6087 5477 6135
rect 5006 6079 5494 6087
rect 5556 6513 5614 6521
rect 5573 6486 5614 6513
rect 5986 6521 6021 6527
rect 6123 6521 6577 6527
rect 6679 6521 6714 6527
rect 5986 6513 6044 6521
rect 5986 6486 6027 6513
rect 5573 6087 5614 6114
rect 5556 6079 5614 6087
rect 4886 6073 4921 6079
rect 5023 6073 5477 6079
rect 5579 6073 5614 6079
rect 5986 6087 6027 6114
rect 5986 6079 6044 6087
rect 6106 6513 6594 6521
rect 6123 6465 6577 6513
rect 6123 6135 6185 6465
rect 6515 6135 6577 6465
rect 6123 6087 6577 6135
rect 6106 6079 6594 6087
rect 6656 6513 6714 6521
rect 6673 6486 6714 6513
rect 7086 6521 7121 6527
rect 7223 6521 7677 6527
rect 7779 6521 7814 6527
rect 7086 6513 7144 6521
rect 7086 6486 7127 6513
rect 6673 6087 6714 6114
rect 6656 6079 6714 6087
rect 5986 6073 6021 6079
rect 6123 6073 6577 6079
rect 6679 6073 6714 6079
rect 7086 6087 7127 6114
rect 7086 6079 7144 6087
rect 7206 6513 7694 6521
rect 7223 6465 7677 6513
rect 7223 6135 7285 6465
rect 7615 6135 7677 6465
rect 7223 6087 7677 6135
rect 7206 6079 7694 6087
rect 7756 6513 7814 6521
rect 7773 6486 7814 6513
rect 8186 6521 8221 6527
rect 8323 6521 8777 6527
rect 8879 6521 8914 6527
rect 8186 6513 8244 6521
rect 8186 6486 8227 6513
rect 7773 6087 7814 6114
rect 7756 6079 7814 6087
rect 7086 6073 7121 6079
rect 7223 6073 7677 6079
rect 7779 6073 7814 6079
rect 8186 6087 8227 6114
rect 8186 6079 8244 6087
rect 8306 6513 8794 6521
rect 8323 6465 8777 6513
rect 8323 6135 8385 6465
rect 8715 6135 8777 6465
rect 8323 6087 8777 6135
rect 8306 6079 8794 6087
rect 8856 6513 8914 6521
rect 8873 6486 8914 6513
rect 9286 6521 9321 6527
rect 9423 6521 9877 6527
rect 9979 6521 10014 6527
rect 9286 6513 9344 6521
rect 9286 6486 9327 6513
rect 8873 6087 8914 6114
rect 8856 6079 8914 6087
rect 8186 6073 8221 6079
rect 8323 6073 8777 6079
rect 8879 6073 8914 6079
rect 9286 6087 9327 6114
rect 9286 6079 9344 6087
rect 9406 6513 9894 6521
rect 9423 6465 9877 6513
rect 9423 6135 9485 6465
rect 9815 6135 9877 6465
rect 9423 6087 9877 6135
rect 9406 6079 9894 6087
rect 9956 6513 10014 6521
rect 9973 6486 10014 6513
rect 10386 6521 10421 6527
rect 10523 6521 10977 6527
rect 11079 6521 11114 6527
rect 10386 6513 10444 6521
rect 10386 6486 10427 6513
rect 9973 6087 10014 6114
rect 9956 6079 10014 6087
rect 9286 6073 9321 6079
rect 9423 6073 9877 6079
rect 9979 6073 10014 6079
rect 10386 6087 10427 6114
rect 10386 6079 10444 6087
rect 10506 6513 10994 6521
rect 10523 6465 10977 6513
rect 10523 6135 10585 6465
rect 10915 6135 10977 6465
rect 10523 6087 10977 6135
rect 10506 6079 10994 6087
rect 11056 6513 11114 6521
rect 11073 6486 11114 6513
rect 11486 6521 11521 6527
rect 11623 6521 12077 6527
rect 12179 6521 12214 6527
rect 11486 6513 11544 6521
rect 11486 6486 11527 6513
rect 11073 6087 11114 6114
rect 11056 6079 11114 6087
rect 10386 6073 10421 6079
rect 10523 6073 10977 6079
rect 11079 6073 11114 6079
rect 11486 6087 11527 6114
rect 11486 6079 11544 6087
rect 11606 6513 12094 6521
rect 11623 6465 12077 6513
rect 11623 6135 11685 6465
rect 12015 6135 12077 6465
rect 11623 6087 12077 6135
rect 11606 6079 12094 6087
rect 12156 6513 12214 6521
rect 12173 6486 12214 6513
rect 12586 6521 12621 6527
rect 12723 6521 13177 6527
rect 13279 6521 13314 6527
rect 12586 6513 12644 6521
rect 12586 6486 12627 6513
rect 12173 6087 12214 6114
rect 12156 6079 12214 6087
rect 11486 6073 11521 6079
rect 11623 6073 12077 6079
rect 12179 6073 12214 6079
rect 12586 6087 12627 6114
rect 12586 6079 12644 6087
rect 12706 6513 13194 6521
rect 12723 6465 13177 6513
rect 12723 6135 12785 6465
rect 13115 6135 13177 6465
rect 12723 6087 13177 6135
rect 12706 6079 13194 6087
rect 13256 6513 13314 6521
rect 13273 6486 13314 6513
rect 13273 6087 13314 6114
rect 13256 6079 13314 6087
rect 12586 6073 12621 6079
rect 12723 6073 13177 6079
rect 13279 6073 13314 6079
rect -1025 6050 -725 6067
rect -471 6056 -463 6073
rect -37 6056 -29 6073
rect 79 6056 87 6073
rect 513 6056 521 6073
rect 629 6056 637 6073
rect 1063 6056 1071 6073
rect 1179 6056 1187 6073
rect 1613 6056 1621 6073
rect 1729 6056 1737 6073
rect 2163 6056 2171 6073
rect 2279 6056 2287 6073
rect 2713 6056 2721 6073
rect 2829 6056 2837 6073
rect 3263 6056 3271 6073
rect 3379 6056 3387 6073
rect 3813 6056 3821 6073
rect 3929 6056 3937 6073
rect 4363 6056 4371 6073
rect 4479 6056 4487 6073
rect 4913 6056 4921 6073
rect 5029 6056 5037 6073
rect 5463 6056 5471 6073
rect 5579 6056 5587 6073
rect 6013 6056 6021 6073
rect 6129 6056 6137 6073
rect 6563 6056 6571 6073
rect 6679 6056 6687 6073
rect 7113 6056 7121 6073
rect 7229 6056 7237 6073
rect 7663 6056 7671 6073
rect 7779 6056 7787 6073
rect 8213 6056 8221 6073
rect 8329 6056 8337 6073
rect 8763 6056 8771 6073
rect 8879 6056 8887 6073
rect 9313 6056 9321 6073
rect 9429 6056 9437 6073
rect 9863 6056 9871 6073
rect 9979 6056 9987 6073
rect 10413 6056 10421 6073
rect 10529 6056 10537 6073
rect 10963 6056 10971 6073
rect 11079 6056 11087 6073
rect 11513 6056 11521 6073
rect 11629 6056 11637 6073
rect 12063 6056 12071 6073
rect 12179 6056 12187 6073
rect 12613 6056 12621 6073
rect 12729 6056 12737 6073
rect 13163 6056 13171 6073
rect 13279 6056 13287 6073
rect 13713 6056 13721 6073
rect 13975 6069 13987 6600
rect 14263 6069 14275 6600
rect 13975 6050 14275 6069
rect -1025 5517 -1013 6050
rect -737 5517 -725 6050
rect -550 6042 -500 6050
rect -550 6008 -542 6042
rect -508 6008 -500 6042
rect -550 6000 -500 6008
rect 0 6042 50 6050
rect 0 6008 8 6042
rect 42 6008 50 6042
rect 0 6000 50 6008
rect 550 6042 600 6050
rect 550 6008 558 6042
rect 592 6008 600 6042
rect 550 6000 600 6008
rect 1100 6042 1150 6050
rect 1100 6008 1108 6042
rect 1142 6008 1150 6042
rect 1100 6000 1150 6008
rect 1650 6042 1700 6050
rect 1650 6008 1658 6042
rect 1692 6008 1700 6042
rect 1650 6000 1700 6008
rect 2200 6042 2250 6050
rect 2200 6008 2208 6042
rect 2242 6008 2250 6042
rect 2200 6000 2250 6008
rect 2750 6042 2800 6050
rect 2750 6008 2758 6042
rect 2792 6008 2800 6042
rect 2750 6000 2800 6008
rect 3300 6042 3350 6050
rect 3300 6008 3308 6042
rect 3342 6008 3350 6042
rect 3300 6000 3350 6008
rect 3850 6042 3900 6050
rect 3850 6008 3858 6042
rect 3892 6008 3900 6042
rect 3850 6000 3900 6008
rect 4400 6042 4450 6050
rect 4400 6008 4408 6042
rect 4442 6008 4450 6042
rect 4400 6000 4450 6008
rect 4950 6042 5000 6050
rect 4950 6008 4958 6042
rect 4992 6008 5000 6042
rect 4950 6000 5000 6008
rect 5500 6042 5550 6050
rect 5500 6008 5508 6042
rect 5542 6008 5550 6042
rect 5500 6000 5550 6008
rect 6050 6042 6100 6050
rect 6050 6008 6058 6042
rect 6092 6008 6100 6042
rect 6050 6000 6100 6008
rect 6600 6042 6650 6050
rect 6600 6008 6608 6042
rect 6642 6008 6650 6042
rect 6600 6000 6650 6008
rect 7150 6042 7200 6050
rect 7150 6008 7158 6042
rect 7192 6008 7200 6042
rect 7150 6000 7200 6008
rect 7700 6042 7750 6050
rect 7700 6008 7708 6042
rect 7742 6008 7750 6042
rect 7700 6000 7750 6008
rect 8250 6042 8300 6050
rect 8250 6008 8258 6042
rect 8292 6008 8300 6042
rect 8250 6000 8300 6008
rect 8800 6042 8850 6050
rect 8800 6008 8808 6042
rect 8842 6008 8850 6042
rect 8800 6000 8850 6008
rect 9350 6042 9400 6050
rect 9350 6008 9358 6042
rect 9392 6008 9400 6042
rect 9350 6000 9400 6008
rect 9900 6042 9950 6050
rect 9900 6008 9908 6042
rect 9942 6008 9950 6042
rect 9900 6000 9950 6008
rect 10450 6042 10500 6050
rect 10450 6008 10458 6042
rect 10492 6008 10500 6042
rect 10450 6000 10500 6008
rect 11000 6042 11050 6050
rect 11000 6008 11008 6042
rect 11042 6008 11050 6042
rect 11000 6000 11050 6008
rect 11550 6042 11600 6050
rect 11550 6008 11558 6042
rect 11592 6008 11600 6042
rect 11550 6000 11600 6008
rect 12100 6042 12150 6050
rect 12100 6008 12108 6042
rect 12142 6008 12150 6042
rect 12100 6000 12150 6008
rect 12650 6042 12700 6050
rect 12650 6008 12658 6042
rect 12692 6008 12700 6042
rect 12650 6000 12700 6008
rect 13200 6042 13250 6050
rect 13200 6008 13208 6042
rect 13242 6008 13250 6042
rect 13200 6000 13250 6008
rect 13750 6042 13800 6050
rect 13750 6008 13758 6042
rect 13792 6008 13800 6042
rect 13750 6000 13800 6008
rect -471 5977 -463 5994
rect -37 5977 -29 5994
rect 79 5977 87 5994
rect 513 5977 521 5994
rect 629 5977 637 5994
rect 1063 5977 1071 5994
rect 1179 5977 1187 5994
rect 1613 5977 1621 5994
rect 1729 5977 1737 5994
rect 2163 5977 2171 5994
rect 2279 5977 2287 5994
rect 2713 5977 2721 5994
rect 2829 5977 2837 5994
rect 3263 5977 3271 5994
rect 3379 5977 3387 5994
rect 3813 5977 3821 5994
rect 3929 5977 3937 5994
rect 4363 5977 4371 5994
rect 4479 5977 4487 5994
rect 4913 5977 4921 5994
rect 5029 5977 5037 5994
rect 5463 5977 5471 5994
rect 5579 5977 5587 5994
rect 6013 5977 6021 5994
rect 6129 5977 6137 5994
rect 6563 5977 6571 5994
rect 6679 5977 6687 5994
rect 7113 5977 7121 5994
rect 7229 5977 7237 5994
rect 7663 5977 7671 5994
rect 7779 5977 7787 5994
rect 8213 5977 8221 5994
rect 8329 5977 8337 5994
rect 8763 5977 8771 5994
rect 8879 5977 8887 5994
rect 9313 5977 9321 5994
rect 9429 5977 9437 5994
rect 9863 5977 9871 5994
rect 9979 5977 9987 5994
rect 10413 5977 10421 5994
rect 10529 5977 10537 5994
rect 10963 5977 10971 5994
rect 11079 5977 11087 5994
rect 11513 5977 11521 5994
rect 11629 5977 11637 5994
rect 12063 5977 12071 5994
rect 12179 5977 12187 5994
rect 12613 5977 12621 5994
rect 12729 5977 12737 5994
rect 13163 5977 13171 5994
rect 13279 5977 13287 5994
rect 13713 5977 13721 5994
rect -64 5971 -29 5977
rect 73 5971 527 5977
rect 629 5971 664 5977
rect -64 5963 -6 5971
rect -64 5936 -23 5963
rect -64 5537 -23 5564
rect -64 5529 -6 5537
rect 56 5963 544 5971
rect 73 5915 527 5963
rect 73 5585 135 5915
rect 465 5585 527 5915
rect 73 5537 527 5585
rect 56 5529 544 5537
rect 606 5963 664 5971
rect 623 5936 664 5963
rect 1036 5971 1071 5977
rect 1173 5971 1627 5977
rect 1729 5971 1764 5977
rect 1036 5963 1094 5971
rect 1036 5936 1077 5963
rect 623 5537 664 5564
rect 606 5529 664 5537
rect -64 5523 -29 5529
rect 73 5523 527 5529
rect 629 5523 664 5529
rect 1036 5537 1077 5564
rect 1036 5529 1094 5537
rect 1156 5963 1644 5971
rect 1173 5915 1627 5963
rect 1173 5585 1235 5915
rect 1565 5585 1627 5915
rect 1173 5537 1627 5585
rect 1156 5529 1644 5537
rect 1706 5963 1764 5971
rect 1723 5936 1764 5963
rect 2136 5971 2171 5977
rect 2273 5971 2727 5977
rect 2829 5971 2864 5977
rect 2136 5963 2194 5971
rect 2136 5936 2177 5963
rect 1723 5537 1764 5564
rect 1706 5529 1764 5537
rect 1036 5523 1071 5529
rect 1173 5523 1627 5529
rect 1729 5523 1764 5529
rect 2136 5537 2177 5564
rect 2136 5529 2194 5537
rect 2256 5963 2744 5971
rect 2273 5915 2727 5963
rect 2273 5585 2335 5915
rect 2665 5585 2727 5915
rect 2273 5537 2727 5585
rect 2256 5529 2744 5537
rect 2806 5963 2864 5971
rect 2823 5936 2864 5963
rect 3236 5971 3271 5977
rect 3373 5971 3827 5977
rect 3929 5971 3964 5977
rect 3236 5963 3294 5971
rect 3236 5936 3277 5963
rect 2823 5537 2864 5564
rect 2806 5529 2864 5537
rect 2136 5523 2171 5529
rect 2273 5523 2727 5529
rect 2829 5523 2864 5529
rect 3236 5537 3277 5564
rect 3236 5529 3294 5537
rect 3356 5963 3844 5971
rect 3373 5915 3827 5963
rect 3373 5585 3435 5915
rect 3765 5585 3827 5915
rect 3373 5537 3827 5585
rect 3356 5529 3844 5537
rect 3906 5963 3964 5971
rect 3923 5936 3964 5963
rect 4336 5971 4371 5977
rect 4473 5971 4927 5977
rect 5029 5971 5064 5977
rect 4336 5963 4394 5971
rect 4336 5936 4377 5963
rect 3923 5537 3964 5564
rect 3906 5529 3964 5537
rect 3236 5523 3271 5529
rect 3373 5523 3827 5529
rect 3929 5523 3964 5529
rect 4336 5537 4377 5564
rect 4336 5529 4394 5537
rect 4456 5963 4944 5971
rect 4473 5915 4927 5963
rect 4473 5585 4535 5915
rect 4865 5585 4927 5915
rect 4473 5537 4927 5585
rect 4456 5529 4944 5537
rect 5006 5963 5064 5971
rect 5023 5936 5064 5963
rect 5436 5971 5471 5977
rect 5573 5971 6027 5977
rect 6129 5971 6164 5977
rect 5436 5963 5494 5971
rect 5436 5936 5477 5963
rect 5023 5537 5064 5564
rect 5006 5529 5064 5537
rect 4336 5523 4371 5529
rect 4473 5523 4927 5529
rect 5029 5523 5064 5529
rect 5436 5537 5477 5564
rect 5436 5529 5494 5537
rect 5556 5963 6044 5971
rect 5573 5915 6027 5963
rect 5573 5585 5635 5915
rect 5965 5585 6027 5915
rect 5573 5537 6027 5585
rect 5556 5529 6044 5537
rect 6106 5963 6164 5971
rect 6123 5936 6164 5963
rect 6536 5971 6571 5977
rect 6673 5971 7127 5977
rect 7229 5971 7264 5977
rect 6536 5963 6594 5971
rect 6536 5936 6577 5963
rect 6123 5537 6164 5564
rect 6106 5529 6164 5537
rect 5436 5523 5471 5529
rect 5573 5523 6027 5529
rect 6129 5523 6164 5529
rect 6536 5537 6577 5564
rect 6536 5529 6594 5537
rect 6656 5963 7144 5971
rect 6673 5915 7127 5963
rect 6673 5585 6735 5915
rect 7065 5585 7127 5915
rect 6673 5537 7127 5585
rect 6656 5529 7144 5537
rect 7206 5963 7264 5971
rect 7223 5936 7264 5963
rect 7636 5971 7671 5977
rect 7773 5971 8227 5977
rect 8329 5971 8364 5977
rect 7636 5963 7694 5971
rect 7636 5936 7677 5963
rect 7223 5537 7264 5564
rect 7206 5529 7264 5537
rect 6536 5523 6571 5529
rect 6673 5523 7127 5529
rect 7229 5523 7264 5529
rect 7636 5537 7677 5564
rect 7636 5529 7694 5537
rect 7756 5963 8244 5971
rect 7773 5915 8227 5963
rect 7773 5585 7835 5915
rect 8165 5585 8227 5915
rect 7773 5537 8227 5585
rect 7756 5529 8244 5537
rect 8306 5963 8364 5971
rect 8323 5936 8364 5963
rect 8736 5971 8771 5977
rect 8873 5971 9327 5977
rect 9429 5971 9464 5977
rect 8736 5963 8794 5971
rect 8736 5936 8777 5963
rect 8323 5537 8364 5564
rect 8306 5529 8364 5537
rect 7636 5523 7671 5529
rect 7773 5523 8227 5529
rect 8329 5523 8364 5529
rect 8736 5537 8777 5564
rect 8736 5529 8794 5537
rect 8856 5963 9344 5971
rect 8873 5915 9327 5963
rect 8873 5585 8935 5915
rect 9265 5585 9327 5915
rect 8873 5537 9327 5585
rect 8856 5529 9344 5537
rect 9406 5963 9464 5971
rect 9423 5936 9464 5963
rect 9836 5971 9871 5977
rect 9973 5971 10427 5977
rect 10529 5971 10564 5977
rect 9836 5963 9894 5971
rect 9836 5936 9877 5963
rect 9423 5537 9464 5564
rect 9406 5529 9464 5537
rect 8736 5523 8771 5529
rect 8873 5523 9327 5529
rect 9429 5523 9464 5529
rect 9836 5537 9877 5564
rect 9836 5529 9894 5537
rect 9956 5963 10444 5971
rect 9973 5915 10427 5963
rect 9973 5585 10035 5915
rect 10365 5585 10427 5915
rect 9973 5537 10427 5585
rect 9956 5529 10444 5537
rect 10506 5963 10564 5971
rect 10523 5936 10564 5963
rect 10936 5971 10971 5977
rect 11073 5971 11527 5977
rect 11629 5971 11664 5977
rect 10936 5963 10994 5971
rect 10936 5936 10977 5963
rect 10523 5537 10564 5564
rect 10506 5529 10564 5537
rect 9836 5523 9871 5529
rect 9973 5523 10427 5529
rect 10529 5523 10564 5529
rect 10936 5537 10977 5564
rect 10936 5529 10994 5537
rect 11056 5963 11544 5971
rect 11073 5915 11527 5963
rect 11073 5585 11135 5915
rect 11465 5585 11527 5915
rect 11073 5537 11527 5585
rect 11056 5529 11544 5537
rect 11606 5963 11664 5971
rect 11623 5936 11664 5963
rect 12036 5971 12071 5977
rect 12173 5971 12627 5977
rect 12729 5971 12764 5977
rect 12036 5963 12094 5971
rect 12036 5936 12077 5963
rect 11623 5537 11664 5564
rect 11606 5529 11664 5537
rect 10936 5523 10971 5529
rect 11073 5523 11527 5529
rect 11629 5523 11664 5529
rect 12036 5537 12077 5564
rect 12036 5529 12094 5537
rect 12156 5963 12644 5971
rect 12173 5915 12627 5963
rect 12173 5585 12235 5915
rect 12565 5585 12627 5915
rect 12173 5537 12627 5585
rect 12156 5529 12644 5537
rect 12706 5963 12764 5971
rect 12723 5936 12764 5963
rect 13136 5971 13171 5977
rect 13273 5971 13727 5977
rect 13136 5963 13194 5971
rect 13136 5936 13177 5963
rect 12723 5537 12764 5564
rect 12706 5529 12764 5537
rect 12036 5523 12071 5529
rect 12173 5523 12627 5529
rect 12729 5523 12764 5529
rect 13136 5537 13177 5564
rect 13136 5529 13194 5537
rect 13256 5963 13727 5971
rect 13273 5915 13727 5963
rect 13273 5585 13335 5915
rect 13665 5585 13727 5915
rect 13273 5537 13727 5585
rect 13256 5529 13727 5537
rect 13136 5523 13171 5529
rect 13273 5523 13727 5529
rect -1025 5500 -725 5517
rect -471 5506 -463 5523
rect -37 5506 -29 5523
rect 79 5506 87 5523
rect 513 5506 521 5523
rect 629 5506 637 5523
rect 1063 5506 1071 5523
rect 1179 5506 1187 5523
rect 1613 5506 1621 5523
rect 1729 5506 1737 5523
rect 2163 5506 2171 5523
rect 2279 5506 2287 5523
rect 2713 5506 2721 5523
rect 2829 5506 2837 5523
rect 3263 5506 3271 5523
rect 3379 5506 3387 5523
rect 3813 5506 3821 5523
rect 3929 5506 3937 5523
rect 4363 5506 4371 5523
rect 4479 5506 4487 5523
rect 4913 5506 4921 5523
rect 5029 5506 5037 5523
rect 5463 5506 5471 5523
rect 5579 5506 5587 5523
rect 6013 5506 6021 5523
rect 6129 5506 6137 5523
rect 6563 5506 6571 5523
rect 6679 5506 6687 5523
rect 7113 5506 7121 5523
rect 7229 5506 7237 5523
rect 7663 5506 7671 5523
rect 7779 5506 7787 5523
rect 8213 5506 8221 5523
rect 8329 5506 8337 5523
rect 8763 5506 8771 5523
rect 8879 5506 8887 5523
rect 9313 5506 9321 5523
rect 9429 5506 9437 5523
rect 9863 5506 9871 5523
rect 9979 5506 9987 5523
rect 10413 5506 10421 5523
rect 10529 5506 10537 5523
rect 10963 5506 10971 5523
rect 11079 5506 11087 5523
rect 11513 5506 11521 5523
rect 11629 5506 11637 5523
rect 12063 5506 12071 5523
rect 12179 5506 12187 5523
rect 12613 5506 12621 5523
rect 12729 5506 12737 5523
rect 13163 5506 13171 5523
rect 13279 5506 13287 5523
rect 13713 5506 13721 5523
rect 13975 5517 13987 6050
rect 14263 5517 14275 6050
rect 13975 5500 14275 5517
rect -1025 4967 -1013 5500
rect -737 4967 -725 5500
rect -550 5492 -500 5500
rect -550 5458 -542 5492
rect -508 5458 -500 5492
rect -550 5450 -500 5458
rect 0 5492 50 5500
rect 0 5458 8 5492
rect 42 5458 50 5492
rect 0 5450 50 5458
rect 550 5492 600 5500
rect 550 5458 558 5492
rect 592 5458 600 5492
rect 550 5450 600 5458
rect 1100 5492 1150 5500
rect 1100 5458 1108 5492
rect 1142 5458 1150 5492
rect 1100 5450 1150 5458
rect 1650 5492 1700 5500
rect 1650 5458 1658 5492
rect 1692 5458 1700 5492
rect 1650 5450 1700 5458
rect 2200 5492 2250 5500
rect 2200 5458 2208 5492
rect 2242 5458 2250 5492
rect 2200 5450 2250 5458
rect 2750 5492 2800 5500
rect 2750 5458 2758 5492
rect 2792 5458 2800 5492
rect 2750 5450 2800 5458
rect 3300 5492 3350 5500
rect 3300 5458 3308 5492
rect 3342 5458 3350 5492
rect 3300 5450 3350 5458
rect 3850 5492 3900 5500
rect 3850 5458 3858 5492
rect 3892 5458 3900 5492
rect 3850 5450 3900 5458
rect 4400 5492 4450 5500
rect 4400 5458 4408 5492
rect 4442 5458 4450 5492
rect 4400 5450 4450 5458
rect 4950 5492 5000 5500
rect 4950 5458 4958 5492
rect 4992 5458 5000 5492
rect 4950 5450 5000 5458
rect 5500 5492 5550 5500
rect 5500 5458 5508 5492
rect 5542 5458 5550 5492
rect 5500 5450 5550 5458
rect 6050 5492 6100 5500
rect 6050 5458 6058 5492
rect 6092 5458 6100 5492
rect 6050 5450 6100 5458
rect 6600 5492 6650 5500
rect 6600 5458 6608 5492
rect 6642 5458 6650 5492
rect 6600 5450 6650 5458
rect 7150 5492 7200 5500
rect 7150 5458 7158 5492
rect 7192 5458 7200 5492
rect 7150 5450 7200 5458
rect 7700 5492 7750 5500
rect 7700 5458 7708 5492
rect 7742 5458 7750 5492
rect 7700 5450 7750 5458
rect 8250 5492 8300 5500
rect 8250 5458 8258 5492
rect 8292 5458 8300 5492
rect 8250 5450 8300 5458
rect 8800 5492 8850 5500
rect 8800 5458 8808 5492
rect 8842 5458 8850 5492
rect 8800 5450 8850 5458
rect 9350 5492 9400 5500
rect 9350 5458 9358 5492
rect 9392 5458 9400 5492
rect 9350 5450 9400 5458
rect 9900 5492 9950 5500
rect 9900 5458 9908 5492
rect 9942 5458 9950 5492
rect 9900 5450 9950 5458
rect 10450 5492 10500 5500
rect 10450 5458 10458 5492
rect 10492 5458 10500 5492
rect 10450 5450 10500 5458
rect 11000 5492 11050 5500
rect 11000 5458 11008 5492
rect 11042 5458 11050 5492
rect 11000 5450 11050 5458
rect 11550 5492 11600 5500
rect 11550 5458 11558 5492
rect 11592 5458 11600 5492
rect 11550 5450 11600 5458
rect 12100 5492 12150 5500
rect 12100 5458 12108 5492
rect 12142 5458 12150 5492
rect 12100 5450 12150 5458
rect 12650 5492 12700 5500
rect 12650 5458 12658 5492
rect 12692 5458 12700 5492
rect 12650 5450 12700 5458
rect 13200 5492 13250 5500
rect 13200 5458 13208 5492
rect 13242 5458 13250 5492
rect 13200 5450 13250 5458
rect 13750 5492 13800 5500
rect 13750 5458 13758 5492
rect 13792 5458 13800 5492
rect 13750 5450 13800 5458
rect -471 5427 -463 5444
rect -37 5427 -29 5444
rect 79 5427 87 5444
rect 513 5427 521 5444
rect 629 5427 637 5444
rect 1063 5427 1071 5444
rect 1179 5427 1187 5444
rect 1613 5427 1621 5444
rect 1729 5427 1737 5444
rect 2163 5427 2171 5444
rect 2279 5427 2287 5444
rect 2713 5427 2721 5444
rect 2829 5427 2837 5444
rect 3263 5427 3271 5444
rect 3379 5427 3387 5444
rect 3813 5427 3821 5444
rect 3929 5427 3937 5444
rect 4363 5427 4371 5444
rect 4479 5427 4487 5444
rect 4913 5427 4921 5444
rect 5029 5427 5037 5444
rect 5463 5427 5471 5444
rect 5579 5427 5587 5444
rect 6013 5427 6021 5444
rect 6129 5427 6137 5444
rect 6563 5427 6571 5444
rect 6679 5427 6687 5444
rect 7113 5427 7121 5444
rect 7229 5427 7237 5444
rect 7663 5427 7671 5444
rect 7779 5427 7787 5444
rect 8213 5427 8221 5444
rect 8329 5427 8337 5444
rect 8763 5427 8771 5444
rect 8879 5427 8887 5444
rect 9313 5427 9321 5444
rect 9429 5427 9437 5444
rect 9863 5427 9871 5444
rect 9979 5427 9987 5444
rect 10413 5427 10421 5444
rect 10529 5427 10537 5444
rect 10963 5427 10971 5444
rect 11079 5427 11087 5444
rect 11513 5427 11521 5444
rect 11629 5427 11637 5444
rect 12063 5427 12071 5444
rect 12179 5427 12187 5444
rect 12613 5427 12621 5444
rect 12729 5427 12737 5444
rect 13163 5427 13171 5444
rect 13279 5427 13287 5444
rect 13713 5427 13721 5444
rect -477 5421 -23 5427
rect 79 5421 114 5427
rect -477 5413 -6 5421
rect -477 5365 -23 5413
rect -477 5035 -415 5365
rect -85 5035 -23 5365
rect -477 4987 -23 5035
rect -477 4979 -6 4987
rect 56 5413 114 5421
rect 73 5386 114 5413
rect 486 5421 521 5427
rect 623 5421 1077 5427
rect 1179 5421 1214 5427
rect 486 5413 544 5421
rect 486 5386 527 5413
rect 73 4987 114 5014
rect 56 4979 114 4987
rect -477 4973 -23 4979
rect 79 4973 114 4979
rect 486 4987 527 5014
rect 486 4979 544 4987
rect 606 5413 1094 5421
rect 623 5365 1077 5413
rect 623 5035 685 5365
rect 1015 5035 1077 5365
rect 623 4987 1077 5035
rect 606 4979 1094 4987
rect 1156 5413 1214 5421
rect 1173 5386 1214 5413
rect 1586 5421 1621 5427
rect 1723 5421 2177 5427
rect 2279 5421 2314 5427
rect 1586 5413 1644 5421
rect 1586 5386 1627 5413
rect 1173 4987 1214 5014
rect 1156 4979 1214 4987
rect 486 4973 521 4979
rect 623 4973 1077 4979
rect 1179 4973 1214 4979
rect 1586 4987 1627 5014
rect 1586 4979 1644 4987
rect 1706 5413 2194 5421
rect 1723 5365 2177 5413
rect 1723 5035 1785 5365
rect 2115 5035 2177 5365
rect 1723 4987 2177 5035
rect 1706 4979 2194 4987
rect 2256 5413 2314 5421
rect 2273 5386 2314 5413
rect 2686 5421 2721 5427
rect 2823 5421 3277 5427
rect 3379 5421 3414 5427
rect 2686 5413 2744 5421
rect 2686 5386 2727 5413
rect 2273 4987 2314 5014
rect 2256 4979 2314 4987
rect 1586 4973 1621 4979
rect 1723 4973 2177 4979
rect 2279 4973 2314 4979
rect 2686 4987 2727 5014
rect 2686 4979 2744 4987
rect 2806 5413 3294 5421
rect 2823 5365 3277 5413
rect 2823 5035 2885 5365
rect 3215 5035 3277 5365
rect 2823 4987 3277 5035
rect 2806 4979 3294 4987
rect 3356 5413 3414 5421
rect 3373 5386 3414 5413
rect 3786 5421 3821 5427
rect 3923 5421 4377 5427
rect 4479 5421 4514 5427
rect 3786 5413 3844 5421
rect 3786 5386 3827 5413
rect 3373 4987 3414 5014
rect 3356 4979 3414 4987
rect 2686 4973 2721 4979
rect 2823 4973 3277 4979
rect 3379 4973 3414 4979
rect 3786 4987 3827 5014
rect 3786 4979 3844 4987
rect 3906 5413 4394 5421
rect 3923 5365 4377 5413
rect 3923 5035 3985 5365
rect 4315 5035 4377 5365
rect 3923 4987 4377 5035
rect 3906 4979 4394 4987
rect 4456 5413 4514 5421
rect 4473 5386 4514 5413
rect 4886 5421 4921 5427
rect 5023 5421 5477 5427
rect 5579 5421 5614 5427
rect 4886 5413 4944 5421
rect 4886 5386 4927 5413
rect 4473 4987 4514 5014
rect 4456 4979 4514 4987
rect 3786 4973 3821 4979
rect 3923 4973 4377 4979
rect 4479 4973 4514 4979
rect 4886 4987 4927 5014
rect 4886 4979 4944 4987
rect 5006 5413 5494 5421
rect 5023 5365 5477 5413
rect 5023 5035 5085 5365
rect 5415 5035 5477 5365
rect 5023 4987 5477 5035
rect 5006 4979 5494 4987
rect 5556 5413 5614 5421
rect 5573 5386 5614 5413
rect 5986 5421 6021 5427
rect 6123 5421 6577 5427
rect 6679 5421 6714 5427
rect 5986 5413 6044 5421
rect 5986 5386 6027 5413
rect 5573 4987 5614 5014
rect 5556 4979 5614 4987
rect 4886 4973 4921 4979
rect 5023 4973 5477 4979
rect 5579 4973 5614 4979
rect 5986 4987 6027 5014
rect 5986 4979 6044 4987
rect 6106 5413 6594 5421
rect 6123 5365 6577 5413
rect 6123 5035 6185 5365
rect 6515 5035 6577 5365
rect 6123 4987 6577 5035
rect 6106 4979 6594 4987
rect 6656 5413 6714 5421
rect 6673 5386 6714 5413
rect 7086 5421 7121 5427
rect 7223 5421 7677 5427
rect 7779 5421 7814 5427
rect 7086 5413 7144 5421
rect 7086 5386 7127 5413
rect 6673 4987 6714 5014
rect 6656 4979 6714 4987
rect 5986 4973 6021 4979
rect 6123 4973 6577 4979
rect 6679 4973 6714 4979
rect 7086 4987 7127 5014
rect 7086 4979 7144 4987
rect 7206 5413 7694 5421
rect 7223 5365 7677 5413
rect 7223 5035 7285 5365
rect 7615 5035 7677 5365
rect 7223 4987 7677 5035
rect 7206 4979 7694 4987
rect 7756 5413 7814 5421
rect 7773 5386 7814 5413
rect 8186 5421 8221 5427
rect 8323 5421 8777 5427
rect 8879 5421 8914 5427
rect 8186 5413 8244 5421
rect 8186 5386 8227 5413
rect 7773 4987 7814 5014
rect 7756 4979 7814 4987
rect 7086 4973 7121 4979
rect 7223 4973 7677 4979
rect 7779 4973 7814 4979
rect 8186 4987 8227 5014
rect 8186 4979 8244 4987
rect 8306 5413 8794 5421
rect 8323 5365 8777 5413
rect 8323 5035 8385 5365
rect 8715 5035 8777 5365
rect 8323 4987 8777 5035
rect 8306 4979 8794 4987
rect 8856 5413 8914 5421
rect 8873 5386 8914 5413
rect 9286 5421 9321 5427
rect 9423 5421 9877 5427
rect 9979 5421 10014 5427
rect 9286 5413 9344 5421
rect 9286 5386 9327 5413
rect 8873 4987 8914 5014
rect 8856 4979 8914 4987
rect 8186 4973 8221 4979
rect 8323 4973 8777 4979
rect 8879 4973 8914 4979
rect 9286 4987 9327 5014
rect 9286 4979 9344 4987
rect 9406 5413 9894 5421
rect 9423 5365 9877 5413
rect 9423 5035 9485 5365
rect 9815 5035 9877 5365
rect 9423 4987 9877 5035
rect 9406 4979 9894 4987
rect 9956 5413 10014 5421
rect 9973 5386 10014 5413
rect 10386 5421 10421 5427
rect 10523 5421 10977 5427
rect 11079 5421 11114 5427
rect 10386 5413 10444 5421
rect 10386 5386 10427 5413
rect 9973 4987 10014 5014
rect 9956 4979 10014 4987
rect 9286 4973 9321 4979
rect 9423 4973 9877 4979
rect 9979 4973 10014 4979
rect 10386 4987 10427 5014
rect 10386 4979 10444 4987
rect 10506 5413 10994 5421
rect 10523 5365 10977 5413
rect 10523 5035 10585 5365
rect 10915 5035 10977 5365
rect 10523 4987 10977 5035
rect 10506 4979 10994 4987
rect 11056 5413 11114 5421
rect 11073 5386 11114 5413
rect 11486 5421 11521 5427
rect 11623 5421 12077 5427
rect 12179 5421 12214 5427
rect 11486 5413 11544 5421
rect 11486 5386 11527 5413
rect 11073 4987 11114 5014
rect 11056 4979 11114 4987
rect 10386 4973 10421 4979
rect 10523 4973 10977 4979
rect 11079 4973 11114 4979
rect 11486 4987 11527 5014
rect 11486 4979 11544 4987
rect 11606 5413 12094 5421
rect 11623 5365 12077 5413
rect 11623 5035 11685 5365
rect 12015 5035 12077 5365
rect 11623 4987 12077 5035
rect 11606 4979 12094 4987
rect 12156 5413 12214 5421
rect 12173 5386 12214 5413
rect 12586 5421 12621 5427
rect 12723 5421 13177 5427
rect 13279 5421 13314 5427
rect 12586 5413 12644 5421
rect 12586 5386 12627 5413
rect 12173 4987 12214 5014
rect 12156 4979 12214 4987
rect 11486 4973 11521 4979
rect 11623 4973 12077 4979
rect 12179 4973 12214 4979
rect 12586 4987 12627 5014
rect 12586 4979 12644 4987
rect 12706 5413 13194 5421
rect 12723 5365 13177 5413
rect 12723 5035 12785 5365
rect 13115 5035 13177 5365
rect 12723 4987 13177 5035
rect 12706 4979 13194 4987
rect 13256 5413 13314 5421
rect 13273 5386 13314 5413
rect 13273 4987 13314 5014
rect 13256 4979 13314 4987
rect 12586 4973 12621 4979
rect 12723 4973 13177 4979
rect 13279 4973 13314 4979
rect -1025 4950 -725 4967
rect -471 4956 -463 4973
rect -37 4956 -29 4973
rect 79 4956 87 4973
rect 513 4956 521 4973
rect 629 4956 637 4973
rect 1063 4956 1071 4973
rect 1179 4956 1187 4973
rect 1613 4956 1621 4973
rect 1729 4956 1737 4973
rect 2163 4956 2171 4973
rect 2279 4956 2287 4973
rect 2713 4956 2721 4973
rect 2829 4956 2837 4973
rect 3263 4956 3271 4973
rect 3379 4956 3387 4973
rect 3813 4956 3821 4973
rect 3929 4956 3937 4973
rect 4363 4956 4371 4973
rect 4479 4956 4487 4973
rect 4913 4956 4921 4973
rect 5029 4956 5037 4973
rect 5463 4956 5471 4973
rect 5579 4956 5587 4973
rect 6013 4956 6021 4973
rect 6129 4956 6137 4973
rect 6563 4956 6571 4973
rect 6679 4956 6687 4973
rect 7113 4956 7121 4973
rect 7229 4956 7237 4973
rect 7663 4956 7671 4973
rect 7779 4956 7787 4973
rect 8213 4956 8221 4973
rect 8329 4956 8337 4973
rect 8763 4956 8771 4973
rect 8879 4956 8887 4973
rect 9313 4956 9321 4973
rect 9429 4956 9437 4973
rect 9863 4956 9871 4973
rect 9979 4956 9987 4973
rect 10413 4956 10421 4973
rect 10529 4956 10537 4973
rect 10963 4956 10971 4973
rect 11079 4956 11087 4973
rect 11513 4956 11521 4973
rect 11629 4956 11637 4973
rect 12063 4956 12071 4973
rect 12179 4956 12187 4973
rect 12613 4956 12621 4973
rect 12729 4956 12737 4973
rect 13163 4956 13171 4973
rect 13279 4956 13287 4973
rect 13713 4956 13721 4973
rect 13975 4969 13987 5500
rect 14263 4969 14275 5500
rect 13975 4950 14275 4969
rect -1025 4417 -1013 4950
rect -737 4417 -725 4950
rect -550 4942 -500 4950
rect -550 4908 -542 4942
rect -508 4908 -500 4942
rect -550 4900 -500 4908
rect 0 4942 50 4950
rect 0 4908 8 4942
rect 42 4908 50 4942
rect 0 4900 50 4908
rect 550 4942 600 4950
rect 550 4908 558 4942
rect 592 4908 600 4942
rect 550 4900 600 4908
rect 1100 4942 1150 4950
rect 1100 4908 1108 4942
rect 1142 4908 1150 4942
rect 1100 4900 1150 4908
rect 1650 4942 1700 4950
rect 1650 4908 1658 4942
rect 1692 4908 1700 4942
rect 1650 4900 1700 4908
rect 2200 4942 2250 4950
rect 2200 4908 2208 4942
rect 2242 4908 2250 4942
rect 2200 4900 2250 4908
rect 2750 4942 2800 4950
rect 2750 4908 2758 4942
rect 2792 4908 2800 4942
rect 2750 4900 2800 4908
rect 3300 4942 3350 4950
rect 3300 4908 3308 4942
rect 3342 4908 3350 4942
rect 3300 4900 3350 4908
rect 3850 4942 3900 4950
rect 3850 4908 3858 4942
rect 3892 4908 3900 4942
rect 3850 4900 3900 4908
rect 4400 4942 4450 4950
rect 4400 4908 4408 4942
rect 4442 4908 4450 4942
rect 4400 4900 4450 4908
rect 4950 4942 5000 4950
rect 4950 4908 4958 4942
rect 4992 4908 5000 4942
rect 4950 4900 5000 4908
rect 5500 4942 5550 4950
rect 5500 4908 5508 4942
rect 5542 4908 5550 4942
rect 5500 4900 5550 4908
rect 6050 4942 6100 4950
rect 6050 4908 6058 4942
rect 6092 4908 6100 4942
rect 6050 4900 6100 4908
rect 6600 4942 6650 4950
rect 6600 4908 6608 4942
rect 6642 4908 6650 4942
rect 6600 4900 6650 4908
rect 7150 4942 7200 4950
rect 7150 4908 7158 4942
rect 7192 4908 7200 4942
rect 7150 4900 7200 4908
rect 7700 4942 7750 4950
rect 7700 4908 7708 4942
rect 7742 4908 7750 4942
rect 7700 4900 7750 4908
rect 8250 4942 8300 4950
rect 8250 4908 8258 4942
rect 8292 4908 8300 4942
rect 8250 4900 8300 4908
rect 8800 4942 8850 4950
rect 8800 4908 8808 4942
rect 8842 4908 8850 4942
rect 8800 4900 8850 4908
rect 9350 4942 9400 4950
rect 9350 4908 9358 4942
rect 9392 4908 9400 4942
rect 9350 4900 9400 4908
rect 9900 4942 9950 4950
rect 9900 4908 9908 4942
rect 9942 4908 9950 4942
rect 9900 4900 9950 4908
rect 10450 4942 10500 4950
rect 10450 4908 10458 4942
rect 10492 4908 10500 4942
rect 10450 4900 10500 4908
rect 11000 4942 11050 4950
rect 11000 4908 11008 4942
rect 11042 4908 11050 4942
rect 11000 4900 11050 4908
rect 11550 4942 11600 4950
rect 11550 4908 11558 4942
rect 11592 4908 11600 4942
rect 11550 4900 11600 4908
rect 12100 4942 12150 4950
rect 12100 4908 12108 4942
rect 12142 4908 12150 4942
rect 12100 4900 12150 4908
rect 12650 4942 12700 4950
rect 12650 4908 12658 4942
rect 12692 4908 12700 4942
rect 12650 4900 12700 4908
rect 13200 4942 13250 4950
rect 13200 4908 13208 4942
rect 13242 4908 13250 4942
rect 13200 4900 13250 4908
rect 13750 4942 13800 4950
rect 13750 4908 13758 4942
rect 13792 4908 13800 4942
rect 13750 4900 13800 4908
rect -471 4877 -463 4894
rect -37 4877 -29 4894
rect 79 4877 87 4894
rect 513 4877 521 4894
rect 629 4877 637 4894
rect 1063 4877 1071 4894
rect 1179 4877 1187 4894
rect 1613 4877 1621 4894
rect 1729 4877 1737 4894
rect 2163 4877 2171 4894
rect 2279 4877 2287 4894
rect 2713 4877 2721 4894
rect 2829 4877 2837 4894
rect 3263 4877 3271 4894
rect 3379 4877 3387 4894
rect 3813 4877 3821 4894
rect 3929 4877 3937 4894
rect 4363 4877 4371 4894
rect 4479 4877 4487 4894
rect 4913 4877 4921 4894
rect 5029 4877 5037 4894
rect 5463 4877 5471 4894
rect 5579 4877 5587 4894
rect 6013 4877 6021 4894
rect 6129 4877 6137 4894
rect 6563 4877 6571 4894
rect 6679 4877 6687 4894
rect 7113 4877 7121 4894
rect 7229 4877 7237 4894
rect 7663 4877 7671 4894
rect 7779 4877 7787 4894
rect 8213 4877 8221 4894
rect 8329 4877 8337 4894
rect 8763 4877 8771 4894
rect 8879 4877 8887 4894
rect 9313 4877 9321 4894
rect 9429 4877 9437 4894
rect 9863 4877 9871 4894
rect 9979 4877 9987 4894
rect 10413 4877 10421 4894
rect 10529 4877 10537 4894
rect 10963 4877 10971 4894
rect 11079 4877 11087 4894
rect 11513 4877 11521 4894
rect 11629 4877 11637 4894
rect 12063 4877 12071 4894
rect 12179 4877 12187 4894
rect 12613 4877 12621 4894
rect 12729 4877 12737 4894
rect 13163 4877 13171 4894
rect 13279 4877 13287 4894
rect 13713 4877 13721 4894
rect -64 4871 -29 4877
rect 73 4871 527 4877
rect 629 4871 664 4877
rect -64 4863 -6 4871
rect -64 4836 -23 4863
rect -64 4437 -23 4464
rect -64 4429 -6 4437
rect 56 4863 544 4871
rect 73 4815 527 4863
rect 73 4485 135 4815
rect 465 4485 527 4815
rect 73 4437 527 4485
rect 56 4429 544 4437
rect 606 4863 664 4871
rect 623 4836 664 4863
rect 1036 4871 1071 4877
rect 1173 4871 1627 4877
rect 1729 4871 1764 4877
rect 1036 4863 1094 4871
rect 1036 4836 1077 4863
rect 623 4437 664 4464
rect 606 4429 664 4437
rect -64 4423 -29 4429
rect 73 4423 527 4429
rect 629 4423 664 4429
rect 1036 4437 1077 4464
rect 1036 4429 1094 4437
rect 1156 4863 1644 4871
rect 1173 4815 1627 4863
rect 1173 4485 1235 4815
rect 1565 4485 1627 4815
rect 1173 4437 1627 4485
rect 1156 4429 1644 4437
rect 1706 4863 1764 4871
rect 1723 4836 1764 4863
rect 2136 4871 2171 4877
rect 2273 4871 2727 4877
rect 2829 4871 2864 4877
rect 2136 4863 2194 4871
rect 2136 4836 2177 4863
rect 1723 4437 1764 4464
rect 1706 4429 1764 4437
rect 1036 4423 1071 4429
rect 1173 4423 1627 4429
rect 1729 4423 1764 4429
rect 2136 4437 2177 4464
rect 2136 4429 2194 4437
rect 2256 4863 2744 4871
rect 2273 4815 2727 4863
rect 2273 4485 2335 4815
rect 2665 4485 2727 4815
rect 2273 4437 2727 4485
rect 2256 4429 2744 4437
rect 2806 4863 2864 4871
rect 2823 4836 2864 4863
rect 3236 4871 3271 4877
rect 3373 4871 3827 4877
rect 3929 4871 3964 4877
rect 3236 4863 3294 4871
rect 3236 4836 3277 4863
rect 2823 4437 2864 4464
rect 2806 4429 2864 4437
rect 2136 4423 2171 4429
rect 2273 4423 2727 4429
rect 2829 4423 2864 4429
rect 3236 4437 3277 4464
rect 3236 4429 3294 4437
rect 3356 4863 3844 4871
rect 3373 4815 3827 4863
rect 3373 4485 3435 4815
rect 3765 4485 3827 4815
rect 3373 4437 3827 4485
rect 3356 4429 3844 4437
rect 3906 4863 3964 4871
rect 3923 4836 3964 4863
rect 4336 4871 4371 4877
rect 4473 4871 4927 4877
rect 5029 4871 5064 4877
rect 4336 4863 4394 4871
rect 4336 4836 4377 4863
rect 3923 4437 3964 4464
rect 3906 4429 3964 4437
rect 3236 4423 3271 4429
rect 3373 4423 3827 4429
rect 3929 4423 3964 4429
rect 4336 4437 4377 4464
rect 4336 4429 4394 4437
rect 4456 4863 4944 4871
rect 4473 4815 4927 4863
rect 4473 4485 4535 4815
rect 4865 4485 4927 4815
rect 4473 4437 4927 4485
rect 4456 4429 4944 4437
rect 5006 4863 5064 4871
rect 5023 4836 5064 4863
rect 5436 4871 5471 4877
rect 5573 4871 6027 4877
rect 6129 4871 6164 4877
rect 5436 4863 5494 4871
rect 5436 4836 5477 4863
rect 5023 4437 5064 4464
rect 5006 4429 5064 4437
rect 4336 4423 4371 4429
rect 4473 4423 4927 4429
rect 5029 4423 5064 4429
rect 5436 4437 5477 4464
rect 5436 4429 5494 4437
rect 5556 4863 6044 4871
rect 5573 4815 6027 4863
rect 5573 4485 5635 4815
rect 5965 4485 6027 4815
rect 5573 4437 6027 4485
rect 5556 4429 6044 4437
rect 6106 4863 6164 4871
rect 6123 4836 6164 4863
rect 6536 4871 6571 4877
rect 6673 4871 7127 4877
rect 7229 4871 7264 4877
rect 6536 4863 6594 4871
rect 6536 4836 6577 4863
rect 6123 4437 6164 4464
rect 6106 4429 6164 4437
rect 5436 4423 5471 4429
rect 5573 4423 6027 4429
rect 6129 4423 6164 4429
rect 6536 4437 6577 4464
rect 6536 4429 6594 4437
rect 6656 4863 7144 4871
rect 6673 4815 7127 4863
rect 6673 4485 6735 4815
rect 7065 4485 7127 4815
rect 6673 4437 7127 4485
rect 6656 4429 7144 4437
rect 7206 4863 7264 4871
rect 7223 4836 7264 4863
rect 7636 4871 7671 4877
rect 7773 4871 8227 4877
rect 8329 4871 8364 4877
rect 7636 4863 7694 4871
rect 7636 4836 7677 4863
rect 7223 4437 7264 4464
rect 7206 4429 7264 4437
rect 6536 4423 6571 4429
rect 6673 4423 7127 4429
rect 7229 4423 7264 4429
rect 7636 4437 7677 4464
rect 7636 4429 7694 4437
rect 7756 4863 8244 4871
rect 7773 4815 8227 4863
rect 7773 4485 7835 4815
rect 8165 4485 8227 4815
rect 7773 4437 8227 4485
rect 7756 4429 8244 4437
rect 8306 4863 8364 4871
rect 8323 4836 8364 4863
rect 8736 4871 8771 4877
rect 8873 4871 9327 4877
rect 9429 4871 9464 4877
rect 8736 4863 8794 4871
rect 8736 4836 8777 4863
rect 8323 4437 8364 4464
rect 8306 4429 8364 4437
rect 7636 4423 7671 4429
rect 7773 4423 8227 4429
rect 8329 4423 8364 4429
rect 8736 4437 8777 4464
rect 8736 4429 8794 4437
rect 8856 4863 9344 4871
rect 8873 4815 9327 4863
rect 8873 4485 8935 4815
rect 9265 4485 9327 4815
rect 8873 4437 9327 4485
rect 8856 4429 9344 4437
rect 9406 4863 9464 4871
rect 9423 4836 9464 4863
rect 9836 4871 9871 4877
rect 9973 4871 10427 4877
rect 10529 4871 10564 4877
rect 9836 4863 9894 4871
rect 9836 4836 9877 4863
rect 9423 4437 9464 4464
rect 9406 4429 9464 4437
rect 8736 4423 8771 4429
rect 8873 4423 9327 4429
rect 9429 4423 9464 4429
rect 9836 4437 9877 4464
rect 9836 4429 9894 4437
rect 9956 4863 10444 4871
rect 9973 4815 10427 4863
rect 9973 4485 10035 4815
rect 10365 4485 10427 4815
rect 9973 4437 10427 4485
rect 9956 4429 10444 4437
rect 10506 4863 10564 4871
rect 10523 4836 10564 4863
rect 10936 4871 10971 4877
rect 11073 4871 11527 4877
rect 11629 4871 11664 4877
rect 10936 4863 10994 4871
rect 10936 4836 10977 4863
rect 10523 4437 10564 4464
rect 10506 4429 10564 4437
rect 9836 4423 9871 4429
rect 9973 4423 10427 4429
rect 10529 4423 10564 4429
rect 10936 4437 10977 4464
rect 10936 4429 10994 4437
rect 11056 4863 11544 4871
rect 11073 4815 11527 4863
rect 11073 4485 11135 4815
rect 11465 4485 11527 4815
rect 11073 4437 11527 4485
rect 11056 4429 11544 4437
rect 11606 4863 11664 4871
rect 11623 4836 11664 4863
rect 12036 4871 12071 4877
rect 12173 4871 12627 4877
rect 12729 4871 12764 4877
rect 12036 4863 12094 4871
rect 12036 4836 12077 4863
rect 11623 4437 11664 4464
rect 11606 4429 11664 4437
rect 10936 4423 10971 4429
rect 11073 4423 11527 4429
rect 11629 4423 11664 4429
rect 12036 4437 12077 4464
rect 12036 4429 12094 4437
rect 12156 4863 12644 4871
rect 12173 4815 12627 4863
rect 12173 4485 12235 4815
rect 12565 4485 12627 4815
rect 12173 4437 12627 4485
rect 12156 4429 12644 4437
rect 12706 4863 12764 4871
rect 12723 4836 12764 4863
rect 13136 4871 13171 4877
rect 13273 4871 13727 4877
rect 13136 4863 13194 4871
rect 13136 4836 13177 4863
rect 12723 4437 12764 4464
rect 12706 4429 12764 4437
rect 12036 4423 12071 4429
rect 12173 4423 12627 4429
rect 12729 4423 12764 4429
rect 13136 4437 13177 4464
rect 13136 4429 13194 4437
rect 13256 4863 13727 4871
rect 13273 4815 13727 4863
rect 13273 4485 13335 4815
rect 13665 4485 13727 4815
rect 13273 4437 13727 4485
rect 13256 4429 13727 4437
rect 13136 4423 13171 4429
rect 13273 4423 13727 4429
rect -1025 4400 -725 4417
rect -471 4406 -463 4423
rect -37 4406 -29 4423
rect 79 4406 87 4423
rect 513 4406 521 4423
rect 629 4406 637 4423
rect 1063 4406 1071 4423
rect 1179 4406 1187 4423
rect 1613 4406 1621 4423
rect 1729 4406 1737 4423
rect 2163 4406 2171 4423
rect 2279 4406 2287 4423
rect 2713 4406 2721 4423
rect 2829 4406 2837 4423
rect 3263 4406 3271 4423
rect 3379 4406 3387 4423
rect 3813 4406 3821 4423
rect 3929 4406 3937 4423
rect 4363 4406 4371 4423
rect 4479 4406 4487 4423
rect 4913 4406 4921 4423
rect 5029 4406 5037 4423
rect 5463 4406 5471 4423
rect 5579 4406 5587 4423
rect 6013 4406 6021 4423
rect 6129 4406 6137 4423
rect 6563 4406 6571 4423
rect 6679 4406 6687 4423
rect 7113 4406 7121 4423
rect 7229 4406 7237 4423
rect 7663 4406 7671 4423
rect 7779 4406 7787 4423
rect 8213 4406 8221 4423
rect 8329 4406 8337 4423
rect 8763 4406 8771 4423
rect 8879 4406 8887 4423
rect 9313 4406 9321 4423
rect 9429 4406 9437 4423
rect 9863 4406 9871 4423
rect 9979 4406 9987 4423
rect 10413 4406 10421 4423
rect 10529 4406 10537 4423
rect 10963 4406 10971 4423
rect 11079 4406 11087 4423
rect 11513 4406 11521 4423
rect 11629 4406 11637 4423
rect 12063 4406 12071 4423
rect 12179 4406 12187 4423
rect 12613 4406 12621 4423
rect 12729 4406 12737 4423
rect 13163 4406 13171 4423
rect 13279 4406 13287 4423
rect 13713 4406 13721 4423
rect 13975 4417 13987 4950
rect 14263 4417 14275 4950
rect 13975 4400 14275 4417
rect -1025 3867 -1013 4400
rect -737 3867 -725 4400
rect -550 4392 -500 4400
rect -550 4358 -542 4392
rect -508 4358 -500 4392
rect -550 4350 -500 4358
rect 0 4392 50 4400
rect 0 4358 8 4392
rect 42 4358 50 4392
rect 0 4350 50 4358
rect 550 4392 600 4400
rect 550 4358 558 4392
rect 592 4358 600 4392
rect 550 4350 600 4358
rect 1100 4392 1150 4400
rect 1100 4358 1108 4392
rect 1142 4358 1150 4392
rect 1100 4350 1150 4358
rect 1650 4392 1700 4400
rect 1650 4358 1658 4392
rect 1692 4358 1700 4392
rect 1650 4350 1700 4358
rect 2200 4392 2250 4400
rect 2200 4358 2208 4392
rect 2242 4358 2250 4392
rect 2200 4350 2250 4358
rect 2750 4392 2800 4400
rect 2750 4358 2758 4392
rect 2792 4358 2800 4392
rect 2750 4350 2800 4358
rect 3300 4392 3350 4400
rect 3300 4358 3308 4392
rect 3342 4358 3350 4392
rect 3300 4350 3350 4358
rect 3850 4392 3900 4400
rect 3850 4358 3858 4392
rect 3892 4358 3900 4392
rect 3850 4350 3900 4358
rect 4400 4392 4450 4400
rect 4400 4358 4408 4392
rect 4442 4358 4450 4392
rect 4400 4350 4450 4358
rect 4950 4392 5000 4400
rect 4950 4358 4958 4392
rect 4992 4358 5000 4392
rect 4950 4350 5000 4358
rect 5500 4392 5550 4400
rect 5500 4358 5508 4392
rect 5542 4358 5550 4392
rect 5500 4350 5550 4358
rect 6050 4392 6100 4400
rect 6050 4358 6058 4392
rect 6092 4358 6100 4392
rect 6050 4350 6100 4358
rect 6600 4392 6650 4400
rect 6600 4358 6608 4392
rect 6642 4358 6650 4392
rect 6600 4350 6650 4358
rect 7150 4392 7200 4400
rect 7150 4358 7158 4392
rect 7192 4358 7200 4392
rect 7150 4350 7200 4358
rect 7700 4392 7750 4400
rect 7700 4358 7708 4392
rect 7742 4358 7750 4392
rect 7700 4350 7750 4358
rect 8250 4392 8300 4400
rect 8250 4358 8258 4392
rect 8292 4358 8300 4392
rect 8250 4350 8300 4358
rect 8800 4392 8850 4400
rect 8800 4358 8808 4392
rect 8842 4358 8850 4392
rect 8800 4350 8850 4358
rect 9350 4392 9400 4400
rect 9350 4358 9358 4392
rect 9392 4358 9400 4392
rect 9350 4350 9400 4358
rect 9900 4392 9950 4400
rect 9900 4358 9908 4392
rect 9942 4358 9950 4392
rect 9900 4350 9950 4358
rect 10450 4392 10500 4400
rect 10450 4358 10458 4392
rect 10492 4358 10500 4392
rect 10450 4350 10500 4358
rect 11000 4392 11050 4400
rect 11000 4358 11008 4392
rect 11042 4358 11050 4392
rect 11000 4350 11050 4358
rect 11550 4392 11600 4400
rect 11550 4358 11558 4392
rect 11592 4358 11600 4392
rect 11550 4350 11600 4358
rect 12100 4392 12150 4400
rect 12100 4358 12108 4392
rect 12142 4358 12150 4392
rect 12100 4350 12150 4358
rect 12650 4392 12700 4400
rect 12650 4358 12658 4392
rect 12692 4358 12700 4392
rect 12650 4350 12700 4358
rect 13200 4392 13250 4400
rect 13200 4358 13208 4392
rect 13242 4358 13250 4392
rect 13200 4350 13250 4358
rect 13750 4392 13800 4400
rect 13750 4358 13758 4392
rect 13792 4358 13800 4392
rect 13750 4350 13800 4358
rect -471 4327 -463 4344
rect -37 4327 -29 4344
rect 79 4327 87 4344
rect 513 4327 521 4344
rect 629 4327 637 4344
rect 1063 4327 1071 4344
rect 1179 4327 1187 4344
rect 1613 4327 1621 4344
rect 1729 4327 1737 4344
rect 2163 4327 2171 4344
rect 2279 4327 2287 4344
rect 2713 4327 2721 4344
rect 2829 4327 2837 4344
rect 3263 4327 3271 4344
rect 3379 4327 3387 4344
rect 3813 4327 3821 4344
rect 3929 4327 3937 4344
rect 4363 4327 4371 4344
rect 4479 4327 4487 4344
rect 4913 4327 4921 4344
rect 5029 4327 5037 4344
rect 5463 4327 5471 4344
rect 5579 4327 5587 4344
rect 6013 4327 6021 4344
rect 6129 4327 6137 4344
rect 6563 4327 6571 4344
rect 6679 4327 6687 4344
rect 7113 4327 7121 4344
rect 7229 4327 7237 4344
rect 7663 4327 7671 4344
rect 7779 4327 7787 4344
rect 8213 4327 8221 4344
rect 8329 4327 8337 4344
rect 8763 4327 8771 4344
rect 8879 4327 8887 4344
rect 9313 4327 9321 4344
rect 9429 4327 9437 4344
rect 9863 4327 9871 4344
rect 9979 4327 9987 4344
rect 10413 4327 10421 4344
rect 10529 4327 10537 4344
rect 10963 4327 10971 4344
rect 11079 4327 11087 4344
rect 11513 4327 11521 4344
rect 11629 4327 11637 4344
rect 12063 4327 12071 4344
rect 12179 4327 12187 4344
rect 12613 4327 12621 4344
rect 12729 4327 12737 4344
rect 13163 4327 13171 4344
rect 13279 4327 13287 4344
rect 13713 4327 13721 4344
rect -477 4321 -23 4327
rect 79 4321 114 4327
rect -477 4313 -6 4321
rect -477 4265 -23 4313
rect -477 3935 -415 4265
rect -85 3935 -23 4265
rect -477 3887 -23 3935
rect -477 3879 -6 3887
rect 56 4313 114 4321
rect 73 4286 114 4313
rect 486 4321 521 4327
rect 623 4321 1077 4327
rect 1179 4321 1214 4327
rect 486 4313 544 4321
rect 486 4286 527 4313
rect 73 3887 114 3914
rect 56 3879 114 3887
rect -477 3873 -23 3879
rect 79 3873 114 3879
rect 486 3887 527 3914
rect 486 3879 544 3887
rect 606 4313 1094 4321
rect 623 4265 1077 4313
rect 623 3935 685 4265
rect 1015 3935 1077 4265
rect 623 3887 1077 3935
rect 606 3879 1094 3887
rect 1156 4313 1214 4321
rect 1173 4286 1214 4313
rect 1586 4321 1621 4327
rect 1723 4321 2177 4327
rect 2279 4321 2314 4327
rect 1586 4313 1644 4321
rect 1586 4286 1627 4313
rect 1173 3887 1214 3914
rect 1156 3879 1214 3887
rect 486 3873 521 3879
rect 623 3873 1077 3879
rect 1179 3873 1214 3879
rect 1586 3887 1627 3914
rect 1586 3879 1644 3887
rect 1706 4313 2194 4321
rect 1723 4265 2177 4313
rect 1723 3935 1785 4265
rect 2115 3935 2177 4265
rect 1723 3887 2177 3935
rect 1706 3879 2194 3887
rect 2256 4313 2314 4321
rect 2273 4286 2314 4313
rect 2686 4321 2721 4327
rect 2823 4321 3277 4327
rect 3379 4321 3414 4327
rect 2686 4313 2744 4321
rect 2686 4286 2727 4313
rect 2273 3887 2314 3914
rect 2256 3879 2314 3887
rect 1586 3873 1621 3879
rect 1723 3873 2177 3879
rect 2279 3873 2314 3879
rect 2686 3887 2727 3914
rect 2686 3879 2744 3887
rect 2806 4313 3294 4321
rect 2823 4265 3277 4313
rect 2823 3935 2885 4265
rect 3215 3935 3277 4265
rect 2823 3887 3277 3935
rect 2806 3879 3294 3887
rect 3356 4313 3414 4321
rect 3373 4286 3414 4313
rect 3786 4321 3821 4327
rect 3923 4321 4377 4327
rect 4479 4321 4514 4327
rect 3786 4313 3844 4321
rect 3786 4286 3827 4313
rect 3373 3887 3414 3914
rect 3356 3879 3414 3887
rect 2686 3873 2721 3879
rect 2823 3873 3277 3879
rect 3379 3873 3414 3879
rect 3786 3887 3827 3914
rect 3786 3879 3844 3887
rect 3906 4313 4394 4321
rect 3923 4265 4377 4313
rect 3923 3935 3985 4265
rect 4315 3935 4377 4265
rect 3923 3887 4377 3935
rect 3906 3879 4394 3887
rect 4456 4313 4514 4321
rect 4473 4286 4514 4313
rect 4886 4321 4921 4327
rect 5023 4321 5477 4327
rect 5579 4321 5614 4327
rect 4886 4313 4944 4321
rect 4886 4286 4927 4313
rect 4473 3887 4514 3914
rect 4456 3879 4514 3887
rect 3786 3873 3821 3879
rect 3923 3873 4377 3879
rect 4479 3873 4514 3879
rect 4886 3887 4927 3914
rect 4886 3879 4944 3887
rect 5006 4313 5494 4321
rect 5023 4265 5477 4313
rect 5023 3935 5085 4265
rect 5415 3935 5477 4265
rect 5023 3887 5477 3935
rect 5006 3879 5494 3887
rect 5556 4313 5614 4321
rect 5573 4286 5614 4313
rect 5986 4321 6021 4327
rect 6123 4321 6577 4327
rect 6679 4321 6714 4327
rect 5986 4313 6044 4321
rect 5986 4286 6027 4313
rect 5573 3887 5614 3914
rect 5556 3879 5614 3887
rect 4886 3873 4921 3879
rect 5023 3873 5477 3879
rect 5579 3873 5614 3879
rect 5986 3887 6027 3914
rect 5986 3879 6044 3887
rect 6106 4313 6594 4321
rect 6123 4265 6577 4313
rect 6123 3935 6185 4265
rect 6515 3935 6577 4265
rect 6123 3887 6577 3935
rect 6106 3879 6594 3887
rect 6656 4313 6714 4321
rect 6673 4286 6714 4313
rect 7086 4321 7121 4327
rect 7223 4321 7677 4327
rect 7779 4321 7814 4327
rect 7086 4313 7144 4321
rect 7086 4286 7127 4313
rect 6673 3887 6714 3914
rect 6656 3879 6714 3887
rect 5986 3873 6021 3879
rect 6123 3873 6577 3879
rect 6679 3873 6714 3879
rect 7086 3887 7127 3914
rect 7086 3879 7144 3887
rect 7206 4313 7694 4321
rect 7223 4265 7677 4313
rect 7223 3935 7285 4265
rect 7615 3935 7677 4265
rect 7223 3887 7677 3935
rect 7206 3879 7694 3887
rect 7756 4313 7814 4321
rect 7773 4286 7814 4313
rect 8186 4321 8221 4327
rect 8323 4321 8777 4327
rect 8879 4321 8914 4327
rect 8186 4313 8244 4321
rect 8186 4286 8227 4313
rect 7773 3887 7814 3914
rect 7756 3879 7814 3887
rect 7086 3873 7121 3879
rect 7223 3873 7677 3879
rect 7779 3873 7814 3879
rect 8186 3887 8227 3914
rect 8186 3879 8244 3887
rect 8306 4313 8794 4321
rect 8323 4265 8777 4313
rect 8323 3935 8385 4265
rect 8715 3935 8777 4265
rect 8323 3887 8777 3935
rect 8306 3879 8794 3887
rect 8856 4313 8914 4321
rect 8873 4286 8914 4313
rect 9286 4321 9321 4327
rect 9423 4321 9877 4327
rect 9979 4321 10014 4327
rect 9286 4313 9344 4321
rect 9286 4286 9327 4313
rect 8873 3887 8914 3914
rect 8856 3879 8914 3887
rect 8186 3873 8221 3879
rect 8323 3873 8777 3879
rect 8879 3873 8914 3879
rect 9286 3887 9327 3914
rect 9286 3879 9344 3887
rect 9406 4313 9894 4321
rect 9423 4265 9877 4313
rect 9423 3935 9485 4265
rect 9815 3935 9877 4265
rect 9423 3887 9877 3935
rect 9406 3879 9894 3887
rect 9956 4313 10014 4321
rect 9973 4286 10014 4313
rect 10386 4321 10421 4327
rect 10523 4321 10977 4327
rect 11079 4321 11114 4327
rect 10386 4313 10444 4321
rect 10386 4286 10427 4313
rect 9973 3887 10014 3914
rect 9956 3879 10014 3887
rect 9286 3873 9321 3879
rect 9423 3873 9877 3879
rect 9979 3873 10014 3879
rect 10386 3887 10427 3914
rect 10386 3879 10444 3887
rect 10506 4313 10994 4321
rect 10523 4265 10977 4313
rect 10523 3935 10585 4265
rect 10915 3935 10977 4265
rect 10523 3887 10977 3935
rect 10506 3879 10994 3887
rect 11056 4313 11114 4321
rect 11073 4286 11114 4313
rect 11486 4321 11521 4327
rect 11623 4321 12077 4327
rect 12179 4321 12214 4327
rect 11486 4313 11544 4321
rect 11486 4286 11527 4313
rect 11073 3887 11114 3914
rect 11056 3879 11114 3887
rect 10386 3873 10421 3879
rect 10523 3873 10977 3879
rect 11079 3873 11114 3879
rect 11486 3887 11527 3914
rect 11486 3879 11544 3887
rect 11606 4313 12094 4321
rect 11623 4265 12077 4313
rect 11623 3935 11685 4265
rect 12015 3935 12077 4265
rect 11623 3887 12077 3935
rect 11606 3879 12094 3887
rect 12156 4313 12214 4321
rect 12173 4286 12214 4313
rect 12586 4321 12621 4327
rect 12723 4321 13177 4327
rect 13279 4321 13314 4327
rect 12586 4313 12644 4321
rect 12586 4286 12627 4313
rect 12173 3887 12214 3914
rect 12156 3879 12214 3887
rect 11486 3873 11521 3879
rect 11623 3873 12077 3879
rect 12179 3873 12214 3879
rect 12586 3887 12627 3914
rect 12586 3879 12644 3887
rect 12706 4313 13194 4321
rect 12723 4265 13177 4313
rect 12723 3935 12785 4265
rect 13115 3935 13177 4265
rect 12723 3887 13177 3935
rect 12706 3879 13194 3887
rect 13256 4313 13314 4321
rect 13273 4286 13314 4313
rect 13273 3887 13314 3914
rect 13256 3879 13314 3887
rect 12586 3873 12621 3879
rect 12723 3873 13177 3879
rect 13279 3873 13314 3879
rect -1025 3850 -725 3867
rect -471 3856 -463 3873
rect -37 3856 -29 3873
rect 79 3856 87 3873
rect 513 3856 521 3873
rect 629 3856 637 3873
rect 1063 3856 1071 3873
rect 1179 3856 1187 3873
rect 1613 3856 1621 3873
rect 1729 3856 1737 3873
rect 2163 3856 2171 3873
rect 2279 3856 2287 3873
rect 2713 3856 2721 3873
rect 2829 3856 2837 3873
rect 3263 3856 3271 3873
rect 3379 3856 3387 3873
rect 3813 3856 3821 3873
rect 3929 3856 3937 3873
rect 4363 3856 4371 3873
rect 4479 3856 4487 3873
rect 4913 3856 4921 3873
rect 5029 3856 5037 3873
rect 5463 3856 5471 3873
rect 5579 3856 5587 3873
rect 6013 3856 6021 3873
rect 6129 3856 6137 3873
rect 6563 3856 6571 3873
rect 6679 3856 6687 3873
rect 7113 3856 7121 3873
rect 7229 3856 7237 3873
rect 7663 3856 7671 3873
rect 7779 3856 7787 3873
rect 8213 3856 8221 3873
rect 8329 3856 8337 3873
rect 8763 3856 8771 3873
rect 8879 3856 8887 3873
rect 9313 3856 9321 3873
rect 9429 3856 9437 3873
rect 9863 3856 9871 3873
rect 9979 3856 9987 3873
rect 10413 3856 10421 3873
rect 10529 3856 10537 3873
rect 10963 3856 10971 3873
rect 11079 3856 11087 3873
rect 11513 3856 11521 3873
rect 11629 3856 11637 3873
rect 12063 3856 12071 3873
rect 12179 3856 12187 3873
rect 12613 3856 12621 3873
rect 12729 3856 12737 3873
rect 13163 3856 13171 3873
rect 13279 3856 13287 3873
rect 13713 3856 13721 3873
rect 13975 3869 13987 4400
rect 14263 3869 14275 4400
rect 13975 3850 14275 3869
rect -1025 3317 -1013 3850
rect -737 3317 -725 3850
rect -550 3842 -500 3850
rect -550 3808 -542 3842
rect -508 3808 -500 3842
rect -550 3800 -500 3808
rect 0 3842 50 3850
rect 0 3808 8 3842
rect 42 3808 50 3842
rect 0 3800 50 3808
rect 550 3842 600 3850
rect 550 3808 558 3842
rect 592 3808 600 3842
rect 550 3800 600 3808
rect 1100 3842 1150 3850
rect 1100 3808 1108 3842
rect 1142 3808 1150 3842
rect 1100 3800 1150 3808
rect 1650 3842 1700 3850
rect 1650 3808 1658 3842
rect 1692 3808 1700 3842
rect 1650 3800 1700 3808
rect 2200 3842 2250 3850
rect 2200 3808 2208 3842
rect 2242 3808 2250 3842
rect 2200 3800 2250 3808
rect 2750 3842 2800 3850
rect 2750 3808 2758 3842
rect 2792 3808 2800 3842
rect 2750 3800 2800 3808
rect 3300 3842 3350 3850
rect 3300 3808 3308 3842
rect 3342 3808 3350 3842
rect 3300 3800 3350 3808
rect 3850 3842 3900 3850
rect 3850 3808 3858 3842
rect 3892 3808 3900 3842
rect 3850 3800 3900 3808
rect 4400 3842 4450 3850
rect 4400 3808 4408 3842
rect 4442 3808 4450 3842
rect 4400 3800 4450 3808
rect 4950 3842 5000 3850
rect 4950 3808 4958 3842
rect 4992 3808 5000 3842
rect 4950 3800 5000 3808
rect 5500 3842 5550 3850
rect 5500 3808 5508 3842
rect 5542 3808 5550 3842
rect 5500 3800 5550 3808
rect 6050 3842 6100 3850
rect 6050 3808 6058 3842
rect 6092 3808 6100 3842
rect 6050 3800 6100 3808
rect 6600 3842 6650 3850
rect 6600 3808 6608 3842
rect 6642 3808 6650 3842
rect 6600 3800 6650 3808
rect 7150 3842 7200 3850
rect 7150 3808 7158 3842
rect 7192 3808 7200 3842
rect 7150 3800 7200 3808
rect 7700 3842 7750 3850
rect 7700 3808 7708 3842
rect 7742 3808 7750 3842
rect 7700 3800 7750 3808
rect 8250 3842 8300 3850
rect 8250 3808 8258 3842
rect 8292 3808 8300 3842
rect 8250 3800 8300 3808
rect 8800 3842 8850 3850
rect 8800 3808 8808 3842
rect 8842 3808 8850 3842
rect 8800 3800 8850 3808
rect 9350 3842 9400 3850
rect 9350 3808 9358 3842
rect 9392 3808 9400 3842
rect 9350 3800 9400 3808
rect 9900 3842 9950 3850
rect 9900 3808 9908 3842
rect 9942 3808 9950 3842
rect 9900 3800 9950 3808
rect 10450 3842 10500 3850
rect 10450 3808 10458 3842
rect 10492 3808 10500 3842
rect 10450 3800 10500 3808
rect 11000 3842 11050 3850
rect 11000 3808 11008 3842
rect 11042 3808 11050 3842
rect 11000 3800 11050 3808
rect 11550 3842 11600 3850
rect 11550 3808 11558 3842
rect 11592 3808 11600 3842
rect 11550 3800 11600 3808
rect 12100 3842 12150 3850
rect 12100 3808 12108 3842
rect 12142 3808 12150 3842
rect 12100 3800 12150 3808
rect 12650 3842 12700 3850
rect 12650 3808 12658 3842
rect 12692 3808 12700 3842
rect 12650 3800 12700 3808
rect 13200 3842 13250 3850
rect 13200 3808 13208 3842
rect 13242 3808 13250 3842
rect 13200 3800 13250 3808
rect 13750 3842 13800 3850
rect 13750 3808 13758 3842
rect 13792 3808 13800 3842
rect 13750 3800 13800 3808
rect -471 3777 -463 3794
rect -37 3777 -29 3794
rect 79 3777 87 3794
rect 513 3777 521 3794
rect 629 3777 637 3794
rect 1063 3777 1071 3794
rect 1179 3777 1187 3794
rect 1613 3777 1621 3794
rect 1729 3777 1737 3794
rect 2163 3777 2171 3794
rect 2279 3777 2287 3794
rect 2713 3777 2721 3794
rect 2829 3777 2837 3794
rect 3263 3777 3271 3794
rect 3379 3777 3387 3794
rect 3813 3777 3821 3794
rect 3929 3777 3937 3794
rect 4363 3777 4371 3794
rect 4479 3777 4487 3794
rect 4913 3777 4921 3794
rect 5029 3777 5037 3794
rect 5463 3777 5471 3794
rect 5579 3777 5587 3794
rect 6013 3777 6021 3794
rect 6129 3777 6137 3794
rect 6563 3777 6571 3794
rect 6679 3777 6687 3794
rect 7113 3777 7121 3794
rect 7229 3777 7237 3794
rect 7663 3777 7671 3794
rect 7779 3777 7787 3794
rect 8213 3777 8221 3794
rect 8329 3777 8337 3794
rect 8763 3777 8771 3794
rect 8879 3777 8887 3794
rect 9313 3777 9321 3794
rect 9429 3777 9437 3794
rect 9863 3777 9871 3794
rect 9979 3777 9987 3794
rect 10413 3777 10421 3794
rect 10529 3777 10537 3794
rect 10963 3777 10971 3794
rect 11079 3777 11087 3794
rect 11513 3777 11521 3794
rect 11629 3777 11637 3794
rect 12063 3777 12071 3794
rect 12179 3777 12187 3794
rect 12613 3777 12621 3794
rect 12729 3777 12737 3794
rect 13163 3777 13171 3794
rect 13279 3777 13287 3794
rect 13713 3777 13721 3794
rect -64 3771 -29 3777
rect 73 3771 527 3777
rect 629 3771 664 3777
rect -64 3763 -6 3771
rect -64 3736 -23 3763
rect -64 3337 -23 3364
rect -64 3329 -6 3337
rect 56 3763 544 3771
rect 73 3715 527 3763
rect 73 3385 135 3715
rect 465 3385 527 3715
rect 73 3337 527 3385
rect 56 3329 544 3337
rect 606 3763 664 3771
rect 623 3736 664 3763
rect 1036 3771 1071 3777
rect 1173 3771 1627 3777
rect 1729 3771 1764 3777
rect 1036 3763 1094 3771
rect 1036 3736 1077 3763
rect 623 3337 664 3364
rect 606 3329 664 3337
rect -64 3323 -29 3329
rect 73 3323 527 3329
rect 629 3323 664 3329
rect 1036 3337 1077 3364
rect 1036 3329 1094 3337
rect 1156 3763 1644 3771
rect 1173 3715 1627 3763
rect 1173 3385 1235 3715
rect 1565 3385 1627 3715
rect 1173 3337 1627 3385
rect 1156 3329 1644 3337
rect 1706 3763 1764 3771
rect 1723 3736 1764 3763
rect 2136 3771 2171 3777
rect 2273 3771 2727 3777
rect 2829 3771 2864 3777
rect 2136 3763 2194 3771
rect 2136 3736 2177 3763
rect 1723 3337 1764 3364
rect 1706 3329 1764 3337
rect 1036 3323 1071 3329
rect 1173 3323 1627 3329
rect 1729 3323 1764 3329
rect 2136 3337 2177 3364
rect 2136 3329 2194 3337
rect 2256 3763 2744 3771
rect 2273 3715 2727 3763
rect 2273 3385 2335 3715
rect 2665 3385 2727 3715
rect 2273 3337 2727 3385
rect 2256 3329 2744 3337
rect 2806 3763 2864 3771
rect 2823 3736 2864 3763
rect 3236 3771 3271 3777
rect 3373 3771 3827 3777
rect 3929 3771 3964 3777
rect 3236 3763 3294 3771
rect 3236 3736 3277 3763
rect 2823 3337 2864 3364
rect 2806 3329 2864 3337
rect 2136 3323 2171 3329
rect 2273 3323 2727 3329
rect 2829 3323 2864 3329
rect 3236 3337 3277 3364
rect 3236 3329 3294 3337
rect 3356 3763 3844 3771
rect 3373 3715 3827 3763
rect 3373 3385 3435 3715
rect 3765 3385 3827 3715
rect 3373 3337 3827 3385
rect 3356 3329 3844 3337
rect 3906 3763 3964 3771
rect 3923 3736 3964 3763
rect 4336 3771 4371 3777
rect 4473 3771 4927 3777
rect 5029 3771 5064 3777
rect 4336 3763 4394 3771
rect 4336 3736 4377 3763
rect 3923 3337 3964 3364
rect 3906 3329 3964 3337
rect 3236 3323 3271 3329
rect 3373 3323 3827 3329
rect 3929 3323 3964 3329
rect 4336 3337 4377 3364
rect 4336 3329 4394 3337
rect 4456 3763 4944 3771
rect 4473 3715 4927 3763
rect 4473 3385 4535 3715
rect 4865 3385 4927 3715
rect 4473 3337 4927 3385
rect 4456 3329 4944 3337
rect 5006 3763 5064 3771
rect 5023 3736 5064 3763
rect 5436 3771 5471 3777
rect 5573 3771 6027 3777
rect 6129 3771 6164 3777
rect 5436 3763 5494 3771
rect 5436 3736 5477 3763
rect 5023 3337 5064 3364
rect 5006 3329 5064 3337
rect 4336 3323 4371 3329
rect 4473 3323 4927 3329
rect 5029 3323 5064 3329
rect 5436 3337 5477 3364
rect 5436 3329 5494 3337
rect 5556 3763 6044 3771
rect 5573 3715 6027 3763
rect 5573 3385 5635 3715
rect 5965 3385 6027 3715
rect 5573 3337 6027 3385
rect 5556 3329 6044 3337
rect 6106 3763 6164 3771
rect 6123 3736 6164 3763
rect 6536 3771 6571 3777
rect 6673 3771 7127 3777
rect 7229 3771 7264 3777
rect 6536 3763 6594 3771
rect 6536 3736 6577 3763
rect 6123 3337 6164 3364
rect 6106 3329 6164 3337
rect 5436 3323 5471 3329
rect 5573 3323 6027 3329
rect 6129 3323 6164 3329
rect 6536 3337 6577 3364
rect 6536 3329 6594 3337
rect 6656 3763 7144 3771
rect 6673 3715 7127 3763
rect 6673 3385 6735 3715
rect 7065 3385 7127 3715
rect 6673 3337 7127 3385
rect 6656 3329 7144 3337
rect 7206 3763 7264 3771
rect 7223 3736 7264 3763
rect 7636 3771 7671 3777
rect 7773 3771 8227 3777
rect 8329 3771 8364 3777
rect 7636 3763 7694 3771
rect 7636 3736 7677 3763
rect 7223 3337 7264 3364
rect 7206 3329 7264 3337
rect 6536 3323 6571 3329
rect 6673 3323 7127 3329
rect 7229 3323 7264 3329
rect 7636 3337 7677 3364
rect 7636 3329 7694 3337
rect 7756 3763 8244 3771
rect 7773 3715 8227 3763
rect 7773 3385 7835 3715
rect 8165 3385 8227 3715
rect 7773 3337 8227 3385
rect 7756 3329 8244 3337
rect 8306 3763 8364 3771
rect 8323 3736 8364 3763
rect 8736 3771 8771 3777
rect 8873 3771 9327 3777
rect 9429 3771 9464 3777
rect 8736 3763 8794 3771
rect 8736 3736 8777 3763
rect 8323 3337 8364 3364
rect 8306 3329 8364 3337
rect 7636 3323 7671 3329
rect 7773 3323 8227 3329
rect 8329 3323 8364 3329
rect 8736 3337 8777 3364
rect 8736 3329 8794 3337
rect 8856 3763 9344 3771
rect 8873 3715 9327 3763
rect 8873 3385 8935 3715
rect 9265 3385 9327 3715
rect 8873 3337 9327 3385
rect 8856 3329 9344 3337
rect 9406 3763 9464 3771
rect 9423 3736 9464 3763
rect 9836 3771 9871 3777
rect 9973 3771 10427 3777
rect 10529 3771 10564 3777
rect 9836 3763 9894 3771
rect 9836 3736 9877 3763
rect 9423 3337 9464 3364
rect 9406 3329 9464 3337
rect 8736 3323 8771 3329
rect 8873 3323 9327 3329
rect 9429 3323 9464 3329
rect 9836 3337 9877 3364
rect 9836 3329 9894 3337
rect 9956 3763 10444 3771
rect 9973 3715 10427 3763
rect 9973 3385 10035 3715
rect 10365 3385 10427 3715
rect 9973 3337 10427 3385
rect 9956 3329 10444 3337
rect 10506 3763 10564 3771
rect 10523 3736 10564 3763
rect 10936 3771 10971 3777
rect 11073 3771 11527 3777
rect 11629 3771 11664 3777
rect 10936 3763 10994 3771
rect 10936 3736 10977 3763
rect 10523 3337 10564 3364
rect 10506 3329 10564 3337
rect 9836 3323 9871 3329
rect 9973 3323 10427 3329
rect 10529 3323 10564 3329
rect 10936 3337 10977 3364
rect 10936 3329 10994 3337
rect 11056 3763 11544 3771
rect 11073 3715 11527 3763
rect 11073 3385 11135 3715
rect 11465 3385 11527 3715
rect 11073 3337 11527 3385
rect 11056 3329 11544 3337
rect 11606 3763 11664 3771
rect 11623 3736 11664 3763
rect 12036 3771 12071 3777
rect 12173 3771 12627 3777
rect 12729 3771 12764 3777
rect 12036 3763 12094 3771
rect 12036 3736 12077 3763
rect 11623 3337 11664 3364
rect 11606 3329 11664 3337
rect 10936 3323 10971 3329
rect 11073 3323 11527 3329
rect 11629 3323 11664 3329
rect 12036 3337 12077 3364
rect 12036 3329 12094 3337
rect 12156 3763 12644 3771
rect 12173 3715 12627 3763
rect 12173 3385 12235 3715
rect 12565 3385 12627 3715
rect 12173 3337 12627 3385
rect 12156 3329 12644 3337
rect 12706 3763 12764 3771
rect 12723 3736 12764 3763
rect 13136 3771 13171 3777
rect 13273 3771 13727 3777
rect 13136 3763 13194 3771
rect 13136 3736 13177 3763
rect 12723 3337 12764 3364
rect 12706 3329 12764 3337
rect 12036 3323 12071 3329
rect 12173 3323 12627 3329
rect 12729 3323 12764 3329
rect 13136 3337 13177 3364
rect 13136 3329 13194 3337
rect 13256 3763 13727 3771
rect 13273 3715 13727 3763
rect 13273 3385 13335 3715
rect 13665 3385 13727 3715
rect 13273 3337 13727 3385
rect 13256 3329 13727 3337
rect 13136 3323 13171 3329
rect 13273 3323 13727 3329
rect -1025 3300 -725 3317
rect -471 3306 -463 3323
rect -37 3306 -29 3323
rect 79 3306 87 3323
rect 513 3306 521 3323
rect 629 3306 637 3323
rect 1063 3306 1071 3323
rect 1179 3306 1187 3323
rect 1613 3306 1621 3323
rect 1729 3306 1737 3323
rect 2163 3306 2171 3323
rect 2279 3306 2287 3323
rect 2713 3306 2721 3323
rect 2829 3306 2837 3323
rect 3263 3306 3271 3323
rect 3379 3306 3387 3323
rect 3813 3306 3821 3323
rect 3929 3306 3937 3323
rect 4363 3306 4371 3323
rect 4479 3306 4487 3323
rect 4913 3306 4921 3323
rect 5029 3306 5037 3323
rect 5463 3306 5471 3323
rect 5579 3306 5587 3323
rect 6013 3306 6021 3323
rect 6129 3306 6137 3323
rect 6563 3306 6571 3323
rect 6679 3306 6687 3323
rect 7113 3306 7121 3323
rect 7229 3306 7237 3323
rect 7663 3306 7671 3323
rect 7779 3306 7787 3323
rect 8213 3306 8221 3323
rect 8329 3306 8337 3323
rect 8763 3306 8771 3323
rect 8879 3306 8887 3323
rect 9313 3306 9321 3323
rect 9429 3306 9437 3323
rect 9863 3306 9871 3323
rect 9979 3306 9987 3323
rect 10413 3306 10421 3323
rect 10529 3306 10537 3323
rect 10963 3306 10971 3323
rect 11079 3306 11087 3323
rect 11513 3306 11521 3323
rect 11629 3306 11637 3323
rect 12063 3306 12071 3323
rect 12179 3306 12187 3323
rect 12613 3306 12621 3323
rect 12729 3306 12737 3323
rect 13163 3306 13171 3323
rect 13279 3306 13287 3323
rect 13713 3306 13721 3323
rect 13975 3317 13987 3850
rect 14263 3317 14275 3850
rect 13975 3300 14275 3317
rect -1025 2767 -1013 3300
rect -737 2767 -725 3300
rect -550 3292 -500 3300
rect -550 3258 -542 3292
rect -508 3258 -500 3292
rect -550 3250 -500 3258
rect 0 3292 50 3300
rect 0 3258 8 3292
rect 42 3258 50 3292
rect 0 3250 50 3258
rect 550 3292 600 3300
rect 550 3258 558 3292
rect 592 3258 600 3292
rect 550 3250 600 3258
rect 1100 3292 1150 3300
rect 1100 3258 1108 3292
rect 1142 3258 1150 3292
rect 1100 3250 1150 3258
rect 1650 3292 1700 3300
rect 1650 3258 1658 3292
rect 1692 3258 1700 3292
rect 1650 3250 1700 3258
rect 2200 3292 2250 3300
rect 2200 3258 2208 3292
rect 2242 3258 2250 3292
rect 2200 3250 2250 3258
rect 2750 3292 2800 3300
rect 2750 3258 2758 3292
rect 2792 3258 2800 3292
rect 2750 3250 2800 3258
rect 3300 3292 3350 3300
rect 3300 3258 3308 3292
rect 3342 3258 3350 3292
rect 3300 3250 3350 3258
rect 3850 3292 3900 3300
rect 3850 3258 3858 3292
rect 3892 3258 3900 3292
rect 3850 3250 3900 3258
rect 4400 3292 4450 3300
rect 4400 3258 4408 3292
rect 4442 3258 4450 3292
rect 4400 3250 4450 3258
rect 4950 3292 5000 3300
rect 4950 3258 4958 3292
rect 4992 3258 5000 3292
rect 4950 3250 5000 3258
rect 5500 3292 5550 3300
rect 5500 3258 5508 3292
rect 5542 3258 5550 3292
rect 5500 3250 5550 3258
rect 6050 3292 6100 3300
rect 6050 3258 6058 3292
rect 6092 3258 6100 3292
rect 6050 3250 6100 3258
rect 6600 3292 6650 3300
rect 6600 3258 6608 3292
rect 6642 3258 6650 3292
rect 6600 3250 6650 3258
rect 7150 3292 7200 3300
rect 7150 3258 7158 3292
rect 7192 3258 7200 3292
rect 7150 3250 7200 3258
rect 7700 3292 7750 3300
rect 7700 3258 7708 3292
rect 7742 3258 7750 3292
rect 7700 3250 7750 3258
rect 8250 3292 8300 3300
rect 8250 3258 8258 3292
rect 8292 3258 8300 3292
rect 8250 3250 8300 3258
rect 8800 3292 8850 3300
rect 8800 3258 8808 3292
rect 8842 3258 8850 3292
rect 8800 3250 8850 3258
rect 9350 3292 9400 3300
rect 9350 3258 9358 3292
rect 9392 3258 9400 3292
rect 9350 3250 9400 3258
rect 9900 3292 9950 3300
rect 9900 3258 9908 3292
rect 9942 3258 9950 3292
rect 9900 3250 9950 3258
rect 10450 3292 10500 3300
rect 10450 3258 10458 3292
rect 10492 3258 10500 3292
rect 10450 3250 10500 3258
rect 11000 3292 11050 3300
rect 11000 3258 11008 3292
rect 11042 3258 11050 3292
rect 11000 3250 11050 3258
rect 11550 3292 11600 3300
rect 11550 3258 11558 3292
rect 11592 3258 11600 3292
rect 11550 3250 11600 3258
rect 12100 3292 12150 3300
rect 12100 3258 12108 3292
rect 12142 3258 12150 3292
rect 12100 3250 12150 3258
rect 12650 3292 12700 3300
rect 12650 3258 12658 3292
rect 12692 3258 12700 3292
rect 12650 3250 12700 3258
rect 13200 3292 13250 3300
rect 13200 3258 13208 3292
rect 13242 3258 13250 3292
rect 13200 3250 13250 3258
rect 13750 3292 13800 3300
rect 13750 3258 13758 3292
rect 13792 3258 13800 3292
rect 13750 3250 13800 3258
rect -471 3227 -463 3244
rect -37 3227 -29 3244
rect 79 3227 87 3244
rect 513 3227 521 3244
rect 629 3227 637 3244
rect 1063 3227 1071 3244
rect 1179 3227 1187 3244
rect 1613 3227 1621 3244
rect 1729 3227 1737 3244
rect 2163 3227 2171 3244
rect 2279 3227 2287 3244
rect 2713 3227 2721 3244
rect 2829 3227 2837 3244
rect 3263 3227 3271 3244
rect 3379 3227 3387 3244
rect 3813 3227 3821 3244
rect 3929 3227 3937 3244
rect 4363 3227 4371 3244
rect 4479 3227 4487 3244
rect 4913 3227 4921 3244
rect 5029 3227 5037 3244
rect 5463 3227 5471 3244
rect 5579 3227 5587 3244
rect 6013 3227 6021 3244
rect 6129 3227 6137 3244
rect 6563 3227 6571 3244
rect 6679 3227 6687 3244
rect 7113 3227 7121 3244
rect 7229 3227 7237 3244
rect 7663 3227 7671 3244
rect 7779 3227 7787 3244
rect 8213 3227 8221 3244
rect 8329 3227 8337 3244
rect 8763 3227 8771 3244
rect 8879 3227 8887 3244
rect 9313 3227 9321 3244
rect 9429 3227 9437 3244
rect 9863 3227 9871 3244
rect 9979 3227 9987 3244
rect 10413 3227 10421 3244
rect 10529 3227 10537 3244
rect 10963 3227 10971 3244
rect 11079 3227 11087 3244
rect 11513 3227 11521 3244
rect 11629 3227 11637 3244
rect 12063 3227 12071 3244
rect 12179 3227 12187 3244
rect 12613 3227 12621 3244
rect 12729 3227 12737 3244
rect 13163 3227 13171 3244
rect 13279 3227 13287 3244
rect 13713 3227 13721 3244
rect -477 3221 -23 3227
rect 79 3221 114 3227
rect -477 3213 -6 3221
rect -477 3165 -23 3213
rect -477 2835 -415 3165
rect -85 2835 -23 3165
rect -477 2787 -23 2835
rect -477 2779 -6 2787
rect 56 3213 114 3221
rect 73 3186 114 3213
rect 486 3221 521 3227
rect 623 3221 1077 3227
rect 1179 3221 1214 3227
rect 486 3213 544 3221
rect 486 3186 527 3213
rect 73 2787 114 2814
rect 56 2779 114 2787
rect -477 2773 -23 2779
rect 79 2773 114 2779
rect 486 2787 527 2814
rect 486 2779 544 2787
rect 606 3213 1094 3221
rect 623 3165 1077 3213
rect 623 2835 685 3165
rect 1015 2835 1077 3165
rect 623 2787 1077 2835
rect 606 2779 1094 2787
rect 1156 3213 1214 3221
rect 1173 3186 1214 3213
rect 1586 3221 1621 3227
rect 1723 3221 2177 3227
rect 2279 3221 2314 3227
rect 1586 3213 1644 3221
rect 1586 3186 1627 3213
rect 1173 2787 1214 2814
rect 1156 2779 1214 2787
rect 486 2773 521 2779
rect 623 2773 1077 2779
rect 1179 2773 1214 2779
rect 1586 2787 1627 2814
rect 1586 2779 1644 2787
rect 1706 3213 2194 3221
rect 1723 3165 2177 3213
rect 1723 2835 1785 3165
rect 2115 2835 2177 3165
rect 1723 2787 2177 2835
rect 1706 2779 2194 2787
rect 2256 3213 2314 3221
rect 2273 3186 2314 3213
rect 2686 3221 2721 3227
rect 2823 3221 3277 3227
rect 3379 3221 3414 3227
rect 2686 3213 2744 3221
rect 2686 3186 2727 3213
rect 2273 2787 2314 2814
rect 2256 2779 2314 2787
rect 1586 2773 1621 2779
rect 1723 2773 2177 2779
rect 2279 2773 2314 2779
rect 2686 2787 2727 2814
rect 2686 2779 2744 2787
rect 2806 3213 3294 3221
rect 2823 3165 3277 3213
rect 2823 2835 2885 3165
rect 3215 2835 3277 3165
rect 2823 2787 3277 2835
rect 2806 2779 3294 2787
rect 3356 3213 3414 3221
rect 3373 3186 3414 3213
rect 3786 3221 3821 3227
rect 3923 3221 4377 3227
rect 4479 3221 4514 3227
rect 3786 3213 3844 3221
rect 3786 3186 3827 3213
rect 3373 2787 3414 2814
rect 3356 2779 3414 2787
rect 2686 2773 2721 2779
rect 2823 2773 3277 2779
rect 3379 2773 3414 2779
rect 3786 2787 3827 2814
rect 3786 2779 3844 2787
rect 3906 3213 4394 3221
rect 3923 3165 4377 3213
rect 3923 2835 3985 3165
rect 4315 2835 4377 3165
rect 3923 2787 4377 2835
rect 3906 2779 4394 2787
rect 4456 3213 4514 3221
rect 4473 3186 4514 3213
rect 4886 3221 4921 3227
rect 5023 3221 5477 3227
rect 5579 3221 5614 3227
rect 4886 3213 4944 3221
rect 4886 3186 4927 3213
rect 4473 2787 4514 2814
rect 4456 2779 4514 2787
rect 3786 2773 3821 2779
rect 3923 2773 4377 2779
rect 4479 2773 4514 2779
rect 4886 2787 4927 2814
rect 4886 2779 4944 2787
rect 5006 3213 5494 3221
rect 5023 3165 5477 3213
rect 5023 2835 5085 3165
rect 5415 2835 5477 3165
rect 5023 2787 5477 2835
rect 5006 2779 5494 2787
rect 5556 3213 5614 3221
rect 5573 3186 5614 3213
rect 5986 3221 6021 3227
rect 6123 3221 6577 3227
rect 6679 3221 6714 3227
rect 5986 3213 6044 3221
rect 5986 3186 6027 3213
rect 5573 2787 5614 2814
rect 5556 2779 5614 2787
rect 4886 2773 4921 2779
rect 5023 2773 5477 2779
rect 5579 2773 5614 2779
rect 5986 2787 6027 2814
rect 5986 2779 6044 2787
rect 6106 3213 6594 3221
rect 6123 3165 6577 3213
rect 6123 2835 6185 3165
rect 6515 2835 6577 3165
rect 6123 2787 6577 2835
rect 6106 2779 6594 2787
rect 6656 3213 6714 3221
rect 6673 3186 6714 3213
rect 7086 3221 7121 3227
rect 7223 3221 7677 3227
rect 7779 3221 7814 3227
rect 7086 3213 7144 3221
rect 7086 3186 7127 3213
rect 6673 2787 6714 2814
rect 6656 2779 6714 2787
rect 5986 2773 6021 2779
rect 6123 2773 6577 2779
rect 6679 2773 6714 2779
rect 7086 2787 7127 2814
rect 7086 2779 7144 2787
rect 7206 3213 7694 3221
rect 7223 3165 7677 3213
rect 7223 2835 7285 3165
rect 7615 2835 7677 3165
rect 7223 2787 7677 2835
rect 7206 2779 7694 2787
rect 7756 3213 7814 3221
rect 7773 3186 7814 3213
rect 8186 3221 8221 3227
rect 8323 3221 8777 3227
rect 8879 3221 8914 3227
rect 8186 3213 8244 3221
rect 8186 3186 8227 3213
rect 7773 2787 7814 2814
rect 7756 2779 7814 2787
rect 7086 2773 7121 2779
rect 7223 2773 7677 2779
rect 7779 2773 7814 2779
rect 8186 2787 8227 2814
rect 8186 2779 8244 2787
rect 8306 3213 8794 3221
rect 8323 3165 8777 3213
rect 8323 2835 8385 3165
rect 8715 2835 8777 3165
rect 8323 2787 8777 2835
rect 8306 2779 8794 2787
rect 8856 3213 8914 3221
rect 8873 3186 8914 3213
rect 9286 3221 9321 3227
rect 9423 3221 9877 3227
rect 9979 3221 10014 3227
rect 9286 3213 9344 3221
rect 9286 3186 9327 3213
rect 8873 2787 8914 2814
rect 8856 2779 8914 2787
rect 8186 2773 8221 2779
rect 8323 2773 8777 2779
rect 8879 2773 8914 2779
rect 9286 2787 9327 2814
rect 9286 2779 9344 2787
rect 9406 3213 9894 3221
rect 9423 3165 9877 3213
rect 9423 2835 9485 3165
rect 9815 2835 9877 3165
rect 9423 2787 9877 2835
rect 9406 2779 9894 2787
rect 9956 3213 10014 3221
rect 9973 3186 10014 3213
rect 10386 3221 10421 3227
rect 10523 3221 10977 3227
rect 11079 3221 11114 3227
rect 10386 3213 10444 3221
rect 10386 3186 10427 3213
rect 9973 2787 10014 2814
rect 9956 2779 10014 2787
rect 9286 2773 9321 2779
rect 9423 2773 9877 2779
rect 9979 2773 10014 2779
rect 10386 2787 10427 2814
rect 10386 2779 10444 2787
rect 10506 3213 10994 3221
rect 10523 3165 10977 3213
rect 10523 2835 10585 3165
rect 10915 2835 10977 3165
rect 10523 2787 10977 2835
rect 10506 2779 10994 2787
rect 11056 3213 11114 3221
rect 11073 3186 11114 3213
rect 11486 3221 11521 3227
rect 11623 3221 12077 3227
rect 12179 3221 12214 3227
rect 11486 3213 11544 3221
rect 11486 3186 11527 3213
rect 11073 2787 11114 2814
rect 11056 2779 11114 2787
rect 10386 2773 10421 2779
rect 10523 2773 10977 2779
rect 11079 2773 11114 2779
rect 11486 2787 11527 2814
rect 11486 2779 11544 2787
rect 11606 3213 12094 3221
rect 11623 3165 12077 3213
rect 11623 2835 11685 3165
rect 12015 2835 12077 3165
rect 11623 2787 12077 2835
rect 11606 2779 12094 2787
rect 12156 3213 12214 3221
rect 12173 3186 12214 3213
rect 12586 3221 12621 3227
rect 12723 3221 13177 3227
rect 13279 3221 13314 3227
rect 12586 3213 12644 3221
rect 12586 3186 12627 3213
rect 12173 2787 12214 2814
rect 12156 2779 12214 2787
rect 11486 2773 11521 2779
rect 11623 2773 12077 2779
rect 12179 2773 12214 2779
rect 12586 2787 12627 2814
rect 12586 2779 12644 2787
rect 12706 3213 13194 3221
rect 12723 3165 13177 3213
rect 12723 2835 12785 3165
rect 13115 2835 13177 3165
rect 12723 2787 13177 2835
rect 12706 2779 13194 2787
rect 13256 3213 13314 3221
rect 13273 3186 13314 3213
rect 13273 2787 13314 2814
rect 13256 2779 13314 2787
rect 12586 2773 12621 2779
rect 12723 2773 13177 2779
rect 13279 2773 13314 2779
rect -1025 2750 -725 2767
rect -471 2756 -463 2773
rect -37 2756 -29 2773
rect 79 2756 87 2773
rect 513 2756 521 2773
rect 629 2756 637 2773
rect 1063 2756 1071 2773
rect 1179 2756 1187 2773
rect 1613 2756 1621 2773
rect 1729 2756 1737 2773
rect 2163 2756 2171 2773
rect 2279 2756 2287 2773
rect 2713 2756 2721 2773
rect 2829 2756 2837 2773
rect 3263 2756 3271 2773
rect 3379 2756 3387 2773
rect 3813 2756 3821 2773
rect 3929 2756 3937 2773
rect 4363 2756 4371 2773
rect 4479 2756 4487 2773
rect 4913 2756 4921 2773
rect 5029 2756 5037 2773
rect 5463 2756 5471 2773
rect 5579 2756 5587 2773
rect 6013 2756 6021 2773
rect 6129 2756 6137 2773
rect 6563 2756 6571 2773
rect 6679 2756 6687 2773
rect 7113 2756 7121 2773
rect 7229 2756 7237 2773
rect 7663 2756 7671 2773
rect 7779 2756 7787 2773
rect 8213 2756 8221 2773
rect 8329 2756 8337 2773
rect 8763 2756 8771 2773
rect 8879 2756 8887 2773
rect 9313 2756 9321 2773
rect 9429 2756 9437 2773
rect 9863 2756 9871 2773
rect 9979 2756 9987 2773
rect 10413 2756 10421 2773
rect 10529 2756 10537 2773
rect 10963 2756 10971 2773
rect 11079 2756 11087 2773
rect 11513 2756 11521 2773
rect 11629 2756 11637 2773
rect 12063 2756 12071 2773
rect 12179 2756 12187 2773
rect 12613 2756 12621 2773
rect 12729 2756 12737 2773
rect 13163 2756 13171 2773
rect 13279 2756 13287 2773
rect 13713 2756 13721 2773
rect 13975 2769 13987 3300
rect 14263 2769 14275 3300
rect 13975 2750 14275 2769
rect -1025 2217 -1013 2750
rect -737 2217 -725 2750
rect -550 2742 -500 2750
rect -550 2708 -542 2742
rect -508 2708 -500 2742
rect -550 2700 -500 2708
rect 0 2742 50 2750
rect 0 2708 8 2742
rect 42 2708 50 2742
rect 0 2700 50 2708
rect 550 2742 600 2750
rect 550 2708 558 2742
rect 592 2708 600 2742
rect 550 2700 600 2708
rect 1100 2742 1150 2750
rect 1100 2708 1108 2742
rect 1142 2708 1150 2742
rect 1100 2700 1150 2708
rect 1650 2742 1700 2750
rect 1650 2708 1658 2742
rect 1692 2708 1700 2742
rect 1650 2700 1700 2708
rect 2200 2742 2250 2750
rect 2200 2708 2208 2742
rect 2242 2708 2250 2742
rect 2200 2700 2250 2708
rect 2750 2742 2800 2750
rect 2750 2708 2758 2742
rect 2792 2708 2800 2742
rect 2750 2700 2800 2708
rect 3300 2742 3350 2750
rect 3300 2708 3308 2742
rect 3342 2708 3350 2742
rect 3300 2700 3350 2708
rect 3850 2742 3900 2750
rect 3850 2708 3858 2742
rect 3892 2708 3900 2742
rect 3850 2700 3900 2708
rect 4400 2742 4450 2750
rect 4400 2708 4408 2742
rect 4442 2708 4450 2742
rect 4400 2700 4450 2708
rect 4950 2742 5000 2750
rect 4950 2708 4958 2742
rect 4992 2708 5000 2742
rect 4950 2700 5000 2708
rect 5500 2742 5550 2750
rect 5500 2708 5508 2742
rect 5542 2708 5550 2742
rect 5500 2700 5550 2708
rect 6050 2742 6100 2750
rect 6050 2708 6058 2742
rect 6092 2708 6100 2742
rect 6050 2700 6100 2708
rect 6600 2742 6650 2750
rect 6600 2708 6608 2742
rect 6642 2708 6650 2742
rect 6600 2700 6650 2708
rect 7150 2742 7200 2750
rect 7150 2708 7158 2742
rect 7192 2708 7200 2742
rect 7150 2700 7200 2708
rect 7700 2742 7750 2750
rect 7700 2708 7708 2742
rect 7742 2708 7750 2742
rect 7700 2700 7750 2708
rect 8250 2742 8300 2750
rect 8250 2708 8258 2742
rect 8292 2708 8300 2742
rect 8250 2700 8300 2708
rect 8800 2742 8850 2750
rect 8800 2708 8808 2742
rect 8842 2708 8850 2742
rect 8800 2700 8850 2708
rect 9350 2742 9400 2750
rect 9350 2708 9358 2742
rect 9392 2708 9400 2742
rect 9350 2700 9400 2708
rect 9900 2742 9950 2750
rect 9900 2708 9908 2742
rect 9942 2708 9950 2742
rect 9900 2700 9950 2708
rect 10450 2742 10500 2750
rect 10450 2708 10458 2742
rect 10492 2708 10500 2742
rect 10450 2700 10500 2708
rect 11000 2742 11050 2750
rect 11000 2708 11008 2742
rect 11042 2708 11050 2742
rect 11000 2700 11050 2708
rect 11550 2742 11600 2750
rect 11550 2708 11558 2742
rect 11592 2708 11600 2742
rect 11550 2700 11600 2708
rect 12100 2742 12150 2750
rect 12100 2708 12108 2742
rect 12142 2708 12150 2742
rect 12100 2700 12150 2708
rect 12650 2742 12700 2750
rect 12650 2708 12658 2742
rect 12692 2708 12700 2742
rect 12650 2700 12700 2708
rect 13200 2742 13250 2750
rect 13200 2708 13208 2742
rect 13242 2708 13250 2742
rect 13200 2700 13250 2708
rect 13750 2742 13800 2750
rect 13750 2708 13758 2742
rect 13792 2708 13800 2742
rect 13750 2700 13800 2708
rect -471 2677 -463 2694
rect -37 2677 -29 2694
rect 79 2677 87 2694
rect 513 2677 521 2694
rect 629 2677 637 2694
rect 1063 2677 1071 2694
rect 1179 2677 1187 2694
rect 1613 2677 1621 2694
rect 1729 2677 1737 2694
rect 2163 2677 2171 2694
rect 2279 2677 2287 2694
rect 2713 2677 2721 2694
rect 2829 2677 2837 2694
rect 3263 2677 3271 2694
rect 3379 2677 3387 2694
rect 3813 2677 3821 2694
rect 3929 2677 3937 2694
rect 4363 2677 4371 2694
rect 4479 2677 4487 2694
rect 4913 2677 4921 2694
rect 5029 2677 5037 2694
rect 5463 2677 5471 2694
rect 5579 2677 5587 2694
rect 6013 2677 6021 2694
rect 6129 2677 6137 2694
rect 6563 2677 6571 2694
rect 6679 2677 6687 2694
rect 7113 2677 7121 2694
rect 7229 2677 7237 2694
rect 7663 2677 7671 2694
rect 7779 2677 7787 2694
rect 8213 2677 8221 2694
rect 8329 2677 8337 2694
rect 8763 2677 8771 2694
rect 8879 2677 8887 2694
rect 9313 2677 9321 2694
rect 9429 2677 9437 2694
rect 9863 2677 9871 2694
rect 9979 2677 9987 2694
rect 10413 2677 10421 2694
rect 10529 2677 10537 2694
rect 10963 2677 10971 2694
rect 11079 2677 11087 2694
rect 11513 2677 11521 2694
rect 11629 2677 11637 2694
rect 12063 2677 12071 2694
rect 12179 2677 12187 2694
rect 12613 2677 12621 2694
rect 12729 2677 12737 2694
rect 13163 2677 13171 2694
rect 13279 2677 13287 2694
rect 13713 2677 13721 2694
rect -64 2671 -29 2677
rect 73 2671 527 2677
rect 629 2671 664 2677
rect -64 2663 -6 2671
rect -64 2636 -23 2663
rect -64 2237 -23 2264
rect -64 2229 -6 2237
rect 56 2663 544 2671
rect 73 2615 527 2663
rect 73 2285 135 2615
rect 465 2285 527 2615
rect 73 2237 527 2285
rect 56 2229 544 2237
rect 606 2663 664 2671
rect 623 2636 664 2663
rect 1036 2671 1071 2677
rect 1173 2671 1627 2677
rect 1729 2671 1764 2677
rect 1036 2663 1094 2671
rect 1036 2636 1077 2663
rect 623 2237 664 2264
rect 606 2229 664 2237
rect -64 2223 -29 2229
rect 73 2223 527 2229
rect 629 2223 664 2229
rect 1036 2237 1077 2264
rect 1036 2229 1094 2237
rect 1156 2663 1644 2671
rect 1173 2615 1627 2663
rect 1173 2285 1235 2615
rect 1565 2285 1627 2615
rect 1173 2237 1627 2285
rect 1156 2229 1644 2237
rect 1706 2663 1764 2671
rect 1723 2636 1764 2663
rect 2136 2671 2171 2677
rect 2273 2671 2727 2677
rect 2829 2671 2864 2677
rect 2136 2663 2194 2671
rect 2136 2636 2177 2663
rect 1723 2237 1764 2264
rect 1706 2229 1764 2237
rect 1036 2223 1071 2229
rect 1173 2223 1627 2229
rect 1729 2223 1764 2229
rect 2136 2237 2177 2264
rect 2136 2229 2194 2237
rect 2256 2663 2744 2671
rect 2273 2615 2727 2663
rect 2273 2285 2335 2615
rect 2665 2285 2727 2615
rect 2273 2237 2727 2285
rect 2256 2229 2744 2237
rect 2806 2663 2864 2671
rect 2823 2636 2864 2663
rect 3236 2671 3271 2677
rect 3373 2671 3827 2677
rect 3929 2671 3964 2677
rect 3236 2663 3294 2671
rect 3236 2636 3277 2663
rect 2823 2237 2864 2264
rect 2806 2229 2864 2237
rect 2136 2223 2171 2229
rect 2273 2223 2727 2229
rect 2829 2223 2864 2229
rect 3236 2237 3277 2264
rect 3236 2229 3294 2237
rect 3356 2663 3844 2671
rect 3373 2615 3827 2663
rect 3373 2285 3435 2615
rect 3765 2285 3827 2615
rect 3373 2237 3827 2285
rect 3356 2229 3844 2237
rect 3906 2663 3964 2671
rect 3923 2636 3964 2663
rect 4336 2671 4371 2677
rect 4473 2671 4927 2677
rect 5029 2671 5064 2677
rect 4336 2663 4394 2671
rect 4336 2636 4377 2663
rect 3923 2237 3964 2264
rect 3906 2229 3964 2237
rect 3236 2223 3271 2229
rect 3373 2223 3827 2229
rect 3929 2223 3964 2229
rect 4336 2237 4377 2264
rect 4336 2229 4394 2237
rect 4456 2663 4944 2671
rect 4473 2615 4927 2663
rect 4473 2285 4535 2615
rect 4865 2285 4927 2615
rect 4473 2237 4927 2285
rect 4456 2229 4944 2237
rect 5006 2663 5064 2671
rect 5023 2636 5064 2663
rect 5436 2671 5471 2677
rect 5573 2671 6027 2677
rect 6129 2671 6164 2677
rect 5436 2663 5494 2671
rect 5436 2636 5477 2663
rect 5023 2237 5064 2264
rect 5006 2229 5064 2237
rect 4336 2223 4371 2229
rect 4473 2223 4927 2229
rect 5029 2223 5064 2229
rect 5436 2237 5477 2264
rect 5436 2229 5494 2237
rect 5556 2663 6044 2671
rect 5573 2615 6027 2663
rect 5573 2285 5635 2615
rect 5965 2285 6027 2615
rect 5573 2237 6027 2285
rect 5556 2229 6044 2237
rect 6106 2663 6164 2671
rect 6123 2636 6164 2663
rect 6536 2671 6571 2677
rect 6673 2671 7127 2677
rect 7229 2671 7264 2677
rect 6536 2663 6594 2671
rect 6536 2636 6577 2663
rect 6123 2237 6164 2264
rect 6106 2229 6164 2237
rect 5436 2223 5471 2229
rect 5573 2223 6027 2229
rect 6129 2223 6164 2229
rect 6536 2237 6577 2264
rect 6536 2229 6594 2237
rect 6656 2663 7144 2671
rect 6673 2615 7127 2663
rect 6673 2285 6735 2615
rect 7065 2285 7127 2615
rect 6673 2237 7127 2285
rect 6656 2229 7144 2237
rect 7206 2663 7264 2671
rect 7223 2636 7264 2663
rect 7636 2671 7671 2677
rect 7773 2671 8227 2677
rect 8329 2671 8364 2677
rect 7636 2663 7694 2671
rect 7636 2636 7677 2663
rect 7223 2237 7264 2264
rect 7206 2229 7264 2237
rect 6536 2223 6571 2229
rect 6673 2223 7127 2229
rect 7229 2223 7264 2229
rect 7636 2237 7677 2264
rect 7636 2229 7694 2237
rect 7756 2663 8244 2671
rect 7773 2615 8227 2663
rect 7773 2285 7835 2615
rect 8165 2285 8227 2615
rect 7773 2237 8227 2285
rect 7756 2229 8244 2237
rect 8306 2663 8364 2671
rect 8323 2636 8364 2663
rect 8736 2671 8771 2677
rect 8873 2671 9327 2677
rect 9429 2671 9464 2677
rect 8736 2663 8794 2671
rect 8736 2636 8777 2663
rect 8323 2237 8364 2264
rect 8306 2229 8364 2237
rect 7636 2223 7671 2229
rect 7773 2223 8227 2229
rect 8329 2223 8364 2229
rect 8736 2237 8777 2264
rect 8736 2229 8794 2237
rect 8856 2663 9344 2671
rect 8873 2615 9327 2663
rect 8873 2285 8935 2615
rect 9265 2285 9327 2615
rect 8873 2237 9327 2285
rect 8856 2229 9344 2237
rect 9406 2663 9464 2671
rect 9423 2636 9464 2663
rect 9836 2671 9871 2677
rect 9973 2671 10427 2677
rect 10529 2671 10564 2677
rect 9836 2663 9894 2671
rect 9836 2636 9877 2663
rect 9423 2237 9464 2264
rect 9406 2229 9464 2237
rect 8736 2223 8771 2229
rect 8873 2223 9327 2229
rect 9429 2223 9464 2229
rect 9836 2237 9877 2264
rect 9836 2229 9894 2237
rect 9956 2663 10444 2671
rect 9973 2615 10427 2663
rect 9973 2285 10035 2615
rect 10365 2285 10427 2615
rect 9973 2237 10427 2285
rect 9956 2229 10444 2237
rect 10506 2663 10564 2671
rect 10523 2636 10564 2663
rect 10936 2671 10971 2677
rect 11073 2671 11527 2677
rect 11629 2671 11664 2677
rect 10936 2663 10994 2671
rect 10936 2636 10977 2663
rect 10523 2237 10564 2264
rect 10506 2229 10564 2237
rect 9836 2223 9871 2229
rect 9973 2223 10427 2229
rect 10529 2223 10564 2229
rect 10936 2237 10977 2264
rect 10936 2229 10994 2237
rect 11056 2663 11544 2671
rect 11073 2615 11527 2663
rect 11073 2285 11135 2615
rect 11465 2285 11527 2615
rect 11073 2237 11527 2285
rect 11056 2229 11544 2237
rect 11606 2663 11664 2671
rect 11623 2636 11664 2663
rect 12036 2671 12071 2677
rect 12173 2671 12627 2677
rect 12729 2671 12764 2677
rect 12036 2663 12094 2671
rect 12036 2636 12077 2663
rect 11623 2237 11664 2264
rect 11606 2229 11664 2237
rect 10936 2223 10971 2229
rect 11073 2223 11527 2229
rect 11629 2223 11664 2229
rect 12036 2237 12077 2264
rect 12036 2229 12094 2237
rect 12156 2663 12644 2671
rect 12173 2615 12627 2663
rect 12173 2285 12235 2615
rect 12565 2285 12627 2615
rect 12173 2237 12627 2285
rect 12156 2229 12644 2237
rect 12706 2663 12764 2671
rect 12723 2636 12764 2663
rect 13136 2671 13171 2677
rect 13273 2671 13727 2677
rect 13136 2663 13194 2671
rect 13136 2636 13177 2663
rect 12723 2237 12764 2264
rect 12706 2229 12764 2237
rect 12036 2223 12071 2229
rect 12173 2223 12627 2229
rect 12729 2223 12764 2229
rect 13136 2237 13177 2264
rect 13136 2229 13194 2237
rect 13256 2663 13727 2671
rect 13273 2615 13727 2663
rect 13273 2285 13335 2615
rect 13665 2285 13727 2615
rect 13273 2237 13727 2285
rect 13256 2229 13727 2237
rect 13136 2223 13171 2229
rect 13273 2223 13727 2229
rect -1025 2200 -725 2217
rect -471 2206 -463 2223
rect -37 2206 -29 2223
rect 79 2206 87 2223
rect 513 2206 521 2223
rect 629 2206 637 2223
rect 1063 2206 1071 2223
rect 1179 2206 1187 2223
rect 1613 2206 1621 2223
rect 1729 2206 1737 2223
rect 2163 2206 2171 2223
rect 2279 2206 2287 2223
rect 2713 2206 2721 2223
rect 2829 2206 2837 2223
rect 3263 2206 3271 2223
rect 3379 2206 3387 2223
rect 3813 2206 3821 2223
rect 3929 2206 3937 2223
rect 4363 2206 4371 2223
rect 4479 2206 4487 2223
rect 4913 2206 4921 2223
rect 5029 2206 5037 2223
rect 5463 2206 5471 2223
rect 5579 2206 5587 2223
rect 6013 2206 6021 2223
rect 6129 2206 6137 2223
rect 6563 2206 6571 2223
rect 6679 2206 6687 2223
rect 7113 2206 7121 2223
rect 7229 2206 7237 2223
rect 7663 2206 7671 2223
rect 7779 2206 7787 2223
rect 8213 2206 8221 2223
rect 8329 2206 8337 2223
rect 8763 2206 8771 2223
rect 8879 2206 8887 2223
rect 9313 2206 9321 2223
rect 9429 2206 9437 2223
rect 9863 2206 9871 2223
rect 9979 2206 9987 2223
rect 10413 2206 10421 2223
rect 10529 2206 10537 2223
rect 10963 2206 10971 2223
rect 11079 2206 11087 2223
rect 11513 2206 11521 2223
rect 11629 2206 11637 2223
rect 12063 2206 12071 2223
rect 12179 2206 12187 2223
rect 12613 2206 12621 2223
rect 12729 2206 12737 2223
rect 13163 2206 13171 2223
rect 13279 2206 13287 2223
rect 13713 2206 13721 2223
rect 13975 2217 13987 2750
rect 14263 2217 14275 2750
rect 13975 2200 14275 2217
rect -1025 1667 -1013 2200
rect -737 1667 -725 2200
rect -550 2192 -500 2200
rect -550 2158 -542 2192
rect -508 2158 -500 2192
rect -550 2150 -500 2158
rect 0 2192 50 2200
rect 0 2158 8 2192
rect 42 2158 50 2192
rect 0 2150 50 2158
rect 550 2192 600 2200
rect 550 2158 558 2192
rect 592 2158 600 2192
rect 550 2150 600 2158
rect 1100 2192 1150 2200
rect 1100 2158 1108 2192
rect 1142 2158 1150 2192
rect 1100 2150 1150 2158
rect 1650 2192 1700 2200
rect 1650 2158 1658 2192
rect 1692 2158 1700 2192
rect 1650 2150 1700 2158
rect 2200 2192 2250 2200
rect 2200 2158 2208 2192
rect 2242 2158 2250 2192
rect 2200 2150 2250 2158
rect 2750 2192 2800 2200
rect 2750 2158 2758 2192
rect 2792 2158 2800 2192
rect 2750 2150 2800 2158
rect 3300 2192 3350 2200
rect 3300 2158 3308 2192
rect 3342 2158 3350 2192
rect 3300 2150 3350 2158
rect 3850 2192 3900 2200
rect 3850 2158 3858 2192
rect 3892 2158 3900 2192
rect 3850 2150 3900 2158
rect 4400 2192 4450 2200
rect 4400 2158 4408 2192
rect 4442 2158 4450 2192
rect 4400 2150 4450 2158
rect 4950 2192 5000 2200
rect 4950 2158 4958 2192
rect 4992 2158 5000 2192
rect 4950 2150 5000 2158
rect 5500 2192 5550 2200
rect 5500 2158 5508 2192
rect 5542 2158 5550 2192
rect 5500 2150 5550 2158
rect 6050 2192 6100 2200
rect 6050 2158 6058 2192
rect 6092 2158 6100 2192
rect 6050 2150 6100 2158
rect 6600 2192 6650 2200
rect 6600 2158 6608 2192
rect 6642 2158 6650 2192
rect 6600 2150 6650 2158
rect 7150 2192 7200 2200
rect 7150 2158 7158 2192
rect 7192 2158 7200 2192
rect 7150 2150 7200 2158
rect 7700 2192 7750 2200
rect 7700 2158 7708 2192
rect 7742 2158 7750 2192
rect 7700 2150 7750 2158
rect 8250 2192 8300 2200
rect 8250 2158 8258 2192
rect 8292 2158 8300 2192
rect 8250 2150 8300 2158
rect 8800 2192 8850 2200
rect 8800 2158 8808 2192
rect 8842 2158 8850 2192
rect 8800 2150 8850 2158
rect 9350 2192 9400 2200
rect 9350 2158 9358 2192
rect 9392 2158 9400 2192
rect 9350 2150 9400 2158
rect 9900 2192 9950 2200
rect 9900 2158 9908 2192
rect 9942 2158 9950 2192
rect 9900 2150 9950 2158
rect 10450 2192 10500 2200
rect 10450 2158 10458 2192
rect 10492 2158 10500 2192
rect 10450 2150 10500 2158
rect 11000 2192 11050 2200
rect 11000 2158 11008 2192
rect 11042 2158 11050 2192
rect 11000 2150 11050 2158
rect 11550 2192 11600 2200
rect 11550 2158 11558 2192
rect 11592 2158 11600 2192
rect 11550 2150 11600 2158
rect 12100 2192 12150 2200
rect 12100 2158 12108 2192
rect 12142 2158 12150 2192
rect 12100 2150 12150 2158
rect 12650 2192 12700 2200
rect 12650 2158 12658 2192
rect 12692 2158 12700 2192
rect 12650 2150 12700 2158
rect 13200 2192 13250 2200
rect 13200 2158 13208 2192
rect 13242 2158 13250 2192
rect 13200 2150 13250 2158
rect 13750 2192 13800 2200
rect 13750 2158 13758 2192
rect 13792 2158 13800 2192
rect 13750 2150 13800 2158
rect -471 2127 -463 2144
rect -37 2127 -29 2144
rect 79 2127 87 2144
rect 513 2127 521 2144
rect 629 2127 637 2144
rect 1063 2127 1071 2144
rect 1179 2127 1187 2144
rect 1613 2127 1621 2144
rect 1729 2127 1737 2144
rect 2163 2127 2171 2144
rect 2279 2127 2287 2144
rect 2713 2127 2721 2144
rect 2829 2127 2837 2144
rect 3263 2127 3271 2144
rect 3379 2127 3387 2144
rect 3813 2127 3821 2144
rect 3929 2127 3937 2144
rect 4363 2127 4371 2144
rect 4479 2127 4487 2144
rect 4913 2127 4921 2144
rect 5029 2127 5037 2144
rect 5463 2127 5471 2144
rect 5579 2127 5587 2144
rect 6013 2127 6021 2144
rect 6129 2127 6137 2144
rect 6563 2127 6571 2144
rect 6679 2127 6687 2144
rect 7113 2127 7121 2144
rect 7229 2127 7237 2144
rect 7663 2127 7671 2144
rect 7779 2127 7787 2144
rect 8213 2127 8221 2144
rect 8329 2127 8337 2144
rect 8763 2127 8771 2144
rect 8879 2127 8887 2144
rect 9313 2127 9321 2144
rect 9429 2127 9437 2144
rect 9863 2127 9871 2144
rect 9979 2127 9987 2144
rect 10413 2127 10421 2144
rect 10529 2127 10537 2144
rect 10963 2127 10971 2144
rect 11079 2127 11087 2144
rect 11513 2127 11521 2144
rect 11629 2127 11637 2144
rect 12063 2127 12071 2144
rect 12179 2127 12187 2144
rect 12613 2127 12621 2144
rect 12729 2127 12737 2144
rect 13163 2127 13171 2144
rect 13279 2127 13287 2144
rect 13713 2127 13721 2144
rect -477 2121 -23 2127
rect 79 2121 114 2127
rect -477 2113 -6 2121
rect -477 2065 -23 2113
rect -477 1735 -415 2065
rect -85 1735 -23 2065
rect -477 1687 -23 1735
rect -477 1679 -6 1687
rect 56 2113 114 2121
rect 73 2086 114 2113
rect 486 2121 521 2127
rect 623 2121 1077 2127
rect 1179 2121 1214 2127
rect 486 2113 544 2121
rect 486 2086 527 2113
rect 73 1687 114 1714
rect 56 1679 114 1687
rect -477 1673 -23 1679
rect 79 1673 114 1679
rect 486 1687 527 1714
rect 486 1679 544 1687
rect 606 2113 1094 2121
rect 623 2065 1077 2113
rect 623 1735 685 2065
rect 1015 1735 1077 2065
rect 623 1687 1077 1735
rect 606 1679 1094 1687
rect 1156 2113 1214 2121
rect 1173 2086 1214 2113
rect 1586 2121 1621 2127
rect 1723 2121 2177 2127
rect 2279 2121 2314 2127
rect 1586 2113 1644 2121
rect 1586 2086 1627 2113
rect 1173 1687 1214 1714
rect 1156 1679 1214 1687
rect 486 1673 521 1679
rect 623 1673 1077 1679
rect 1179 1673 1214 1679
rect 1586 1687 1627 1714
rect 1586 1679 1644 1687
rect 1706 2113 2194 2121
rect 1723 2065 2177 2113
rect 1723 1735 1785 2065
rect 2115 1735 2177 2065
rect 1723 1687 2177 1735
rect 1706 1679 2194 1687
rect 2256 2113 2314 2121
rect 2273 2086 2314 2113
rect 2686 2121 2721 2127
rect 2823 2121 3277 2127
rect 3379 2121 3414 2127
rect 2686 2113 2744 2121
rect 2686 2086 2727 2113
rect 2273 1687 2314 1714
rect 2256 1679 2314 1687
rect 1586 1673 1621 1679
rect 1723 1673 2177 1679
rect 2279 1673 2314 1679
rect 2686 1687 2727 1714
rect 2686 1679 2744 1687
rect 2806 2113 3294 2121
rect 2823 2065 3277 2113
rect 2823 1735 2885 2065
rect 3215 1735 3277 2065
rect 2823 1687 3277 1735
rect 2806 1679 3294 1687
rect 3356 2113 3414 2121
rect 3373 2086 3414 2113
rect 3786 2121 3821 2127
rect 3923 2121 4377 2127
rect 4479 2121 4514 2127
rect 3786 2113 3844 2121
rect 3786 2086 3827 2113
rect 3373 1687 3414 1714
rect 3356 1679 3414 1687
rect 2686 1673 2721 1679
rect 2823 1673 3277 1679
rect 3379 1673 3414 1679
rect 3786 1687 3827 1714
rect 3786 1679 3844 1687
rect 3906 2113 4394 2121
rect 3923 2065 4377 2113
rect 3923 1735 3985 2065
rect 4315 1735 4377 2065
rect 3923 1687 4377 1735
rect 3906 1679 4394 1687
rect 4456 2113 4514 2121
rect 4473 2086 4514 2113
rect 4886 2121 4921 2127
rect 5023 2121 5477 2127
rect 5579 2121 5614 2127
rect 4886 2113 4944 2121
rect 4886 2086 4927 2113
rect 4473 1687 4514 1714
rect 4456 1679 4514 1687
rect 3786 1673 3821 1679
rect 3923 1673 4377 1679
rect 4479 1673 4514 1679
rect 4886 1687 4927 1714
rect 4886 1679 4944 1687
rect 5006 2113 5494 2121
rect 5023 2065 5477 2113
rect 5023 1735 5085 2065
rect 5415 1735 5477 2065
rect 5023 1687 5477 1735
rect 5006 1679 5494 1687
rect 5556 2113 5614 2121
rect 5573 2086 5614 2113
rect 5986 2121 6021 2127
rect 6123 2121 6577 2127
rect 6679 2121 6714 2127
rect 5986 2113 6044 2121
rect 5986 2086 6027 2113
rect 5573 1687 5614 1714
rect 5556 1679 5614 1687
rect 4886 1673 4921 1679
rect 5023 1673 5477 1679
rect 5579 1673 5614 1679
rect 5986 1687 6027 1714
rect 5986 1679 6044 1687
rect 6106 2113 6594 2121
rect 6123 2065 6577 2113
rect 6123 1735 6185 2065
rect 6515 1735 6577 2065
rect 6123 1687 6577 1735
rect 6106 1679 6594 1687
rect 6656 2113 6714 2121
rect 6673 2086 6714 2113
rect 7086 2121 7121 2127
rect 7223 2121 7677 2127
rect 7779 2121 7814 2127
rect 7086 2113 7144 2121
rect 7086 2086 7127 2113
rect 6673 1687 6714 1714
rect 6656 1679 6714 1687
rect 5986 1673 6021 1679
rect 6123 1673 6577 1679
rect 6679 1673 6714 1679
rect 7086 1687 7127 1714
rect 7086 1679 7144 1687
rect 7206 2113 7694 2121
rect 7223 2065 7677 2113
rect 7223 1735 7285 2065
rect 7615 1735 7677 2065
rect 7223 1687 7677 1735
rect 7206 1679 7694 1687
rect 7756 2113 7814 2121
rect 7773 2086 7814 2113
rect 8186 2121 8221 2127
rect 8323 2121 8777 2127
rect 8879 2121 8914 2127
rect 8186 2113 8244 2121
rect 8186 2086 8227 2113
rect 7773 1687 7814 1714
rect 7756 1679 7814 1687
rect 7086 1673 7121 1679
rect 7223 1673 7677 1679
rect 7779 1673 7814 1679
rect 8186 1687 8227 1714
rect 8186 1679 8244 1687
rect 8306 2113 8794 2121
rect 8323 2065 8777 2113
rect 8323 1735 8385 2065
rect 8715 1735 8777 2065
rect 8323 1687 8777 1735
rect 8306 1679 8794 1687
rect 8856 2113 8914 2121
rect 8873 2086 8914 2113
rect 9286 2121 9321 2127
rect 9423 2121 9877 2127
rect 9979 2121 10014 2127
rect 9286 2113 9344 2121
rect 9286 2086 9327 2113
rect 8873 1687 8914 1714
rect 8856 1679 8914 1687
rect 8186 1673 8221 1679
rect 8323 1673 8777 1679
rect 8879 1673 8914 1679
rect 9286 1687 9327 1714
rect 9286 1679 9344 1687
rect 9406 2113 9894 2121
rect 9423 2065 9877 2113
rect 9423 1735 9485 2065
rect 9815 1735 9877 2065
rect 9423 1687 9877 1735
rect 9406 1679 9894 1687
rect 9956 2113 10014 2121
rect 9973 2086 10014 2113
rect 10386 2121 10421 2127
rect 10523 2121 10977 2127
rect 11079 2121 11114 2127
rect 10386 2113 10444 2121
rect 10386 2086 10427 2113
rect 9973 1687 10014 1714
rect 9956 1679 10014 1687
rect 9286 1673 9321 1679
rect 9423 1673 9877 1679
rect 9979 1673 10014 1679
rect 10386 1687 10427 1714
rect 10386 1679 10444 1687
rect 10506 2113 10994 2121
rect 10523 2065 10977 2113
rect 10523 1735 10585 2065
rect 10915 1735 10977 2065
rect 10523 1687 10977 1735
rect 10506 1679 10994 1687
rect 11056 2113 11114 2121
rect 11073 2086 11114 2113
rect 11486 2121 11521 2127
rect 11623 2121 12077 2127
rect 12179 2121 12214 2127
rect 11486 2113 11544 2121
rect 11486 2086 11527 2113
rect 11073 1687 11114 1714
rect 11056 1679 11114 1687
rect 10386 1673 10421 1679
rect 10523 1673 10977 1679
rect 11079 1673 11114 1679
rect 11486 1687 11527 1714
rect 11486 1679 11544 1687
rect 11606 2113 12094 2121
rect 11623 2065 12077 2113
rect 11623 1735 11685 2065
rect 12015 1735 12077 2065
rect 11623 1687 12077 1735
rect 11606 1679 12094 1687
rect 12156 2113 12214 2121
rect 12173 2086 12214 2113
rect 12586 2121 12621 2127
rect 12723 2121 13177 2127
rect 13279 2121 13314 2127
rect 12586 2113 12644 2121
rect 12586 2086 12627 2113
rect 12173 1687 12214 1714
rect 12156 1679 12214 1687
rect 11486 1673 11521 1679
rect 11623 1673 12077 1679
rect 12179 1673 12214 1679
rect 12586 1687 12627 1714
rect 12586 1679 12644 1687
rect 12706 2113 13194 2121
rect 12723 2065 13177 2113
rect 12723 1735 12785 2065
rect 13115 1735 13177 2065
rect 12723 1687 13177 1735
rect 12706 1679 13194 1687
rect 13256 2113 13314 2121
rect 13273 2086 13314 2113
rect 13273 1687 13314 1714
rect 13256 1679 13314 1687
rect 12586 1673 12621 1679
rect 12723 1673 13177 1679
rect 13279 1673 13314 1679
rect -1025 1650 -725 1667
rect -471 1656 -463 1673
rect -37 1656 -29 1673
rect 79 1656 87 1673
rect 513 1656 521 1673
rect 629 1656 637 1673
rect 1063 1656 1071 1673
rect 1179 1656 1187 1673
rect 1613 1656 1621 1673
rect 1729 1656 1737 1673
rect 2163 1656 2171 1673
rect 2279 1656 2287 1673
rect 2713 1656 2721 1673
rect 2829 1656 2837 1673
rect 3263 1656 3271 1673
rect 3379 1656 3387 1673
rect 3813 1656 3821 1673
rect 3929 1656 3937 1673
rect 4363 1656 4371 1673
rect 4479 1656 4487 1673
rect 4913 1656 4921 1673
rect 5029 1656 5037 1673
rect 5463 1656 5471 1673
rect 5579 1656 5587 1673
rect 6013 1656 6021 1673
rect 6129 1656 6137 1673
rect 6563 1656 6571 1673
rect 6679 1656 6687 1673
rect 7113 1656 7121 1673
rect 7229 1656 7237 1673
rect 7663 1656 7671 1673
rect 7779 1656 7787 1673
rect 8213 1656 8221 1673
rect 8329 1656 8337 1673
rect 8763 1656 8771 1673
rect 8879 1656 8887 1673
rect 9313 1656 9321 1673
rect 9429 1656 9437 1673
rect 9863 1656 9871 1673
rect 9979 1656 9987 1673
rect 10413 1656 10421 1673
rect 10529 1656 10537 1673
rect 10963 1656 10971 1673
rect 11079 1656 11087 1673
rect 11513 1656 11521 1673
rect 11629 1656 11637 1673
rect 12063 1656 12071 1673
rect 12179 1656 12187 1673
rect 12613 1656 12621 1673
rect 12729 1656 12737 1673
rect 13163 1656 13171 1673
rect 13279 1656 13287 1673
rect 13713 1656 13721 1673
rect 13975 1669 13987 2200
rect 14263 1669 14275 2200
rect 13975 1650 14275 1669
rect -1025 1117 -1013 1650
rect -737 1117 -725 1650
rect -550 1642 -500 1650
rect -550 1608 -542 1642
rect -508 1608 -500 1642
rect -550 1600 -500 1608
rect 0 1642 50 1650
rect 0 1608 8 1642
rect 42 1608 50 1642
rect 0 1600 50 1608
rect 550 1642 600 1650
rect 550 1608 558 1642
rect 592 1608 600 1642
rect 550 1600 600 1608
rect 1100 1642 1150 1650
rect 1100 1608 1108 1642
rect 1142 1608 1150 1642
rect 1100 1600 1150 1608
rect 1650 1642 1700 1650
rect 1650 1608 1658 1642
rect 1692 1608 1700 1642
rect 1650 1600 1700 1608
rect 2200 1642 2250 1650
rect 2200 1608 2208 1642
rect 2242 1608 2250 1642
rect 2200 1600 2250 1608
rect 2750 1642 2800 1650
rect 2750 1608 2758 1642
rect 2792 1608 2800 1642
rect 2750 1600 2800 1608
rect 3300 1642 3350 1650
rect 3300 1608 3308 1642
rect 3342 1608 3350 1642
rect 3300 1600 3350 1608
rect 3850 1642 3900 1650
rect 3850 1608 3858 1642
rect 3892 1608 3900 1642
rect 3850 1600 3900 1608
rect 4400 1642 4450 1650
rect 4400 1608 4408 1642
rect 4442 1608 4450 1642
rect 4400 1600 4450 1608
rect 4950 1642 5000 1650
rect 4950 1608 4958 1642
rect 4992 1608 5000 1642
rect 4950 1600 5000 1608
rect 5500 1642 5550 1650
rect 5500 1608 5508 1642
rect 5542 1608 5550 1642
rect 5500 1600 5550 1608
rect 6050 1642 6100 1650
rect 6050 1608 6058 1642
rect 6092 1608 6100 1642
rect 6050 1600 6100 1608
rect 6600 1642 6650 1650
rect 6600 1608 6608 1642
rect 6642 1608 6650 1642
rect 6600 1600 6650 1608
rect 7150 1642 7200 1650
rect 7150 1608 7158 1642
rect 7192 1608 7200 1642
rect 7150 1600 7200 1608
rect 7700 1642 7750 1650
rect 7700 1608 7708 1642
rect 7742 1608 7750 1642
rect 7700 1600 7750 1608
rect 8250 1642 8300 1650
rect 8250 1608 8258 1642
rect 8292 1608 8300 1642
rect 8250 1600 8300 1608
rect 8800 1642 8850 1650
rect 8800 1608 8808 1642
rect 8842 1608 8850 1642
rect 8800 1600 8850 1608
rect 9350 1642 9400 1650
rect 9350 1608 9358 1642
rect 9392 1608 9400 1642
rect 9350 1600 9400 1608
rect 9900 1642 9950 1650
rect 9900 1608 9908 1642
rect 9942 1608 9950 1642
rect 9900 1600 9950 1608
rect 10450 1642 10500 1650
rect 10450 1608 10458 1642
rect 10492 1608 10500 1642
rect 10450 1600 10500 1608
rect 11000 1642 11050 1650
rect 11000 1608 11008 1642
rect 11042 1608 11050 1642
rect 11000 1600 11050 1608
rect 11550 1642 11600 1650
rect 11550 1608 11558 1642
rect 11592 1608 11600 1642
rect 11550 1600 11600 1608
rect 12100 1642 12150 1650
rect 12100 1608 12108 1642
rect 12142 1608 12150 1642
rect 12100 1600 12150 1608
rect 12650 1642 12700 1650
rect 12650 1608 12658 1642
rect 12692 1608 12700 1642
rect 12650 1600 12700 1608
rect 13200 1642 13250 1650
rect 13200 1608 13208 1642
rect 13242 1608 13250 1642
rect 13200 1600 13250 1608
rect 13750 1642 13800 1650
rect 13750 1608 13758 1642
rect 13792 1608 13800 1642
rect 13750 1600 13800 1608
rect -471 1577 -463 1594
rect -37 1577 -29 1594
rect 79 1577 87 1594
rect 513 1577 521 1594
rect 629 1577 637 1594
rect 1063 1577 1071 1594
rect 1179 1577 1187 1594
rect 1613 1577 1621 1594
rect 1729 1577 1737 1594
rect 2163 1577 2171 1594
rect 2279 1577 2287 1594
rect 2713 1577 2721 1594
rect 2829 1577 2837 1594
rect 3263 1577 3271 1594
rect 3379 1577 3387 1594
rect 3813 1577 3821 1594
rect 3929 1577 3937 1594
rect 4363 1577 4371 1594
rect 4479 1577 4487 1594
rect 4913 1577 4921 1594
rect 5029 1577 5037 1594
rect 5463 1577 5471 1594
rect 5579 1577 5587 1594
rect 6013 1577 6021 1594
rect 6129 1577 6137 1594
rect 6563 1577 6571 1594
rect 6679 1577 6687 1594
rect 7113 1577 7121 1594
rect 7229 1577 7237 1594
rect 7663 1577 7671 1594
rect 7779 1577 7787 1594
rect 8213 1577 8221 1594
rect 8329 1577 8337 1594
rect 8763 1577 8771 1594
rect 8879 1577 8887 1594
rect 9313 1577 9321 1594
rect 9429 1577 9437 1594
rect 9863 1577 9871 1594
rect 9979 1577 9987 1594
rect 10413 1577 10421 1594
rect 10529 1577 10537 1594
rect 10963 1577 10971 1594
rect 11079 1577 11087 1594
rect 11513 1577 11521 1594
rect 11629 1577 11637 1594
rect 12063 1577 12071 1594
rect 12179 1577 12187 1594
rect 12613 1577 12621 1594
rect 12729 1577 12737 1594
rect 13163 1577 13171 1594
rect 13279 1577 13287 1594
rect 13713 1577 13721 1594
rect -64 1571 -29 1577
rect 73 1571 527 1577
rect 629 1571 664 1577
rect -64 1563 -6 1571
rect -64 1536 -23 1563
rect -64 1137 -23 1164
rect -64 1129 -6 1137
rect 56 1563 544 1571
rect 73 1515 527 1563
rect 73 1185 135 1515
rect 465 1185 527 1515
rect 73 1137 527 1185
rect 56 1129 544 1137
rect 606 1563 664 1571
rect 623 1536 664 1563
rect 1036 1571 1071 1577
rect 1173 1571 1627 1577
rect 1729 1571 1764 1577
rect 1036 1563 1094 1571
rect 1036 1536 1077 1563
rect 623 1137 664 1164
rect 606 1129 664 1137
rect -64 1123 -29 1129
rect 73 1123 527 1129
rect 629 1123 664 1129
rect 1036 1137 1077 1164
rect 1036 1129 1094 1137
rect 1156 1563 1644 1571
rect 1173 1515 1627 1563
rect 1173 1185 1235 1515
rect 1565 1185 1627 1515
rect 1173 1137 1627 1185
rect 1156 1129 1644 1137
rect 1706 1563 1764 1571
rect 1723 1536 1764 1563
rect 2136 1571 2171 1577
rect 2273 1571 2727 1577
rect 2829 1571 2864 1577
rect 2136 1563 2194 1571
rect 2136 1536 2177 1563
rect 1723 1137 1764 1164
rect 1706 1129 1764 1137
rect 1036 1123 1071 1129
rect 1173 1123 1627 1129
rect 1729 1123 1764 1129
rect 2136 1137 2177 1164
rect 2136 1129 2194 1137
rect 2256 1563 2744 1571
rect 2273 1515 2727 1563
rect 2273 1185 2335 1515
rect 2665 1185 2727 1515
rect 2273 1137 2727 1185
rect 2256 1129 2744 1137
rect 2806 1563 2864 1571
rect 2823 1536 2864 1563
rect 3236 1571 3271 1577
rect 3373 1571 3827 1577
rect 3929 1571 3964 1577
rect 3236 1563 3294 1571
rect 3236 1536 3277 1563
rect 2823 1137 2864 1164
rect 2806 1129 2864 1137
rect 2136 1123 2171 1129
rect 2273 1123 2727 1129
rect 2829 1123 2864 1129
rect 3236 1137 3277 1164
rect 3236 1129 3294 1137
rect 3356 1563 3844 1571
rect 3373 1515 3827 1563
rect 3373 1185 3435 1515
rect 3765 1185 3827 1515
rect 3373 1137 3827 1185
rect 3356 1129 3844 1137
rect 3906 1563 3964 1571
rect 3923 1536 3964 1563
rect 4336 1571 4371 1577
rect 4473 1571 4927 1577
rect 5029 1571 5064 1577
rect 4336 1563 4394 1571
rect 4336 1536 4377 1563
rect 3923 1137 3964 1164
rect 3906 1129 3964 1137
rect 3236 1123 3271 1129
rect 3373 1123 3827 1129
rect 3929 1123 3964 1129
rect 4336 1137 4377 1164
rect 4336 1129 4394 1137
rect 4456 1563 4944 1571
rect 4473 1515 4927 1563
rect 4473 1185 4535 1515
rect 4865 1185 4927 1515
rect 4473 1137 4927 1185
rect 4456 1129 4944 1137
rect 5006 1563 5064 1571
rect 5023 1536 5064 1563
rect 5436 1571 5471 1577
rect 5573 1571 6027 1577
rect 6129 1571 6164 1577
rect 5436 1563 5494 1571
rect 5436 1536 5477 1563
rect 5023 1137 5064 1164
rect 5006 1129 5064 1137
rect 4336 1123 4371 1129
rect 4473 1123 4927 1129
rect 5029 1123 5064 1129
rect 5436 1137 5477 1164
rect 5436 1129 5494 1137
rect 5556 1563 6044 1571
rect 5573 1515 6027 1563
rect 5573 1185 5635 1515
rect 5965 1185 6027 1515
rect 5573 1137 6027 1185
rect 5556 1129 6044 1137
rect 6106 1563 6164 1571
rect 6123 1536 6164 1563
rect 6536 1571 6571 1577
rect 6673 1571 7127 1577
rect 7229 1571 7264 1577
rect 6536 1563 6594 1571
rect 6536 1536 6577 1563
rect 6123 1137 6164 1164
rect 6106 1129 6164 1137
rect 5436 1123 5471 1129
rect 5573 1123 6027 1129
rect 6129 1123 6164 1129
rect 6536 1137 6577 1164
rect 6536 1129 6594 1137
rect 6656 1563 7144 1571
rect 6673 1515 7127 1563
rect 6673 1185 6735 1515
rect 7065 1185 7127 1515
rect 6673 1137 7127 1185
rect 6656 1129 7144 1137
rect 7206 1563 7264 1571
rect 7223 1536 7264 1563
rect 7636 1571 7671 1577
rect 7773 1571 8227 1577
rect 8329 1571 8364 1577
rect 7636 1563 7694 1571
rect 7636 1536 7677 1563
rect 7223 1137 7264 1164
rect 7206 1129 7264 1137
rect 6536 1123 6571 1129
rect 6673 1123 7127 1129
rect 7229 1123 7264 1129
rect 7636 1137 7677 1164
rect 7636 1129 7694 1137
rect 7756 1563 8244 1571
rect 7773 1515 8227 1563
rect 7773 1185 7835 1515
rect 8165 1185 8227 1515
rect 7773 1137 8227 1185
rect 7756 1129 8244 1137
rect 8306 1563 8364 1571
rect 8323 1536 8364 1563
rect 8736 1571 8771 1577
rect 8873 1571 9327 1577
rect 9429 1571 9464 1577
rect 8736 1563 8794 1571
rect 8736 1536 8777 1563
rect 8323 1137 8364 1164
rect 8306 1129 8364 1137
rect 7636 1123 7671 1129
rect 7773 1123 8227 1129
rect 8329 1123 8364 1129
rect 8736 1137 8777 1164
rect 8736 1129 8794 1137
rect 8856 1563 9344 1571
rect 8873 1515 9327 1563
rect 8873 1185 8935 1515
rect 9265 1185 9327 1515
rect 8873 1137 9327 1185
rect 8856 1129 9344 1137
rect 9406 1563 9464 1571
rect 9423 1536 9464 1563
rect 9836 1571 9871 1577
rect 9973 1571 10427 1577
rect 10529 1571 10564 1577
rect 9836 1563 9894 1571
rect 9836 1536 9877 1563
rect 9423 1137 9464 1164
rect 9406 1129 9464 1137
rect 8736 1123 8771 1129
rect 8873 1123 9327 1129
rect 9429 1123 9464 1129
rect 9836 1137 9877 1164
rect 9836 1129 9894 1137
rect 9956 1563 10444 1571
rect 9973 1515 10427 1563
rect 9973 1185 10035 1515
rect 10365 1185 10427 1515
rect 9973 1137 10427 1185
rect 9956 1129 10444 1137
rect 10506 1563 10564 1571
rect 10523 1536 10564 1563
rect 10936 1571 10971 1577
rect 11073 1571 11527 1577
rect 11629 1571 11664 1577
rect 10936 1563 10994 1571
rect 10936 1536 10977 1563
rect 10523 1137 10564 1164
rect 10506 1129 10564 1137
rect 9836 1123 9871 1129
rect 9973 1123 10427 1129
rect 10529 1123 10564 1129
rect 10936 1137 10977 1164
rect 10936 1129 10994 1137
rect 11056 1563 11544 1571
rect 11073 1515 11527 1563
rect 11073 1185 11135 1515
rect 11465 1185 11527 1515
rect 11073 1137 11527 1185
rect 11056 1129 11544 1137
rect 11606 1563 11664 1571
rect 11623 1536 11664 1563
rect 12036 1571 12071 1577
rect 12173 1571 12627 1577
rect 12729 1571 12764 1577
rect 12036 1563 12094 1571
rect 12036 1536 12077 1563
rect 11623 1137 11664 1164
rect 11606 1129 11664 1137
rect 10936 1123 10971 1129
rect 11073 1123 11527 1129
rect 11629 1123 11664 1129
rect 12036 1137 12077 1164
rect 12036 1129 12094 1137
rect 12156 1563 12644 1571
rect 12173 1515 12627 1563
rect 12173 1185 12235 1515
rect 12565 1185 12627 1515
rect 12173 1137 12627 1185
rect 12156 1129 12644 1137
rect 12706 1563 12764 1571
rect 12723 1536 12764 1563
rect 13136 1571 13171 1577
rect 13273 1571 13727 1577
rect 13136 1563 13194 1571
rect 13136 1536 13177 1563
rect 12723 1137 12764 1164
rect 12706 1129 12764 1137
rect 12036 1123 12071 1129
rect 12173 1123 12627 1129
rect 12729 1123 12764 1129
rect 13136 1137 13177 1164
rect 13136 1129 13194 1137
rect 13256 1563 13727 1571
rect 13273 1515 13727 1563
rect 13273 1185 13335 1515
rect 13665 1185 13727 1515
rect 13273 1137 13727 1185
rect 13256 1129 13727 1137
rect 13136 1123 13171 1129
rect 13273 1123 13727 1129
rect -1025 1100 -725 1117
rect -471 1106 -463 1123
rect -37 1106 -29 1123
rect 79 1106 87 1123
rect 513 1106 521 1123
rect 629 1106 637 1123
rect 1063 1106 1071 1123
rect 1179 1106 1187 1123
rect 1613 1106 1621 1123
rect 1729 1106 1737 1123
rect 2163 1106 2171 1123
rect 2279 1106 2287 1123
rect 2713 1106 2721 1123
rect 2829 1106 2837 1123
rect 3263 1106 3271 1123
rect 3379 1106 3387 1123
rect 3813 1106 3821 1123
rect 3929 1106 3937 1123
rect 4363 1106 4371 1123
rect 4479 1106 4487 1123
rect 4913 1106 4921 1123
rect 5029 1106 5037 1123
rect 5463 1106 5471 1123
rect 5579 1106 5587 1123
rect 6013 1106 6021 1123
rect 6129 1106 6137 1123
rect 6563 1106 6571 1123
rect 6679 1106 6687 1123
rect 7113 1106 7121 1123
rect 7229 1106 7237 1123
rect 7663 1106 7671 1123
rect 7779 1106 7787 1123
rect 8213 1106 8221 1123
rect 8329 1106 8337 1123
rect 8763 1106 8771 1123
rect 8879 1106 8887 1123
rect 9313 1106 9321 1123
rect 9429 1106 9437 1123
rect 9863 1106 9871 1123
rect 9979 1106 9987 1123
rect 10413 1106 10421 1123
rect 10529 1106 10537 1123
rect 10963 1106 10971 1123
rect 11079 1106 11087 1123
rect 11513 1106 11521 1123
rect 11629 1106 11637 1123
rect 12063 1106 12071 1123
rect 12179 1106 12187 1123
rect 12613 1106 12621 1123
rect 12729 1106 12737 1123
rect 13163 1106 13171 1123
rect 13279 1106 13287 1123
rect 13713 1106 13721 1123
rect 13975 1117 13987 1650
rect 14263 1117 14275 1650
rect 13975 1100 14275 1117
rect -1025 567 -1013 1100
rect -737 567 -725 1100
rect -550 1092 -500 1100
rect -550 1058 -542 1092
rect -508 1058 -500 1092
rect -550 1050 -500 1058
rect 0 1092 50 1100
rect 0 1058 8 1092
rect 42 1058 50 1092
rect 0 1050 50 1058
rect 550 1092 600 1100
rect 550 1058 558 1092
rect 592 1058 600 1092
rect 550 1050 600 1058
rect 1100 1092 1150 1100
rect 1100 1058 1108 1092
rect 1142 1058 1150 1092
rect 1100 1050 1150 1058
rect 1650 1092 1700 1100
rect 1650 1058 1658 1092
rect 1692 1058 1700 1092
rect 1650 1050 1700 1058
rect 2200 1092 2250 1100
rect 2200 1058 2208 1092
rect 2242 1058 2250 1092
rect 2200 1050 2250 1058
rect 2750 1092 2800 1100
rect 2750 1058 2758 1092
rect 2792 1058 2800 1092
rect 2750 1050 2800 1058
rect 3300 1092 3350 1100
rect 3300 1058 3308 1092
rect 3342 1058 3350 1092
rect 3300 1050 3350 1058
rect 3850 1092 3900 1100
rect 3850 1058 3858 1092
rect 3892 1058 3900 1092
rect 3850 1050 3900 1058
rect 4400 1092 4450 1100
rect 4400 1058 4408 1092
rect 4442 1058 4450 1092
rect 4400 1050 4450 1058
rect 4950 1092 5000 1100
rect 4950 1058 4958 1092
rect 4992 1058 5000 1092
rect 4950 1050 5000 1058
rect 5500 1092 5550 1100
rect 5500 1058 5508 1092
rect 5542 1058 5550 1092
rect 5500 1050 5550 1058
rect 6050 1092 6100 1100
rect 6050 1058 6058 1092
rect 6092 1058 6100 1092
rect 6050 1050 6100 1058
rect 6600 1092 6650 1100
rect 6600 1058 6608 1092
rect 6642 1058 6650 1092
rect 6600 1050 6650 1058
rect 7150 1092 7200 1100
rect 7150 1058 7158 1092
rect 7192 1058 7200 1092
rect 7150 1050 7200 1058
rect 7700 1092 7750 1100
rect 7700 1058 7708 1092
rect 7742 1058 7750 1092
rect 7700 1050 7750 1058
rect 8250 1092 8300 1100
rect 8250 1058 8258 1092
rect 8292 1058 8300 1092
rect 8250 1050 8300 1058
rect 8800 1092 8850 1100
rect 8800 1058 8808 1092
rect 8842 1058 8850 1092
rect 8800 1050 8850 1058
rect 9350 1092 9400 1100
rect 9350 1058 9358 1092
rect 9392 1058 9400 1092
rect 9350 1050 9400 1058
rect 9900 1092 9950 1100
rect 9900 1058 9908 1092
rect 9942 1058 9950 1092
rect 9900 1050 9950 1058
rect 10450 1092 10500 1100
rect 10450 1058 10458 1092
rect 10492 1058 10500 1092
rect 10450 1050 10500 1058
rect 11000 1092 11050 1100
rect 11000 1058 11008 1092
rect 11042 1058 11050 1092
rect 11000 1050 11050 1058
rect 11550 1092 11600 1100
rect 11550 1058 11558 1092
rect 11592 1058 11600 1092
rect 11550 1050 11600 1058
rect 12100 1092 12150 1100
rect 12100 1058 12108 1092
rect 12142 1058 12150 1092
rect 12100 1050 12150 1058
rect 12650 1092 12700 1100
rect 12650 1058 12658 1092
rect 12692 1058 12700 1092
rect 12650 1050 12700 1058
rect 13200 1092 13250 1100
rect 13200 1058 13208 1092
rect 13242 1058 13250 1092
rect 13200 1050 13250 1058
rect 13750 1092 13800 1100
rect 13750 1058 13758 1092
rect 13792 1058 13800 1092
rect 13750 1050 13800 1058
rect -471 1027 -463 1044
rect -37 1027 -29 1044
rect 79 1027 87 1044
rect 513 1027 521 1044
rect 629 1027 637 1044
rect 1063 1027 1071 1044
rect 1179 1027 1187 1044
rect 1613 1027 1621 1044
rect 1729 1027 1737 1044
rect 2163 1027 2171 1044
rect 2279 1027 2287 1044
rect 2713 1027 2721 1044
rect 2829 1027 2837 1044
rect 3263 1027 3271 1044
rect 3379 1027 3387 1044
rect 3813 1027 3821 1044
rect 3929 1027 3937 1044
rect 4363 1027 4371 1044
rect 4479 1027 4487 1044
rect 4913 1027 4921 1044
rect 5029 1027 5037 1044
rect 5463 1027 5471 1044
rect 5579 1027 5587 1044
rect 6013 1027 6021 1044
rect 6129 1027 6137 1044
rect 6563 1027 6571 1044
rect 6679 1027 6687 1044
rect 7113 1027 7121 1044
rect 7229 1027 7237 1044
rect 7663 1027 7671 1044
rect 7779 1027 7787 1044
rect 8213 1027 8221 1044
rect 8329 1027 8337 1044
rect 8763 1027 8771 1044
rect 8879 1027 8887 1044
rect 9313 1027 9321 1044
rect 9429 1027 9437 1044
rect 9863 1027 9871 1044
rect 9979 1027 9987 1044
rect 10413 1027 10421 1044
rect 10529 1027 10537 1044
rect 10963 1027 10971 1044
rect 11079 1027 11087 1044
rect 11513 1027 11521 1044
rect 11629 1027 11637 1044
rect 12063 1027 12071 1044
rect 12179 1027 12187 1044
rect 12613 1027 12621 1044
rect 12729 1027 12737 1044
rect 13163 1027 13171 1044
rect 13279 1027 13287 1044
rect 13713 1027 13721 1044
rect -477 1021 -23 1027
rect 79 1021 114 1027
rect -477 1013 -6 1021
rect -477 965 -23 1013
rect -477 635 -415 965
rect -85 635 -23 965
rect -477 587 -23 635
rect -477 579 -6 587
rect 56 1013 114 1021
rect 73 986 114 1013
rect 486 1021 521 1027
rect 623 1021 1077 1027
rect 1179 1021 1214 1027
rect 486 1013 544 1021
rect 486 986 527 1013
rect 73 587 114 614
rect 56 579 114 587
rect -477 573 -23 579
rect 79 573 114 579
rect 486 587 527 614
rect 486 579 544 587
rect 606 1013 1094 1021
rect 623 965 1077 1013
rect 623 635 685 965
rect 1015 635 1077 965
rect 623 587 1077 635
rect 606 579 1094 587
rect 1156 1013 1214 1021
rect 1173 986 1214 1013
rect 1586 1021 1621 1027
rect 1723 1021 2177 1027
rect 2279 1021 2314 1027
rect 1586 1013 1644 1021
rect 1586 986 1627 1013
rect 1173 587 1214 614
rect 1156 579 1214 587
rect 486 573 521 579
rect 623 573 1077 579
rect 1179 573 1214 579
rect 1586 587 1627 614
rect 1586 579 1644 587
rect 1706 1013 2194 1021
rect 1723 965 2177 1013
rect 1723 635 1785 965
rect 2115 635 2177 965
rect 1723 587 2177 635
rect 1706 579 2194 587
rect 2256 1013 2314 1021
rect 2273 986 2314 1013
rect 2686 1021 2721 1027
rect 2823 1021 3277 1027
rect 3379 1021 3414 1027
rect 2686 1013 2744 1021
rect 2686 986 2727 1013
rect 2273 587 2314 614
rect 2256 579 2314 587
rect 1586 573 1621 579
rect 1723 573 2177 579
rect 2279 573 2314 579
rect 2686 587 2727 614
rect 2686 579 2744 587
rect 2806 1013 3294 1021
rect 2823 965 3277 1013
rect 2823 635 2885 965
rect 3215 635 3277 965
rect 2823 587 3277 635
rect 2806 579 3294 587
rect 3356 1013 3414 1021
rect 3373 986 3414 1013
rect 3786 1021 3821 1027
rect 3923 1021 4377 1027
rect 4479 1021 4514 1027
rect 3786 1013 3844 1021
rect 3786 986 3827 1013
rect 3373 587 3414 614
rect 3356 579 3414 587
rect 2686 573 2721 579
rect 2823 573 3277 579
rect 3379 573 3414 579
rect 3786 587 3827 614
rect 3786 579 3844 587
rect 3906 1013 4394 1021
rect 3923 965 4377 1013
rect 3923 635 3985 965
rect 4315 635 4377 965
rect 3923 587 4377 635
rect 3906 579 4394 587
rect 4456 1013 4514 1021
rect 4473 986 4514 1013
rect 4886 1021 4921 1027
rect 5023 1021 5477 1027
rect 5579 1021 5614 1027
rect 4886 1013 4944 1021
rect 4886 986 4927 1013
rect 4473 587 4514 614
rect 4456 579 4514 587
rect 3786 573 3821 579
rect 3923 573 4377 579
rect 4479 573 4514 579
rect 4886 587 4927 614
rect 4886 579 4944 587
rect 5006 1013 5494 1021
rect 5023 965 5477 1013
rect 5023 635 5085 965
rect 5415 635 5477 965
rect 5023 587 5477 635
rect 5006 579 5494 587
rect 5556 1013 5614 1021
rect 5573 986 5614 1013
rect 5986 1021 6021 1027
rect 6123 1021 6577 1027
rect 6679 1021 6714 1027
rect 5986 1013 6044 1021
rect 5986 986 6027 1013
rect 5573 587 5614 614
rect 5556 579 5614 587
rect 4886 573 4921 579
rect 5023 573 5477 579
rect 5579 573 5614 579
rect 5986 587 6027 614
rect 5986 579 6044 587
rect 6106 1013 6594 1021
rect 6123 965 6577 1013
rect 6123 635 6185 965
rect 6515 635 6577 965
rect 6123 587 6577 635
rect 6106 579 6594 587
rect 6656 1013 6714 1021
rect 6673 986 6714 1013
rect 7086 1021 7121 1027
rect 7223 1021 7677 1027
rect 7779 1021 7814 1027
rect 7086 1013 7144 1021
rect 7086 986 7127 1013
rect 6673 587 6714 614
rect 6656 579 6714 587
rect 5986 573 6021 579
rect 6123 573 6577 579
rect 6679 573 6714 579
rect 7086 587 7127 614
rect 7086 579 7144 587
rect 7206 1013 7694 1021
rect 7223 965 7677 1013
rect 7223 635 7285 965
rect 7615 635 7677 965
rect 7223 587 7677 635
rect 7206 579 7694 587
rect 7756 1013 7814 1021
rect 7773 986 7814 1013
rect 8186 1021 8221 1027
rect 8323 1021 8777 1027
rect 8879 1021 8914 1027
rect 8186 1013 8244 1021
rect 8186 986 8227 1013
rect 7773 587 7814 614
rect 7756 579 7814 587
rect 7086 573 7121 579
rect 7223 573 7677 579
rect 7779 573 7814 579
rect 8186 587 8227 614
rect 8186 579 8244 587
rect 8306 1013 8794 1021
rect 8323 965 8777 1013
rect 8323 635 8385 965
rect 8715 635 8777 965
rect 8323 587 8777 635
rect 8306 579 8794 587
rect 8856 1013 8914 1021
rect 8873 986 8914 1013
rect 9286 1021 9321 1027
rect 9423 1021 9877 1027
rect 9979 1021 10014 1027
rect 9286 1013 9344 1021
rect 9286 986 9327 1013
rect 8873 587 8914 614
rect 8856 579 8914 587
rect 8186 573 8221 579
rect 8323 573 8777 579
rect 8879 573 8914 579
rect 9286 587 9327 614
rect 9286 579 9344 587
rect 9406 1013 9894 1021
rect 9423 965 9877 1013
rect 9423 635 9485 965
rect 9815 635 9877 965
rect 9423 587 9877 635
rect 9406 579 9894 587
rect 9956 1013 10014 1021
rect 9973 986 10014 1013
rect 10386 1021 10421 1027
rect 10523 1021 10977 1027
rect 11079 1021 11114 1027
rect 10386 1013 10444 1021
rect 10386 986 10427 1013
rect 9973 587 10014 614
rect 9956 579 10014 587
rect 9286 573 9321 579
rect 9423 573 9877 579
rect 9979 573 10014 579
rect 10386 587 10427 614
rect 10386 579 10444 587
rect 10506 1013 10994 1021
rect 10523 965 10977 1013
rect 10523 635 10585 965
rect 10915 635 10977 965
rect 10523 587 10977 635
rect 10506 579 10994 587
rect 11056 1013 11114 1021
rect 11073 986 11114 1013
rect 11486 1021 11521 1027
rect 11623 1021 12077 1027
rect 12179 1021 12214 1027
rect 11486 1013 11544 1021
rect 11486 986 11527 1013
rect 11073 587 11114 614
rect 11056 579 11114 587
rect 10386 573 10421 579
rect 10523 573 10977 579
rect 11079 573 11114 579
rect 11486 587 11527 614
rect 11486 579 11544 587
rect 11606 1013 12094 1021
rect 11623 965 12077 1013
rect 11623 635 11685 965
rect 12015 635 12077 965
rect 11623 587 12077 635
rect 11606 579 12094 587
rect 12156 1013 12214 1021
rect 12173 986 12214 1013
rect 12586 1021 12621 1027
rect 12723 1021 13177 1027
rect 13279 1021 13314 1027
rect 12586 1013 12644 1021
rect 12586 986 12627 1013
rect 12173 587 12214 614
rect 12156 579 12214 587
rect 11486 573 11521 579
rect 11623 573 12077 579
rect 12179 573 12214 579
rect 12586 587 12627 614
rect 12586 579 12644 587
rect 12706 1013 13194 1021
rect 12723 965 13177 1013
rect 12723 635 12785 965
rect 13115 635 13177 965
rect 12723 587 13177 635
rect 12706 579 13194 587
rect 13256 1013 13314 1021
rect 13273 986 13314 1013
rect 13273 587 13314 614
rect 13256 579 13314 587
rect 12586 573 12621 579
rect 12723 573 13177 579
rect 13279 573 13314 579
rect -1025 550 -725 567
rect -471 556 -463 573
rect -37 556 -29 573
rect 79 556 87 573
rect 513 556 521 573
rect 629 556 637 573
rect 1063 556 1071 573
rect 1179 556 1187 573
rect 1613 556 1621 573
rect 1729 556 1737 573
rect 2163 556 2171 573
rect 2279 556 2287 573
rect 2713 556 2721 573
rect 2829 556 2837 573
rect 3263 556 3271 573
rect 3379 556 3387 573
rect 3813 556 3821 573
rect 3929 556 3937 573
rect 4363 556 4371 573
rect 4479 556 4487 573
rect 4913 556 4921 573
rect 5029 556 5037 573
rect 5463 556 5471 573
rect 5579 556 5587 573
rect 6013 556 6021 573
rect 6129 556 6137 573
rect 6563 556 6571 573
rect 6679 556 6687 573
rect 7113 556 7121 573
rect 7229 556 7237 573
rect 7663 556 7671 573
rect 7779 556 7787 573
rect 8213 556 8221 573
rect 8329 556 8337 573
rect 8763 556 8771 573
rect 8879 556 8887 573
rect 9313 556 9321 573
rect 9429 556 9437 573
rect 9863 556 9871 573
rect 9979 556 9987 573
rect 10413 556 10421 573
rect 10529 556 10537 573
rect 10963 556 10971 573
rect 11079 556 11087 573
rect 11513 556 11521 573
rect 11629 556 11637 573
rect 12063 556 12071 573
rect 12179 556 12187 573
rect 12613 556 12621 573
rect 12729 556 12737 573
rect 13163 556 13171 573
rect 13279 556 13287 573
rect 13713 556 13721 573
rect 13975 569 13987 1100
rect 14263 569 14275 1100
rect 13975 550 14275 569
rect -1025 17 -1013 550
rect -737 17 -725 550
rect -550 542 -500 550
rect -550 508 -542 542
rect -508 508 -500 542
rect -550 500 -500 508
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 550 542 600 550
rect 550 508 558 542
rect 592 508 600 542
rect 550 500 600 508
rect 1100 542 1150 550
rect 1100 508 1108 542
rect 1142 508 1150 542
rect 1100 500 1150 508
rect 1650 542 1700 550
rect 1650 508 1658 542
rect 1692 508 1700 542
rect 1650 500 1700 508
rect 2200 542 2250 550
rect 2200 508 2208 542
rect 2242 508 2250 542
rect 2200 500 2250 508
rect 2750 542 2800 550
rect 2750 508 2758 542
rect 2792 508 2800 542
rect 2750 500 2800 508
rect 3300 542 3350 550
rect 3300 508 3308 542
rect 3342 508 3350 542
rect 3300 500 3350 508
rect 3850 542 3900 550
rect 3850 508 3858 542
rect 3892 508 3900 542
rect 3850 500 3900 508
rect 4400 542 4450 550
rect 4400 508 4408 542
rect 4442 508 4450 542
rect 4400 500 4450 508
rect 4950 542 5000 550
rect 4950 508 4958 542
rect 4992 508 5000 542
rect 4950 500 5000 508
rect 5500 542 5550 550
rect 5500 508 5508 542
rect 5542 508 5550 542
rect 5500 500 5550 508
rect 6050 542 6100 550
rect 6050 508 6058 542
rect 6092 508 6100 542
rect 6050 500 6100 508
rect 6600 542 6650 550
rect 6600 508 6608 542
rect 6642 508 6650 542
rect 6600 500 6650 508
rect 7150 542 7200 550
rect 7150 508 7158 542
rect 7192 508 7200 542
rect 7150 500 7200 508
rect 7700 542 7750 550
rect 7700 508 7708 542
rect 7742 508 7750 542
rect 7700 500 7750 508
rect 8250 542 8300 550
rect 8250 508 8258 542
rect 8292 508 8300 542
rect 8250 500 8300 508
rect 8800 542 8850 550
rect 8800 508 8808 542
rect 8842 508 8850 542
rect 8800 500 8850 508
rect 9350 542 9400 550
rect 9350 508 9358 542
rect 9392 508 9400 542
rect 9350 500 9400 508
rect 9900 542 9950 550
rect 9900 508 9908 542
rect 9942 508 9950 542
rect 9900 500 9950 508
rect 10450 542 10500 550
rect 10450 508 10458 542
rect 10492 508 10500 542
rect 10450 500 10500 508
rect 11000 542 11050 550
rect 11000 508 11008 542
rect 11042 508 11050 542
rect 11000 500 11050 508
rect 11550 542 11600 550
rect 11550 508 11558 542
rect 11592 508 11600 542
rect 11550 500 11600 508
rect 12100 542 12150 550
rect 12100 508 12108 542
rect 12142 508 12150 542
rect 12100 500 12150 508
rect 12650 542 12700 550
rect 12650 508 12658 542
rect 12692 508 12700 542
rect 12650 500 12700 508
rect 13200 542 13250 550
rect 13200 508 13208 542
rect 13242 508 13250 542
rect 13200 500 13250 508
rect 13750 542 13800 550
rect 13750 508 13758 542
rect 13792 508 13800 542
rect 13750 500 13800 508
rect -471 477 -463 494
rect -37 477 -29 494
rect 79 477 87 494
rect 513 477 521 494
rect 629 477 637 494
rect 1063 477 1071 494
rect 1179 477 1187 494
rect 1613 477 1621 494
rect 1729 477 1737 494
rect 2163 477 2171 494
rect 2279 477 2287 494
rect 2713 477 2721 494
rect 2829 477 2837 494
rect 3263 477 3271 494
rect 3379 477 3387 494
rect 3813 477 3821 494
rect 3929 477 3937 494
rect 4363 477 4371 494
rect 4479 477 4487 494
rect 4913 477 4921 494
rect 5029 477 5037 494
rect 5463 477 5471 494
rect 5579 477 5587 494
rect 6013 477 6021 494
rect 6129 477 6137 494
rect 6563 477 6571 494
rect 6679 477 6687 494
rect 7113 477 7121 494
rect 7229 477 7237 494
rect 7663 477 7671 494
rect 7779 477 7787 494
rect 8213 477 8221 494
rect 8329 477 8337 494
rect 8763 477 8771 494
rect 8879 477 8887 494
rect 9313 477 9321 494
rect 9429 477 9437 494
rect 9863 477 9871 494
rect 9979 477 9987 494
rect 10413 477 10421 494
rect 10529 477 10537 494
rect 10963 477 10971 494
rect 11079 477 11087 494
rect 11513 477 11521 494
rect 11629 477 11637 494
rect 12063 477 12071 494
rect 12179 477 12187 494
rect 12613 477 12621 494
rect 12729 477 12737 494
rect 13163 477 13171 494
rect 13279 477 13287 494
rect 13713 477 13721 494
rect -64 471 -29 477
rect 73 471 527 477
rect 629 471 664 477
rect -64 463 -6 471
rect -64 436 -23 463
rect -64 37 -23 64
rect -64 29 -6 37
rect 56 463 544 471
rect 73 415 527 463
rect 73 85 135 415
rect 465 85 527 415
rect 73 37 527 85
rect 56 29 544 37
rect 606 463 664 471
rect 623 436 664 463
rect 1036 471 1071 477
rect 1173 471 1627 477
rect 1729 471 1764 477
rect 1036 463 1094 471
rect 1036 436 1077 463
rect 623 37 664 64
rect 606 29 664 37
rect -64 23 -29 29
rect 73 23 527 29
rect 629 23 664 29
rect 1036 37 1077 64
rect 1036 29 1094 37
rect 1156 463 1644 471
rect 1173 415 1627 463
rect 1173 85 1235 415
rect 1565 85 1627 415
rect 1173 37 1627 85
rect 1156 29 1644 37
rect 1706 463 1764 471
rect 1723 436 1764 463
rect 2136 471 2171 477
rect 2273 471 2727 477
rect 2829 471 2864 477
rect 2136 463 2194 471
rect 2136 436 2177 463
rect 1723 37 1764 64
rect 1706 29 1764 37
rect 1036 23 1071 29
rect 1173 23 1627 29
rect 1729 23 1764 29
rect 2136 37 2177 64
rect 2136 29 2194 37
rect 2256 463 2744 471
rect 2273 415 2727 463
rect 2273 85 2335 415
rect 2665 85 2727 415
rect 2273 37 2727 85
rect 2256 29 2744 37
rect 2806 463 2864 471
rect 2823 436 2864 463
rect 3236 471 3271 477
rect 3373 471 3827 477
rect 3929 471 3964 477
rect 3236 463 3294 471
rect 3236 436 3277 463
rect 2823 37 2864 64
rect 2806 29 2864 37
rect 2136 23 2171 29
rect 2273 23 2727 29
rect 2829 23 2864 29
rect 3236 37 3277 64
rect 3236 29 3294 37
rect 3356 463 3844 471
rect 3373 415 3827 463
rect 3373 85 3435 415
rect 3765 85 3827 415
rect 3373 37 3827 85
rect 3356 29 3844 37
rect 3906 463 3964 471
rect 3923 436 3964 463
rect 4336 471 4371 477
rect 4473 471 4927 477
rect 5029 471 5064 477
rect 4336 463 4394 471
rect 4336 436 4377 463
rect 3923 37 3964 64
rect 3906 29 3964 37
rect 3236 23 3271 29
rect 3373 23 3827 29
rect 3929 23 3964 29
rect 4336 37 4377 64
rect 4336 29 4394 37
rect 4456 463 4944 471
rect 4473 415 4927 463
rect 4473 85 4535 415
rect 4865 85 4927 415
rect 4473 37 4927 85
rect 4456 29 4944 37
rect 5006 463 5064 471
rect 5023 436 5064 463
rect 5436 471 5471 477
rect 5573 471 6027 477
rect 6129 471 6164 477
rect 5436 463 5494 471
rect 5436 436 5477 463
rect 5023 37 5064 64
rect 5006 29 5064 37
rect 4336 23 4371 29
rect 4473 23 4927 29
rect 5029 23 5064 29
rect 5436 37 5477 64
rect 5436 29 5494 37
rect 5556 463 6044 471
rect 5573 415 6027 463
rect 5573 85 5635 415
rect 5965 85 6027 415
rect 5573 37 6027 85
rect 5556 29 6044 37
rect 6106 463 6164 471
rect 6123 436 6164 463
rect 6536 471 6571 477
rect 6673 471 7127 477
rect 7229 471 7264 477
rect 6536 463 6594 471
rect 6536 436 6577 463
rect 6123 37 6164 64
rect 6106 29 6164 37
rect 5436 23 5471 29
rect 5573 23 6027 29
rect 6129 23 6164 29
rect 6536 37 6577 64
rect 6536 29 6594 37
rect 6656 463 7144 471
rect 6673 415 7127 463
rect 6673 85 6735 415
rect 7065 85 7127 415
rect 6673 37 7127 85
rect 6656 29 7144 37
rect 7206 463 7264 471
rect 7223 436 7264 463
rect 7636 471 7671 477
rect 7773 471 8227 477
rect 8329 471 8364 477
rect 7636 463 7694 471
rect 7636 436 7677 463
rect 7223 37 7264 64
rect 7206 29 7264 37
rect 6536 23 6571 29
rect 6673 23 7127 29
rect 7229 23 7264 29
rect 7636 37 7677 64
rect 7636 29 7694 37
rect 7756 463 8244 471
rect 7773 415 8227 463
rect 7773 85 7835 415
rect 8165 85 8227 415
rect 7773 37 8227 85
rect 7756 29 8244 37
rect 8306 463 8364 471
rect 8323 436 8364 463
rect 8736 471 8771 477
rect 8873 471 9327 477
rect 9429 471 9464 477
rect 8736 463 8794 471
rect 8736 436 8777 463
rect 8323 37 8364 64
rect 8306 29 8364 37
rect 7636 23 7671 29
rect 7773 23 8227 29
rect 8329 23 8364 29
rect 8736 37 8777 64
rect 8736 29 8794 37
rect 8856 463 9344 471
rect 8873 415 9327 463
rect 8873 85 8935 415
rect 9265 85 9327 415
rect 8873 37 9327 85
rect 8856 29 9344 37
rect 9406 463 9464 471
rect 9423 436 9464 463
rect 9836 471 9871 477
rect 9973 471 10427 477
rect 10529 471 10564 477
rect 9836 463 9894 471
rect 9836 436 9877 463
rect 9423 37 9464 64
rect 9406 29 9464 37
rect 8736 23 8771 29
rect 8873 23 9327 29
rect 9429 23 9464 29
rect 9836 37 9877 64
rect 9836 29 9894 37
rect 9956 463 10444 471
rect 9973 415 10427 463
rect 9973 85 10035 415
rect 10365 85 10427 415
rect 9973 37 10427 85
rect 9956 29 10444 37
rect 10506 463 10564 471
rect 10523 436 10564 463
rect 10936 471 10971 477
rect 11073 471 11527 477
rect 11629 471 11664 477
rect 10936 463 10994 471
rect 10936 436 10977 463
rect 10523 37 10564 64
rect 10506 29 10564 37
rect 9836 23 9871 29
rect 9973 23 10427 29
rect 10529 23 10564 29
rect 10936 37 10977 64
rect 10936 29 10994 37
rect 11056 463 11544 471
rect 11073 415 11527 463
rect 11073 85 11135 415
rect 11465 85 11527 415
rect 11073 37 11527 85
rect 11056 29 11544 37
rect 11606 463 11664 471
rect 11623 436 11664 463
rect 12036 471 12071 477
rect 12173 471 12627 477
rect 12729 471 12764 477
rect 12036 463 12094 471
rect 12036 436 12077 463
rect 11623 37 11664 64
rect 11606 29 11664 37
rect 10936 23 10971 29
rect 11073 23 11527 29
rect 11629 23 11664 29
rect 12036 37 12077 64
rect 12036 29 12094 37
rect 12156 463 12644 471
rect 12173 415 12627 463
rect 12173 85 12235 415
rect 12565 85 12627 415
rect 12173 37 12627 85
rect 12156 29 12644 37
rect 12706 463 12764 471
rect 12723 436 12764 463
rect 13136 471 13171 477
rect 13273 471 13727 477
rect 13136 463 13194 471
rect 13136 436 13177 463
rect 12723 37 12764 64
rect 12706 29 12764 37
rect 12036 23 12071 29
rect 12173 23 12627 29
rect 12729 23 12764 29
rect 13136 37 13177 64
rect 13136 29 13194 37
rect 13256 463 13727 471
rect 13273 415 13727 463
rect 13273 85 13335 415
rect 13665 85 13727 415
rect 13273 37 13727 85
rect 13256 29 13727 37
rect 13136 23 13171 29
rect 13273 23 13727 29
rect -1025 0 -725 17
rect -471 6 -463 23
rect -37 6 -29 23
rect 79 6 87 23
rect 513 6 521 23
rect 629 6 637 23
rect 1063 6 1071 23
rect 1179 6 1187 23
rect 1613 6 1621 23
rect 1729 6 1737 23
rect 2163 6 2171 23
rect 2279 6 2287 23
rect 2713 6 2721 23
rect 2829 6 2837 23
rect 3263 6 3271 23
rect 3379 6 3387 23
rect 3813 6 3821 23
rect 3929 6 3937 23
rect 4363 6 4371 23
rect 4479 6 4487 23
rect 4913 6 4921 23
rect 5029 6 5037 23
rect 5463 6 5471 23
rect 5579 6 5587 23
rect 6013 6 6021 23
rect 6129 6 6137 23
rect 6563 6 6571 23
rect 6679 6 6687 23
rect 7113 6 7121 23
rect 7229 6 7237 23
rect 7663 6 7671 23
rect 7779 6 7787 23
rect 8213 6 8221 23
rect 8329 6 8337 23
rect 8763 6 8771 23
rect 8879 6 8887 23
rect 9313 6 9321 23
rect 9429 6 9437 23
rect 9863 6 9871 23
rect 9979 6 9987 23
rect 10413 6 10421 23
rect 10529 6 10537 23
rect 10963 6 10971 23
rect 11079 6 11087 23
rect 11513 6 11521 23
rect 11629 6 11637 23
rect 12063 6 12071 23
rect 12179 6 12187 23
rect 12613 6 12621 23
rect 12729 6 12737 23
rect 13163 6 13171 23
rect 13279 6 13287 23
rect 13713 6 13721 23
rect 13975 17 13987 550
rect 14263 17 14275 550
rect 13975 0 14275 17
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 0 -8 50 0
rect 0 -42 8 -8
rect 42 -42 50 -8
rect 0 -50 50 -42
rect 550 -8 600 0
rect 550 -42 558 -8
rect 592 -42 600 -8
rect 550 -50 600 -42
rect 1100 -8 1150 0
rect 1100 -42 1108 -8
rect 1142 -42 1150 -8
rect 1100 -50 1150 -42
rect 1650 -8 1700 0
rect 1650 -42 1658 -8
rect 1692 -42 1700 -8
rect 1650 -50 1700 -42
rect 2200 -8 2250 0
rect 2200 -42 2208 -8
rect 2242 -42 2250 -8
rect 2200 -50 2250 -42
rect 2750 -8 2800 0
rect 2750 -42 2758 -8
rect 2792 -42 2800 -8
rect 2750 -50 2800 -42
rect 3300 -8 3350 0
rect 3300 -42 3308 -8
rect 3342 -42 3350 -8
rect 3300 -50 3350 -42
rect 3850 -8 3900 0
rect 3850 -42 3858 -8
rect 3892 -42 3900 -8
rect 3850 -50 3900 -42
rect 4400 -8 4450 0
rect 4400 -42 4408 -8
rect 4442 -42 4450 -8
rect 4400 -50 4450 -42
rect 4950 -8 5000 0
rect 4950 -42 4958 -8
rect 4992 -42 5000 -8
rect 4950 -50 5000 -42
rect 5500 -8 5550 0
rect 5500 -42 5508 -8
rect 5542 -42 5550 -8
rect 5500 -50 5550 -42
rect 6050 -8 6100 0
rect 6050 -42 6058 -8
rect 6092 -42 6100 -8
rect 6050 -50 6100 -42
rect 6600 -8 6650 0
rect 6600 -42 6608 -8
rect 6642 -42 6650 -8
rect 6600 -50 6650 -42
rect 7150 -8 7200 0
rect 7150 -42 7158 -8
rect 7192 -42 7200 -8
rect 7150 -50 7200 -42
rect 7700 -8 7750 0
rect 7700 -42 7708 -8
rect 7742 -42 7750 -8
rect 7700 -50 7750 -42
rect 8250 -8 8300 0
rect 8250 -42 8258 -8
rect 8292 -42 8300 -8
rect 8250 -50 8300 -42
rect 8800 -8 8850 0
rect 8800 -42 8808 -8
rect 8842 -42 8850 -8
rect 8800 -50 8850 -42
rect 9350 -8 9400 0
rect 9350 -42 9358 -8
rect 9392 -42 9400 -8
rect 9350 -50 9400 -42
rect 9900 -8 9950 0
rect 9900 -42 9908 -8
rect 9942 -42 9950 -8
rect 9900 -50 9950 -42
rect 10450 -8 10500 0
rect 10450 -42 10458 -8
rect 10492 -42 10500 -8
rect 10450 -50 10500 -42
rect 11000 -8 11050 0
rect 11000 -42 11008 -8
rect 11042 -42 11050 -8
rect 11000 -50 11050 -42
rect 11550 -8 11600 0
rect 11550 -42 11558 -8
rect 11592 -42 11600 -8
rect 11550 -50 11600 -42
rect 12100 -8 12150 0
rect 12100 -42 12108 -8
rect 12142 -42 12150 -8
rect 12100 -50 12150 -42
rect 12650 -8 12700 0
rect 12650 -42 12658 -8
rect 12692 -42 12700 -8
rect 12650 -50 12700 -42
rect 13200 -8 13250 0
rect 13200 -42 13208 -8
rect 13242 -42 13250 -8
rect 13200 -50 13250 -42
rect 13750 -8 13800 0
rect 13750 -42 13758 -8
rect 13792 -42 13800 -8
rect 13750 -50 13800 -42
rect -471 -73 -463 -56
rect -37 -73 -29 -56
rect 79 -73 87 -56
rect 513 -73 521 -56
rect 629 -73 637 -56
rect 1063 -73 1071 -56
rect 1179 -73 1187 -56
rect 1613 -73 1621 -56
rect 1729 -73 1737 -56
rect 2163 -73 2171 -56
rect 2279 -73 2287 -56
rect 2713 -73 2721 -56
rect 2829 -73 2837 -56
rect 3263 -73 3271 -56
rect 3379 -73 3387 -56
rect 3813 -73 3821 -56
rect 3929 -73 3937 -56
rect 4363 -73 4371 -56
rect 4479 -73 4487 -56
rect 4913 -73 4921 -56
rect 5029 -73 5037 -56
rect 5463 -73 5471 -56
rect 5579 -73 5587 -56
rect 6013 -73 6021 -56
rect 6129 -73 6137 -56
rect 6563 -73 6571 -56
rect 6679 -73 6687 -56
rect 7113 -73 7121 -56
rect 7229 -73 7237 -56
rect 7663 -73 7671 -56
rect 7779 -73 7787 -56
rect 8213 -73 8221 -56
rect 8329 -73 8337 -56
rect 8763 -73 8771 -56
rect 8879 -73 8887 -56
rect 9313 -73 9321 -56
rect 9429 -73 9437 -56
rect 9863 -73 9871 -56
rect 9979 -73 9987 -56
rect 10413 -73 10421 -56
rect 10529 -73 10537 -56
rect 10963 -73 10971 -56
rect 11079 -73 11087 -56
rect 11513 -73 11521 -56
rect 11629 -73 11637 -56
rect 12063 -73 12071 -56
rect 12179 -73 12187 -56
rect 12613 -73 12621 -56
rect 12729 -73 12737 -56
rect 13163 -73 13171 -56
rect 13279 -73 13287 -56
rect 13713 -73 13721 -56
rect -477 -79 -23 -73
rect 79 -79 114 -73
rect -477 -87 -6 -79
rect -477 -135 -23 -87
rect -477 -465 -415 -135
rect -85 -465 -23 -135
rect -477 -513 -23 -465
rect -477 -521 -6 -513
rect 56 -87 114 -79
rect 73 -114 114 -87
rect 486 -79 521 -73
rect 623 -79 1077 -73
rect 1179 -79 1214 -73
rect 486 -87 544 -79
rect 486 -114 527 -87
rect 56 -521 73 -513
rect 527 -521 544 -513
rect 606 -87 1094 -79
rect 623 -135 1077 -87
rect 623 -465 685 -135
rect 1015 -465 1077 -135
rect 623 -513 1077 -465
rect 606 -521 1094 -513
rect 1156 -87 1214 -79
rect 1173 -114 1214 -87
rect 1586 -79 1621 -73
rect 1723 -79 2177 -73
rect 2279 -79 2314 -73
rect 1586 -87 1644 -79
rect 1586 -114 1627 -87
rect 1156 -521 1173 -513
rect 1627 -521 1644 -513
rect 1706 -87 2194 -79
rect 1723 -135 2177 -87
rect 1723 -465 1785 -135
rect 2115 -465 2177 -135
rect 1723 -513 2177 -465
rect 1706 -521 2194 -513
rect 2256 -87 2314 -79
rect 2273 -114 2314 -87
rect 2686 -79 2721 -73
rect 2823 -79 3277 -73
rect 3379 -79 3414 -73
rect 2686 -87 2744 -79
rect 2686 -114 2727 -87
rect 2256 -521 2273 -513
rect 2727 -521 2744 -513
rect 2806 -87 3294 -79
rect 2823 -135 3277 -87
rect 2823 -465 2885 -135
rect 3215 -465 3277 -135
rect 2823 -513 3277 -465
rect 2806 -521 3294 -513
rect 3356 -87 3414 -79
rect 3373 -114 3414 -87
rect 3786 -79 3821 -73
rect 3923 -79 4377 -73
rect 4479 -79 4514 -73
rect 3786 -87 3844 -79
rect 3786 -114 3827 -87
rect 3356 -521 3373 -513
rect 3827 -521 3844 -513
rect 3906 -87 4394 -79
rect 3923 -135 4377 -87
rect 3923 -465 3985 -135
rect 4315 -465 4377 -135
rect 3923 -513 4377 -465
rect 3906 -521 4394 -513
rect 4456 -87 4514 -79
rect 4473 -114 4514 -87
rect 4886 -79 4921 -73
rect 5023 -79 5477 -73
rect 5579 -79 5614 -73
rect 4886 -87 4944 -79
rect 4886 -114 4927 -87
rect 4456 -521 4473 -513
rect 4927 -521 4944 -513
rect 5006 -87 5494 -79
rect 5023 -135 5477 -87
rect 5023 -465 5085 -135
rect 5415 -465 5477 -135
rect 5023 -513 5477 -465
rect 5006 -521 5494 -513
rect 5556 -87 5614 -79
rect 5573 -114 5614 -87
rect 5986 -79 6021 -73
rect 6123 -79 6577 -73
rect 6679 -79 6714 -73
rect 5986 -87 6044 -79
rect 5986 -114 6027 -87
rect 5556 -521 5573 -513
rect 6027 -521 6044 -513
rect 6106 -87 6594 -79
rect 6123 -135 6577 -87
rect 6123 -465 6185 -135
rect 6515 -465 6577 -135
rect 6123 -513 6577 -465
rect 6106 -521 6594 -513
rect 6656 -87 6714 -79
rect 6673 -114 6714 -87
rect 7086 -79 7121 -73
rect 7223 -79 7677 -73
rect 7779 -79 7814 -73
rect 7086 -87 7144 -79
rect 7086 -114 7127 -87
rect 6656 -521 6673 -513
rect 7127 -521 7144 -513
rect 7206 -87 7694 -79
rect 7223 -135 7677 -87
rect 7223 -465 7285 -135
rect 7615 -465 7677 -135
rect 7223 -513 7677 -465
rect 7206 -521 7694 -513
rect 7756 -87 7814 -79
rect 7773 -114 7814 -87
rect 8186 -79 8221 -73
rect 8323 -79 8777 -73
rect 8879 -79 8914 -73
rect 8186 -87 8244 -79
rect 8186 -114 8227 -87
rect 7756 -521 7773 -513
rect 8227 -521 8244 -513
rect 8306 -87 8794 -79
rect 8323 -135 8777 -87
rect 8323 -465 8385 -135
rect 8715 -465 8777 -135
rect 8323 -513 8777 -465
rect 8306 -521 8794 -513
rect 8856 -87 8914 -79
rect 8873 -114 8914 -87
rect 9286 -79 9321 -73
rect 9423 -79 9877 -73
rect 9979 -79 10014 -73
rect 9286 -87 9344 -79
rect 9286 -114 9327 -87
rect 8856 -521 8873 -513
rect 9327 -521 9344 -513
rect 9406 -87 9894 -79
rect 9423 -135 9877 -87
rect 9423 -465 9485 -135
rect 9815 -465 9877 -135
rect 9423 -513 9877 -465
rect 9406 -521 9894 -513
rect 9956 -87 10014 -79
rect 9973 -114 10014 -87
rect 10386 -79 10421 -73
rect 10523 -79 10977 -73
rect 11079 -79 11114 -73
rect 10386 -87 10444 -79
rect 10386 -114 10427 -87
rect 9956 -521 9973 -513
rect 10427 -521 10444 -513
rect 10506 -87 10994 -79
rect 10523 -135 10977 -87
rect 10523 -465 10585 -135
rect 10915 -465 10977 -135
rect 10523 -513 10977 -465
rect 10506 -521 10994 -513
rect 11056 -87 11114 -79
rect 11073 -114 11114 -87
rect 11486 -79 11521 -73
rect 11623 -79 12077 -73
rect 12179 -79 12214 -73
rect 11486 -87 11544 -79
rect 11486 -114 11527 -87
rect 11056 -521 11073 -513
rect 11527 -521 11544 -513
rect 11606 -87 12094 -79
rect 11623 -135 12077 -87
rect 11623 -465 11685 -135
rect 12015 -465 12077 -135
rect 11623 -513 12077 -465
rect 11606 -521 12094 -513
rect 12156 -87 12214 -79
rect 12173 -114 12214 -87
rect 12586 -79 12621 -73
rect 12723 -79 13177 -73
rect 13279 -79 13314 -73
rect 12586 -87 12644 -79
rect 12586 -114 12627 -87
rect 12156 -521 12173 -513
rect 12627 -521 12644 -513
rect 12706 -87 13194 -79
rect 12723 -135 13177 -87
rect 12723 -465 12785 -135
rect 13115 -465 13177 -135
rect 12723 -513 13177 -465
rect 12706 -521 13194 -513
rect 13256 -87 13314 -79
rect 13273 -114 13314 -87
rect 13256 -521 13273 -513
rect -477 -527 -23 -521
rect 623 -527 1077 -521
rect 1723 -527 2177 -521
rect 2823 -527 3277 -521
rect 3923 -527 4377 -521
rect 5023 -527 5477 -521
rect 6123 -527 6577 -521
rect 7223 -527 7677 -521
rect 8323 -527 8777 -521
rect 9423 -527 9877 -521
rect 10523 -527 10977 -521
rect 11623 -527 12077 -521
rect 12723 -527 13177 -521
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 0 -558 50 -550
rect 0 -592 8 -558
rect 42 -592 50 -558
rect 0 -600 50 -592
rect 550 -558 600 -550
rect 550 -592 558 -558
rect 592 -592 600 -558
rect 550 -600 600 -592
rect 1100 -558 1150 -550
rect 1100 -592 1108 -558
rect 1142 -592 1150 -558
rect 1100 -600 1150 -592
rect 1650 -558 1700 -550
rect 1650 -592 1658 -558
rect 1692 -592 1700 -558
rect 1650 -600 1700 -592
rect 2200 -558 2250 -550
rect 2200 -592 2208 -558
rect 2242 -592 2250 -558
rect 2200 -600 2250 -592
rect 2750 -558 2800 -550
rect 2750 -592 2758 -558
rect 2792 -592 2800 -558
rect 2750 -600 2800 -592
rect 3300 -558 3350 -550
rect 3300 -592 3308 -558
rect 3342 -592 3350 -558
rect 3300 -600 3350 -592
rect 3850 -558 3900 -550
rect 3850 -592 3858 -558
rect 3892 -592 3900 -558
rect 3850 -600 3900 -592
rect 4400 -558 4450 -550
rect 4400 -592 4408 -558
rect 4442 -592 4450 -558
rect 4400 -600 4450 -592
rect 4950 -558 5000 -550
rect 4950 -592 4958 -558
rect 4992 -592 5000 -558
rect 4950 -600 5000 -592
rect 5500 -558 5550 -550
rect 5500 -592 5508 -558
rect 5542 -592 5550 -558
rect 5500 -600 5550 -592
rect 6050 -558 6100 -550
rect 6050 -592 6058 -558
rect 6092 -592 6100 -558
rect 6050 -600 6100 -592
rect 6600 -558 6650 -550
rect 6600 -592 6608 -558
rect 6642 -592 6650 -558
rect 6600 -600 6650 -592
rect 7150 -558 7200 -550
rect 7150 -592 7158 -558
rect 7192 -592 7200 -558
rect 7150 -600 7200 -592
rect 7700 -558 7750 -550
rect 7700 -592 7708 -558
rect 7742 -592 7750 -558
rect 7700 -600 7750 -592
rect 8250 -558 8300 -550
rect 8250 -592 8258 -558
rect 8292 -592 8300 -558
rect 8250 -600 8300 -592
rect 8800 -558 8850 -550
rect 8800 -592 8808 -558
rect 8842 -592 8850 -558
rect 8800 -600 8850 -592
rect 9350 -558 9400 -550
rect 9350 -592 9358 -558
rect 9392 -592 9400 -558
rect 9350 -600 9400 -592
rect 9900 -558 9950 -550
rect 9900 -592 9908 -558
rect 9942 -592 9950 -558
rect 9900 -600 9950 -592
rect 10450 -558 10500 -550
rect 10450 -592 10458 -558
rect 10492 -592 10500 -558
rect 10450 -600 10500 -592
rect 11000 -558 11050 -550
rect 11000 -592 11008 -558
rect 11042 -592 11050 -558
rect 11000 -600 11050 -592
rect 11550 -558 11600 -550
rect 11550 -592 11558 -558
rect 11592 -592 11600 -558
rect 11550 -600 11600 -592
rect 12100 -558 12150 -550
rect 12100 -592 12108 -558
rect 12142 -592 12150 -558
rect 12100 -600 12150 -592
rect 12650 -558 12700 -550
rect 12650 -592 12658 -558
rect 12692 -592 12700 -558
rect 12650 -600 12700 -592
rect 13200 -558 13250 -550
rect 13200 -592 13208 -558
rect 13242 -592 13250 -558
rect 13200 -600 13250 -592
rect 13750 -558 13800 -550
rect 13750 -592 13758 -558
rect 13792 -592 13800 -558
rect 13750 -600 13800 -592
rect 13975 -775 13987 0
rect -737 -787 13987 -775
rect -17 -1063 0 -787
rect 531 -1063 550 -787
rect 1083 -1063 1100 -787
rect 1631 -1063 1650 -787
rect 2183 -1063 2200 -787
rect 2731 -1063 2750 -787
rect 3283 -1063 3300 -787
rect 3831 -1063 3850 -787
rect 4383 -1063 4400 -787
rect 4931 -1063 4950 -787
rect 5483 -1063 5500 -787
rect 6031 -1063 6050 -787
rect 6583 -1063 6600 -787
rect 7131 -1063 7150 -787
rect 7683 -1063 7700 -787
rect 8231 -1063 8250 -787
rect 8783 -1063 8800 -787
rect 9331 -1063 9350 -787
rect 9883 -1063 9900 -787
rect 10431 -1063 10450 -787
rect 10983 -1063 11000 -787
rect 11531 -1063 11550 -787
rect 12083 -1063 12100 -787
rect 12631 -1063 12650 -787
rect 13183 -1063 13200 -787
rect 14263 -1063 14275 0
rect -1025 -1075 14275 -1063
rect 14775 -1575 14787 14725
rect -1537 -1587 14787 -1575
rect 18763 -5563 18775 18713
rect -5525 -5575 18775 -5563
<< viali >>
rect -5513 14737 18763 18713
rect -5513 -1587 -1537 14737
rect -1013 13937 -19 14213
rect 0 13937 531 14213
rect 550 13937 1081 14213
rect 1100 13937 1631 14213
rect 1650 13937 2181 14213
rect 2200 13937 2731 14213
rect 2750 13937 3281 14213
rect 3300 13937 3831 14213
rect 3850 13937 4381 14213
rect 4400 13937 4931 14213
rect 4950 13937 5481 14213
rect 5500 13937 6031 14213
rect 6050 13937 6581 14213
rect 6600 13937 7131 14213
rect 7150 13937 7681 14213
rect 7700 13937 8231 14213
rect 8250 13937 8781 14213
rect 8800 13937 9331 14213
rect 9350 13937 9881 14213
rect 9900 13937 10431 14213
rect 10450 13937 10981 14213
rect 11000 13937 11531 14213
rect 11550 13937 12081 14213
rect 12100 13937 12631 14213
rect 12650 13937 13181 14213
rect 13200 13937 14263 14213
rect -1013 13219 -737 13937
rect -542 13708 -508 13742
rect 8 13708 42 13742
rect 558 13708 592 13742
rect 1108 13708 1142 13742
rect 1658 13708 1692 13742
rect 2208 13708 2242 13742
rect 2758 13708 2792 13742
rect 3308 13708 3342 13742
rect 3858 13708 3892 13742
rect 4408 13708 4442 13742
rect 4958 13708 4992 13742
rect 5508 13708 5542 13742
rect 6058 13708 6092 13742
rect 6608 13708 6642 13742
rect 7158 13708 7192 13742
rect 7708 13708 7742 13742
rect 8258 13708 8292 13742
rect 8808 13708 8842 13742
rect 9358 13708 9392 13742
rect 9908 13708 9942 13742
rect 10458 13708 10492 13742
rect 11008 13708 11042 13742
rect 11558 13708 11592 13742
rect 12108 13708 12142 13742
rect 12658 13708 12692 13742
rect 13208 13708 13242 13742
rect 13758 13708 13792 13742
rect -23 13237 -6 13663
rect 56 13237 73 13663
rect 135 13603 465 13615
rect 135 13297 147 13603
rect 147 13297 453 13603
rect 453 13297 465 13603
rect 135 13285 465 13297
rect 527 13237 544 13663
rect 606 13237 623 13663
rect 1077 13237 1094 13663
rect 1156 13237 1173 13663
rect 1235 13603 1565 13615
rect 1235 13297 1247 13603
rect 1247 13297 1553 13603
rect 1553 13297 1565 13603
rect 1235 13285 1565 13297
rect 1627 13237 1644 13663
rect 1706 13237 1723 13663
rect 2177 13237 2194 13663
rect 2256 13237 2273 13663
rect 2335 13603 2665 13615
rect 2335 13297 2347 13603
rect 2347 13297 2653 13603
rect 2653 13297 2665 13603
rect 2335 13285 2665 13297
rect 2727 13237 2744 13663
rect 2806 13237 2823 13663
rect 3277 13237 3294 13663
rect 3356 13237 3373 13663
rect 3435 13603 3765 13615
rect 3435 13297 3447 13603
rect 3447 13297 3753 13603
rect 3753 13297 3765 13603
rect 3435 13285 3765 13297
rect 3827 13237 3844 13663
rect 3906 13237 3923 13663
rect 4377 13237 4394 13663
rect 4456 13237 4473 13663
rect 4535 13603 4865 13615
rect 4535 13297 4547 13603
rect 4547 13297 4853 13603
rect 4853 13297 4865 13603
rect 4535 13285 4865 13297
rect 4927 13237 4944 13663
rect 5006 13237 5023 13663
rect 5477 13237 5494 13663
rect 5556 13237 5573 13663
rect 5635 13603 5965 13615
rect 5635 13297 5647 13603
rect 5647 13297 5953 13603
rect 5953 13297 5965 13603
rect 5635 13285 5965 13297
rect 6027 13237 6044 13663
rect 6106 13237 6123 13663
rect 6577 13237 6594 13663
rect 6656 13237 6673 13663
rect 6735 13603 7065 13615
rect 6735 13297 6747 13603
rect 6747 13297 7053 13603
rect 7053 13297 7065 13603
rect 6735 13285 7065 13297
rect 7127 13237 7144 13663
rect 7206 13237 7223 13663
rect 7677 13237 7694 13663
rect 7756 13237 7773 13663
rect 7835 13603 8165 13615
rect 7835 13297 7847 13603
rect 7847 13297 8153 13603
rect 8153 13297 8165 13603
rect 7835 13285 8165 13297
rect 8227 13237 8244 13663
rect 8306 13237 8323 13663
rect 8777 13237 8794 13663
rect 8856 13237 8873 13663
rect 8935 13603 9265 13615
rect 8935 13297 8947 13603
rect 8947 13297 9253 13603
rect 9253 13297 9265 13603
rect 8935 13285 9265 13297
rect 9327 13237 9344 13663
rect 9406 13237 9423 13663
rect 9877 13237 9894 13663
rect 9956 13237 9973 13663
rect 10035 13603 10365 13615
rect 10035 13297 10047 13603
rect 10047 13297 10353 13603
rect 10353 13297 10365 13603
rect 10035 13285 10365 13297
rect 10427 13237 10444 13663
rect 10506 13237 10523 13663
rect 10977 13237 10994 13663
rect 11056 13237 11073 13663
rect 11135 13603 11465 13615
rect 11135 13297 11147 13603
rect 11147 13297 11453 13603
rect 11453 13297 11465 13603
rect 11135 13285 11465 13297
rect 11527 13237 11544 13663
rect 11606 13237 11623 13663
rect 12077 13237 12094 13663
rect 12156 13237 12173 13663
rect 12235 13603 12565 13615
rect 12235 13297 12247 13603
rect 12247 13297 12553 13603
rect 12553 13297 12565 13603
rect 12235 13285 12565 13297
rect 12627 13237 12644 13663
rect 12706 13237 12723 13663
rect 13177 13237 13194 13663
rect 13256 13237 13273 13663
rect 13335 13603 13665 13615
rect 13335 13297 13347 13603
rect 13347 13297 13653 13603
rect 13653 13297 13665 13603
rect 13335 13285 13665 13297
rect -463 13206 -37 13223
rect 87 13206 513 13223
rect 637 13206 1063 13223
rect 1187 13206 1613 13223
rect 1737 13206 2163 13223
rect 2287 13206 2713 13223
rect 2837 13206 3263 13223
rect 3387 13206 3813 13223
rect 3937 13206 4363 13223
rect 4487 13206 4913 13223
rect 5037 13206 5463 13223
rect 5587 13206 6013 13223
rect 6137 13206 6563 13223
rect 6687 13206 7113 13223
rect 7237 13206 7663 13223
rect 7787 13206 8213 13223
rect 8337 13206 8763 13223
rect 8887 13206 9313 13223
rect 9437 13206 9863 13223
rect 9987 13206 10413 13223
rect 10537 13206 10963 13223
rect 11087 13206 11513 13223
rect 11637 13206 12063 13223
rect 12187 13206 12613 13223
rect 12737 13206 13163 13223
rect 13287 13206 13713 13223
rect 13987 13219 14263 13937
rect -1013 12669 -737 13200
rect -542 13158 -508 13192
rect 8 13158 42 13192
rect 558 13158 592 13192
rect 1108 13158 1142 13192
rect 1658 13158 1692 13192
rect 2208 13158 2242 13192
rect 2758 13158 2792 13192
rect 3308 13158 3342 13192
rect 3858 13158 3892 13192
rect 4408 13158 4442 13192
rect 4958 13158 4992 13192
rect 5508 13158 5542 13192
rect 6058 13158 6092 13192
rect 6608 13158 6642 13192
rect 7158 13158 7192 13192
rect 7708 13158 7742 13192
rect 8258 13158 8292 13192
rect 8808 13158 8842 13192
rect 9358 13158 9392 13192
rect 9908 13158 9942 13192
rect 10458 13158 10492 13192
rect 11008 13158 11042 13192
rect 11558 13158 11592 13192
rect 12108 13158 12142 13192
rect 12658 13158 12692 13192
rect 13208 13158 13242 13192
rect 13758 13158 13792 13192
rect -463 13127 -37 13144
rect 87 13127 513 13144
rect 637 13127 1063 13144
rect 1187 13127 1613 13144
rect 1737 13127 2163 13144
rect 2287 13127 2713 13144
rect 2837 13127 3263 13144
rect 3387 13127 3813 13144
rect 3937 13127 4363 13144
rect 4487 13127 4913 13144
rect 5037 13127 5463 13144
rect 5587 13127 6013 13144
rect 6137 13127 6563 13144
rect 6687 13127 7113 13144
rect 7237 13127 7663 13144
rect 7787 13127 8213 13144
rect 8337 13127 8763 13144
rect 8887 13127 9313 13144
rect 9437 13127 9863 13144
rect 9987 13127 10413 13144
rect 10537 13127 10963 13144
rect 11087 13127 11513 13144
rect 11637 13127 12063 13144
rect 12187 13127 12613 13144
rect 12737 13127 13163 13144
rect 13287 13127 13713 13144
rect -415 13053 -85 13065
rect -415 12747 -403 13053
rect -403 12747 -97 13053
rect -97 12747 -85 13053
rect -415 12735 -85 12747
rect -23 12687 -6 13113
rect 56 12687 73 13113
rect 527 12687 544 13113
rect 606 12687 623 13113
rect 685 13053 1015 13065
rect 685 12747 697 13053
rect 697 12747 1003 13053
rect 1003 12747 1015 13053
rect 685 12735 1015 12747
rect 1077 12687 1094 13113
rect 1156 12687 1173 13113
rect 1627 12687 1644 13113
rect 1706 12687 1723 13113
rect 1785 13053 2115 13065
rect 1785 12747 1797 13053
rect 1797 12747 2103 13053
rect 2103 12747 2115 13053
rect 1785 12735 2115 12747
rect 2177 12687 2194 13113
rect 2256 12687 2273 13113
rect 2727 12687 2744 13113
rect 2806 12687 2823 13113
rect 2885 13053 3215 13065
rect 2885 12747 2897 13053
rect 2897 12747 3203 13053
rect 3203 12747 3215 13053
rect 2885 12735 3215 12747
rect 3277 12687 3294 13113
rect 3356 12687 3373 13113
rect 3827 12687 3844 13113
rect 3906 12687 3923 13113
rect 3985 13053 4315 13065
rect 3985 12747 3997 13053
rect 3997 12747 4303 13053
rect 4303 12747 4315 13053
rect 3985 12735 4315 12747
rect 4377 12687 4394 13113
rect 4456 12687 4473 13113
rect 4927 12687 4944 13113
rect 5006 12687 5023 13113
rect 5085 13053 5415 13065
rect 5085 12747 5097 13053
rect 5097 12747 5403 13053
rect 5403 12747 5415 13053
rect 5085 12735 5415 12747
rect 5477 12687 5494 13113
rect 5556 12687 5573 13113
rect 6027 12687 6044 13113
rect 6106 12687 6123 13113
rect 6185 13053 6515 13065
rect 6185 12747 6197 13053
rect 6197 12747 6503 13053
rect 6503 12747 6515 13053
rect 6185 12735 6515 12747
rect 6577 12687 6594 13113
rect 6656 12687 6673 13113
rect 7127 12687 7144 13113
rect 7206 12687 7223 13113
rect 7285 13053 7615 13065
rect 7285 12747 7297 13053
rect 7297 12747 7603 13053
rect 7603 12747 7615 13053
rect 7285 12735 7615 12747
rect 7677 12687 7694 13113
rect 7756 12687 7773 13113
rect 8227 12687 8244 13113
rect 8306 12687 8323 13113
rect 8385 13053 8715 13065
rect 8385 12747 8397 13053
rect 8397 12747 8703 13053
rect 8703 12747 8715 13053
rect 8385 12735 8715 12747
rect 8777 12687 8794 13113
rect 8856 12687 8873 13113
rect 9327 12687 9344 13113
rect 9406 12687 9423 13113
rect 9485 13053 9815 13065
rect 9485 12747 9497 13053
rect 9497 12747 9803 13053
rect 9803 12747 9815 13053
rect 9485 12735 9815 12747
rect 9877 12687 9894 13113
rect 9956 12687 9973 13113
rect 10427 12687 10444 13113
rect 10506 12687 10523 13113
rect 10585 13053 10915 13065
rect 10585 12747 10597 13053
rect 10597 12747 10903 13053
rect 10903 12747 10915 13053
rect 10585 12735 10915 12747
rect 10977 12687 10994 13113
rect 11056 12687 11073 13113
rect 11527 12687 11544 13113
rect 11606 12687 11623 13113
rect 11685 13053 12015 13065
rect 11685 12747 11697 13053
rect 11697 12747 12003 13053
rect 12003 12747 12015 13053
rect 11685 12735 12015 12747
rect 12077 12687 12094 13113
rect 12156 12687 12173 13113
rect 12627 12687 12644 13113
rect 12706 12687 12723 13113
rect 12785 13053 13115 13065
rect 12785 12747 12797 13053
rect 12797 12747 13103 13053
rect 13103 12747 13115 13053
rect 12785 12735 13115 12747
rect 13177 12687 13194 13113
rect 13256 12687 13273 13113
rect -463 12656 -37 12673
rect 87 12656 513 12673
rect 637 12656 1063 12673
rect 1187 12656 1613 12673
rect 1737 12656 2163 12673
rect 2287 12656 2713 12673
rect 2837 12656 3263 12673
rect 3387 12656 3813 12673
rect 3937 12656 4363 12673
rect 4487 12656 4913 12673
rect 5037 12656 5463 12673
rect 5587 12656 6013 12673
rect 6137 12656 6563 12673
rect 6687 12656 7113 12673
rect 7237 12656 7663 12673
rect 7787 12656 8213 12673
rect 8337 12656 8763 12673
rect 8887 12656 9313 12673
rect 9437 12656 9863 12673
rect 9987 12656 10413 12673
rect 10537 12656 10963 12673
rect 11087 12656 11513 12673
rect 11637 12656 12063 12673
rect 12187 12656 12613 12673
rect 12737 12656 13163 12673
rect 13287 12656 13713 12673
rect 13987 12669 14263 13200
rect -1013 12119 -737 12650
rect -542 12608 -508 12642
rect 8 12608 42 12642
rect 558 12608 592 12642
rect 1108 12608 1142 12642
rect 1658 12608 1692 12642
rect 2208 12608 2242 12642
rect 2758 12608 2792 12642
rect 3308 12608 3342 12642
rect 3858 12608 3892 12642
rect 4408 12608 4442 12642
rect 4958 12608 4992 12642
rect 5508 12608 5542 12642
rect 6058 12608 6092 12642
rect 6608 12608 6642 12642
rect 7158 12608 7192 12642
rect 7708 12608 7742 12642
rect 8258 12608 8292 12642
rect 8808 12608 8842 12642
rect 9358 12608 9392 12642
rect 9908 12608 9942 12642
rect 10458 12608 10492 12642
rect 11008 12608 11042 12642
rect 11558 12608 11592 12642
rect 12108 12608 12142 12642
rect 12658 12608 12692 12642
rect 13208 12608 13242 12642
rect 13758 12608 13792 12642
rect -463 12577 -37 12594
rect 87 12577 513 12594
rect 637 12577 1063 12594
rect 1187 12577 1613 12594
rect 1737 12577 2163 12594
rect 2287 12577 2713 12594
rect 2837 12577 3263 12594
rect 3387 12577 3813 12594
rect 3937 12577 4363 12594
rect 4487 12577 4913 12594
rect 5037 12577 5463 12594
rect 5587 12577 6013 12594
rect 6137 12577 6563 12594
rect 6687 12577 7113 12594
rect 7237 12577 7663 12594
rect 7787 12577 8213 12594
rect 8337 12577 8763 12594
rect 8887 12577 9313 12594
rect 9437 12577 9863 12594
rect 9987 12577 10413 12594
rect 10537 12577 10963 12594
rect 11087 12577 11513 12594
rect 11637 12577 12063 12594
rect 12187 12577 12613 12594
rect 12737 12577 13163 12594
rect 13287 12577 13713 12594
rect -23 12137 -6 12563
rect 56 12137 73 12563
rect 135 12503 465 12515
rect 135 12197 147 12503
rect 147 12197 453 12503
rect 453 12197 465 12503
rect 135 12185 465 12197
rect 527 12137 544 12563
rect 606 12137 623 12563
rect 1077 12137 1094 12563
rect 1156 12137 1173 12563
rect 1235 12503 1565 12515
rect 1235 12197 1247 12503
rect 1247 12197 1553 12503
rect 1553 12197 1565 12503
rect 1235 12185 1565 12197
rect 1627 12137 1644 12563
rect 1706 12137 1723 12563
rect 2177 12137 2194 12563
rect 2256 12137 2273 12563
rect 2335 12503 2665 12515
rect 2335 12197 2347 12503
rect 2347 12197 2653 12503
rect 2653 12197 2665 12503
rect 2335 12185 2665 12197
rect 2727 12137 2744 12563
rect 2806 12137 2823 12563
rect 3277 12137 3294 12563
rect 3356 12137 3373 12563
rect 3435 12503 3765 12515
rect 3435 12197 3447 12503
rect 3447 12197 3753 12503
rect 3753 12197 3765 12503
rect 3435 12185 3765 12197
rect 3827 12137 3844 12563
rect 3906 12137 3923 12563
rect 4377 12137 4394 12563
rect 4456 12137 4473 12563
rect 4535 12503 4865 12515
rect 4535 12197 4547 12503
rect 4547 12197 4853 12503
rect 4853 12197 4865 12503
rect 4535 12185 4865 12197
rect 4927 12137 4944 12563
rect 5006 12137 5023 12563
rect 5477 12137 5494 12563
rect 5556 12137 5573 12563
rect 5635 12503 5965 12515
rect 5635 12197 5647 12503
rect 5647 12197 5953 12503
rect 5953 12197 5965 12503
rect 5635 12185 5965 12197
rect 6027 12137 6044 12563
rect 6106 12137 6123 12563
rect 6577 12137 6594 12563
rect 6656 12137 6673 12563
rect 6735 12503 7065 12515
rect 6735 12197 6747 12503
rect 6747 12197 7053 12503
rect 7053 12197 7065 12503
rect 6735 12185 7065 12197
rect 7127 12137 7144 12563
rect 7206 12137 7223 12563
rect 7677 12137 7694 12563
rect 7756 12137 7773 12563
rect 7835 12503 8165 12515
rect 7835 12197 7847 12503
rect 7847 12197 8153 12503
rect 8153 12197 8165 12503
rect 7835 12185 8165 12197
rect 8227 12137 8244 12563
rect 8306 12137 8323 12563
rect 8777 12137 8794 12563
rect 8856 12137 8873 12563
rect 8935 12503 9265 12515
rect 8935 12197 8947 12503
rect 8947 12197 9253 12503
rect 9253 12197 9265 12503
rect 8935 12185 9265 12197
rect 9327 12137 9344 12563
rect 9406 12137 9423 12563
rect 9877 12137 9894 12563
rect 9956 12137 9973 12563
rect 10035 12503 10365 12515
rect 10035 12197 10047 12503
rect 10047 12197 10353 12503
rect 10353 12197 10365 12503
rect 10035 12185 10365 12197
rect 10427 12137 10444 12563
rect 10506 12137 10523 12563
rect 10977 12137 10994 12563
rect 11056 12137 11073 12563
rect 11135 12503 11465 12515
rect 11135 12197 11147 12503
rect 11147 12197 11453 12503
rect 11453 12197 11465 12503
rect 11135 12185 11465 12197
rect 11527 12137 11544 12563
rect 11606 12137 11623 12563
rect 12077 12137 12094 12563
rect 12156 12137 12173 12563
rect 12235 12503 12565 12515
rect 12235 12197 12247 12503
rect 12247 12197 12553 12503
rect 12553 12197 12565 12503
rect 12235 12185 12565 12197
rect 12627 12137 12644 12563
rect 12706 12137 12723 12563
rect 13177 12137 13194 12563
rect 13256 12137 13273 12563
rect 13335 12503 13665 12515
rect 13335 12197 13347 12503
rect 13347 12197 13653 12503
rect 13653 12197 13665 12503
rect 13335 12185 13665 12197
rect -463 12106 -37 12123
rect 87 12106 513 12123
rect 637 12106 1063 12123
rect 1187 12106 1613 12123
rect 1737 12106 2163 12123
rect 2287 12106 2713 12123
rect 2837 12106 3263 12123
rect 3387 12106 3813 12123
rect 3937 12106 4363 12123
rect 4487 12106 4913 12123
rect 5037 12106 5463 12123
rect 5587 12106 6013 12123
rect 6137 12106 6563 12123
rect 6687 12106 7113 12123
rect 7237 12106 7663 12123
rect 7787 12106 8213 12123
rect 8337 12106 8763 12123
rect 8887 12106 9313 12123
rect 9437 12106 9863 12123
rect 9987 12106 10413 12123
rect 10537 12106 10963 12123
rect 11087 12106 11513 12123
rect 11637 12106 12063 12123
rect 12187 12106 12613 12123
rect 12737 12106 13163 12123
rect 13287 12106 13713 12123
rect 13987 12119 14263 12650
rect -1013 11569 -737 12100
rect -542 12058 -508 12092
rect 8 12058 42 12092
rect 558 12058 592 12092
rect 1108 12058 1142 12092
rect 1658 12058 1692 12092
rect 2208 12058 2242 12092
rect 2758 12058 2792 12092
rect 3308 12058 3342 12092
rect 3858 12058 3892 12092
rect 4408 12058 4442 12092
rect 4958 12058 4992 12092
rect 5508 12058 5542 12092
rect 6058 12058 6092 12092
rect 6608 12058 6642 12092
rect 7158 12058 7192 12092
rect 7708 12058 7742 12092
rect 8258 12058 8292 12092
rect 8808 12058 8842 12092
rect 9358 12058 9392 12092
rect 9908 12058 9942 12092
rect 10458 12058 10492 12092
rect 11008 12058 11042 12092
rect 11558 12058 11592 12092
rect 12108 12058 12142 12092
rect 12658 12058 12692 12092
rect 13208 12058 13242 12092
rect 13758 12058 13792 12092
rect -463 12027 -37 12044
rect 87 12027 513 12044
rect 637 12027 1063 12044
rect 1187 12027 1613 12044
rect 1737 12027 2163 12044
rect 2287 12027 2713 12044
rect 2837 12027 3263 12044
rect 3387 12027 3813 12044
rect 3937 12027 4363 12044
rect 4487 12027 4913 12044
rect 5037 12027 5463 12044
rect 5587 12027 6013 12044
rect 6137 12027 6563 12044
rect 6687 12027 7113 12044
rect 7237 12027 7663 12044
rect 7787 12027 8213 12044
rect 8337 12027 8763 12044
rect 8887 12027 9313 12044
rect 9437 12027 9863 12044
rect 9987 12027 10413 12044
rect 10537 12027 10963 12044
rect 11087 12027 11513 12044
rect 11637 12027 12063 12044
rect 12187 12027 12613 12044
rect 12737 12027 13163 12044
rect 13287 12027 13713 12044
rect -415 11953 -85 11965
rect -415 11647 -403 11953
rect -403 11647 -97 11953
rect -97 11647 -85 11953
rect -415 11635 -85 11647
rect -23 11587 -6 12013
rect 56 11587 73 12013
rect 527 11587 544 12013
rect 606 11587 623 12013
rect 685 11953 1015 11965
rect 685 11647 697 11953
rect 697 11647 1003 11953
rect 1003 11647 1015 11953
rect 685 11635 1015 11647
rect 1077 11587 1094 12013
rect 1156 11587 1173 12013
rect 1627 11587 1644 12013
rect 1706 11587 1723 12013
rect 1785 11953 2115 11965
rect 1785 11647 1797 11953
rect 1797 11647 2103 11953
rect 2103 11647 2115 11953
rect 1785 11635 2115 11647
rect 2177 11587 2194 12013
rect 2256 11587 2273 12013
rect 2727 11587 2744 12013
rect 2806 11587 2823 12013
rect 2885 11953 3215 11965
rect 2885 11647 2897 11953
rect 2897 11647 3203 11953
rect 3203 11647 3215 11953
rect 2885 11635 3215 11647
rect 3277 11587 3294 12013
rect 3356 11587 3373 12013
rect 3827 11587 3844 12013
rect 3906 11587 3923 12013
rect 3985 11953 4315 11965
rect 3985 11647 3997 11953
rect 3997 11647 4303 11953
rect 4303 11647 4315 11953
rect 3985 11635 4315 11647
rect 4377 11587 4394 12013
rect 4456 11587 4473 12013
rect 4927 11587 4944 12013
rect 5006 11587 5023 12013
rect 5085 11953 5415 11965
rect 5085 11647 5097 11953
rect 5097 11647 5403 11953
rect 5403 11647 5415 11953
rect 5085 11635 5415 11647
rect 5477 11587 5494 12013
rect 5556 11587 5573 12013
rect 6027 11587 6044 12013
rect 6106 11587 6123 12013
rect 6185 11953 6515 11965
rect 6185 11647 6197 11953
rect 6197 11647 6503 11953
rect 6503 11647 6515 11953
rect 6185 11635 6515 11647
rect 6577 11587 6594 12013
rect 6656 11587 6673 12013
rect 7127 11587 7144 12013
rect 7206 11587 7223 12013
rect 7285 11953 7615 11965
rect 7285 11647 7297 11953
rect 7297 11647 7603 11953
rect 7603 11647 7615 11953
rect 7285 11635 7615 11647
rect 7677 11587 7694 12013
rect 7756 11587 7773 12013
rect 8227 11587 8244 12013
rect 8306 11587 8323 12013
rect 8385 11953 8715 11965
rect 8385 11647 8397 11953
rect 8397 11647 8703 11953
rect 8703 11647 8715 11953
rect 8385 11635 8715 11647
rect 8777 11587 8794 12013
rect 8856 11587 8873 12013
rect 9327 11587 9344 12013
rect 9406 11587 9423 12013
rect 9485 11953 9815 11965
rect 9485 11647 9497 11953
rect 9497 11647 9803 11953
rect 9803 11647 9815 11953
rect 9485 11635 9815 11647
rect 9877 11587 9894 12013
rect 9956 11587 9973 12013
rect 10427 11587 10444 12013
rect 10506 11587 10523 12013
rect 10585 11953 10915 11965
rect 10585 11647 10597 11953
rect 10597 11647 10903 11953
rect 10903 11647 10915 11953
rect 10585 11635 10915 11647
rect 10977 11587 10994 12013
rect 11056 11587 11073 12013
rect 11527 11587 11544 12013
rect 11606 11587 11623 12013
rect 11685 11953 12015 11965
rect 11685 11647 11697 11953
rect 11697 11647 12003 11953
rect 12003 11647 12015 11953
rect 11685 11635 12015 11647
rect 12077 11587 12094 12013
rect 12156 11587 12173 12013
rect 12627 11587 12644 12013
rect 12706 11587 12723 12013
rect 12785 11953 13115 11965
rect 12785 11647 12797 11953
rect 12797 11647 13103 11953
rect 13103 11647 13115 11953
rect 12785 11635 13115 11647
rect 13177 11587 13194 12013
rect 13256 11587 13273 12013
rect -463 11556 -37 11573
rect 87 11556 513 11573
rect 637 11556 1063 11573
rect 1187 11556 1613 11573
rect 1737 11556 2163 11573
rect 2287 11556 2713 11573
rect 2837 11556 3263 11573
rect 3387 11556 3813 11573
rect 3937 11556 4363 11573
rect 4487 11556 4913 11573
rect 5037 11556 5463 11573
rect 5587 11556 6013 11573
rect 6137 11556 6563 11573
rect 6687 11556 7113 11573
rect 7237 11556 7663 11573
rect 7787 11556 8213 11573
rect 8337 11556 8763 11573
rect 8887 11556 9313 11573
rect 9437 11556 9863 11573
rect 9987 11556 10413 11573
rect 10537 11556 10963 11573
rect 11087 11556 11513 11573
rect 11637 11556 12063 11573
rect 12187 11556 12613 11573
rect 12737 11556 13163 11573
rect 13287 11556 13713 11573
rect 13987 11569 14263 12100
rect -1013 11019 -737 11550
rect -542 11508 -508 11542
rect 8 11508 42 11542
rect 558 11508 592 11542
rect 1108 11508 1142 11542
rect 1658 11508 1692 11542
rect 2208 11508 2242 11542
rect 2758 11508 2792 11542
rect 3308 11508 3342 11542
rect 3858 11508 3892 11542
rect 4408 11508 4442 11542
rect 4958 11508 4992 11542
rect 5508 11508 5542 11542
rect 6058 11508 6092 11542
rect 6608 11508 6642 11542
rect 7158 11508 7192 11542
rect 7708 11508 7742 11542
rect 8258 11508 8292 11542
rect 8808 11508 8842 11542
rect 9358 11508 9392 11542
rect 9908 11508 9942 11542
rect 10458 11508 10492 11542
rect 11008 11508 11042 11542
rect 11558 11508 11592 11542
rect 12108 11508 12142 11542
rect 12658 11508 12692 11542
rect 13208 11508 13242 11542
rect 13758 11508 13792 11542
rect -463 11477 -37 11494
rect 87 11477 513 11494
rect 637 11477 1063 11494
rect 1187 11477 1613 11494
rect 1737 11477 2163 11494
rect 2287 11477 2713 11494
rect 2837 11477 3263 11494
rect 3387 11477 3813 11494
rect 3937 11477 4363 11494
rect 4487 11477 4913 11494
rect 5037 11477 5463 11494
rect 5587 11477 6013 11494
rect 6137 11477 6563 11494
rect 6687 11477 7113 11494
rect 7237 11477 7663 11494
rect 7787 11477 8213 11494
rect 8337 11477 8763 11494
rect 8887 11477 9313 11494
rect 9437 11477 9863 11494
rect 9987 11477 10413 11494
rect 10537 11477 10963 11494
rect 11087 11477 11513 11494
rect 11637 11477 12063 11494
rect 12187 11477 12613 11494
rect 12737 11477 13163 11494
rect 13287 11477 13713 11494
rect -23 11037 -6 11463
rect 56 11037 73 11463
rect 135 11403 465 11415
rect 135 11097 147 11403
rect 147 11097 453 11403
rect 453 11097 465 11403
rect 135 11085 465 11097
rect 527 11037 544 11463
rect 606 11037 623 11463
rect 1077 11037 1094 11463
rect 1156 11037 1173 11463
rect 1235 11403 1565 11415
rect 1235 11097 1247 11403
rect 1247 11097 1553 11403
rect 1553 11097 1565 11403
rect 1235 11085 1565 11097
rect 1627 11037 1644 11463
rect 1706 11037 1723 11463
rect 2177 11037 2194 11463
rect 2256 11037 2273 11463
rect 2335 11403 2665 11415
rect 2335 11097 2347 11403
rect 2347 11097 2653 11403
rect 2653 11097 2665 11403
rect 2335 11085 2665 11097
rect 2727 11037 2744 11463
rect 2806 11037 2823 11463
rect 3277 11037 3294 11463
rect 3356 11037 3373 11463
rect 3435 11403 3765 11415
rect 3435 11097 3447 11403
rect 3447 11097 3753 11403
rect 3753 11097 3765 11403
rect 3435 11085 3765 11097
rect 3827 11037 3844 11463
rect 3906 11037 3923 11463
rect 4377 11037 4394 11463
rect 4456 11037 4473 11463
rect 4535 11403 4865 11415
rect 4535 11097 4547 11403
rect 4547 11097 4853 11403
rect 4853 11097 4865 11403
rect 4535 11085 4865 11097
rect 4927 11037 4944 11463
rect 5006 11037 5023 11463
rect 5477 11037 5494 11463
rect 5556 11037 5573 11463
rect 5635 11403 5965 11415
rect 5635 11097 5647 11403
rect 5647 11097 5953 11403
rect 5953 11097 5965 11403
rect 5635 11085 5965 11097
rect 6027 11037 6044 11463
rect 6106 11037 6123 11463
rect 6577 11037 6594 11463
rect 6656 11037 6673 11463
rect 6735 11403 7065 11415
rect 6735 11097 6747 11403
rect 6747 11097 7053 11403
rect 7053 11097 7065 11403
rect 6735 11085 7065 11097
rect 7127 11037 7144 11463
rect 7206 11037 7223 11463
rect 7677 11037 7694 11463
rect 7756 11037 7773 11463
rect 7835 11403 8165 11415
rect 7835 11097 7847 11403
rect 7847 11097 8153 11403
rect 8153 11097 8165 11403
rect 7835 11085 8165 11097
rect 8227 11037 8244 11463
rect 8306 11037 8323 11463
rect 8777 11037 8794 11463
rect 8856 11037 8873 11463
rect 8935 11403 9265 11415
rect 8935 11097 8947 11403
rect 8947 11097 9253 11403
rect 9253 11097 9265 11403
rect 8935 11085 9265 11097
rect 9327 11037 9344 11463
rect 9406 11037 9423 11463
rect 9877 11037 9894 11463
rect 9956 11037 9973 11463
rect 10035 11403 10365 11415
rect 10035 11097 10047 11403
rect 10047 11097 10353 11403
rect 10353 11097 10365 11403
rect 10035 11085 10365 11097
rect 10427 11037 10444 11463
rect 10506 11037 10523 11463
rect 10977 11037 10994 11463
rect 11056 11037 11073 11463
rect 11135 11403 11465 11415
rect 11135 11097 11147 11403
rect 11147 11097 11453 11403
rect 11453 11097 11465 11403
rect 11135 11085 11465 11097
rect 11527 11037 11544 11463
rect 11606 11037 11623 11463
rect 12077 11037 12094 11463
rect 12156 11037 12173 11463
rect 12235 11403 12565 11415
rect 12235 11097 12247 11403
rect 12247 11097 12553 11403
rect 12553 11097 12565 11403
rect 12235 11085 12565 11097
rect 12627 11037 12644 11463
rect 12706 11037 12723 11463
rect 13177 11037 13194 11463
rect 13256 11037 13273 11463
rect 13335 11403 13665 11415
rect 13335 11097 13347 11403
rect 13347 11097 13653 11403
rect 13653 11097 13665 11403
rect 13335 11085 13665 11097
rect -463 11006 -37 11023
rect 87 11006 513 11023
rect 637 11006 1063 11023
rect 1187 11006 1613 11023
rect 1737 11006 2163 11023
rect 2287 11006 2713 11023
rect 2837 11006 3263 11023
rect 3387 11006 3813 11023
rect 3937 11006 4363 11023
rect 4487 11006 4913 11023
rect 5037 11006 5463 11023
rect 5587 11006 6013 11023
rect 6137 11006 6563 11023
rect 6687 11006 7113 11023
rect 7237 11006 7663 11023
rect 7787 11006 8213 11023
rect 8337 11006 8763 11023
rect 8887 11006 9313 11023
rect 9437 11006 9863 11023
rect 9987 11006 10413 11023
rect 10537 11006 10963 11023
rect 11087 11006 11513 11023
rect 11637 11006 12063 11023
rect 12187 11006 12613 11023
rect 12737 11006 13163 11023
rect 13287 11006 13713 11023
rect 13987 11019 14263 11550
rect -1013 10469 -737 11000
rect -542 10958 -508 10992
rect 8 10958 42 10992
rect 558 10958 592 10992
rect 1108 10958 1142 10992
rect 1658 10958 1692 10992
rect 2208 10958 2242 10992
rect 2758 10958 2792 10992
rect 3308 10958 3342 10992
rect 3858 10958 3892 10992
rect 4408 10958 4442 10992
rect 4958 10958 4992 10992
rect 5508 10958 5542 10992
rect 6058 10958 6092 10992
rect 6608 10958 6642 10992
rect 7158 10958 7192 10992
rect 7708 10958 7742 10992
rect 8258 10958 8292 10992
rect 8808 10958 8842 10992
rect 9358 10958 9392 10992
rect 9908 10958 9942 10992
rect 10458 10958 10492 10992
rect 11008 10958 11042 10992
rect 11558 10958 11592 10992
rect 12108 10958 12142 10992
rect 12658 10958 12692 10992
rect 13208 10958 13242 10992
rect 13758 10958 13792 10992
rect -463 10927 -37 10944
rect 87 10927 513 10944
rect 637 10927 1063 10944
rect 1187 10927 1613 10944
rect 1737 10927 2163 10944
rect 2287 10927 2713 10944
rect 2837 10927 3263 10944
rect 3387 10927 3813 10944
rect 3937 10927 4363 10944
rect 4487 10927 4913 10944
rect 5037 10927 5463 10944
rect 5587 10927 6013 10944
rect 6137 10927 6563 10944
rect 6687 10927 7113 10944
rect 7237 10927 7663 10944
rect 7787 10927 8213 10944
rect 8337 10927 8763 10944
rect 8887 10927 9313 10944
rect 9437 10927 9863 10944
rect 9987 10927 10413 10944
rect 10537 10927 10963 10944
rect 11087 10927 11513 10944
rect 11637 10927 12063 10944
rect 12187 10927 12613 10944
rect 12737 10927 13163 10944
rect 13287 10927 13713 10944
rect -415 10853 -85 10865
rect -415 10547 -403 10853
rect -403 10547 -97 10853
rect -97 10547 -85 10853
rect -415 10535 -85 10547
rect -23 10487 -6 10913
rect 56 10487 73 10913
rect 527 10487 544 10913
rect 606 10487 623 10913
rect 685 10853 1015 10865
rect 685 10547 697 10853
rect 697 10547 1003 10853
rect 1003 10547 1015 10853
rect 685 10535 1015 10547
rect 1077 10487 1094 10913
rect 1156 10487 1173 10913
rect 1627 10487 1644 10913
rect 1706 10487 1723 10913
rect 1785 10853 2115 10865
rect 1785 10547 1797 10853
rect 1797 10547 2103 10853
rect 2103 10547 2115 10853
rect 1785 10535 2115 10547
rect 2177 10487 2194 10913
rect 2256 10487 2273 10913
rect 2727 10487 2744 10913
rect 2806 10487 2823 10913
rect 2885 10853 3215 10865
rect 2885 10547 2897 10853
rect 2897 10547 3203 10853
rect 3203 10547 3215 10853
rect 2885 10535 3215 10547
rect 3277 10487 3294 10913
rect 3356 10487 3373 10913
rect 3827 10487 3844 10913
rect 3906 10487 3923 10913
rect 3985 10853 4315 10865
rect 3985 10547 3997 10853
rect 3997 10547 4303 10853
rect 4303 10547 4315 10853
rect 3985 10535 4315 10547
rect 4377 10487 4394 10913
rect 4456 10487 4473 10913
rect 4927 10487 4944 10913
rect 5006 10487 5023 10913
rect 5085 10853 5415 10865
rect 5085 10547 5097 10853
rect 5097 10547 5403 10853
rect 5403 10547 5415 10853
rect 5085 10535 5415 10547
rect 5477 10487 5494 10913
rect 5556 10487 5573 10913
rect 6027 10487 6044 10913
rect 6106 10487 6123 10913
rect 6185 10853 6515 10865
rect 6185 10547 6197 10853
rect 6197 10547 6503 10853
rect 6503 10547 6515 10853
rect 6185 10535 6515 10547
rect 6577 10487 6594 10913
rect 6656 10487 6673 10913
rect 7127 10487 7144 10913
rect 7206 10487 7223 10913
rect 7285 10853 7615 10865
rect 7285 10547 7297 10853
rect 7297 10547 7603 10853
rect 7603 10547 7615 10853
rect 7285 10535 7615 10547
rect 7677 10487 7694 10913
rect 7756 10487 7773 10913
rect 8227 10487 8244 10913
rect 8306 10487 8323 10913
rect 8385 10853 8715 10865
rect 8385 10547 8397 10853
rect 8397 10547 8703 10853
rect 8703 10547 8715 10853
rect 8385 10535 8715 10547
rect 8777 10487 8794 10913
rect 8856 10487 8873 10913
rect 9327 10487 9344 10913
rect 9406 10487 9423 10913
rect 9485 10853 9815 10865
rect 9485 10547 9497 10853
rect 9497 10547 9803 10853
rect 9803 10547 9815 10853
rect 9485 10535 9815 10547
rect 9877 10487 9894 10913
rect 9956 10487 9973 10913
rect 10427 10487 10444 10913
rect 10506 10487 10523 10913
rect 10585 10853 10915 10865
rect 10585 10547 10597 10853
rect 10597 10547 10903 10853
rect 10903 10547 10915 10853
rect 10585 10535 10915 10547
rect 10977 10487 10994 10913
rect 11056 10487 11073 10913
rect 11527 10487 11544 10913
rect 11606 10487 11623 10913
rect 11685 10853 12015 10865
rect 11685 10547 11697 10853
rect 11697 10547 12003 10853
rect 12003 10547 12015 10853
rect 11685 10535 12015 10547
rect 12077 10487 12094 10913
rect 12156 10487 12173 10913
rect 12627 10487 12644 10913
rect 12706 10487 12723 10913
rect 12785 10853 13115 10865
rect 12785 10547 12797 10853
rect 12797 10547 13103 10853
rect 13103 10547 13115 10853
rect 12785 10535 13115 10547
rect 13177 10487 13194 10913
rect 13256 10487 13273 10913
rect -463 10456 -37 10473
rect 87 10456 513 10473
rect 637 10456 1063 10473
rect 1187 10456 1613 10473
rect 1737 10456 2163 10473
rect 2287 10456 2713 10473
rect 2837 10456 3263 10473
rect 3387 10456 3813 10473
rect 3937 10456 4363 10473
rect 4487 10456 4913 10473
rect 5037 10456 5463 10473
rect 5587 10456 6013 10473
rect 6137 10456 6563 10473
rect 6687 10456 7113 10473
rect 7237 10456 7663 10473
rect 7787 10456 8213 10473
rect 8337 10456 8763 10473
rect 8887 10456 9313 10473
rect 9437 10456 9863 10473
rect 9987 10456 10413 10473
rect 10537 10456 10963 10473
rect 11087 10456 11513 10473
rect 11637 10456 12063 10473
rect 12187 10456 12613 10473
rect 12737 10456 13163 10473
rect 13287 10456 13713 10473
rect 13987 10469 14263 11000
rect -1013 9919 -737 10450
rect -542 10408 -508 10442
rect 8 10408 42 10442
rect 558 10408 592 10442
rect 1108 10408 1142 10442
rect 1658 10408 1692 10442
rect 2208 10408 2242 10442
rect 2758 10408 2792 10442
rect 3308 10408 3342 10442
rect 3858 10408 3892 10442
rect 4408 10408 4442 10442
rect 4958 10408 4992 10442
rect 5508 10408 5542 10442
rect 6058 10408 6092 10442
rect 6608 10408 6642 10442
rect 7158 10408 7192 10442
rect 7708 10408 7742 10442
rect 8258 10408 8292 10442
rect 8808 10408 8842 10442
rect 9358 10408 9392 10442
rect 9908 10408 9942 10442
rect 10458 10408 10492 10442
rect 11008 10408 11042 10442
rect 11558 10408 11592 10442
rect 12108 10408 12142 10442
rect 12658 10408 12692 10442
rect 13208 10408 13242 10442
rect 13758 10408 13792 10442
rect -463 10377 -37 10394
rect 87 10377 513 10394
rect 637 10377 1063 10394
rect 1187 10377 1613 10394
rect 1737 10377 2163 10394
rect 2287 10377 2713 10394
rect 2837 10377 3263 10394
rect 3387 10377 3813 10394
rect 3937 10377 4363 10394
rect 4487 10377 4913 10394
rect 5037 10377 5463 10394
rect 5587 10377 6013 10394
rect 6137 10377 6563 10394
rect 6687 10377 7113 10394
rect 7237 10377 7663 10394
rect 7787 10377 8213 10394
rect 8337 10377 8763 10394
rect 8887 10377 9313 10394
rect 9437 10377 9863 10394
rect 9987 10377 10413 10394
rect 10537 10377 10963 10394
rect 11087 10377 11513 10394
rect 11637 10377 12063 10394
rect 12187 10377 12613 10394
rect 12737 10377 13163 10394
rect 13287 10377 13713 10394
rect -23 9937 -6 10363
rect 56 9937 73 10363
rect 135 10303 465 10315
rect 135 9997 147 10303
rect 147 9997 453 10303
rect 453 9997 465 10303
rect 135 9985 465 9997
rect 527 9937 544 10363
rect 606 9937 623 10363
rect 1077 9937 1094 10363
rect 1156 9937 1173 10363
rect 1235 10303 1565 10315
rect 1235 9997 1247 10303
rect 1247 9997 1553 10303
rect 1553 9997 1565 10303
rect 1235 9985 1565 9997
rect 1627 9937 1644 10363
rect 1706 9937 1723 10363
rect 2177 9937 2194 10363
rect 2256 9937 2273 10363
rect 2335 10303 2665 10315
rect 2335 9997 2347 10303
rect 2347 9997 2653 10303
rect 2653 9997 2665 10303
rect 2335 9985 2665 9997
rect 2727 9937 2744 10363
rect 2806 9937 2823 10363
rect 3277 9937 3294 10363
rect 3356 9937 3373 10363
rect 3435 10303 3765 10315
rect 3435 9997 3447 10303
rect 3447 9997 3753 10303
rect 3753 9997 3765 10303
rect 3435 9985 3765 9997
rect 3827 9937 3844 10363
rect 3906 9937 3923 10363
rect 4377 9937 4394 10363
rect 4456 9937 4473 10363
rect 4535 10303 4865 10315
rect 4535 9997 4547 10303
rect 4547 9997 4853 10303
rect 4853 9997 4865 10303
rect 4535 9985 4865 9997
rect 4927 9937 4944 10363
rect 5006 9937 5023 10363
rect 5477 9937 5494 10363
rect 5556 9937 5573 10363
rect 5635 10303 5965 10315
rect 5635 9997 5647 10303
rect 5647 9997 5953 10303
rect 5953 9997 5965 10303
rect 5635 9985 5965 9997
rect 6027 9937 6044 10363
rect 6106 9937 6123 10363
rect 6577 9937 6594 10363
rect 6656 9937 6673 10363
rect 6735 10303 7065 10315
rect 6735 9997 6747 10303
rect 6747 9997 7053 10303
rect 7053 9997 7065 10303
rect 6735 9985 7065 9997
rect 7127 9937 7144 10363
rect 7206 9937 7223 10363
rect 7677 9937 7694 10363
rect 7756 9937 7773 10363
rect 7835 10303 8165 10315
rect 7835 9997 7847 10303
rect 7847 9997 8153 10303
rect 8153 9997 8165 10303
rect 7835 9985 8165 9997
rect 8227 9937 8244 10363
rect 8306 9937 8323 10363
rect 8777 9937 8794 10363
rect 8856 9937 8873 10363
rect 8935 10303 9265 10315
rect 8935 9997 8947 10303
rect 8947 9997 9253 10303
rect 9253 9997 9265 10303
rect 8935 9985 9265 9997
rect 9327 9937 9344 10363
rect 9406 9937 9423 10363
rect 9877 9937 9894 10363
rect 9956 9937 9973 10363
rect 10035 10303 10365 10315
rect 10035 9997 10047 10303
rect 10047 9997 10353 10303
rect 10353 9997 10365 10303
rect 10035 9985 10365 9997
rect 10427 9937 10444 10363
rect 10506 9937 10523 10363
rect 10977 9937 10994 10363
rect 11056 9937 11073 10363
rect 11135 10303 11465 10315
rect 11135 9997 11147 10303
rect 11147 9997 11453 10303
rect 11453 9997 11465 10303
rect 11135 9985 11465 9997
rect 11527 9937 11544 10363
rect 11606 9937 11623 10363
rect 12077 9937 12094 10363
rect 12156 9937 12173 10363
rect 12235 10303 12565 10315
rect 12235 9997 12247 10303
rect 12247 9997 12553 10303
rect 12553 9997 12565 10303
rect 12235 9985 12565 9997
rect 12627 9937 12644 10363
rect 12706 9937 12723 10363
rect 13177 9937 13194 10363
rect 13256 9937 13273 10363
rect 13335 10303 13665 10315
rect 13335 9997 13347 10303
rect 13347 9997 13653 10303
rect 13653 9997 13665 10303
rect 13335 9985 13665 9997
rect -463 9906 -37 9923
rect 87 9906 513 9923
rect 637 9906 1063 9923
rect 1187 9906 1613 9923
rect 1737 9906 2163 9923
rect 2287 9906 2713 9923
rect 2837 9906 3263 9923
rect 3387 9906 3813 9923
rect 3937 9906 4363 9923
rect 4487 9906 4913 9923
rect 5037 9906 5463 9923
rect 5587 9906 6013 9923
rect 6137 9906 6563 9923
rect 6687 9906 7113 9923
rect 7237 9906 7663 9923
rect 7787 9906 8213 9923
rect 8337 9906 8763 9923
rect 8887 9906 9313 9923
rect 9437 9906 9863 9923
rect 9987 9906 10413 9923
rect 10537 9906 10963 9923
rect 11087 9906 11513 9923
rect 11637 9906 12063 9923
rect 12187 9906 12613 9923
rect 12737 9906 13163 9923
rect 13287 9906 13713 9923
rect 13987 9919 14263 10450
rect -1013 9369 -737 9900
rect -542 9858 -508 9892
rect 8 9858 42 9892
rect 558 9858 592 9892
rect 1108 9858 1142 9892
rect 1658 9858 1692 9892
rect 2208 9858 2242 9892
rect 2758 9858 2792 9892
rect 3308 9858 3342 9892
rect 3858 9858 3892 9892
rect 4408 9858 4442 9892
rect 4958 9858 4992 9892
rect 5508 9858 5542 9892
rect 6058 9858 6092 9892
rect 6608 9858 6642 9892
rect 7158 9858 7192 9892
rect 7708 9858 7742 9892
rect 8258 9858 8292 9892
rect 8808 9858 8842 9892
rect 9358 9858 9392 9892
rect 9908 9858 9942 9892
rect 10458 9858 10492 9892
rect 11008 9858 11042 9892
rect 11558 9858 11592 9892
rect 12108 9858 12142 9892
rect 12658 9858 12692 9892
rect 13208 9858 13242 9892
rect 13758 9858 13792 9892
rect -463 9827 -37 9844
rect 87 9827 513 9844
rect 637 9827 1063 9844
rect 1187 9827 1613 9844
rect 1737 9827 2163 9844
rect 2287 9827 2713 9844
rect 2837 9827 3263 9844
rect 3387 9827 3813 9844
rect 3937 9827 4363 9844
rect 4487 9827 4913 9844
rect 5037 9827 5463 9844
rect 5587 9827 6013 9844
rect 6137 9827 6563 9844
rect 6687 9827 7113 9844
rect 7237 9827 7663 9844
rect 7787 9827 8213 9844
rect 8337 9827 8763 9844
rect 8887 9827 9313 9844
rect 9437 9827 9863 9844
rect 9987 9827 10413 9844
rect 10537 9827 10963 9844
rect 11087 9827 11513 9844
rect 11637 9827 12063 9844
rect 12187 9827 12613 9844
rect 12737 9827 13163 9844
rect 13287 9827 13713 9844
rect -415 9753 -85 9765
rect -415 9447 -403 9753
rect -403 9447 -97 9753
rect -97 9447 -85 9753
rect -415 9435 -85 9447
rect -23 9387 -6 9813
rect 56 9387 73 9813
rect 527 9387 544 9813
rect 606 9387 623 9813
rect 685 9753 1015 9765
rect 685 9447 697 9753
rect 697 9447 1003 9753
rect 1003 9447 1015 9753
rect 685 9435 1015 9447
rect 1077 9387 1094 9813
rect 1156 9387 1173 9813
rect 1627 9387 1644 9813
rect 1706 9387 1723 9813
rect 1785 9753 2115 9765
rect 1785 9447 1797 9753
rect 1797 9447 2103 9753
rect 2103 9447 2115 9753
rect 1785 9435 2115 9447
rect 2177 9387 2194 9813
rect 2256 9387 2273 9813
rect 2727 9387 2744 9813
rect 2806 9387 2823 9813
rect 2885 9753 3215 9765
rect 2885 9447 2897 9753
rect 2897 9447 3203 9753
rect 3203 9447 3215 9753
rect 2885 9435 3215 9447
rect 3277 9387 3294 9813
rect 3356 9387 3373 9813
rect 3827 9387 3844 9813
rect 3906 9387 3923 9813
rect 3985 9753 4315 9765
rect 3985 9447 3997 9753
rect 3997 9447 4303 9753
rect 4303 9447 4315 9753
rect 3985 9435 4315 9447
rect 4377 9387 4394 9813
rect 4456 9387 4473 9813
rect 4927 9387 4944 9813
rect 5006 9387 5023 9813
rect 5085 9753 5415 9765
rect 5085 9447 5097 9753
rect 5097 9447 5403 9753
rect 5403 9447 5415 9753
rect 5085 9435 5415 9447
rect 5477 9387 5494 9813
rect 5556 9387 5573 9813
rect 6027 9387 6044 9813
rect 6106 9387 6123 9813
rect 6185 9753 6515 9765
rect 6185 9447 6197 9753
rect 6197 9447 6503 9753
rect 6503 9447 6515 9753
rect 6185 9435 6515 9447
rect 6577 9387 6594 9813
rect 6656 9387 6673 9813
rect 7127 9387 7144 9813
rect 7206 9387 7223 9813
rect 7285 9753 7615 9765
rect 7285 9447 7297 9753
rect 7297 9447 7603 9753
rect 7603 9447 7615 9753
rect 7285 9435 7615 9447
rect 7677 9387 7694 9813
rect 7756 9387 7773 9813
rect 8227 9387 8244 9813
rect 8306 9387 8323 9813
rect 8385 9753 8715 9765
rect 8385 9447 8397 9753
rect 8397 9447 8703 9753
rect 8703 9447 8715 9753
rect 8385 9435 8715 9447
rect 8777 9387 8794 9813
rect 8856 9387 8873 9813
rect 9327 9387 9344 9813
rect 9406 9387 9423 9813
rect 9485 9753 9815 9765
rect 9485 9447 9497 9753
rect 9497 9447 9803 9753
rect 9803 9447 9815 9753
rect 9485 9435 9815 9447
rect 9877 9387 9894 9813
rect 9956 9387 9973 9813
rect 10427 9387 10444 9813
rect 10506 9387 10523 9813
rect 10585 9753 10915 9765
rect 10585 9447 10597 9753
rect 10597 9447 10903 9753
rect 10903 9447 10915 9753
rect 10585 9435 10915 9447
rect 10977 9387 10994 9813
rect 11056 9387 11073 9813
rect 11527 9387 11544 9813
rect 11606 9387 11623 9813
rect 11685 9753 12015 9765
rect 11685 9447 11697 9753
rect 11697 9447 12003 9753
rect 12003 9447 12015 9753
rect 11685 9435 12015 9447
rect 12077 9387 12094 9813
rect 12156 9387 12173 9813
rect 12627 9387 12644 9813
rect 12706 9387 12723 9813
rect 12785 9753 13115 9765
rect 12785 9447 12797 9753
rect 12797 9447 13103 9753
rect 13103 9447 13115 9753
rect 12785 9435 13115 9447
rect 13177 9387 13194 9813
rect 13256 9387 13273 9813
rect -463 9356 -37 9373
rect 87 9356 513 9373
rect 637 9356 1063 9373
rect 1187 9356 1613 9373
rect 1737 9356 2163 9373
rect 2287 9356 2713 9373
rect 2837 9356 3263 9373
rect 3387 9356 3813 9373
rect 3937 9356 4363 9373
rect 4487 9356 4913 9373
rect 5037 9356 5463 9373
rect 5587 9356 6013 9373
rect 6137 9356 6563 9373
rect 6687 9356 7113 9373
rect 7237 9356 7663 9373
rect 7787 9356 8213 9373
rect 8337 9356 8763 9373
rect 8887 9356 9313 9373
rect 9437 9356 9863 9373
rect 9987 9356 10413 9373
rect 10537 9356 10963 9373
rect 11087 9356 11513 9373
rect 11637 9356 12063 9373
rect 12187 9356 12613 9373
rect 12737 9356 13163 9373
rect 13287 9356 13713 9373
rect 13987 9369 14263 9900
rect -1013 8819 -737 9350
rect -542 9308 -508 9342
rect 8 9308 42 9342
rect 558 9308 592 9342
rect 1108 9308 1142 9342
rect 1658 9308 1692 9342
rect 2208 9308 2242 9342
rect 2758 9308 2792 9342
rect 3308 9308 3342 9342
rect 3858 9308 3892 9342
rect 4408 9308 4442 9342
rect 4958 9308 4992 9342
rect 5508 9308 5542 9342
rect 6058 9308 6092 9342
rect 6608 9308 6642 9342
rect 7158 9308 7192 9342
rect 7708 9308 7742 9342
rect 8258 9308 8292 9342
rect 8808 9308 8842 9342
rect 9358 9308 9392 9342
rect 9908 9308 9942 9342
rect 10458 9308 10492 9342
rect 11008 9308 11042 9342
rect 11558 9308 11592 9342
rect 12108 9308 12142 9342
rect 12658 9308 12692 9342
rect 13208 9308 13242 9342
rect 13758 9308 13792 9342
rect -463 9277 -37 9294
rect 87 9277 513 9294
rect 637 9277 1063 9294
rect 1187 9277 1613 9294
rect 1737 9277 2163 9294
rect 2287 9277 2713 9294
rect 2837 9277 3263 9294
rect 3387 9277 3813 9294
rect 3937 9277 4363 9294
rect 4487 9277 4913 9294
rect 5037 9277 5463 9294
rect 5587 9277 6013 9294
rect 6137 9277 6563 9294
rect 6687 9277 7113 9294
rect 7237 9277 7663 9294
rect 7787 9277 8213 9294
rect 8337 9277 8763 9294
rect 8887 9277 9313 9294
rect 9437 9277 9863 9294
rect 9987 9277 10413 9294
rect 10537 9277 10963 9294
rect 11087 9277 11513 9294
rect 11637 9277 12063 9294
rect 12187 9277 12613 9294
rect 12737 9277 13163 9294
rect 13287 9277 13713 9294
rect -23 8837 -6 9263
rect 56 8837 73 9263
rect 135 9203 465 9215
rect 135 8897 147 9203
rect 147 8897 453 9203
rect 453 8897 465 9203
rect 135 8885 465 8897
rect 527 8837 544 9263
rect 606 8837 623 9263
rect 1077 8837 1094 9263
rect 1156 8837 1173 9263
rect 1235 9203 1565 9215
rect 1235 8897 1247 9203
rect 1247 8897 1553 9203
rect 1553 8897 1565 9203
rect 1235 8885 1565 8897
rect 1627 8837 1644 9263
rect 1706 8837 1723 9263
rect 2177 8837 2194 9263
rect 2256 8837 2273 9263
rect 2335 9203 2665 9215
rect 2335 8897 2347 9203
rect 2347 8897 2653 9203
rect 2653 8897 2665 9203
rect 2335 8885 2665 8897
rect 2727 8837 2744 9263
rect 2806 8837 2823 9263
rect 3277 8837 3294 9263
rect 3356 8837 3373 9263
rect 3435 9203 3765 9215
rect 3435 8897 3447 9203
rect 3447 8897 3753 9203
rect 3753 8897 3765 9203
rect 3435 8885 3765 8897
rect 3827 8837 3844 9263
rect 3906 8837 3923 9263
rect 4377 8837 4394 9263
rect 4456 8837 4473 9263
rect 4535 9203 4865 9215
rect 4535 8897 4547 9203
rect 4547 8897 4853 9203
rect 4853 8897 4865 9203
rect 4535 8885 4865 8897
rect 4927 8837 4944 9263
rect 5006 8837 5023 9263
rect 5477 8837 5494 9263
rect 5556 8837 5573 9263
rect 5635 9203 5965 9215
rect 5635 8897 5647 9203
rect 5647 8897 5953 9203
rect 5953 8897 5965 9203
rect 5635 8885 5965 8897
rect 6027 8837 6044 9263
rect 6106 8837 6123 9263
rect 6577 8837 6594 9263
rect 6656 8837 6673 9263
rect 6735 9203 7065 9215
rect 6735 8897 6747 9203
rect 6747 8897 7053 9203
rect 7053 8897 7065 9203
rect 6735 8885 7065 8897
rect 7127 8837 7144 9263
rect 7206 8837 7223 9263
rect 7677 8837 7694 9263
rect 7756 8837 7773 9263
rect 7835 9203 8165 9215
rect 7835 8897 7847 9203
rect 7847 8897 8153 9203
rect 8153 8897 8165 9203
rect 7835 8885 8165 8897
rect 8227 8837 8244 9263
rect 8306 8837 8323 9263
rect 8777 8837 8794 9263
rect 8856 8837 8873 9263
rect 8935 9203 9265 9215
rect 8935 8897 8947 9203
rect 8947 8897 9253 9203
rect 9253 8897 9265 9203
rect 8935 8885 9265 8897
rect 9327 8837 9344 9263
rect 9406 8837 9423 9263
rect 9877 8837 9894 9263
rect 9956 8837 9973 9263
rect 10035 9203 10365 9215
rect 10035 8897 10047 9203
rect 10047 8897 10353 9203
rect 10353 8897 10365 9203
rect 10035 8885 10365 8897
rect 10427 8837 10444 9263
rect 10506 8837 10523 9263
rect 10977 8837 10994 9263
rect 11056 8837 11073 9263
rect 11135 9203 11465 9215
rect 11135 8897 11147 9203
rect 11147 8897 11453 9203
rect 11453 8897 11465 9203
rect 11135 8885 11465 8897
rect 11527 8837 11544 9263
rect 11606 8837 11623 9263
rect 12077 8837 12094 9263
rect 12156 8837 12173 9263
rect 12235 9203 12565 9215
rect 12235 8897 12247 9203
rect 12247 8897 12553 9203
rect 12553 8897 12565 9203
rect 12235 8885 12565 8897
rect 12627 8837 12644 9263
rect 12706 8837 12723 9263
rect 13177 8837 13194 9263
rect 13256 8837 13273 9263
rect 13335 9203 13665 9215
rect 13335 8897 13347 9203
rect 13347 8897 13653 9203
rect 13653 8897 13665 9203
rect 13335 8885 13665 8897
rect -463 8806 -37 8823
rect 87 8806 513 8823
rect 637 8806 1063 8823
rect 1187 8806 1613 8823
rect 1737 8806 2163 8823
rect 2287 8806 2713 8823
rect 2837 8806 3263 8823
rect 3387 8806 3813 8823
rect 3937 8806 4363 8823
rect 4487 8806 4913 8823
rect 5037 8806 5463 8823
rect 5587 8806 6013 8823
rect 6137 8806 6563 8823
rect 6687 8806 7113 8823
rect 7237 8806 7663 8823
rect 7787 8806 8213 8823
rect 8337 8806 8763 8823
rect 8887 8806 9313 8823
rect 9437 8806 9863 8823
rect 9987 8806 10413 8823
rect 10537 8806 10963 8823
rect 11087 8806 11513 8823
rect 11637 8806 12063 8823
rect 12187 8806 12613 8823
rect 12737 8806 13163 8823
rect 13287 8806 13713 8823
rect 13987 8819 14263 9350
rect -1013 8269 -737 8800
rect -542 8758 -508 8792
rect 8 8758 42 8792
rect 558 8758 592 8792
rect 1108 8758 1142 8792
rect 1658 8758 1692 8792
rect 2208 8758 2242 8792
rect 2758 8758 2792 8792
rect 3308 8758 3342 8792
rect 3858 8758 3892 8792
rect 4408 8758 4442 8792
rect 4958 8758 4992 8792
rect 5508 8758 5542 8792
rect 6058 8758 6092 8792
rect 6608 8758 6642 8792
rect 7158 8758 7192 8792
rect 7708 8758 7742 8792
rect 8258 8758 8292 8792
rect 8808 8758 8842 8792
rect 9358 8758 9392 8792
rect 9908 8758 9942 8792
rect 10458 8758 10492 8792
rect 11008 8758 11042 8792
rect 11558 8758 11592 8792
rect 12108 8758 12142 8792
rect 12658 8758 12692 8792
rect 13208 8758 13242 8792
rect 13758 8758 13792 8792
rect -463 8727 -37 8744
rect 87 8727 513 8744
rect 637 8727 1063 8744
rect 1187 8727 1613 8744
rect 1737 8727 2163 8744
rect 2287 8727 2713 8744
rect 2837 8727 3263 8744
rect 3387 8727 3813 8744
rect 3937 8727 4363 8744
rect 4487 8727 4913 8744
rect 5037 8727 5463 8744
rect 5587 8727 6013 8744
rect 6137 8727 6563 8744
rect 6687 8727 7113 8744
rect 7237 8727 7663 8744
rect 7787 8727 8213 8744
rect 8337 8727 8763 8744
rect 8887 8727 9313 8744
rect 9437 8727 9863 8744
rect 9987 8727 10413 8744
rect 10537 8727 10963 8744
rect 11087 8727 11513 8744
rect 11637 8727 12063 8744
rect 12187 8727 12613 8744
rect 12737 8727 13163 8744
rect 13287 8727 13713 8744
rect -415 8653 -85 8665
rect -415 8347 -403 8653
rect -403 8347 -97 8653
rect -97 8347 -85 8653
rect -415 8335 -85 8347
rect -23 8287 -6 8713
rect 56 8287 73 8713
rect 527 8287 544 8713
rect 606 8287 623 8713
rect 685 8653 1015 8665
rect 685 8347 697 8653
rect 697 8347 1003 8653
rect 1003 8347 1015 8653
rect 685 8335 1015 8347
rect 1077 8287 1094 8713
rect 1156 8287 1173 8713
rect 1627 8287 1644 8713
rect 1706 8287 1723 8713
rect 1785 8653 2115 8665
rect 1785 8347 1797 8653
rect 1797 8347 2103 8653
rect 2103 8347 2115 8653
rect 1785 8335 2115 8347
rect 2177 8287 2194 8713
rect 2256 8287 2273 8713
rect 2727 8287 2744 8713
rect 2806 8287 2823 8713
rect 2885 8653 3215 8665
rect 2885 8347 2897 8653
rect 2897 8347 3203 8653
rect 3203 8347 3215 8653
rect 2885 8335 3215 8347
rect 3277 8287 3294 8713
rect 3356 8287 3373 8713
rect 3827 8287 3844 8713
rect 3906 8287 3923 8713
rect 3985 8653 4315 8665
rect 3985 8347 3997 8653
rect 3997 8347 4303 8653
rect 4303 8347 4315 8653
rect 3985 8335 4315 8347
rect 4377 8287 4394 8713
rect 4456 8287 4473 8713
rect 4927 8287 4944 8713
rect 5006 8287 5023 8713
rect 5085 8653 5415 8665
rect 5085 8347 5097 8653
rect 5097 8347 5403 8653
rect 5403 8347 5415 8653
rect 5085 8335 5415 8347
rect 5477 8287 5494 8713
rect 5556 8287 5573 8713
rect 6027 8287 6044 8713
rect 6106 8287 6123 8713
rect 6185 8653 6515 8665
rect 6185 8347 6197 8653
rect 6197 8347 6503 8653
rect 6503 8347 6515 8653
rect 6185 8335 6515 8347
rect 6577 8287 6594 8713
rect 6656 8287 6673 8713
rect 7127 8287 7144 8713
rect 7206 8287 7223 8713
rect 7285 8653 7615 8665
rect 7285 8347 7297 8653
rect 7297 8347 7603 8653
rect 7603 8347 7615 8653
rect 7285 8335 7615 8347
rect 7677 8287 7694 8713
rect 7756 8287 7773 8713
rect 8227 8287 8244 8713
rect 8306 8287 8323 8713
rect 8385 8653 8715 8665
rect 8385 8347 8397 8653
rect 8397 8347 8703 8653
rect 8703 8347 8715 8653
rect 8385 8335 8715 8347
rect 8777 8287 8794 8713
rect 8856 8287 8873 8713
rect 9327 8287 9344 8713
rect 9406 8287 9423 8713
rect 9485 8653 9815 8665
rect 9485 8347 9497 8653
rect 9497 8347 9803 8653
rect 9803 8347 9815 8653
rect 9485 8335 9815 8347
rect 9877 8287 9894 8713
rect 9956 8287 9973 8713
rect 10427 8287 10444 8713
rect 10506 8287 10523 8713
rect 10585 8653 10915 8665
rect 10585 8347 10597 8653
rect 10597 8347 10903 8653
rect 10903 8347 10915 8653
rect 10585 8335 10915 8347
rect 10977 8287 10994 8713
rect 11056 8287 11073 8713
rect 11527 8287 11544 8713
rect 11606 8287 11623 8713
rect 11685 8653 12015 8665
rect 11685 8347 11697 8653
rect 11697 8347 12003 8653
rect 12003 8347 12015 8653
rect 11685 8335 12015 8347
rect 12077 8287 12094 8713
rect 12156 8287 12173 8713
rect 12627 8287 12644 8713
rect 12706 8287 12723 8713
rect 12785 8653 13115 8665
rect 12785 8347 12797 8653
rect 12797 8347 13103 8653
rect 13103 8347 13115 8653
rect 12785 8335 13115 8347
rect 13177 8287 13194 8713
rect 13256 8287 13273 8713
rect -463 8256 -37 8273
rect 87 8256 513 8273
rect 637 8256 1063 8273
rect 1187 8256 1613 8273
rect 1737 8256 2163 8273
rect 2287 8256 2713 8273
rect 2837 8256 3263 8273
rect 3387 8256 3813 8273
rect 3937 8256 4363 8273
rect 4487 8256 4913 8273
rect 5037 8256 5463 8273
rect 5587 8256 6013 8273
rect 6137 8256 6563 8273
rect 6687 8256 7113 8273
rect 7237 8256 7663 8273
rect 7787 8256 8213 8273
rect 8337 8256 8763 8273
rect 8887 8256 9313 8273
rect 9437 8256 9863 8273
rect 9987 8256 10413 8273
rect 10537 8256 10963 8273
rect 11087 8256 11513 8273
rect 11637 8256 12063 8273
rect 12187 8256 12613 8273
rect 12737 8256 13163 8273
rect 13287 8256 13713 8273
rect 13987 8269 14263 8800
rect -1013 7719 -737 8250
rect -542 8208 -508 8242
rect 8 8208 42 8242
rect 558 8208 592 8242
rect 1108 8208 1142 8242
rect 1658 8208 1692 8242
rect 2208 8208 2242 8242
rect 2758 8208 2792 8242
rect 3308 8208 3342 8242
rect 3858 8208 3892 8242
rect 4408 8208 4442 8242
rect 4958 8208 4992 8242
rect 5508 8208 5542 8242
rect 6058 8208 6092 8242
rect 6608 8208 6642 8242
rect 7158 8208 7192 8242
rect 7708 8208 7742 8242
rect 8258 8208 8292 8242
rect 8808 8208 8842 8242
rect 9358 8208 9392 8242
rect 9908 8208 9942 8242
rect 10458 8208 10492 8242
rect 11008 8208 11042 8242
rect 11558 8208 11592 8242
rect 12108 8208 12142 8242
rect 12658 8208 12692 8242
rect 13208 8208 13242 8242
rect 13758 8208 13792 8242
rect -463 8177 -37 8194
rect 87 8177 513 8194
rect 637 8177 1063 8194
rect 1187 8177 1613 8194
rect 1737 8177 2163 8194
rect 2287 8177 2713 8194
rect 2837 8177 3263 8194
rect 3387 8177 3813 8194
rect 3937 8177 4363 8194
rect 4487 8177 4913 8194
rect 5037 8177 5463 8194
rect 5587 8177 6013 8194
rect 6137 8177 6563 8194
rect 6687 8177 7113 8194
rect 7237 8177 7663 8194
rect 7787 8177 8213 8194
rect 8337 8177 8763 8194
rect 8887 8177 9313 8194
rect 9437 8177 9863 8194
rect 9987 8177 10413 8194
rect 10537 8177 10963 8194
rect 11087 8177 11513 8194
rect 11637 8177 12063 8194
rect 12187 8177 12613 8194
rect 12737 8177 13163 8194
rect 13287 8177 13713 8194
rect -23 7737 -6 8163
rect 56 7737 73 8163
rect 135 8103 465 8115
rect 135 7797 147 8103
rect 147 7797 453 8103
rect 453 7797 465 8103
rect 135 7785 465 7797
rect 527 7737 544 8163
rect 606 7737 623 8163
rect 1077 7737 1094 8163
rect 1156 7737 1173 8163
rect 1235 8103 1565 8115
rect 1235 7797 1247 8103
rect 1247 7797 1553 8103
rect 1553 7797 1565 8103
rect 1235 7785 1565 7797
rect 1627 7737 1644 8163
rect 1706 7737 1723 8163
rect 2177 7737 2194 8163
rect 2256 7737 2273 8163
rect 2335 8103 2665 8115
rect 2335 7797 2347 8103
rect 2347 7797 2653 8103
rect 2653 7797 2665 8103
rect 2335 7785 2665 7797
rect 2727 7737 2744 8163
rect 2806 7737 2823 8163
rect 3277 7737 3294 8163
rect 3356 7737 3373 8163
rect 3435 8103 3765 8115
rect 3435 7797 3447 8103
rect 3447 7797 3753 8103
rect 3753 7797 3765 8103
rect 3435 7785 3765 7797
rect 3827 7737 3844 8163
rect 3906 7737 3923 8163
rect 4377 7737 4394 8163
rect 4456 7737 4473 8163
rect 4535 8103 4865 8115
rect 4535 7797 4547 8103
rect 4547 7797 4853 8103
rect 4853 7797 4865 8103
rect 4535 7785 4865 7797
rect 4927 7737 4944 8163
rect 5006 7737 5023 8163
rect 5477 7737 5494 8163
rect 5556 7737 5573 8163
rect 5635 8103 5965 8115
rect 5635 7797 5647 8103
rect 5647 7797 5953 8103
rect 5953 7797 5965 8103
rect 5635 7785 5965 7797
rect 6027 7737 6044 8163
rect 6106 7737 6123 8163
rect 6577 7737 6594 8163
rect 6656 7737 6673 8163
rect 6735 8103 7065 8115
rect 6735 7797 6747 8103
rect 6747 7797 7053 8103
rect 7053 7797 7065 8103
rect 6735 7785 7065 7797
rect 7127 7737 7144 8163
rect 7206 7737 7223 8163
rect 7677 7737 7694 8163
rect 7756 7737 7773 8163
rect 7835 8103 8165 8115
rect 7835 7797 7847 8103
rect 7847 7797 8153 8103
rect 8153 7797 8165 8103
rect 7835 7785 8165 7797
rect 8227 7737 8244 8163
rect 8306 7737 8323 8163
rect 8777 7737 8794 8163
rect 8856 7737 8873 8163
rect 8935 8103 9265 8115
rect 8935 7797 8947 8103
rect 8947 7797 9253 8103
rect 9253 7797 9265 8103
rect 8935 7785 9265 7797
rect 9327 7737 9344 8163
rect 9406 7737 9423 8163
rect 9877 7737 9894 8163
rect 9956 7737 9973 8163
rect 10035 8103 10365 8115
rect 10035 7797 10047 8103
rect 10047 7797 10353 8103
rect 10353 7797 10365 8103
rect 10035 7785 10365 7797
rect 10427 7737 10444 8163
rect 10506 7737 10523 8163
rect 10977 7737 10994 8163
rect 11056 7737 11073 8163
rect 11135 8103 11465 8115
rect 11135 7797 11147 8103
rect 11147 7797 11453 8103
rect 11453 7797 11465 8103
rect 11135 7785 11465 7797
rect 11527 7737 11544 8163
rect 11606 7737 11623 8163
rect 12077 7737 12094 8163
rect 12156 7737 12173 8163
rect 12235 8103 12565 8115
rect 12235 7797 12247 8103
rect 12247 7797 12553 8103
rect 12553 7797 12565 8103
rect 12235 7785 12565 7797
rect 12627 7737 12644 8163
rect 12706 7737 12723 8163
rect 13177 7737 13194 8163
rect 13256 7737 13273 8163
rect 13335 8103 13665 8115
rect 13335 7797 13347 8103
rect 13347 7797 13653 8103
rect 13653 7797 13665 8103
rect 13335 7785 13665 7797
rect -463 7706 -37 7723
rect 87 7706 513 7723
rect 637 7706 1063 7723
rect 1187 7706 1613 7723
rect 1737 7706 2163 7723
rect 2287 7706 2713 7723
rect 2837 7706 3263 7723
rect 3387 7706 3813 7723
rect 3937 7706 4363 7723
rect 4487 7706 4913 7723
rect 5037 7706 5463 7723
rect 5587 7706 6013 7723
rect 6137 7706 6563 7723
rect 6687 7706 7113 7723
rect 7237 7706 7663 7723
rect 7787 7706 8213 7723
rect 8337 7706 8763 7723
rect 8887 7706 9313 7723
rect 9437 7706 9863 7723
rect 9987 7706 10413 7723
rect 10537 7706 10963 7723
rect 11087 7706 11513 7723
rect 11637 7706 12063 7723
rect 12187 7706 12613 7723
rect 12737 7706 13163 7723
rect 13287 7706 13713 7723
rect 13987 7719 14263 8250
rect -1013 7169 -737 7700
rect -542 7658 -508 7692
rect 8 7658 42 7692
rect 558 7658 592 7692
rect 1108 7658 1142 7692
rect 1658 7658 1692 7692
rect 2208 7658 2242 7692
rect 2758 7658 2792 7692
rect 3308 7658 3342 7692
rect 3858 7658 3892 7692
rect 4408 7658 4442 7692
rect 4958 7658 4992 7692
rect 5508 7658 5542 7692
rect 6058 7658 6092 7692
rect 6608 7658 6642 7692
rect 7158 7658 7192 7692
rect 7708 7658 7742 7692
rect 8258 7658 8292 7692
rect 8808 7658 8842 7692
rect 9358 7658 9392 7692
rect 9908 7658 9942 7692
rect 10458 7658 10492 7692
rect 11008 7658 11042 7692
rect 11558 7658 11592 7692
rect 12108 7658 12142 7692
rect 12658 7658 12692 7692
rect 13208 7658 13242 7692
rect 13758 7658 13792 7692
rect -463 7627 -37 7644
rect 87 7627 513 7644
rect 637 7627 1063 7644
rect 1187 7627 1613 7644
rect 1737 7627 2163 7644
rect 2287 7627 2713 7644
rect 2837 7627 3263 7644
rect 3387 7627 3813 7644
rect 3937 7627 4363 7644
rect 4487 7627 4913 7644
rect 5037 7627 5463 7644
rect 5587 7627 6013 7644
rect 6137 7627 6563 7644
rect 6687 7627 7113 7644
rect 7237 7627 7663 7644
rect 7787 7627 8213 7644
rect 8337 7627 8763 7644
rect 8887 7627 9313 7644
rect 9437 7627 9863 7644
rect 9987 7627 10413 7644
rect 10537 7627 10963 7644
rect 11087 7627 11513 7644
rect 11637 7627 12063 7644
rect 12187 7627 12613 7644
rect 12737 7627 13163 7644
rect 13287 7627 13713 7644
rect -415 7553 -85 7565
rect -415 7247 -403 7553
rect -403 7247 -97 7553
rect -97 7247 -85 7553
rect -415 7235 -85 7247
rect -23 7187 -6 7613
rect 56 7187 73 7613
rect 527 7187 544 7613
rect 606 7187 623 7613
rect 685 7553 1015 7565
rect 685 7247 697 7553
rect 697 7247 1003 7553
rect 1003 7247 1015 7553
rect 685 7235 1015 7247
rect 1077 7187 1094 7613
rect 1156 7187 1173 7613
rect 1627 7187 1644 7613
rect 1706 7187 1723 7613
rect 1785 7553 2115 7565
rect 1785 7247 1797 7553
rect 1797 7247 2103 7553
rect 2103 7247 2115 7553
rect 1785 7235 2115 7247
rect 2177 7187 2194 7613
rect 2256 7187 2273 7613
rect 2727 7187 2744 7613
rect 2806 7187 2823 7613
rect 2885 7553 3215 7565
rect 2885 7247 2897 7553
rect 2897 7247 3203 7553
rect 3203 7247 3215 7553
rect 2885 7235 3215 7247
rect 3277 7187 3294 7613
rect 3356 7187 3373 7613
rect 3827 7187 3844 7613
rect 3906 7187 3923 7613
rect 3985 7553 4315 7565
rect 3985 7247 3997 7553
rect 3997 7247 4303 7553
rect 4303 7247 4315 7553
rect 3985 7235 4315 7247
rect 4377 7187 4394 7613
rect 4456 7187 4473 7613
rect 4927 7187 4944 7613
rect 5006 7187 5023 7613
rect 5085 7553 5415 7565
rect 5085 7247 5097 7553
rect 5097 7247 5403 7553
rect 5403 7247 5415 7553
rect 5085 7235 5415 7247
rect 5477 7187 5494 7613
rect 5556 7187 5573 7613
rect 6027 7187 6044 7613
rect 6106 7187 6123 7613
rect 6185 7553 6515 7565
rect 6185 7247 6197 7553
rect 6197 7247 6503 7553
rect 6503 7247 6515 7553
rect 6185 7235 6515 7247
rect 6577 7187 6594 7613
rect 6656 7187 6673 7613
rect 7127 7187 7144 7613
rect 7206 7187 7223 7613
rect 7285 7553 7615 7565
rect 7285 7247 7297 7553
rect 7297 7247 7603 7553
rect 7603 7247 7615 7553
rect 7285 7235 7615 7247
rect 7677 7187 7694 7613
rect 7756 7187 7773 7613
rect 8227 7187 8244 7613
rect 8306 7187 8323 7613
rect 8385 7553 8715 7565
rect 8385 7247 8397 7553
rect 8397 7247 8703 7553
rect 8703 7247 8715 7553
rect 8385 7235 8715 7247
rect 8777 7187 8794 7613
rect 8856 7187 8873 7613
rect 9327 7187 9344 7613
rect 9406 7187 9423 7613
rect 9485 7553 9815 7565
rect 9485 7247 9497 7553
rect 9497 7247 9803 7553
rect 9803 7247 9815 7553
rect 9485 7235 9815 7247
rect 9877 7187 9894 7613
rect 9956 7187 9973 7613
rect 10427 7187 10444 7613
rect 10506 7187 10523 7613
rect 10585 7553 10915 7565
rect 10585 7247 10597 7553
rect 10597 7247 10903 7553
rect 10903 7247 10915 7553
rect 10585 7235 10915 7247
rect 10977 7187 10994 7613
rect 11056 7187 11073 7613
rect 11527 7187 11544 7613
rect 11606 7187 11623 7613
rect 11685 7553 12015 7565
rect 11685 7247 11697 7553
rect 11697 7247 12003 7553
rect 12003 7247 12015 7553
rect 11685 7235 12015 7247
rect 12077 7187 12094 7613
rect 12156 7187 12173 7613
rect 12627 7187 12644 7613
rect 12706 7187 12723 7613
rect 12785 7553 13115 7565
rect 12785 7247 12797 7553
rect 12797 7247 13103 7553
rect 13103 7247 13115 7553
rect 12785 7235 13115 7247
rect 13177 7187 13194 7613
rect 13256 7187 13273 7613
rect -463 7156 -37 7173
rect 87 7156 513 7173
rect 637 7156 1063 7173
rect 1187 7156 1613 7173
rect 1737 7156 2163 7173
rect 2287 7156 2713 7173
rect 2837 7156 3263 7173
rect 3387 7156 3813 7173
rect 3937 7156 4363 7173
rect 4487 7156 4913 7173
rect 5037 7156 5463 7173
rect 5587 7156 6013 7173
rect 6137 7156 6563 7173
rect 6687 7156 7113 7173
rect 7237 7156 7663 7173
rect 7787 7156 8213 7173
rect 8337 7156 8763 7173
rect 8887 7156 9313 7173
rect 9437 7156 9863 7173
rect 9987 7156 10413 7173
rect 10537 7156 10963 7173
rect 11087 7156 11513 7173
rect 11637 7156 12063 7173
rect 12187 7156 12613 7173
rect 12737 7156 13163 7173
rect 13287 7156 13713 7173
rect 13987 7169 14263 7700
rect -1013 6619 -737 7150
rect -542 7108 -508 7142
rect 8 7108 42 7142
rect 558 7108 592 7142
rect 1108 7108 1142 7142
rect 1658 7108 1692 7142
rect 2208 7108 2242 7142
rect 2758 7108 2792 7142
rect 3308 7108 3342 7142
rect 3858 7108 3892 7142
rect 4408 7108 4442 7142
rect 4958 7108 4992 7142
rect 5508 7108 5542 7142
rect 6058 7108 6092 7142
rect 6608 7108 6642 7142
rect 7158 7108 7192 7142
rect 7708 7108 7742 7142
rect 8258 7108 8292 7142
rect 8808 7108 8842 7142
rect 9358 7108 9392 7142
rect 9908 7108 9942 7142
rect 10458 7108 10492 7142
rect 11008 7108 11042 7142
rect 11558 7108 11592 7142
rect 12108 7108 12142 7142
rect 12658 7108 12692 7142
rect 13208 7108 13242 7142
rect 13758 7108 13792 7142
rect -463 7077 -37 7094
rect 87 7077 513 7094
rect 637 7077 1063 7094
rect 1187 7077 1613 7094
rect 1737 7077 2163 7094
rect 2287 7077 2713 7094
rect 2837 7077 3263 7094
rect 3387 7077 3813 7094
rect 3937 7077 4363 7094
rect 4487 7077 4913 7094
rect 5037 7077 5463 7094
rect 5587 7077 6013 7094
rect 6137 7077 6563 7094
rect 6687 7077 7113 7094
rect 7237 7077 7663 7094
rect 7787 7077 8213 7094
rect 8337 7077 8763 7094
rect 8887 7077 9313 7094
rect 9437 7077 9863 7094
rect 9987 7077 10413 7094
rect 10537 7077 10963 7094
rect 11087 7077 11513 7094
rect 11637 7077 12063 7094
rect 12187 7077 12613 7094
rect 12737 7077 13163 7094
rect 13287 7077 13713 7094
rect -23 6637 -6 7063
rect 56 6637 73 7063
rect 135 7003 465 7015
rect 135 6697 147 7003
rect 147 6697 453 7003
rect 453 6697 465 7003
rect 135 6685 465 6697
rect 527 6637 544 7063
rect 606 6637 623 7063
rect 1077 6637 1094 7063
rect 1156 6637 1173 7063
rect 1235 7003 1565 7015
rect 1235 6697 1247 7003
rect 1247 6697 1553 7003
rect 1553 6697 1565 7003
rect 1235 6685 1565 6697
rect 1627 6637 1644 7063
rect 1706 6637 1723 7063
rect 2177 6637 2194 7063
rect 2256 6637 2273 7063
rect 2335 7003 2665 7015
rect 2335 6697 2347 7003
rect 2347 6697 2653 7003
rect 2653 6697 2665 7003
rect 2335 6685 2665 6697
rect 2727 6637 2744 7063
rect 2806 6637 2823 7063
rect 3277 6637 3294 7063
rect 3356 6637 3373 7063
rect 3435 7003 3765 7015
rect 3435 6697 3447 7003
rect 3447 6697 3753 7003
rect 3753 6697 3765 7003
rect 3435 6685 3765 6697
rect 3827 6637 3844 7063
rect 3906 6637 3923 7063
rect 4377 6637 4394 7063
rect 4456 6637 4473 7063
rect 4535 7003 4865 7015
rect 4535 6697 4547 7003
rect 4547 6697 4853 7003
rect 4853 6697 4865 7003
rect 4535 6685 4865 6697
rect 4927 6637 4944 7063
rect 5006 6637 5023 7063
rect 5477 6637 5494 7063
rect 5556 6637 5573 7063
rect 5635 7003 5965 7015
rect 5635 6697 5647 7003
rect 5647 6697 5953 7003
rect 5953 6697 5965 7003
rect 5635 6685 5965 6697
rect 6027 6637 6044 7063
rect 6106 6637 6123 7063
rect 6577 6637 6594 7063
rect 6656 6637 6673 7063
rect 6735 7003 7065 7015
rect 6735 6697 6747 7003
rect 6747 6697 7053 7003
rect 7053 6697 7065 7003
rect 6735 6685 7065 6697
rect 7127 6637 7144 7063
rect 7206 6637 7223 7063
rect 7677 6637 7694 7063
rect 7756 6637 7773 7063
rect 7835 7003 8165 7015
rect 7835 6697 7847 7003
rect 7847 6697 8153 7003
rect 8153 6697 8165 7003
rect 7835 6685 8165 6697
rect 8227 6637 8244 7063
rect 8306 6637 8323 7063
rect 8777 6637 8794 7063
rect 8856 6637 8873 7063
rect 8935 7003 9265 7015
rect 8935 6697 8947 7003
rect 8947 6697 9253 7003
rect 9253 6697 9265 7003
rect 8935 6685 9265 6697
rect 9327 6637 9344 7063
rect 9406 6637 9423 7063
rect 9877 6637 9894 7063
rect 9956 6637 9973 7063
rect 10035 7003 10365 7015
rect 10035 6697 10047 7003
rect 10047 6697 10353 7003
rect 10353 6697 10365 7003
rect 10035 6685 10365 6697
rect 10427 6637 10444 7063
rect 10506 6637 10523 7063
rect 10977 6637 10994 7063
rect 11056 6637 11073 7063
rect 11135 7003 11465 7015
rect 11135 6697 11147 7003
rect 11147 6697 11453 7003
rect 11453 6697 11465 7003
rect 11135 6685 11465 6697
rect 11527 6637 11544 7063
rect 11606 6637 11623 7063
rect 12077 6637 12094 7063
rect 12156 6637 12173 7063
rect 12235 7003 12565 7015
rect 12235 6697 12247 7003
rect 12247 6697 12553 7003
rect 12553 6697 12565 7003
rect 12235 6685 12565 6697
rect 12627 6637 12644 7063
rect 12706 6637 12723 7063
rect 13177 6637 13194 7063
rect 13256 6637 13273 7063
rect 13335 7003 13665 7015
rect 13335 6697 13347 7003
rect 13347 6697 13653 7003
rect 13653 6697 13665 7003
rect 13335 6685 13665 6697
rect -463 6606 -37 6623
rect 87 6606 513 6623
rect 637 6606 1063 6623
rect 1187 6606 1613 6623
rect 1737 6606 2163 6623
rect 2287 6606 2713 6623
rect 2837 6606 3263 6623
rect 3387 6606 3813 6623
rect 3937 6606 4363 6623
rect 4487 6606 4913 6623
rect 5037 6606 5463 6623
rect 5587 6606 6013 6623
rect 6137 6606 6563 6623
rect 6687 6606 7113 6623
rect 7237 6606 7663 6623
rect 7787 6606 8213 6623
rect 8337 6606 8763 6623
rect 8887 6606 9313 6623
rect 9437 6606 9863 6623
rect 9987 6606 10413 6623
rect 10537 6606 10963 6623
rect 11087 6606 11513 6623
rect 11637 6606 12063 6623
rect 12187 6606 12613 6623
rect 12737 6606 13163 6623
rect 13287 6606 13713 6623
rect 13987 6619 14263 7150
rect -1013 6069 -737 6600
rect -542 6558 -508 6592
rect 8 6558 42 6592
rect 558 6558 592 6592
rect 1108 6558 1142 6592
rect 1658 6558 1692 6592
rect 2208 6558 2242 6592
rect 2758 6558 2792 6592
rect 3308 6558 3342 6592
rect 3858 6558 3892 6592
rect 4408 6558 4442 6592
rect 4958 6558 4992 6592
rect 5508 6558 5542 6592
rect 6058 6558 6092 6592
rect 6608 6558 6642 6592
rect 7158 6558 7192 6592
rect 7708 6558 7742 6592
rect 8258 6558 8292 6592
rect 8808 6558 8842 6592
rect 9358 6558 9392 6592
rect 9908 6558 9942 6592
rect 10458 6558 10492 6592
rect 11008 6558 11042 6592
rect 11558 6558 11592 6592
rect 12108 6558 12142 6592
rect 12658 6558 12692 6592
rect 13208 6558 13242 6592
rect 13758 6558 13792 6592
rect -463 6527 -37 6544
rect 87 6527 513 6544
rect 637 6527 1063 6544
rect 1187 6527 1613 6544
rect 1737 6527 2163 6544
rect 2287 6527 2713 6544
rect 2837 6527 3263 6544
rect 3387 6527 3813 6544
rect 3937 6527 4363 6544
rect 4487 6527 4913 6544
rect 5037 6527 5463 6544
rect 5587 6527 6013 6544
rect 6137 6527 6563 6544
rect 6687 6527 7113 6544
rect 7237 6527 7663 6544
rect 7787 6527 8213 6544
rect 8337 6527 8763 6544
rect 8887 6527 9313 6544
rect 9437 6527 9863 6544
rect 9987 6527 10413 6544
rect 10537 6527 10963 6544
rect 11087 6527 11513 6544
rect 11637 6527 12063 6544
rect 12187 6527 12613 6544
rect 12737 6527 13163 6544
rect 13287 6527 13713 6544
rect -415 6453 -85 6465
rect -415 6147 -403 6453
rect -403 6147 -97 6453
rect -97 6147 -85 6453
rect -415 6135 -85 6147
rect -23 6087 -6 6513
rect 56 6087 73 6513
rect 527 6087 544 6513
rect 606 6087 623 6513
rect 685 6453 1015 6465
rect 685 6147 697 6453
rect 697 6147 1003 6453
rect 1003 6147 1015 6453
rect 685 6135 1015 6147
rect 1077 6087 1094 6513
rect 1156 6087 1173 6513
rect 1627 6087 1644 6513
rect 1706 6087 1723 6513
rect 1785 6453 2115 6465
rect 1785 6147 1797 6453
rect 1797 6147 2103 6453
rect 2103 6147 2115 6453
rect 1785 6135 2115 6147
rect 2177 6087 2194 6513
rect 2256 6087 2273 6513
rect 2727 6087 2744 6513
rect 2806 6087 2823 6513
rect 2885 6453 3215 6465
rect 2885 6147 2897 6453
rect 2897 6147 3203 6453
rect 3203 6147 3215 6453
rect 2885 6135 3215 6147
rect 3277 6087 3294 6513
rect 3356 6087 3373 6513
rect 3827 6087 3844 6513
rect 3906 6087 3923 6513
rect 3985 6453 4315 6465
rect 3985 6147 3997 6453
rect 3997 6147 4303 6453
rect 4303 6147 4315 6453
rect 3985 6135 4315 6147
rect 4377 6087 4394 6513
rect 4456 6087 4473 6513
rect 4927 6087 4944 6513
rect 5006 6087 5023 6513
rect 5085 6453 5415 6465
rect 5085 6147 5097 6453
rect 5097 6147 5403 6453
rect 5403 6147 5415 6453
rect 5085 6135 5415 6147
rect 5477 6087 5494 6513
rect 5556 6087 5573 6513
rect 6027 6087 6044 6513
rect 6106 6087 6123 6513
rect 6185 6453 6515 6465
rect 6185 6147 6197 6453
rect 6197 6147 6503 6453
rect 6503 6147 6515 6453
rect 6185 6135 6515 6147
rect 6577 6087 6594 6513
rect 6656 6087 6673 6513
rect 7127 6087 7144 6513
rect 7206 6087 7223 6513
rect 7285 6453 7615 6465
rect 7285 6147 7297 6453
rect 7297 6147 7603 6453
rect 7603 6147 7615 6453
rect 7285 6135 7615 6147
rect 7677 6087 7694 6513
rect 7756 6087 7773 6513
rect 8227 6087 8244 6513
rect 8306 6087 8323 6513
rect 8385 6453 8715 6465
rect 8385 6147 8397 6453
rect 8397 6147 8703 6453
rect 8703 6147 8715 6453
rect 8385 6135 8715 6147
rect 8777 6087 8794 6513
rect 8856 6087 8873 6513
rect 9327 6087 9344 6513
rect 9406 6087 9423 6513
rect 9485 6453 9815 6465
rect 9485 6147 9497 6453
rect 9497 6147 9803 6453
rect 9803 6147 9815 6453
rect 9485 6135 9815 6147
rect 9877 6087 9894 6513
rect 9956 6087 9973 6513
rect 10427 6087 10444 6513
rect 10506 6087 10523 6513
rect 10585 6453 10915 6465
rect 10585 6147 10597 6453
rect 10597 6147 10903 6453
rect 10903 6147 10915 6453
rect 10585 6135 10915 6147
rect 10977 6087 10994 6513
rect 11056 6087 11073 6513
rect 11527 6087 11544 6513
rect 11606 6087 11623 6513
rect 11685 6453 12015 6465
rect 11685 6147 11697 6453
rect 11697 6147 12003 6453
rect 12003 6147 12015 6453
rect 11685 6135 12015 6147
rect 12077 6087 12094 6513
rect 12156 6087 12173 6513
rect 12627 6087 12644 6513
rect 12706 6087 12723 6513
rect 12785 6453 13115 6465
rect 12785 6147 12797 6453
rect 12797 6147 13103 6453
rect 13103 6147 13115 6453
rect 12785 6135 13115 6147
rect 13177 6087 13194 6513
rect 13256 6087 13273 6513
rect -463 6056 -37 6073
rect 87 6056 513 6073
rect 637 6056 1063 6073
rect 1187 6056 1613 6073
rect 1737 6056 2163 6073
rect 2287 6056 2713 6073
rect 2837 6056 3263 6073
rect 3387 6056 3813 6073
rect 3937 6056 4363 6073
rect 4487 6056 4913 6073
rect 5037 6056 5463 6073
rect 5587 6056 6013 6073
rect 6137 6056 6563 6073
rect 6687 6056 7113 6073
rect 7237 6056 7663 6073
rect 7787 6056 8213 6073
rect 8337 6056 8763 6073
rect 8887 6056 9313 6073
rect 9437 6056 9863 6073
rect 9987 6056 10413 6073
rect 10537 6056 10963 6073
rect 11087 6056 11513 6073
rect 11637 6056 12063 6073
rect 12187 6056 12613 6073
rect 12737 6056 13163 6073
rect 13287 6056 13713 6073
rect 13987 6069 14263 6600
rect -1013 5519 -737 6050
rect -542 6008 -508 6042
rect 8 6008 42 6042
rect 558 6008 592 6042
rect 1108 6008 1142 6042
rect 1658 6008 1692 6042
rect 2208 6008 2242 6042
rect 2758 6008 2792 6042
rect 3308 6008 3342 6042
rect 3858 6008 3892 6042
rect 4408 6008 4442 6042
rect 4958 6008 4992 6042
rect 5508 6008 5542 6042
rect 6058 6008 6092 6042
rect 6608 6008 6642 6042
rect 7158 6008 7192 6042
rect 7708 6008 7742 6042
rect 8258 6008 8292 6042
rect 8808 6008 8842 6042
rect 9358 6008 9392 6042
rect 9908 6008 9942 6042
rect 10458 6008 10492 6042
rect 11008 6008 11042 6042
rect 11558 6008 11592 6042
rect 12108 6008 12142 6042
rect 12658 6008 12692 6042
rect 13208 6008 13242 6042
rect 13758 6008 13792 6042
rect -463 5977 -37 5994
rect 87 5977 513 5994
rect 637 5977 1063 5994
rect 1187 5977 1613 5994
rect 1737 5977 2163 5994
rect 2287 5977 2713 5994
rect 2837 5977 3263 5994
rect 3387 5977 3813 5994
rect 3937 5977 4363 5994
rect 4487 5977 4913 5994
rect 5037 5977 5463 5994
rect 5587 5977 6013 5994
rect 6137 5977 6563 5994
rect 6687 5977 7113 5994
rect 7237 5977 7663 5994
rect 7787 5977 8213 5994
rect 8337 5977 8763 5994
rect 8887 5977 9313 5994
rect 9437 5977 9863 5994
rect 9987 5977 10413 5994
rect 10537 5977 10963 5994
rect 11087 5977 11513 5994
rect 11637 5977 12063 5994
rect 12187 5977 12613 5994
rect 12737 5977 13163 5994
rect 13287 5977 13713 5994
rect -23 5537 -6 5963
rect 56 5537 73 5963
rect 135 5903 465 5915
rect 135 5597 147 5903
rect 147 5597 453 5903
rect 453 5597 465 5903
rect 135 5585 465 5597
rect 527 5537 544 5963
rect 606 5537 623 5963
rect 1077 5537 1094 5963
rect 1156 5537 1173 5963
rect 1235 5903 1565 5915
rect 1235 5597 1247 5903
rect 1247 5597 1553 5903
rect 1553 5597 1565 5903
rect 1235 5585 1565 5597
rect 1627 5537 1644 5963
rect 1706 5537 1723 5963
rect 2177 5537 2194 5963
rect 2256 5537 2273 5963
rect 2335 5903 2665 5915
rect 2335 5597 2347 5903
rect 2347 5597 2653 5903
rect 2653 5597 2665 5903
rect 2335 5585 2665 5597
rect 2727 5537 2744 5963
rect 2806 5537 2823 5963
rect 3277 5537 3294 5963
rect 3356 5537 3373 5963
rect 3435 5903 3765 5915
rect 3435 5597 3447 5903
rect 3447 5597 3753 5903
rect 3753 5597 3765 5903
rect 3435 5585 3765 5597
rect 3827 5537 3844 5963
rect 3906 5537 3923 5963
rect 4377 5537 4394 5963
rect 4456 5537 4473 5963
rect 4535 5903 4865 5915
rect 4535 5597 4547 5903
rect 4547 5597 4853 5903
rect 4853 5597 4865 5903
rect 4535 5585 4865 5597
rect 4927 5537 4944 5963
rect 5006 5537 5023 5963
rect 5477 5537 5494 5963
rect 5556 5537 5573 5963
rect 5635 5903 5965 5915
rect 5635 5597 5647 5903
rect 5647 5597 5953 5903
rect 5953 5597 5965 5903
rect 5635 5585 5965 5597
rect 6027 5537 6044 5963
rect 6106 5537 6123 5963
rect 6577 5537 6594 5963
rect 6656 5537 6673 5963
rect 6735 5903 7065 5915
rect 6735 5597 6747 5903
rect 6747 5597 7053 5903
rect 7053 5597 7065 5903
rect 6735 5585 7065 5597
rect 7127 5537 7144 5963
rect 7206 5537 7223 5963
rect 7677 5537 7694 5963
rect 7756 5537 7773 5963
rect 7835 5903 8165 5915
rect 7835 5597 7847 5903
rect 7847 5597 8153 5903
rect 8153 5597 8165 5903
rect 7835 5585 8165 5597
rect 8227 5537 8244 5963
rect 8306 5537 8323 5963
rect 8777 5537 8794 5963
rect 8856 5537 8873 5963
rect 8935 5903 9265 5915
rect 8935 5597 8947 5903
rect 8947 5597 9253 5903
rect 9253 5597 9265 5903
rect 8935 5585 9265 5597
rect 9327 5537 9344 5963
rect 9406 5537 9423 5963
rect 9877 5537 9894 5963
rect 9956 5537 9973 5963
rect 10035 5903 10365 5915
rect 10035 5597 10047 5903
rect 10047 5597 10353 5903
rect 10353 5597 10365 5903
rect 10035 5585 10365 5597
rect 10427 5537 10444 5963
rect 10506 5537 10523 5963
rect 10977 5537 10994 5963
rect 11056 5537 11073 5963
rect 11135 5903 11465 5915
rect 11135 5597 11147 5903
rect 11147 5597 11453 5903
rect 11453 5597 11465 5903
rect 11135 5585 11465 5597
rect 11527 5537 11544 5963
rect 11606 5537 11623 5963
rect 12077 5537 12094 5963
rect 12156 5537 12173 5963
rect 12235 5903 12565 5915
rect 12235 5597 12247 5903
rect 12247 5597 12553 5903
rect 12553 5597 12565 5903
rect 12235 5585 12565 5597
rect 12627 5537 12644 5963
rect 12706 5537 12723 5963
rect 13177 5537 13194 5963
rect 13256 5537 13273 5963
rect 13335 5903 13665 5915
rect 13335 5597 13347 5903
rect 13347 5597 13653 5903
rect 13653 5597 13665 5903
rect 13335 5585 13665 5597
rect -463 5506 -37 5523
rect 87 5506 513 5523
rect 637 5506 1063 5523
rect 1187 5506 1613 5523
rect 1737 5506 2163 5523
rect 2287 5506 2713 5523
rect 2837 5506 3263 5523
rect 3387 5506 3813 5523
rect 3937 5506 4363 5523
rect 4487 5506 4913 5523
rect 5037 5506 5463 5523
rect 5587 5506 6013 5523
rect 6137 5506 6563 5523
rect 6687 5506 7113 5523
rect 7237 5506 7663 5523
rect 7787 5506 8213 5523
rect 8337 5506 8763 5523
rect 8887 5506 9313 5523
rect 9437 5506 9863 5523
rect 9987 5506 10413 5523
rect 10537 5506 10963 5523
rect 11087 5506 11513 5523
rect 11637 5506 12063 5523
rect 12187 5506 12613 5523
rect 12737 5506 13163 5523
rect 13287 5506 13713 5523
rect 13987 5519 14263 6050
rect -1013 4969 -737 5500
rect -542 5458 -508 5492
rect 8 5458 42 5492
rect 558 5458 592 5492
rect 1108 5458 1142 5492
rect 1658 5458 1692 5492
rect 2208 5458 2242 5492
rect 2758 5458 2792 5492
rect 3308 5458 3342 5492
rect 3858 5458 3892 5492
rect 4408 5458 4442 5492
rect 4958 5458 4992 5492
rect 5508 5458 5542 5492
rect 6058 5458 6092 5492
rect 6608 5458 6642 5492
rect 7158 5458 7192 5492
rect 7708 5458 7742 5492
rect 8258 5458 8292 5492
rect 8808 5458 8842 5492
rect 9358 5458 9392 5492
rect 9908 5458 9942 5492
rect 10458 5458 10492 5492
rect 11008 5458 11042 5492
rect 11558 5458 11592 5492
rect 12108 5458 12142 5492
rect 12658 5458 12692 5492
rect 13208 5458 13242 5492
rect 13758 5458 13792 5492
rect -463 5427 -37 5444
rect 87 5427 513 5444
rect 637 5427 1063 5444
rect 1187 5427 1613 5444
rect 1737 5427 2163 5444
rect 2287 5427 2713 5444
rect 2837 5427 3263 5444
rect 3387 5427 3813 5444
rect 3937 5427 4363 5444
rect 4487 5427 4913 5444
rect 5037 5427 5463 5444
rect 5587 5427 6013 5444
rect 6137 5427 6563 5444
rect 6687 5427 7113 5444
rect 7237 5427 7663 5444
rect 7787 5427 8213 5444
rect 8337 5427 8763 5444
rect 8887 5427 9313 5444
rect 9437 5427 9863 5444
rect 9987 5427 10413 5444
rect 10537 5427 10963 5444
rect 11087 5427 11513 5444
rect 11637 5427 12063 5444
rect 12187 5427 12613 5444
rect 12737 5427 13163 5444
rect 13287 5427 13713 5444
rect -415 5353 -85 5365
rect -415 5047 -403 5353
rect -403 5047 -97 5353
rect -97 5047 -85 5353
rect -415 5035 -85 5047
rect -23 4987 -6 5413
rect 56 4987 73 5413
rect 527 4987 544 5413
rect 606 4987 623 5413
rect 685 5353 1015 5365
rect 685 5047 697 5353
rect 697 5047 1003 5353
rect 1003 5047 1015 5353
rect 685 5035 1015 5047
rect 1077 4987 1094 5413
rect 1156 4987 1173 5413
rect 1627 4987 1644 5413
rect 1706 4987 1723 5413
rect 1785 5353 2115 5365
rect 1785 5047 1797 5353
rect 1797 5047 2103 5353
rect 2103 5047 2115 5353
rect 1785 5035 2115 5047
rect 2177 4987 2194 5413
rect 2256 4987 2273 5413
rect 2727 4987 2744 5413
rect 2806 4987 2823 5413
rect 2885 5353 3215 5365
rect 2885 5047 2897 5353
rect 2897 5047 3203 5353
rect 3203 5047 3215 5353
rect 2885 5035 3215 5047
rect 3277 4987 3294 5413
rect 3356 4987 3373 5413
rect 3827 4987 3844 5413
rect 3906 4987 3923 5413
rect 3985 5353 4315 5365
rect 3985 5047 3997 5353
rect 3997 5047 4303 5353
rect 4303 5047 4315 5353
rect 3985 5035 4315 5047
rect 4377 4987 4394 5413
rect 4456 4987 4473 5413
rect 4927 4987 4944 5413
rect 5006 4987 5023 5413
rect 5085 5353 5415 5365
rect 5085 5047 5097 5353
rect 5097 5047 5403 5353
rect 5403 5047 5415 5353
rect 5085 5035 5415 5047
rect 5477 4987 5494 5413
rect 5556 4987 5573 5413
rect 6027 4987 6044 5413
rect 6106 4987 6123 5413
rect 6185 5353 6515 5365
rect 6185 5047 6197 5353
rect 6197 5047 6503 5353
rect 6503 5047 6515 5353
rect 6185 5035 6515 5047
rect 6577 4987 6594 5413
rect 6656 4987 6673 5413
rect 7127 4987 7144 5413
rect 7206 4987 7223 5413
rect 7285 5353 7615 5365
rect 7285 5047 7297 5353
rect 7297 5047 7603 5353
rect 7603 5047 7615 5353
rect 7285 5035 7615 5047
rect 7677 4987 7694 5413
rect 7756 4987 7773 5413
rect 8227 4987 8244 5413
rect 8306 4987 8323 5413
rect 8385 5353 8715 5365
rect 8385 5047 8397 5353
rect 8397 5047 8703 5353
rect 8703 5047 8715 5353
rect 8385 5035 8715 5047
rect 8777 4987 8794 5413
rect 8856 4987 8873 5413
rect 9327 4987 9344 5413
rect 9406 4987 9423 5413
rect 9485 5353 9815 5365
rect 9485 5047 9497 5353
rect 9497 5047 9803 5353
rect 9803 5047 9815 5353
rect 9485 5035 9815 5047
rect 9877 4987 9894 5413
rect 9956 4987 9973 5413
rect 10427 4987 10444 5413
rect 10506 4987 10523 5413
rect 10585 5353 10915 5365
rect 10585 5047 10597 5353
rect 10597 5047 10903 5353
rect 10903 5047 10915 5353
rect 10585 5035 10915 5047
rect 10977 4987 10994 5413
rect 11056 4987 11073 5413
rect 11527 4987 11544 5413
rect 11606 4987 11623 5413
rect 11685 5353 12015 5365
rect 11685 5047 11697 5353
rect 11697 5047 12003 5353
rect 12003 5047 12015 5353
rect 11685 5035 12015 5047
rect 12077 4987 12094 5413
rect 12156 4987 12173 5413
rect 12627 4987 12644 5413
rect 12706 4987 12723 5413
rect 12785 5353 13115 5365
rect 12785 5047 12797 5353
rect 12797 5047 13103 5353
rect 13103 5047 13115 5353
rect 12785 5035 13115 5047
rect 13177 4987 13194 5413
rect 13256 4987 13273 5413
rect -463 4956 -37 4973
rect 87 4956 513 4973
rect 637 4956 1063 4973
rect 1187 4956 1613 4973
rect 1737 4956 2163 4973
rect 2287 4956 2713 4973
rect 2837 4956 3263 4973
rect 3387 4956 3813 4973
rect 3937 4956 4363 4973
rect 4487 4956 4913 4973
rect 5037 4956 5463 4973
rect 5587 4956 6013 4973
rect 6137 4956 6563 4973
rect 6687 4956 7113 4973
rect 7237 4956 7663 4973
rect 7787 4956 8213 4973
rect 8337 4956 8763 4973
rect 8887 4956 9313 4973
rect 9437 4956 9863 4973
rect 9987 4956 10413 4973
rect 10537 4956 10963 4973
rect 11087 4956 11513 4973
rect 11637 4956 12063 4973
rect 12187 4956 12613 4973
rect 12737 4956 13163 4973
rect 13287 4956 13713 4973
rect 13987 4969 14263 5500
rect -1013 4419 -737 4950
rect -542 4908 -508 4942
rect 8 4908 42 4942
rect 558 4908 592 4942
rect 1108 4908 1142 4942
rect 1658 4908 1692 4942
rect 2208 4908 2242 4942
rect 2758 4908 2792 4942
rect 3308 4908 3342 4942
rect 3858 4908 3892 4942
rect 4408 4908 4442 4942
rect 4958 4908 4992 4942
rect 5508 4908 5542 4942
rect 6058 4908 6092 4942
rect 6608 4908 6642 4942
rect 7158 4908 7192 4942
rect 7708 4908 7742 4942
rect 8258 4908 8292 4942
rect 8808 4908 8842 4942
rect 9358 4908 9392 4942
rect 9908 4908 9942 4942
rect 10458 4908 10492 4942
rect 11008 4908 11042 4942
rect 11558 4908 11592 4942
rect 12108 4908 12142 4942
rect 12658 4908 12692 4942
rect 13208 4908 13242 4942
rect 13758 4908 13792 4942
rect -463 4877 -37 4894
rect 87 4877 513 4894
rect 637 4877 1063 4894
rect 1187 4877 1613 4894
rect 1737 4877 2163 4894
rect 2287 4877 2713 4894
rect 2837 4877 3263 4894
rect 3387 4877 3813 4894
rect 3937 4877 4363 4894
rect 4487 4877 4913 4894
rect 5037 4877 5463 4894
rect 5587 4877 6013 4894
rect 6137 4877 6563 4894
rect 6687 4877 7113 4894
rect 7237 4877 7663 4894
rect 7787 4877 8213 4894
rect 8337 4877 8763 4894
rect 8887 4877 9313 4894
rect 9437 4877 9863 4894
rect 9987 4877 10413 4894
rect 10537 4877 10963 4894
rect 11087 4877 11513 4894
rect 11637 4877 12063 4894
rect 12187 4877 12613 4894
rect 12737 4877 13163 4894
rect 13287 4877 13713 4894
rect -23 4437 -6 4863
rect 56 4437 73 4863
rect 135 4803 465 4815
rect 135 4497 147 4803
rect 147 4497 453 4803
rect 453 4497 465 4803
rect 135 4485 465 4497
rect 527 4437 544 4863
rect 606 4437 623 4863
rect 1077 4437 1094 4863
rect 1156 4437 1173 4863
rect 1235 4803 1565 4815
rect 1235 4497 1247 4803
rect 1247 4497 1553 4803
rect 1553 4497 1565 4803
rect 1235 4485 1565 4497
rect 1627 4437 1644 4863
rect 1706 4437 1723 4863
rect 2177 4437 2194 4863
rect 2256 4437 2273 4863
rect 2335 4803 2665 4815
rect 2335 4497 2347 4803
rect 2347 4497 2653 4803
rect 2653 4497 2665 4803
rect 2335 4485 2665 4497
rect 2727 4437 2744 4863
rect 2806 4437 2823 4863
rect 3277 4437 3294 4863
rect 3356 4437 3373 4863
rect 3435 4803 3765 4815
rect 3435 4497 3447 4803
rect 3447 4497 3753 4803
rect 3753 4497 3765 4803
rect 3435 4485 3765 4497
rect 3827 4437 3844 4863
rect 3906 4437 3923 4863
rect 4377 4437 4394 4863
rect 4456 4437 4473 4863
rect 4535 4803 4865 4815
rect 4535 4497 4547 4803
rect 4547 4497 4853 4803
rect 4853 4497 4865 4803
rect 4535 4485 4865 4497
rect 4927 4437 4944 4863
rect 5006 4437 5023 4863
rect 5477 4437 5494 4863
rect 5556 4437 5573 4863
rect 5635 4803 5965 4815
rect 5635 4497 5647 4803
rect 5647 4497 5953 4803
rect 5953 4497 5965 4803
rect 5635 4485 5965 4497
rect 6027 4437 6044 4863
rect 6106 4437 6123 4863
rect 6577 4437 6594 4863
rect 6656 4437 6673 4863
rect 6735 4803 7065 4815
rect 6735 4497 6747 4803
rect 6747 4497 7053 4803
rect 7053 4497 7065 4803
rect 6735 4485 7065 4497
rect 7127 4437 7144 4863
rect 7206 4437 7223 4863
rect 7677 4437 7694 4863
rect 7756 4437 7773 4863
rect 7835 4803 8165 4815
rect 7835 4497 7847 4803
rect 7847 4497 8153 4803
rect 8153 4497 8165 4803
rect 7835 4485 8165 4497
rect 8227 4437 8244 4863
rect 8306 4437 8323 4863
rect 8777 4437 8794 4863
rect 8856 4437 8873 4863
rect 8935 4803 9265 4815
rect 8935 4497 8947 4803
rect 8947 4497 9253 4803
rect 9253 4497 9265 4803
rect 8935 4485 9265 4497
rect 9327 4437 9344 4863
rect 9406 4437 9423 4863
rect 9877 4437 9894 4863
rect 9956 4437 9973 4863
rect 10035 4803 10365 4815
rect 10035 4497 10047 4803
rect 10047 4497 10353 4803
rect 10353 4497 10365 4803
rect 10035 4485 10365 4497
rect 10427 4437 10444 4863
rect 10506 4437 10523 4863
rect 10977 4437 10994 4863
rect 11056 4437 11073 4863
rect 11135 4803 11465 4815
rect 11135 4497 11147 4803
rect 11147 4497 11453 4803
rect 11453 4497 11465 4803
rect 11135 4485 11465 4497
rect 11527 4437 11544 4863
rect 11606 4437 11623 4863
rect 12077 4437 12094 4863
rect 12156 4437 12173 4863
rect 12235 4803 12565 4815
rect 12235 4497 12247 4803
rect 12247 4497 12553 4803
rect 12553 4497 12565 4803
rect 12235 4485 12565 4497
rect 12627 4437 12644 4863
rect 12706 4437 12723 4863
rect 13177 4437 13194 4863
rect 13256 4437 13273 4863
rect 13335 4803 13665 4815
rect 13335 4497 13347 4803
rect 13347 4497 13653 4803
rect 13653 4497 13665 4803
rect 13335 4485 13665 4497
rect -463 4406 -37 4423
rect 87 4406 513 4423
rect 637 4406 1063 4423
rect 1187 4406 1613 4423
rect 1737 4406 2163 4423
rect 2287 4406 2713 4423
rect 2837 4406 3263 4423
rect 3387 4406 3813 4423
rect 3937 4406 4363 4423
rect 4487 4406 4913 4423
rect 5037 4406 5463 4423
rect 5587 4406 6013 4423
rect 6137 4406 6563 4423
rect 6687 4406 7113 4423
rect 7237 4406 7663 4423
rect 7787 4406 8213 4423
rect 8337 4406 8763 4423
rect 8887 4406 9313 4423
rect 9437 4406 9863 4423
rect 9987 4406 10413 4423
rect 10537 4406 10963 4423
rect 11087 4406 11513 4423
rect 11637 4406 12063 4423
rect 12187 4406 12613 4423
rect 12737 4406 13163 4423
rect 13287 4406 13713 4423
rect 13987 4419 14263 4950
rect -1013 3869 -737 4400
rect -542 4358 -508 4392
rect 8 4358 42 4392
rect 558 4358 592 4392
rect 1108 4358 1142 4392
rect 1658 4358 1692 4392
rect 2208 4358 2242 4392
rect 2758 4358 2792 4392
rect 3308 4358 3342 4392
rect 3858 4358 3892 4392
rect 4408 4358 4442 4392
rect 4958 4358 4992 4392
rect 5508 4358 5542 4392
rect 6058 4358 6092 4392
rect 6608 4358 6642 4392
rect 7158 4358 7192 4392
rect 7708 4358 7742 4392
rect 8258 4358 8292 4392
rect 8808 4358 8842 4392
rect 9358 4358 9392 4392
rect 9908 4358 9942 4392
rect 10458 4358 10492 4392
rect 11008 4358 11042 4392
rect 11558 4358 11592 4392
rect 12108 4358 12142 4392
rect 12658 4358 12692 4392
rect 13208 4358 13242 4392
rect 13758 4358 13792 4392
rect -463 4327 -37 4344
rect 87 4327 513 4344
rect 637 4327 1063 4344
rect 1187 4327 1613 4344
rect 1737 4327 2163 4344
rect 2287 4327 2713 4344
rect 2837 4327 3263 4344
rect 3387 4327 3813 4344
rect 3937 4327 4363 4344
rect 4487 4327 4913 4344
rect 5037 4327 5463 4344
rect 5587 4327 6013 4344
rect 6137 4327 6563 4344
rect 6687 4327 7113 4344
rect 7237 4327 7663 4344
rect 7787 4327 8213 4344
rect 8337 4327 8763 4344
rect 8887 4327 9313 4344
rect 9437 4327 9863 4344
rect 9987 4327 10413 4344
rect 10537 4327 10963 4344
rect 11087 4327 11513 4344
rect 11637 4327 12063 4344
rect 12187 4327 12613 4344
rect 12737 4327 13163 4344
rect 13287 4327 13713 4344
rect -415 4253 -85 4265
rect -415 3947 -403 4253
rect -403 3947 -97 4253
rect -97 3947 -85 4253
rect -415 3935 -85 3947
rect -23 3887 -6 4313
rect 56 3887 73 4313
rect 527 3887 544 4313
rect 606 3887 623 4313
rect 685 4253 1015 4265
rect 685 3947 697 4253
rect 697 3947 1003 4253
rect 1003 3947 1015 4253
rect 685 3935 1015 3947
rect 1077 3887 1094 4313
rect 1156 3887 1173 4313
rect 1627 3887 1644 4313
rect 1706 3887 1723 4313
rect 1785 4253 2115 4265
rect 1785 3947 1797 4253
rect 1797 3947 2103 4253
rect 2103 3947 2115 4253
rect 1785 3935 2115 3947
rect 2177 3887 2194 4313
rect 2256 3887 2273 4313
rect 2727 3887 2744 4313
rect 2806 3887 2823 4313
rect 2885 4253 3215 4265
rect 2885 3947 2897 4253
rect 2897 3947 3203 4253
rect 3203 3947 3215 4253
rect 2885 3935 3215 3947
rect 3277 3887 3294 4313
rect 3356 3887 3373 4313
rect 3827 3887 3844 4313
rect 3906 3887 3923 4313
rect 3985 4253 4315 4265
rect 3985 3947 3997 4253
rect 3997 3947 4303 4253
rect 4303 3947 4315 4253
rect 3985 3935 4315 3947
rect 4377 3887 4394 4313
rect 4456 3887 4473 4313
rect 4927 3887 4944 4313
rect 5006 3887 5023 4313
rect 5085 4253 5415 4265
rect 5085 3947 5097 4253
rect 5097 3947 5403 4253
rect 5403 3947 5415 4253
rect 5085 3935 5415 3947
rect 5477 3887 5494 4313
rect 5556 3887 5573 4313
rect 6027 3887 6044 4313
rect 6106 3887 6123 4313
rect 6185 4253 6515 4265
rect 6185 3947 6197 4253
rect 6197 3947 6503 4253
rect 6503 3947 6515 4253
rect 6185 3935 6515 3947
rect 6577 3887 6594 4313
rect 6656 3887 6673 4313
rect 7127 3887 7144 4313
rect 7206 3887 7223 4313
rect 7285 4253 7615 4265
rect 7285 3947 7297 4253
rect 7297 3947 7603 4253
rect 7603 3947 7615 4253
rect 7285 3935 7615 3947
rect 7677 3887 7694 4313
rect 7756 3887 7773 4313
rect 8227 3887 8244 4313
rect 8306 3887 8323 4313
rect 8385 4253 8715 4265
rect 8385 3947 8397 4253
rect 8397 3947 8703 4253
rect 8703 3947 8715 4253
rect 8385 3935 8715 3947
rect 8777 3887 8794 4313
rect 8856 3887 8873 4313
rect 9327 3887 9344 4313
rect 9406 3887 9423 4313
rect 9485 4253 9815 4265
rect 9485 3947 9497 4253
rect 9497 3947 9803 4253
rect 9803 3947 9815 4253
rect 9485 3935 9815 3947
rect 9877 3887 9894 4313
rect 9956 3887 9973 4313
rect 10427 3887 10444 4313
rect 10506 3887 10523 4313
rect 10585 4253 10915 4265
rect 10585 3947 10597 4253
rect 10597 3947 10903 4253
rect 10903 3947 10915 4253
rect 10585 3935 10915 3947
rect 10977 3887 10994 4313
rect 11056 3887 11073 4313
rect 11527 3887 11544 4313
rect 11606 3887 11623 4313
rect 11685 4253 12015 4265
rect 11685 3947 11697 4253
rect 11697 3947 12003 4253
rect 12003 3947 12015 4253
rect 11685 3935 12015 3947
rect 12077 3887 12094 4313
rect 12156 3887 12173 4313
rect 12627 3887 12644 4313
rect 12706 3887 12723 4313
rect 12785 4253 13115 4265
rect 12785 3947 12797 4253
rect 12797 3947 13103 4253
rect 13103 3947 13115 4253
rect 12785 3935 13115 3947
rect 13177 3887 13194 4313
rect 13256 3887 13273 4313
rect -463 3856 -37 3873
rect 87 3856 513 3873
rect 637 3856 1063 3873
rect 1187 3856 1613 3873
rect 1737 3856 2163 3873
rect 2287 3856 2713 3873
rect 2837 3856 3263 3873
rect 3387 3856 3813 3873
rect 3937 3856 4363 3873
rect 4487 3856 4913 3873
rect 5037 3856 5463 3873
rect 5587 3856 6013 3873
rect 6137 3856 6563 3873
rect 6687 3856 7113 3873
rect 7237 3856 7663 3873
rect 7787 3856 8213 3873
rect 8337 3856 8763 3873
rect 8887 3856 9313 3873
rect 9437 3856 9863 3873
rect 9987 3856 10413 3873
rect 10537 3856 10963 3873
rect 11087 3856 11513 3873
rect 11637 3856 12063 3873
rect 12187 3856 12613 3873
rect 12737 3856 13163 3873
rect 13287 3856 13713 3873
rect 13987 3869 14263 4400
rect -1013 3319 -737 3850
rect -542 3808 -508 3842
rect 8 3808 42 3842
rect 558 3808 592 3842
rect 1108 3808 1142 3842
rect 1658 3808 1692 3842
rect 2208 3808 2242 3842
rect 2758 3808 2792 3842
rect 3308 3808 3342 3842
rect 3858 3808 3892 3842
rect 4408 3808 4442 3842
rect 4958 3808 4992 3842
rect 5508 3808 5542 3842
rect 6058 3808 6092 3842
rect 6608 3808 6642 3842
rect 7158 3808 7192 3842
rect 7708 3808 7742 3842
rect 8258 3808 8292 3842
rect 8808 3808 8842 3842
rect 9358 3808 9392 3842
rect 9908 3808 9942 3842
rect 10458 3808 10492 3842
rect 11008 3808 11042 3842
rect 11558 3808 11592 3842
rect 12108 3808 12142 3842
rect 12658 3808 12692 3842
rect 13208 3808 13242 3842
rect 13758 3808 13792 3842
rect -463 3777 -37 3794
rect 87 3777 513 3794
rect 637 3777 1063 3794
rect 1187 3777 1613 3794
rect 1737 3777 2163 3794
rect 2287 3777 2713 3794
rect 2837 3777 3263 3794
rect 3387 3777 3813 3794
rect 3937 3777 4363 3794
rect 4487 3777 4913 3794
rect 5037 3777 5463 3794
rect 5587 3777 6013 3794
rect 6137 3777 6563 3794
rect 6687 3777 7113 3794
rect 7237 3777 7663 3794
rect 7787 3777 8213 3794
rect 8337 3777 8763 3794
rect 8887 3777 9313 3794
rect 9437 3777 9863 3794
rect 9987 3777 10413 3794
rect 10537 3777 10963 3794
rect 11087 3777 11513 3794
rect 11637 3777 12063 3794
rect 12187 3777 12613 3794
rect 12737 3777 13163 3794
rect 13287 3777 13713 3794
rect -23 3337 -6 3763
rect 56 3337 73 3763
rect 135 3703 465 3715
rect 135 3397 147 3703
rect 147 3397 453 3703
rect 453 3397 465 3703
rect 135 3385 465 3397
rect 527 3337 544 3763
rect 606 3337 623 3763
rect 1077 3337 1094 3763
rect 1156 3337 1173 3763
rect 1235 3703 1565 3715
rect 1235 3397 1247 3703
rect 1247 3397 1553 3703
rect 1553 3397 1565 3703
rect 1235 3385 1565 3397
rect 1627 3337 1644 3763
rect 1706 3337 1723 3763
rect 2177 3337 2194 3763
rect 2256 3337 2273 3763
rect 2335 3703 2665 3715
rect 2335 3397 2347 3703
rect 2347 3397 2653 3703
rect 2653 3397 2665 3703
rect 2335 3385 2665 3397
rect 2727 3337 2744 3763
rect 2806 3337 2823 3763
rect 3277 3337 3294 3763
rect 3356 3337 3373 3763
rect 3435 3703 3765 3715
rect 3435 3397 3447 3703
rect 3447 3397 3753 3703
rect 3753 3397 3765 3703
rect 3435 3385 3765 3397
rect 3827 3337 3844 3763
rect 3906 3337 3923 3763
rect 4377 3337 4394 3763
rect 4456 3337 4473 3763
rect 4535 3703 4865 3715
rect 4535 3397 4547 3703
rect 4547 3397 4853 3703
rect 4853 3397 4865 3703
rect 4535 3385 4865 3397
rect 4927 3337 4944 3763
rect 5006 3337 5023 3763
rect 5477 3337 5494 3763
rect 5556 3337 5573 3763
rect 5635 3703 5965 3715
rect 5635 3397 5647 3703
rect 5647 3397 5953 3703
rect 5953 3397 5965 3703
rect 5635 3385 5965 3397
rect 6027 3337 6044 3763
rect 6106 3337 6123 3763
rect 6577 3337 6594 3763
rect 6656 3337 6673 3763
rect 6735 3703 7065 3715
rect 6735 3397 6747 3703
rect 6747 3397 7053 3703
rect 7053 3397 7065 3703
rect 6735 3385 7065 3397
rect 7127 3337 7144 3763
rect 7206 3337 7223 3763
rect 7677 3337 7694 3763
rect 7756 3337 7773 3763
rect 7835 3703 8165 3715
rect 7835 3397 7847 3703
rect 7847 3397 8153 3703
rect 8153 3397 8165 3703
rect 7835 3385 8165 3397
rect 8227 3337 8244 3763
rect 8306 3337 8323 3763
rect 8777 3337 8794 3763
rect 8856 3337 8873 3763
rect 8935 3703 9265 3715
rect 8935 3397 8947 3703
rect 8947 3397 9253 3703
rect 9253 3397 9265 3703
rect 8935 3385 9265 3397
rect 9327 3337 9344 3763
rect 9406 3337 9423 3763
rect 9877 3337 9894 3763
rect 9956 3337 9973 3763
rect 10035 3703 10365 3715
rect 10035 3397 10047 3703
rect 10047 3397 10353 3703
rect 10353 3397 10365 3703
rect 10035 3385 10365 3397
rect 10427 3337 10444 3763
rect 10506 3337 10523 3763
rect 10977 3337 10994 3763
rect 11056 3337 11073 3763
rect 11135 3703 11465 3715
rect 11135 3397 11147 3703
rect 11147 3397 11453 3703
rect 11453 3397 11465 3703
rect 11135 3385 11465 3397
rect 11527 3337 11544 3763
rect 11606 3337 11623 3763
rect 12077 3337 12094 3763
rect 12156 3337 12173 3763
rect 12235 3703 12565 3715
rect 12235 3397 12247 3703
rect 12247 3397 12553 3703
rect 12553 3397 12565 3703
rect 12235 3385 12565 3397
rect 12627 3337 12644 3763
rect 12706 3337 12723 3763
rect 13177 3337 13194 3763
rect 13256 3337 13273 3763
rect 13335 3703 13665 3715
rect 13335 3397 13347 3703
rect 13347 3397 13653 3703
rect 13653 3397 13665 3703
rect 13335 3385 13665 3397
rect -463 3306 -37 3323
rect 87 3306 513 3323
rect 637 3306 1063 3323
rect 1187 3306 1613 3323
rect 1737 3306 2163 3323
rect 2287 3306 2713 3323
rect 2837 3306 3263 3323
rect 3387 3306 3813 3323
rect 3937 3306 4363 3323
rect 4487 3306 4913 3323
rect 5037 3306 5463 3323
rect 5587 3306 6013 3323
rect 6137 3306 6563 3323
rect 6687 3306 7113 3323
rect 7237 3306 7663 3323
rect 7787 3306 8213 3323
rect 8337 3306 8763 3323
rect 8887 3306 9313 3323
rect 9437 3306 9863 3323
rect 9987 3306 10413 3323
rect 10537 3306 10963 3323
rect 11087 3306 11513 3323
rect 11637 3306 12063 3323
rect 12187 3306 12613 3323
rect 12737 3306 13163 3323
rect 13287 3306 13713 3323
rect 13987 3319 14263 3850
rect -1013 2769 -737 3300
rect -542 3258 -508 3292
rect 8 3258 42 3292
rect 558 3258 592 3292
rect 1108 3258 1142 3292
rect 1658 3258 1692 3292
rect 2208 3258 2242 3292
rect 2758 3258 2792 3292
rect 3308 3258 3342 3292
rect 3858 3258 3892 3292
rect 4408 3258 4442 3292
rect 4958 3258 4992 3292
rect 5508 3258 5542 3292
rect 6058 3258 6092 3292
rect 6608 3258 6642 3292
rect 7158 3258 7192 3292
rect 7708 3258 7742 3292
rect 8258 3258 8292 3292
rect 8808 3258 8842 3292
rect 9358 3258 9392 3292
rect 9908 3258 9942 3292
rect 10458 3258 10492 3292
rect 11008 3258 11042 3292
rect 11558 3258 11592 3292
rect 12108 3258 12142 3292
rect 12658 3258 12692 3292
rect 13208 3258 13242 3292
rect 13758 3258 13792 3292
rect -463 3227 -37 3244
rect 87 3227 513 3244
rect 637 3227 1063 3244
rect 1187 3227 1613 3244
rect 1737 3227 2163 3244
rect 2287 3227 2713 3244
rect 2837 3227 3263 3244
rect 3387 3227 3813 3244
rect 3937 3227 4363 3244
rect 4487 3227 4913 3244
rect 5037 3227 5463 3244
rect 5587 3227 6013 3244
rect 6137 3227 6563 3244
rect 6687 3227 7113 3244
rect 7237 3227 7663 3244
rect 7787 3227 8213 3244
rect 8337 3227 8763 3244
rect 8887 3227 9313 3244
rect 9437 3227 9863 3244
rect 9987 3227 10413 3244
rect 10537 3227 10963 3244
rect 11087 3227 11513 3244
rect 11637 3227 12063 3244
rect 12187 3227 12613 3244
rect 12737 3227 13163 3244
rect 13287 3227 13713 3244
rect -415 3153 -85 3165
rect -415 2847 -403 3153
rect -403 2847 -97 3153
rect -97 2847 -85 3153
rect -415 2835 -85 2847
rect -23 2787 -6 3213
rect 56 2787 73 3213
rect 527 2787 544 3213
rect 606 2787 623 3213
rect 685 3153 1015 3165
rect 685 2847 697 3153
rect 697 2847 1003 3153
rect 1003 2847 1015 3153
rect 685 2835 1015 2847
rect 1077 2787 1094 3213
rect 1156 2787 1173 3213
rect 1627 2787 1644 3213
rect 1706 2787 1723 3213
rect 1785 3153 2115 3165
rect 1785 2847 1797 3153
rect 1797 2847 2103 3153
rect 2103 2847 2115 3153
rect 1785 2835 2115 2847
rect 2177 2787 2194 3213
rect 2256 2787 2273 3213
rect 2727 2787 2744 3213
rect 2806 2787 2823 3213
rect 2885 3153 3215 3165
rect 2885 2847 2897 3153
rect 2897 2847 3203 3153
rect 3203 2847 3215 3153
rect 2885 2835 3215 2847
rect 3277 2787 3294 3213
rect 3356 2787 3373 3213
rect 3827 2787 3844 3213
rect 3906 2787 3923 3213
rect 3985 3153 4315 3165
rect 3985 2847 3997 3153
rect 3997 2847 4303 3153
rect 4303 2847 4315 3153
rect 3985 2835 4315 2847
rect 4377 2787 4394 3213
rect 4456 2787 4473 3213
rect 4927 2787 4944 3213
rect 5006 2787 5023 3213
rect 5085 3153 5415 3165
rect 5085 2847 5097 3153
rect 5097 2847 5403 3153
rect 5403 2847 5415 3153
rect 5085 2835 5415 2847
rect 5477 2787 5494 3213
rect 5556 2787 5573 3213
rect 6027 2787 6044 3213
rect 6106 2787 6123 3213
rect 6185 3153 6515 3165
rect 6185 2847 6197 3153
rect 6197 2847 6503 3153
rect 6503 2847 6515 3153
rect 6185 2835 6515 2847
rect 6577 2787 6594 3213
rect 6656 2787 6673 3213
rect 7127 2787 7144 3213
rect 7206 2787 7223 3213
rect 7285 3153 7615 3165
rect 7285 2847 7297 3153
rect 7297 2847 7603 3153
rect 7603 2847 7615 3153
rect 7285 2835 7615 2847
rect 7677 2787 7694 3213
rect 7756 2787 7773 3213
rect 8227 2787 8244 3213
rect 8306 2787 8323 3213
rect 8385 3153 8715 3165
rect 8385 2847 8397 3153
rect 8397 2847 8703 3153
rect 8703 2847 8715 3153
rect 8385 2835 8715 2847
rect 8777 2787 8794 3213
rect 8856 2787 8873 3213
rect 9327 2787 9344 3213
rect 9406 2787 9423 3213
rect 9485 3153 9815 3165
rect 9485 2847 9497 3153
rect 9497 2847 9803 3153
rect 9803 2847 9815 3153
rect 9485 2835 9815 2847
rect 9877 2787 9894 3213
rect 9956 2787 9973 3213
rect 10427 2787 10444 3213
rect 10506 2787 10523 3213
rect 10585 3153 10915 3165
rect 10585 2847 10597 3153
rect 10597 2847 10903 3153
rect 10903 2847 10915 3153
rect 10585 2835 10915 2847
rect 10977 2787 10994 3213
rect 11056 2787 11073 3213
rect 11527 2787 11544 3213
rect 11606 2787 11623 3213
rect 11685 3153 12015 3165
rect 11685 2847 11697 3153
rect 11697 2847 12003 3153
rect 12003 2847 12015 3153
rect 11685 2835 12015 2847
rect 12077 2787 12094 3213
rect 12156 2787 12173 3213
rect 12627 2787 12644 3213
rect 12706 2787 12723 3213
rect 12785 3153 13115 3165
rect 12785 2847 12797 3153
rect 12797 2847 13103 3153
rect 13103 2847 13115 3153
rect 12785 2835 13115 2847
rect 13177 2787 13194 3213
rect 13256 2787 13273 3213
rect -463 2756 -37 2773
rect 87 2756 513 2773
rect 637 2756 1063 2773
rect 1187 2756 1613 2773
rect 1737 2756 2163 2773
rect 2287 2756 2713 2773
rect 2837 2756 3263 2773
rect 3387 2756 3813 2773
rect 3937 2756 4363 2773
rect 4487 2756 4913 2773
rect 5037 2756 5463 2773
rect 5587 2756 6013 2773
rect 6137 2756 6563 2773
rect 6687 2756 7113 2773
rect 7237 2756 7663 2773
rect 7787 2756 8213 2773
rect 8337 2756 8763 2773
rect 8887 2756 9313 2773
rect 9437 2756 9863 2773
rect 9987 2756 10413 2773
rect 10537 2756 10963 2773
rect 11087 2756 11513 2773
rect 11637 2756 12063 2773
rect 12187 2756 12613 2773
rect 12737 2756 13163 2773
rect 13287 2756 13713 2773
rect 13987 2769 14263 3300
rect -1013 2219 -737 2750
rect -542 2708 -508 2742
rect 8 2708 42 2742
rect 558 2708 592 2742
rect 1108 2708 1142 2742
rect 1658 2708 1692 2742
rect 2208 2708 2242 2742
rect 2758 2708 2792 2742
rect 3308 2708 3342 2742
rect 3858 2708 3892 2742
rect 4408 2708 4442 2742
rect 4958 2708 4992 2742
rect 5508 2708 5542 2742
rect 6058 2708 6092 2742
rect 6608 2708 6642 2742
rect 7158 2708 7192 2742
rect 7708 2708 7742 2742
rect 8258 2708 8292 2742
rect 8808 2708 8842 2742
rect 9358 2708 9392 2742
rect 9908 2708 9942 2742
rect 10458 2708 10492 2742
rect 11008 2708 11042 2742
rect 11558 2708 11592 2742
rect 12108 2708 12142 2742
rect 12658 2708 12692 2742
rect 13208 2708 13242 2742
rect 13758 2708 13792 2742
rect -463 2677 -37 2694
rect 87 2677 513 2694
rect 637 2677 1063 2694
rect 1187 2677 1613 2694
rect 1737 2677 2163 2694
rect 2287 2677 2713 2694
rect 2837 2677 3263 2694
rect 3387 2677 3813 2694
rect 3937 2677 4363 2694
rect 4487 2677 4913 2694
rect 5037 2677 5463 2694
rect 5587 2677 6013 2694
rect 6137 2677 6563 2694
rect 6687 2677 7113 2694
rect 7237 2677 7663 2694
rect 7787 2677 8213 2694
rect 8337 2677 8763 2694
rect 8887 2677 9313 2694
rect 9437 2677 9863 2694
rect 9987 2677 10413 2694
rect 10537 2677 10963 2694
rect 11087 2677 11513 2694
rect 11637 2677 12063 2694
rect 12187 2677 12613 2694
rect 12737 2677 13163 2694
rect 13287 2677 13713 2694
rect -23 2237 -6 2663
rect 56 2237 73 2663
rect 135 2603 465 2615
rect 135 2297 147 2603
rect 147 2297 453 2603
rect 453 2297 465 2603
rect 135 2285 465 2297
rect 527 2237 544 2663
rect 606 2237 623 2663
rect 1077 2237 1094 2663
rect 1156 2237 1173 2663
rect 1235 2603 1565 2615
rect 1235 2297 1247 2603
rect 1247 2297 1553 2603
rect 1553 2297 1565 2603
rect 1235 2285 1565 2297
rect 1627 2237 1644 2663
rect 1706 2237 1723 2663
rect 2177 2237 2194 2663
rect 2256 2237 2273 2663
rect 2335 2603 2665 2615
rect 2335 2297 2347 2603
rect 2347 2297 2653 2603
rect 2653 2297 2665 2603
rect 2335 2285 2665 2297
rect 2727 2237 2744 2663
rect 2806 2237 2823 2663
rect 3277 2237 3294 2663
rect 3356 2237 3373 2663
rect 3435 2603 3765 2615
rect 3435 2297 3447 2603
rect 3447 2297 3753 2603
rect 3753 2297 3765 2603
rect 3435 2285 3765 2297
rect 3827 2237 3844 2663
rect 3906 2237 3923 2663
rect 4377 2237 4394 2663
rect 4456 2237 4473 2663
rect 4535 2603 4865 2615
rect 4535 2297 4547 2603
rect 4547 2297 4853 2603
rect 4853 2297 4865 2603
rect 4535 2285 4865 2297
rect 4927 2237 4944 2663
rect 5006 2237 5023 2663
rect 5477 2237 5494 2663
rect 5556 2237 5573 2663
rect 5635 2603 5965 2615
rect 5635 2297 5647 2603
rect 5647 2297 5953 2603
rect 5953 2297 5965 2603
rect 5635 2285 5965 2297
rect 6027 2237 6044 2663
rect 6106 2237 6123 2663
rect 6577 2237 6594 2663
rect 6656 2237 6673 2663
rect 6735 2603 7065 2615
rect 6735 2297 6747 2603
rect 6747 2297 7053 2603
rect 7053 2297 7065 2603
rect 6735 2285 7065 2297
rect 7127 2237 7144 2663
rect 7206 2237 7223 2663
rect 7677 2237 7694 2663
rect 7756 2237 7773 2663
rect 7835 2603 8165 2615
rect 7835 2297 7847 2603
rect 7847 2297 8153 2603
rect 8153 2297 8165 2603
rect 7835 2285 8165 2297
rect 8227 2237 8244 2663
rect 8306 2237 8323 2663
rect 8777 2237 8794 2663
rect 8856 2237 8873 2663
rect 8935 2603 9265 2615
rect 8935 2297 8947 2603
rect 8947 2297 9253 2603
rect 9253 2297 9265 2603
rect 8935 2285 9265 2297
rect 9327 2237 9344 2663
rect 9406 2237 9423 2663
rect 9877 2237 9894 2663
rect 9956 2237 9973 2663
rect 10035 2603 10365 2615
rect 10035 2297 10047 2603
rect 10047 2297 10353 2603
rect 10353 2297 10365 2603
rect 10035 2285 10365 2297
rect 10427 2237 10444 2663
rect 10506 2237 10523 2663
rect 10977 2237 10994 2663
rect 11056 2237 11073 2663
rect 11135 2603 11465 2615
rect 11135 2297 11147 2603
rect 11147 2297 11453 2603
rect 11453 2297 11465 2603
rect 11135 2285 11465 2297
rect 11527 2237 11544 2663
rect 11606 2237 11623 2663
rect 12077 2237 12094 2663
rect 12156 2237 12173 2663
rect 12235 2603 12565 2615
rect 12235 2297 12247 2603
rect 12247 2297 12553 2603
rect 12553 2297 12565 2603
rect 12235 2285 12565 2297
rect 12627 2237 12644 2663
rect 12706 2237 12723 2663
rect 13177 2237 13194 2663
rect 13256 2237 13273 2663
rect 13335 2603 13665 2615
rect 13335 2297 13347 2603
rect 13347 2297 13653 2603
rect 13653 2297 13665 2603
rect 13335 2285 13665 2297
rect -463 2206 -37 2223
rect 87 2206 513 2223
rect 637 2206 1063 2223
rect 1187 2206 1613 2223
rect 1737 2206 2163 2223
rect 2287 2206 2713 2223
rect 2837 2206 3263 2223
rect 3387 2206 3813 2223
rect 3937 2206 4363 2223
rect 4487 2206 4913 2223
rect 5037 2206 5463 2223
rect 5587 2206 6013 2223
rect 6137 2206 6563 2223
rect 6687 2206 7113 2223
rect 7237 2206 7663 2223
rect 7787 2206 8213 2223
rect 8337 2206 8763 2223
rect 8887 2206 9313 2223
rect 9437 2206 9863 2223
rect 9987 2206 10413 2223
rect 10537 2206 10963 2223
rect 11087 2206 11513 2223
rect 11637 2206 12063 2223
rect 12187 2206 12613 2223
rect 12737 2206 13163 2223
rect 13287 2206 13713 2223
rect 13987 2219 14263 2750
rect -1013 1669 -737 2200
rect -542 2158 -508 2192
rect 8 2158 42 2192
rect 558 2158 592 2192
rect 1108 2158 1142 2192
rect 1658 2158 1692 2192
rect 2208 2158 2242 2192
rect 2758 2158 2792 2192
rect 3308 2158 3342 2192
rect 3858 2158 3892 2192
rect 4408 2158 4442 2192
rect 4958 2158 4992 2192
rect 5508 2158 5542 2192
rect 6058 2158 6092 2192
rect 6608 2158 6642 2192
rect 7158 2158 7192 2192
rect 7708 2158 7742 2192
rect 8258 2158 8292 2192
rect 8808 2158 8842 2192
rect 9358 2158 9392 2192
rect 9908 2158 9942 2192
rect 10458 2158 10492 2192
rect 11008 2158 11042 2192
rect 11558 2158 11592 2192
rect 12108 2158 12142 2192
rect 12658 2158 12692 2192
rect 13208 2158 13242 2192
rect 13758 2158 13792 2192
rect -463 2127 -37 2144
rect 87 2127 513 2144
rect 637 2127 1063 2144
rect 1187 2127 1613 2144
rect 1737 2127 2163 2144
rect 2287 2127 2713 2144
rect 2837 2127 3263 2144
rect 3387 2127 3813 2144
rect 3937 2127 4363 2144
rect 4487 2127 4913 2144
rect 5037 2127 5463 2144
rect 5587 2127 6013 2144
rect 6137 2127 6563 2144
rect 6687 2127 7113 2144
rect 7237 2127 7663 2144
rect 7787 2127 8213 2144
rect 8337 2127 8763 2144
rect 8887 2127 9313 2144
rect 9437 2127 9863 2144
rect 9987 2127 10413 2144
rect 10537 2127 10963 2144
rect 11087 2127 11513 2144
rect 11637 2127 12063 2144
rect 12187 2127 12613 2144
rect 12737 2127 13163 2144
rect 13287 2127 13713 2144
rect -415 2053 -85 2065
rect -415 1747 -403 2053
rect -403 1747 -97 2053
rect -97 1747 -85 2053
rect -415 1735 -85 1747
rect -23 1687 -6 2113
rect 56 1687 73 2113
rect 527 1687 544 2113
rect 606 1687 623 2113
rect 685 2053 1015 2065
rect 685 1747 697 2053
rect 697 1747 1003 2053
rect 1003 1747 1015 2053
rect 685 1735 1015 1747
rect 1077 1687 1094 2113
rect 1156 1687 1173 2113
rect 1627 1687 1644 2113
rect 1706 1687 1723 2113
rect 1785 2053 2115 2065
rect 1785 1747 1797 2053
rect 1797 1747 2103 2053
rect 2103 1747 2115 2053
rect 1785 1735 2115 1747
rect 2177 1687 2194 2113
rect 2256 1687 2273 2113
rect 2727 1687 2744 2113
rect 2806 1687 2823 2113
rect 2885 2053 3215 2065
rect 2885 1747 2897 2053
rect 2897 1747 3203 2053
rect 3203 1747 3215 2053
rect 2885 1735 3215 1747
rect 3277 1687 3294 2113
rect 3356 1687 3373 2113
rect 3827 1687 3844 2113
rect 3906 1687 3923 2113
rect 3985 2053 4315 2065
rect 3985 1747 3997 2053
rect 3997 1747 4303 2053
rect 4303 1747 4315 2053
rect 3985 1735 4315 1747
rect 4377 1687 4394 2113
rect 4456 1687 4473 2113
rect 4927 1687 4944 2113
rect 5006 1687 5023 2113
rect 5085 2053 5415 2065
rect 5085 1747 5097 2053
rect 5097 1747 5403 2053
rect 5403 1747 5415 2053
rect 5085 1735 5415 1747
rect 5477 1687 5494 2113
rect 5556 1687 5573 2113
rect 6027 1687 6044 2113
rect 6106 1687 6123 2113
rect 6185 2053 6515 2065
rect 6185 1747 6197 2053
rect 6197 1747 6503 2053
rect 6503 1747 6515 2053
rect 6185 1735 6515 1747
rect 6577 1687 6594 2113
rect 6656 1687 6673 2113
rect 7127 1687 7144 2113
rect 7206 1687 7223 2113
rect 7285 2053 7615 2065
rect 7285 1747 7297 2053
rect 7297 1747 7603 2053
rect 7603 1747 7615 2053
rect 7285 1735 7615 1747
rect 7677 1687 7694 2113
rect 7756 1687 7773 2113
rect 8227 1687 8244 2113
rect 8306 1687 8323 2113
rect 8385 2053 8715 2065
rect 8385 1747 8397 2053
rect 8397 1747 8703 2053
rect 8703 1747 8715 2053
rect 8385 1735 8715 1747
rect 8777 1687 8794 2113
rect 8856 1687 8873 2113
rect 9327 1687 9344 2113
rect 9406 1687 9423 2113
rect 9485 2053 9815 2065
rect 9485 1747 9497 2053
rect 9497 1747 9803 2053
rect 9803 1747 9815 2053
rect 9485 1735 9815 1747
rect 9877 1687 9894 2113
rect 9956 1687 9973 2113
rect 10427 1687 10444 2113
rect 10506 1687 10523 2113
rect 10585 2053 10915 2065
rect 10585 1747 10597 2053
rect 10597 1747 10903 2053
rect 10903 1747 10915 2053
rect 10585 1735 10915 1747
rect 10977 1687 10994 2113
rect 11056 1687 11073 2113
rect 11527 1687 11544 2113
rect 11606 1687 11623 2113
rect 11685 2053 12015 2065
rect 11685 1747 11697 2053
rect 11697 1747 12003 2053
rect 12003 1747 12015 2053
rect 11685 1735 12015 1747
rect 12077 1687 12094 2113
rect 12156 1687 12173 2113
rect 12627 1687 12644 2113
rect 12706 1687 12723 2113
rect 12785 2053 13115 2065
rect 12785 1747 12797 2053
rect 12797 1747 13103 2053
rect 13103 1747 13115 2053
rect 12785 1735 13115 1747
rect 13177 1687 13194 2113
rect 13256 1687 13273 2113
rect -463 1656 -37 1673
rect 87 1656 513 1673
rect 637 1656 1063 1673
rect 1187 1656 1613 1673
rect 1737 1656 2163 1673
rect 2287 1656 2713 1673
rect 2837 1656 3263 1673
rect 3387 1656 3813 1673
rect 3937 1656 4363 1673
rect 4487 1656 4913 1673
rect 5037 1656 5463 1673
rect 5587 1656 6013 1673
rect 6137 1656 6563 1673
rect 6687 1656 7113 1673
rect 7237 1656 7663 1673
rect 7787 1656 8213 1673
rect 8337 1656 8763 1673
rect 8887 1656 9313 1673
rect 9437 1656 9863 1673
rect 9987 1656 10413 1673
rect 10537 1656 10963 1673
rect 11087 1656 11513 1673
rect 11637 1656 12063 1673
rect 12187 1656 12613 1673
rect 12737 1656 13163 1673
rect 13287 1656 13713 1673
rect 13987 1669 14263 2200
rect -1013 1119 -737 1650
rect -542 1608 -508 1642
rect 8 1608 42 1642
rect 558 1608 592 1642
rect 1108 1608 1142 1642
rect 1658 1608 1692 1642
rect 2208 1608 2242 1642
rect 2758 1608 2792 1642
rect 3308 1608 3342 1642
rect 3858 1608 3892 1642
rect 4408 1608 4442 1642
rect 4958 1608 4992 1642
rect 5508 1608 5542 1642
rect 6058 1608 6092 1642
rect 6608 1608 6642 1642
rect 7158 1608 7192 1642
rect 7708 1608 7742 1642
rect 8258 1608 8292 1642
rect 8808 1608 8842 1642
rect 9358 1608 9392 1642
rect 9908 1608 9942 1642
rect 10458 1608 10492 1642
rect 11008 1608 11042 1642
rect 11558 1608 11592 1642
rect 12108 1608 12142 1642
rect 12658 1608 12692 1642
rect 13208 1608 13242 1642
rect 13758 1608 13792 1642
rect -463 1577 -37 1594
rect 87 1577 513 1594
rect 637 1577 1063 1594
rect 1187 1577 1613 1594
rect 1737 1577 2163 1594
rect 2287 1577 2713 1594
rect 2837 1577 3263 1594
rect 3387 1577 3813 1594
rect 3937 1577 4363 1594
rect 4487 1577 4913 1594
rect 5037 1577 5463 1594
rect 5587 1577 6013 1594
rect 6137 1577 6563 1594
rect 6687 1577 7113 1594
rect 7237 1577 7663 1594
rect 7787 1577 8213 1594
rect 8337 1577 8763 1594
rect 8887 1577 9313 1594
rect 9437 1577 9863 1594
rect 9987 1577 10413 1594
rect 10537 1577 10963 1594
rect 11087 1577 11513 1594
rect 11637 1577 12063 1594
rect 12187 1577 12613 1594
rect 12737 1577 13163 1594
rect 13287 1577 13713 1594
rect -23 1137 -6 1563
rect 56 1137 73 1563
rect 135 1503 465 1515
rect 135 1197 147 1503
rect 147 1197 453 1503
rect 453 1197 465 1503
rect 135 1185 465 1197
rect 527 1137 544 1563
rect 606 1137 623 1563
rect 1077 1137 1094 1563
rect 1156 1137 1173 1563
rect 1235 1503 1565 1515
rect 1235 1197 1247 1503
rect 1247 1197 1553 1503
rect 1553 1197 1565 1503
rect 1235 1185 1565 1197
rect 1627 1137 1644 1563
rect 1706 1137 1723 1563
rect 2177 1137 2194 1563
rect 2256 1137 2273 1563
rect 2335 1503 2665 1515
rect 2335 1197 2347 1503
rect 2347 1197 2653 1503
rect 2653 1197 2665 1503
rect 2335 1185 2665 1197
rect 2727 1137 2744 1563
rect 2806 1137 2823 1563
rect 3277 1137 3294 1563
rect 3356 1137 3373 1563
rect 3435 1503 3765 1515
rect 3435 1197 3447 1503
rect 3447 1197 3753 1503
rect 3753 1197 3765 1503
rect 3435 1185 3765 1197
rect 3827 1137 3844 1563
rect 3906 1137 3923 1563
rect 4377 1137 4394 1563
rect 4456 1137 4473 1563
rect 4535 1503 4865 1515
rect 4535 1197 4547 1503
rect 4547 1197 4853 1503
rect 4853 1197 4865 1503
rect 4535 1185 4865 1197
rect 4927 1137 4944 1563
rect 5006 1137 5023 1563
rect 5477 1137 5494 1563
rect 5556 1137 5573 1563
rect 5635 1503 5965 1515
rect 5635 1197 5647 1503
rect 5647 1197 5953 1503
rect 5953 1197 5965 1503
rect 5635 1185 5965 1197
rect 6027 1137 6044 1563
rect 6106 1137 6123 1563
rect 6577 1137 6594 1563
rect 6656 1137 6673 1563
rect 6735 1503 7065 1515
rect 6735 1197 6747 1503
rect 6747 1197 7053 1503
rect 7053 1197 7065 1503
rect 6735 1185 7065 1197
rect 7127 1137 7144 1563
rect 7206 1137 7223 1563
rect 7677 1137 7694 1563
rect 7756 1137 7773 1563
rect 7835 1503 8165 1515
rect 7835 1197 7847 1503
rect 7847 1197 8153 1503
rect 8153 1197 8165 1503
rect 7835 1185 8165 1197
rect 8227 1137 8244 1563
rect 8306 1137 8323 1563
rect 8777 1137 8794 1563
rect 8856 1137 8873 1563
rect 8935 1503 9265 1515
rect 8935 1197 8947 1503
rect 8947 1197 9253 1503
rect 9253 1197 9265 1503
rect 8935 1185 9265 1197
rect 9327 1137 9344 1563
rect 9406 1137 9423 1563
rect 9877 1137 9894 1563
rect 9956 1137 9973 1563
rect 10035 1503 10365 1515
rect 10035 1197 10047 1503
rect 10047 1197 10353 1503
rect 10353 1197 10365 1503
rect 10035 1185 10365 1197
rect 10427 1137 10444 1563
rect 10506 1137 10523 1563
rect 10977 1137 10994 1563
rect 11056 1137 11073 1563
rect 11135 1503 11465 1515
rect 11135 1197 11147 1503
rect 11147 1197 11453 1503
rect 11453 1197 11465 1503
rect 11135 1185 11465 1197
rect 11527 1137 11544 1563
rect 11606 1137 11623 1563
rect 12077 1137 12094 1563
rect 12156 1137 12173 1563
rect 12235 1503 12565 1515
rect 12235 1197 12247 1503
rect 12247 1197 12553 1503
rect 12553 1197 12565 1503
rect 12235 1185 12565 1197
rect 12627 1137 12644 1563
rect 12706 1137 12723 1563
rect 13177 1137 13194 1563
rect 13256 1137 13273 1563
rect 13335 1503 13665 1515
rect 13335 1197 13347 1503
rect 13347 1197 13653 1503
rect 13653 1197 13665 1503
rect 13335 1185 13665 1197
rect -463 1106 -37 1123
rect 87 1106 513 1123
rect 637 1106 1063 1123
rect 1187 1106 1613 1123
rect 1737 1106 2163 1123
rect 2287 1106 2713 1123
rect 2837 1106 3263 1123
rect 3387 1106 3813 1123
rect 3937 1106 4363 1123
rect 4487 1106 4913 1123
rect 5037 1106 5463 1123
rect 5587 1106 6013 1123
rect 6137 1106 6563 1123
rect 6687 1106 7113 1123
rect 7237 1106 7663 1123
rect 7787 1106 8213 1123
rect 8337 1106 8763 1123
rect 8887 1106 9313 1123
rect 9437 1106 9863 1123
rect 9987 1106 10413 1123
rect 10537 1106 10963 1123
rect 11087 1106 11513 1123
rect 11637 1106 12063 1123
rect 12187 1106 12613 1123
rect 12737 1106 13163 1123
rect 13287 1106 13713 1123
rect 13987 1119 14263 1650
rect -1013 569 -737 1100
rect -542 1058 -508 1092
rect 8 1058 42 1092
rect 558 1058 592 1092
rect 1108 1058 1142 1092
rect 1658 1058 1692 1092
rect 2208 1058 2242 1092
rect 2758 1058 2792 1092
rect 3308 1058 3342 1092
rect 3858 1058 3892 1092
rect 4408 1058 4442 1092
rect 4958 1058 4992 1092
rect 5508 1058 5542 1092
rect 6058 1058 6092 1092
rect 6608 1058 6642 1092
rect 7158 1058 7192 1092
rect 7708 1058 7742 1092
rect 8258 1058 8292 1092
rect 8808 1058 8842 1092
rect 9358 1058 9392 1092
rect 9908 1058 9942 1092
rect 10458 1058 10492 1092
rect 11008 1058 11042 1092
rect 11558 1058 11592 1092
rect 12108 1058 12142 1092
rect 12658 1058 12692 1092
rect 13208 1058 13242 1092
rect 13758 1058 13792 1092
rect -463 1027 -37 1044
rect 87 1027 513 1044
rect 637 1027 1063 1044
rect 1187 1027 1613 1044
rect 1737 1027 2163 1044
rect 2287 1027 2713 1044
rect 2837 1027 3263 1044
rect 3387 1027 3813 1044
rect 3937 1027 4363 1044
rect 4487 1027 4913 1044
rect 5037 1027 5463 1044
rect 5587 1027 6013 1044
rect 6137 1027 6563 1044
rect 6687 1027 7113 1044
rect 7237 1027 7663 1044
rect 7787 1027 8213 1044
rect 8337 1027 8763 1044
rect 8887 1027 9313 1044
rect 9437 1027 9863 1044
rect 9987 1027 10413 1044
rect 10537 1027 10963 1044
rect 11087 1027 11513 1044
rect 11637 1027 12063 1044
rect 12187 1027 12613 1044
rect 12737 1027 13163 1044
rect 13287 1027 13713 1044
rect -415 953 -85 965
rect -415 647 -403 953
rect -403 647 -97 953
rect -97 647 -85 953
rect -415 635 -85 647
rect -23 587 -6 1013
rect 56 587 73 1013
rect 527 587 544 1013
rect 606 587 623 1013
rect 685 953 1015 965
rect 685 647 697 953
rect 697 647 1003 953
rect 1003 647 1015 953
rect 685 635 1015 647
rect 1077 587 1094 1013
rect 1156 587 1173 1013
rect 1627 587 1644 1013
rect 1706 587 1723 1013
rect 1785 953 2115 965
rect 1785 647 1797 953
rect 1797 647 2103 953
rect 2103 647 2115 953
rect 1785 635 2115 647
rect 2177 587 2194 1013
rect 2256 587 2273 1013
rect 2727 587 2744 1013
rect 2806 587 2823 1013
rect 2885 953 3215 965
rect 2885 647 2897 953
rect 2897 647 3203 953
rect 3203 647 3215 953
rect 2885 635 3215 647
rect 3277 587 3294 1013
rect 3356 587 3373 1013
rect 3827 587 3844 1013
rect 3906 587 3923 1013
rect 3985 953 4315 965
rect 3985 647 3997 953
rect 3997 647 4303 953
rect 4303 647 4315 953
rect 3985 635 4315 647
rect 4377 587 4394 1013
rect 4456 587 4473 1013
rect 4927 587 4944 1013
rect 5006 587 5023 1013
rect 5085 953 5415 965
rect 5085 647 5097 953
rect 5097 647 5403 953
rect 5403 647 5415 953
rect 5085 635 5415 647
rect 5477 587 5494 1013
rect 5556 587 5573 1013
rect 6027 587 6044 1013
rect 6106 587 6123 1013
rect 6185 953 6515 965
rect 6185 647 6197 953
rect 6197 647 6503 953
rect 6503 647 6515 953
rect 6185 635 6515 647
rect 6577 587 6594 1013
rect 6656 587 6673 1013
rect 7127 587 7144 1013
rect 7206 587 7223 1013
rect 7285 953 7615 965
rect 7285 647 7297 953
rect 7297 647 7603 953
rect 7603 647 7615 953
rect 7285 635 7615 647
rect 7677 587 7694 1013
rect 7756 587 7773 1013
rect 8227 587 8244 1013
rect 8306 587 8323 1013
rect 8385 953 8715 965
rect 8385 647 8397 953
rect 8397 647 8703 953
rect 8703 647 8715 953
rect 8385 635 8715 647
rect 8777 587 8794 1013
rect 8856 587 8873 1013
rect 9327 587 9344 1013
rect 9406 587 9423 1013
rect 9485 953 9815 965
rect 9485 647 9497 953
rect 9497 647 9803 953
rect 9803 647 9815 953
rect 9485 635 9815 647
rect 9877 587 9894 1013
rect 9956 587 9973 1013
rect 10427 587 10444 1013
rect 10506 587 10523 1013
rect 10585 953 10915 965
rect 10585 647 10597 953
rect 10597 647 10903 953
rect 10903 647 10915 953
rect 10585 635 10915 647
rect 10977 587 10994 1013
rect 11056 587 11073 1013
rect 11527 587 11544 1013
rect 11606 587 11623 1013
rect 11685 953 12015 965
rect 11685 647 11697 953
rect 11697 647 12003 953
rect 12003 647 12015 953
rect 11685 635 12015 647
rect 12077 587 12094 1013
rect 12156 587 12173 1013
rect 12627 587 12644 1013
rect 12706 587 12723 1013
rect 12785 953 13115 965
rect 12785 647 12797 953
rect 12797 647 13103 953
rect 13103 647 13115 953
rect 12785 635 13115 647
rect 13177 587 13194 1013
rect 13256 587 13273 1013
rect -463 556 -37 573
rect 87 556 513 573
rect 637 556 1063 573
rect 1187 556 1613 573
rect 1737 556 2163 573
rect 2287 556 2713 573
rect 2837 556 3263 573
rect 3387 556 3813 573
rect 3937 556 4363 573
rect 4487 556 4913 573
rect 5037 556 5463 573
rect 5587 556 6013 573
rect 6137 556 6563 573
rect 6687 556 7113 573
rect 7237 556 7663 573
rect 7787 556 8213 573
rect 8337 556 8763 573
rect 8887 556 9313 573
rect 9437 556 9863 573
rect 9987 556 10413 573
rect 10537 556 10963 573
rect 11087 556 11513 573
rect 11637 556 12063 573
rect 12187 556 12613 573
rect 12737 556 13163 573
rect 13287 556 13713 573
rect 13987 569 14263 1100
rect -1013 19 -737 550
rect -542 508 -508 542
rect 8 508 42 542
rect 558 508 592 542
rect 1108 508 1142 542
rect 1658 508 1692 542
rect 2208 508 2242 542
rect 2758 508 2792 542
rect 3308 508 3342 542
rect 3858 508 3892 542
rect 4408 508 4442 542
rect 4958 508 4992 542
rect 5508 508 5542 542
rect 6058 508 6092 542
rect 6608 508 6642 542
rect 7158 508 7192 542
rect 7708 508 7742 542
rect 8258 508 8292 542
rect 8808 508 8842 542
rect 9358 508 9392 542
rect 9908 508 9942 542
rect 10458 508 10492 542
rect 11008 508 11042 542
rect 11558 508 11592 542
rect 12108 508 12142 542
rect 12658 508 12692 542
rect 13208 508 13242 542
rect 13758 508 13792 542
rect -463 477 -37 494
rect 87 477 513 494
rect 637 477 1063 494
rect 1187 477 1613 494
rect 1737 477 2163 494
rect 2287 477 2713 494
rect 2837 477 3263 494
rect 3387 477 3813 494
rect 3937 477 4363 494
rect 4487 477 4913 494
rect 5037 477 5463 494
rect 5587 477 6013 494
rect 6137 477 6563 494
rect 6687 477 7113 494
rect 7237 477 7663 494
rect 7787 477 8213 494
rect 8337 477 8763 494
rect 8887 477 9313 494
rect 9437 477 9863 494
rect 9987 477 10413 494
rect 10537 477 10963 494
rect 11087 477 11513 494
rect 11637 477 12063 494
rect 12187 477 12613 494
rect 12737 477 13163 494
rect 13287 477 13713 494
rect -23 37 -6 463
rect 56 37 73 463
rect 135 403 465 415
rect 135 97 147 403
rect 147 97 453 403
rect 453 97 465 403
rect 135 85 465 97
rect 527 37 544 463
rect 606 37 623 463
rect 1077 37 1094 463
rect 1156 37 1173 463
rect 1235 403 1565 415
rect 1235 97 1247 403
rect 1247 97 1553 403
rect 1553 97 1565 403
rect 1235 85 1565 97
rect 1627 37 1644 463
rect 1706 37 1723 463
rect 2177 37 2194 463
rect 2256 37 2273 463
rect 2335 403 2665 415
rect 2335 97 2347 403
rect 2347 97 2653 403
rect 2653 97 2665 403
rect 2335 85 2665 97
rect 2727 37 2744 463
rect 2806 37 2823 463
rect 3277 37 3294 463
rect 3356 37 3373 463
rect 3435 403 3765 415
rect 3435 97 3447 403
rect 3447 97 3753 403
rect 3753 97 3765 403
rect 3435 85 3765 97
rect 3827 37 3844 463
rect 3906 37 3923 463
rect 4377 37 4394 463
rect 4456 37 4473 463
rect 4535 403 4865 415
rect 4535 97 4547 403
rect 4547 97 4853 403
rect 4853 97 4865 403
rect 4535 85 4865 97
rect 4927 37 4944 463
rect 5006 37 5023 463
rect 5477 37 5494 463
rect 5556 37 5573 463
rect 5635 403 5965 415
rect 5635 97 5647 403
rect 5647 97 5953 403
rect 5953 97 5965 403
rect 5635 85 5965 97
rect 6027 37 6044 463
rect 6106 37 6123 463
rect 6577 37 6594 463
rect 6656 37 6673 463
rect 6735 403 7065 415
rect 6735 97 6747 403
rect 6747 97 7053 403
rect 7053 97 7065 403
rect 6735 85 7065 97
rect 7127 37 7144 463
rect 7206 37 7223 463
rect 7677 37 7694 463
rect 7756 37 7773 463
rect 7835 403 8165 415
rect 7835 97 7847 403
rect 7847 97 8153 403
rect 8153 97 8165 403
rect 7835 85 8165 97
rect 8227 37 8244 463
rect 8306 37 8323 463
rect 8777 37 8794 463
rect 8856 37 8873 463
rect 8935 403 9265 415
rect 8935 97 8947 403
rect 8947 97 9253 403
rect 9253 97 9265 403
rect 8935 85 9265 97
rect 9327 37 9344 463
rect 9406 37 9423 463
rect 9877 37 9894 463
rect 9956 37 9973 463
rect 10035 403 10365 415
rect 10035 97 10047 403
rect 10047 97 10353 403
rect 10353 97 10365 403
rect 10035 85 10365 97
rect 10427 37 10444 463
rect 10506 37 10523 463
rect 10977 37 10994 463
rect 11056 37 11073 463
rect 11135 403 11465 415
rect 11135 97 11147 403
rect 11147 97 11453 403
rect 11453 97 11465 403
rect 11135 85 11465 97
rect 11527 37 11544 463
rect 11606 37 11623 463
rect 12077 37 12094 463
rect 12156 37 12173 463
rect 12235 403 12565 415
rect 12235 97 12247 403
rect 12247 97 12553 403
rect 12553 97 12565 403
rect 12235 85 12565 97
rect 12627 37 12644 463
rect 12706 37 12723 463
rect 13177 37 13194 463
rect 13256 37 13273 463
rect 13335 403 13665 415
rect 13335 97 13347 403
rect 13347 97 13653 403
rect 13653 97 13665 403
rect 13335 85 13665 97
rect -463 6 -37 23
rect 87 6 513 23
rect 637 6 1063 23
rect 1187 6 1613 23
rect 1737 6 2163 23
rect 2287 6 2713 23
rect 2837 6 3263 23
rect 3387 6 3813 23
rect 3937 6 4363 23
rect 4487 6 4913 23
rect 5037 6 5463 23
rect 5587 6 6013 23
rect 6137 6 6563 23
rect 6687 6 7113 23
rect 7237 6 7663 23
rect 7787 6 8213 23
rect 8337 6 8763 23
rect 8887 6 9313 23
rect 9437 6 9863 23
rect 9987 6 10413 23
rect 10537 6 10963 23
rect 11087 6 11513 23
rect 11637 6 12063 23
rect 12187 6 12613 23
rect 12737 6 13163 23
rect 13287 6 13713 23
rect 13987 19 14263 550
rect -1013 -787 -737 0
rect -542 -42 -508 -8
rect 8 -42 42 -8
rect 558 -42 592 -8
rect 1108 -42 1142 -8
rect 1658 -42 1692 -8
rect 2208 -42 2242 -8
rect 2758 -42 2792 -8
rect 3308 -42 3342 -8
rect 3858 -42 3892 -8
rect 4408 -42 4442 -8
rect 4958 -42 4992 -8
rect 5508 -42 5542 -8
rect 6058 -42 6092 -8
rect 6608 -42 6642 -8
rect 7158 -42 7192 -8
rect 7708 -42 7742 -8
rect 8258 -42 8292 -8
rect 8808 -42 8842 -8
rect 9358 -42 9392 -8
rect 9908 -42 9942 -8
rect 10458 -42 10492 -8
rect 11008 -42 11042 -8
rect 11558 -42 11592 -8
rect 12108 -42 12142 -8
rect 12658 -42 12692 -8
rect 13208 -42 13242 -8
rect 13758 -42 13792 -8
rect -463 -73 -37 -56
rect 87 -73 513 -56
rect 637 -73 1063 -56
rect 1187 -73 1613 -56
rect 1737 -73 2163 -56
rect 2287 -73 2713 -56
rect 2837 -73 3263 -56
rect 3387 -73 3813 -56
rect 3937 -73 4363 -56
rect 4487 -73 4913 -56
rect 5037 -73 5463 -56
rect 5587 -73 6013 -56
rect 6137 -73 6563 -56
rect 6687 -73 7113 -56
rect 7237 -73 7663 -56
rect 7787 -73 8213 -56
rect 8337 -73 8763 -56
rect 8887 -73 9313 -56
rect 9437 -73 9863 -56
rect 9987 -73 10413 -56
rect 10537 -73 10963 -56
rect 11087 -73 11513 -56
rect 11637 -73 12063 -56
rect 12187 -73 12613 -56
rect 12737 -73 13163 -56
rect 13287 -73 13713 -56
rect -415 -147 -85 -135
rect -415 -453 -403 -147
rect -403 -453 -97 -147
rect -97 -453 -85 -147
rect -415 -465 -85 -453
rect -23 -513 -6 -87
rect 56 -513 73 -87
rect 527 -513 544 -87
rect 606 -513 623 -87
rect 685 -147 1015 -135
rect 685 -453 697 -147
rect 697 -453 1003 -147
rect 1003 -453 1015 -147
rect 685 -465 1015 -453
rect 1077 -513 1094 -87
rect 1156 -513 1173 -87
rect 1627 -513 1644 -87
rect 1706 -513 1723 -87
rect 1785 -147 2115 -135
rect 1785 -453 1797 -147
rect 1797 -453 2103 -147
rect 2103 -453 2115 -147
rect 1785 -465 2115 -453
rect 2177 -513 2194 -87
rect 2256 -513 2273 -87
rect 2727 -513 2744 -87
rect 2806 -513 2823 -87
rect 2885 -147 3215 -135
rect 2885 -453 2897 -147
rect 2897 -453 3203 -147
rect 3203 -453 3215 -147
rect 2885 -465 3215 -453
rect 3277 -513 3294 -87
rect 3356 -513 3373 -87
rect 3827 -513 3844 -87
rect 3906 -513 3923 -87
rect 3985 -147 4315 -135
rect 3985 -453 3997 -147
rect 3997 -453 4303 -147
rect 4303 -453 4315 -147
rect 3985 -465 4315 -453
rect 4377 -513 4394 -87
rect 4456 -513 4473 -87
rect 4927 -513 4944 -87
rect 5006 -513 5023 -87
rect 5085 -147 5415 -135
rect 5085 -453 5097 -147
rect 5097 -453 5403 -147
rect 5403 -453 5415 -147
rect 5085 -465 5415 -453
rect 5477 -513 5494 -87
rect 5556 -513 5573 -87
rect 6027 -513 6044 -87
rect 6106 -513 6123 -87
rect 6185 -147 6515 -135
rect 6185 -453 6197 -147
rect 6197 -453 6503 -147
rect 6503 -453 6515 -147
rect 6185 -465 6515 -453
rect 6577 -513 6594 -87
rect 6656 -513 6673 -87
rect 7127 -513 7144 -87
rect 7206 -513 7223 -87
rect 7285 -147 7615 -135
rect 7285 -453 7297 -147
rect 7297 -453 7603 -147
rect 7603 -453 7615 -147
rect 7285 -465 7615 -453
rect 7677 -513 7694 -87
rect 7756 -513 7773 -87
rect 8227 -513 8244 -87
rect 8306 -513 8323 -87
rect 8385 -147 8715 -135
rect 8385 -453 8397 -147
rect 8397 -453 8703 -147
rect 8703 -453 8715 -147
rect 8385 -465 8715 -453
rect 8777 -513 8794 -87
rect 8856 -513 8873 -87
rect 9327 -513 9344 -87
rect 9406 -513 9423 -87
rect 9485 -147 9815 -135
rect 9485 -453 9497 -147
rect 9497 -453 9803 -147
rect 9803 -453 9815 -147
rect 9485 -465 9815 -453
rect 9877 -513 9894 -87
rect 9956 -513 9973 -87
rect 10427 -513 10444 -87
rect 10506 -513 10523 -87
rect 10585 -147 10915 -135
rect 10585 -453 10597 -147
rect 10597 -453 10903 -147
rect 10903 -453 10915 -147
rect 10585 -465 10915 -453
rect 10977 -513 10994 -87
rect 11056 -513 11073 -87
rect 11527 -513 11544 -87
rect 11606 -513 11623 -87
rect 11685 -147 12015 -135
rect 11685 -453 11697 -147
rect 11697 -453 12003 -147
rect 12003 -453 12015 -147
rect 11685 -465 12015 -453
rect 12077 -513 12094 -87
rect 12156 -513 12173 -87
rect 12627 -513 12644 -87
rect 12706 -513 12723 -87
rect 12785 -147 13115 -135
rect 12785 -453 12797 -147
rect 12797 -453 13103 -147
rect 13103 -453 13115 -147
rect 12785 -465 13115 -453
rect 13177 -513 13194 -87
rect 13256 -513 13273 -87
rect -542 -592 -508 -558
rect 8 -592 42 -558
rect 558 -592 592 -558
rect 1108 -592 1142 -558
rect 1658 -592 1692 -558
rect 2208 -592 2242 -558
rect 2758 -592 2792 -558
rect 3308 -592 3342 -558
rect 3858 -592 3892 -558
rect 4408 -592 4442 -558
rect 4958 -592 4992 -558
rect 5508 -592 5542 -558
rect 6058 -592 6092 -558
rect 6608 -592 6642 -558
rect 7158 -592 7192 -558
rect 7708 -592 7742 -558
rect 8258 -592 8292 -558
rect 8808 -592 8842 -558
rect 9358 -592 9392 -558
rect 9908 -592 9942 -558
rect 10458 -592 10492 -558
rect 11008 -592 11042 -558
rect 11558 -592 11592 -558
rect 12108 -592 12142 -558
rect 12658 -592 12692 -558
rect 13208 -592 13242 -558
rect 13758 -592 13792 -558
rect 13987 -787 14263 0
rect -1013 -1063 -19 -787
rect 0 -1063 531 -787
rect 550 -1063 1081 -787
rect 1100 -1063 1631 -787
rect 1650 -1063 2181 -787
rect 2200 -1063 2731 -787
rect 2750 -1063 3281 -787
rect 3300 -1063 3831 -787
rect 3850 -1063 4381 -787
rect 4400 -1063 4931 -787
rect 4950 -1063 5481 -787
rect 5500 -1063 6031 -787
rect 6050 -1063 6581 -787
rect 6600 -1063 7131 -787
rect 7150 -1063 7681 -787
rect 7700 -1063 8231 -787
rect 8250 -1063 8781 -787
rect 8800 -1063 9331 -787
rect 9350 -1063 9881 -787
rect 9900 -1063 10431 -787
rect 10450 -1063 10981 -787
rect 11000 -1063 11531 -787
rect 11550 -1063 12081 -787
rect 12100 -1063 12631 -787
rect 12650 -1063 13181 -787
rect 13200 -1063 14263 -787
rect 14787 -1587 18763 14737
rect -5513 -5563 18763 -1587
<< metal1 >>
rect -5525 18713 18775 18725
rect -5525 -5563 -5513 18713
rect -1537 14725 14787 14737
rect -1537 -1575 -1525 14725
rect -1025 14213 14275 14225
rect -1025 13219 -1013 14213
rect -19 13937 0 14213
rect 531 13937 550 14213
rect 1081 13937 1100 14213
rect 1631 13937 1650 14213
rect 2181 13937 2200 14213
rect 2731 13937 2750 14213
rect 3281 13937 3300 14213
rect 3831 13937 3850 14213
rect 4381 13937 4400 14213
rect 4931 13937 4950 14213
rect 5481 13937 5500 14213
rect 6031 13937 6050 14213
rect 6581 13937 6600 14213
rect 7131 13937 7150 14213
rect 7681 13937 7700 14213
rect 8231 13937 8250 14213
rect 8781 13937 8800 14213
rect 9331 13937 9350 14213
rect 9881 13937 9900 14213
rect 10431 13937 10450 14213
rect 10981 13937 11000 14213
rect 11531 13937 11550 14213
rect 12081 13937 12100 14213
rect 12631 13937 12650 14213
rect 13181 13937 13200 14213
rect -737 13925 13987 13937
rect -737 13219 -725 13925
rect -550 13742 -500 13750
rect -550 13708 -542 13742
rect -508 13708 -500 13742
rect -550 13700 -500 13708
rect 0 13742 50 13750
rect 0 13708 8 13742
rect 42 13708 50 13742
rect 0 13700 50 13708
rect 550 13742 600 13750
rect 550 13708 558 13742
rect 592 13708 600 13742
rect 550 13700 600 13708
rect 1100 13742 1150 13750
rect 1100 13708 1108 13742
rect 1142 13708 1150 13742
rect 1100 13700 1150 13708
rect 1650 13742 1700 13750
rect 1650 13708 1658 13742
rect 1692 13708 1700 13742
rect 1650 13700 1700 13708
rect 2200 13742 2250 13750
rect 2200 13708 2208 13742
rect 2242 13708 2250 13742
rect 2200 13700 2250 13708
rect 2750 13742 2800 13750
rect 2750 13708 2758 13742
rect 2792 13708 2800 13742
rect 2750 13700 2800 13708
rect 3300 13742 3350 13750
rect 3300 13708 3308 13742
rect 3342 13708 3350 13742
rect 3300 13700 3350 13708
rect 3850 13742 3900 13750
rect 3850 13708 3858 13742
rect 3892 13708 3900 13742
rect 3850 13700 3900 13708
rect 4400 13742 4450 13750
rect 4400 13708 4408 13742
rect 4442 13708 4450 13742
rect 4400 13700 4450 13708
rect 4950 13742 5000 13750
rect 4950 13708 4958 13742
rect 4992 13708 5000 13742
rect 4950 13700 5000 13708
rect 5500 13742 5550 13750
rect 5500 13708 5508 13742
rect 5542 13708 5550 13742
rect 5500 13700 5550 13708
rect 6050 13742 6100 13750
rect 6050 13708 6058 13742
rect 6092 13708 6100 13742
rect 6050 13700 6100 13708
rect 6600 13742 6650 13750
rect 6600 13708 6608 13742
rect 6642 13708 6650 13742
rect 6600 13700 6650 13708
rect 7150 13742 7200 13750
rect 7150 13708 7158 13742
rect 7192 13708 7200 13742
rect 7150 13700 7200 13708
rect 7700 13742 7750 13750
rect 7700 13708 7708 13742
rect 7742 13708 7750 13742
rect 7700 13700 7750 13708
rect 8250 13742 8300 13750
rect 8250 13708 8258 13742
rect 8292 13708 8300 13742
rect 8250 13700 8300 13708
rect 8800 13742 8850 13750
rect 8800 13708 8808 13742
rect 8842 13708 8850 13742
rect 8800 13700 8850 13708
rect 9350 13742 9400 13750
rect 9350 13708 9358 13742
rect 9392 13708 9400 13742
rect 9350 13700 9400 13708
rect 9900 13742 9950 13750
rect 9900 13708 9908 13742
rect 9942 13708 9950 13742
rect 9900 13700 9950 13708
rect 10450 13742 10500 13750
rect 10450 13708 10458 13742
rect 10492 13708 10500 13742
rect 10450 13700 10500 13708
rect 11000 13742 11050 13750
rect 11000 13708 11008 13742
rect 11042 13708 11050 13742
rect 11000 13700 11050 13708
rect 11550 13742 11600 13750
rect 11550 13708 11558 13742
rect 11592 13708 11600 13742
rect 11550 13700 11600 13708
rect 12100 13742 12150 13750
rect 12100 13708 12108 13742
rect 12142 13708 12150 13742
rect 12100 13700 12150 13708
rect 12650 13742 12700 13750
rect 12650 13708 12658 13742
rect 12692 13708 12700 13742
rect 12650 13700 12700 13708
rect 13200 13742 13250 13750
rect 13200 13708 13208 13742
rect 13242 13708 13250 13742
rect 13200 13700 13250 13708
rect 13750 13742 13800 13750
rect 13750 13708 13758 13742
rect 13792 13708 13800 13742
rect 13750 13700 13800 13708
rect -474 13669 -26 13674
rect 76 13669 524 13674
rect 626 13669 1074 13674
rect 1176 13669 1624 13674
rect 1726 13669 2174 13674
rect 2276 13669 2724 13674
rect 2826 13669 3274 13674
rect 3376 13669 3824 13674
rect 3926 13669 4374 13674
rect 4476 13669 4924 13674
rect 5026 13669 5474 13674
rect 5576 13669 6024 13674
rect 6126 13669 6574 13674
rect 6676 13669 7124 13674
rect 7226 13669 7674 13674
rect 7776 13669 8224 13674
rect 8326 13669 8774 13674
rect 8876 13669 9324 13674
rect 9426 13669 9874 13674
rect 9976 13669 10424 13674
rect 10526 13669 10974 13674
rect 11076 13669 11524 13674
rect 11626 13669 12074 13674
rect 12176 13669 12624 13674
rect 12726 13669 13174 13674
rect 13276 13669 13724 13674
rect -474 13663 -3 13669
rect -474 13615 -23 13663
rect -474 13285 -415 13615
rect -85 13285 -23 13615
rect -474 13237 -23 13285
rect -6 13237 -3 13663
rect -474 13231 -3 13237
rect 53 13663 547 13669
rect 53 13237 56 13663
rect 73 13615 527 13663
rect 73 13285 135 13615
rect 465 13285 527 13615
rect 73 13237 527 13285
rect 544 13237 547 13663
rect 53 13231 547 13237
rect 603 13663 1097 13669
rect 603 13237 606 13663
rect 623 13615 1077 13663
rect 623 13285 685 13615
rect 1015 13285 1077 13615
rect 623 13237 1077 13285
rect 1094 13237 1097 13663
rect 603 13231 1097 13237
rect 1153 13663 1647 13669
rect 1153 13237 1156 13663
rect 1173 13615 1627 13663
rect 1173 13285 1235 13615
rect 1565 13285 1627 13615
rect 1173 13237 1627 13285
rect 1644 13237 1647 13663
rect 1153 13231 1647 13237
rect 1703 13663 2197 13669
rect 1703 13237 1706 13663
rect 1723 13615 2177 13663
rect 1723 13285 1785 13615
rect 2115 13285 2177 13615
rect 1723 13237 2177 13285
rect 2194 13237 2197 13663
rect 1703 13231 2197 13237
rect 2253 13663 2747 13669
rect 2253 13237 2256 13663
rect 2273 13615 2727 13663
rect 2273 13285 2335 13615
rect 2665 13285 2727 13615
rect 2273 13237 2727 13285
rect 2744 13237 2747 13663
rect 2253 13231 2747 13237
rect 2803 13663 3297 13669
rect 2803 13237 2806 13663
rect 2823 13615 3277 13663
rect 2823 13285 2885 13615
rect 3215 13285 3277 13615
rect 2823 13237 3277 13285
rect 3294 13237 3297 13663
rect 2803 13231 3297 13237
rect 3353 13663 3847 13669
rect 3353 13237 3356 13663
rect 3373 13615 3827 13663
rect 3373 13285 3435 13615
rect 3765 13285 3827 13615
rect 3373 13237 3827 13285
rect 3844 13237 3847 13663
rect 3353 13231 3847 13237
rect 3903 13663 4397 13669
rect 3903 13237 3906 13663
rect 3923 13615 4377 13663
rect 3923 13285 3985 13615
rect 4315 13285 4377 13615
rect 3923 13237 4377 13285
rect 4394 13237 4397 13663
rect 3903 13231 4397 13237
rect 4453 13663 4947 13669
rect 4453 13237 4456 13663
rect 4473 13615 4927 13663
rect 4473 13285 4535 13615
rect 4865 13285 4927 13615
rect 4473 13237 4927 13285
rect 4944 13237 4947 13663
rect 4453 13231 4947 13237
rect 5003 13663 5497 13669
rect 5003 13237 5006 13663
rect 5023 13615 5477 13663
rect 5023 13285 5085 13615
rect 5415 13285 5477 13615
rect 5023 13237 5477 13285
rect 5494 13237 5497 13663
rect 5003 13231 5497 13237
rect 5553 13663 6047 13669
rect 5553 13237 5556 13663
rect 5573 13615 6027 13663
rect 5573 13285 5635 13615
rect 5965 13285 6027 13615
rect 5573 13237 6027 13285
rect 6044 13237 6047 13663
rect 5553 13231 6047 13237
rect 6103 13663 6597 13669
rect 6103 13237 6106 13663
rect 6123 13615 6577 13663
rect 6123 13285 6185 13615
rect 6515 13285 6577 13615
rect 6123 13237 6577 13285
rect 6594 13237 6597 13663
rect 6103 13231 6597 13237
rect 6653 13663 7147 13669
rect 6653 13237 6656 13663
rect 6673 13615 7127 13663
rect 6673 13285 6735 13615
rect 7065 13285 7127 13615
rect 6673 13237 7127 13285
rect 7144 13237 7147 13663
rect 6653 13231 7147 13237
rect 7203 13663 7697 13669
rect 7203 13237 7206 13663
rect 7223 13615 7677 13663
rect 7223 13285 7285 13615
rect 7615 13285 7677 13615
rect 7223 13237 7677 13285
rect 7694 13237 7697 13663
rect 7203 13231 7697 13237
rect 7753 13663 8247 13669
rect 7753 13237 7756 13663
rect 7773 13615 8227 13663
rect 7773 13285 7835 13615
rect 8165 13285 8227 13615
rect 7773 13237 8227 13285
rect 8244 13237 8247 13663
rect 7753 13231 8247 13237
rect 8303 13663 8797 13669
rect 8303 13237 8306 13663
rect 8323 13615 8777 13663
rect 8323 13285 8385 13615
rect 8715 13285 8777 13615
rect 8323 13237 8777 13285
rect 8794 13237 8797 13663
rect 8303 13231 8797 13237
rect 8853 13663 9347 13669
rect 8853 13237 8856 13663
rect 8873 13615 9327 13663
rect 8873 13285 8935 13615
rect 9265 13285 9327 13615
rect 8873 13237 9327 13285
rect 9344 13237 9347 13663
rect 8853 13231 9347 13237
rect 9403 13663 9897 13669
rect 9403 13237 9406 13663
rect 9423 13615 9877 13663
rect 9423 13285 9485 13615
rect 9815 13285 9877 13615
rect 9423 13237 9877 13285
rect 9894 13237 9897 13663
rect 9403 13231 9897 13237
rect 9953 13663 10447 13669
rect 9953 13237 9956 13663
rect 9973 13615 10427 13663
rect 9973 13285 10035 13615
rect 10365 13285 10427 13615
rect 9973 13237 10427 13285
rect 10444 13237 10447 13663
rect 9953 13231 10447 13237
rect 10503 13663 10997 13669
rect 10503 13237 10506 13663
rect 10523 13615 10977 13663
rect 10523 13285 10585 13615
rect 10915 13285 10977 13615
rect 10523 13237 10977 13285
rect 10994 13237 10997 13663
rect 10503 13231 10997 13237
rect 11053 13663 11547 13669
rect 11053 13237 11056 13663
rect 11073 13615 11527 13663
rect 11073 13285 11135 13615
rect 11465 13285 11527 13615
rect 11073 13237 11527 13285
rect 11544 13237 11547 13663
rect 11053 13231 11547 13237
rect 11603 13663 12097 13669
rect 11603 13237 11606 13663
rect 11623 13615 12077 13663
rect 11623 13285 11685 13615
rect 12015 13285 12077 13615
rect 11623 13237 12077 13285
rect 12094 13237 12097 13663
rect 11603 13231 12097 13237
rect 12153 13663 12647 13669
rect 12153 13237 12156 13663
rect 12173 13615 12627 13663
rect 12173 13285 12235 13615
rect 12565 13285 12627 13615
rect 12173 13237 12627 13285
rect 12644 13237 12647 13663
rect 12153 13231 12647 13237
rect 12703 13663 13197 13669
rect 12703 13237 12706 13663
rect 12723 13615 13177 13663
rect 12723 13285 12785 13615
rect 13115 13285 13177 13615
rect 12723 13237 13177 13285
rect 13194 13237 13197 13663
rect 12703 13231 13197 13237
rect 13253 13663 13724 13669
rect 13253 13237 13256 13663
rect 13273 13615 13724 13663
rect 13273 13285 13335 13615
rect 13665 13285 13724 13615
rect 13273 13237 13724 13285
rect 13253 13231 13724 13237
rect -474 13226 -26 13231
rect 76 13226 524 13231
rect 626 13226 1074 13231
rect 1176 13226 1624 13231
rect 1726 13226 2174 13231
rect 2276 13226 2724 13231
rect 2826 13226 3274 13231
rect 3376 13226 3824 13231
rect 3926 13226 4374 13231
rect 4476 13226 4924 13231
rect 5026 13226 5474 13231
rect 5576 13226 6024 13231
rect 6126 13226 6574 13231
rect 6676 13226 7124 13231
rect 7226 13226 7674 13231
rect 7776 13226 8224 13231
rect 8326 13226 8774 13231
rect 8876 13226 9324 13231
rect 9426 13226 9874 13231
rect 9976 13226 10424 13231
rect 10526 13226 10974 13231
rect 11076 13226 11524 13231
rect 11626 13226 12074 13231
rect 12176 13226 12624 13231
rect 12726 13226 13174 13231
rect 13276 13226 13724 13231
rect -1025 13200 -725 13219
rect -469 13223 -31 13226
rect -469 13206 -463 13223
rect -37 13206 -31 13223
rect -469 13203 -31 13206
rect 81 13223 519 13226
rect 81 13206 87 13223
rect 513 13206 519 13223
rect 81 13203 519 13206
rect 631 13223 1069 13226
rect 631 13206 637 13223
rect 1063 13206 1069 13223
rect 631 13203 1069 13206
rect 1181 13223 1619 13226
rect 1181 13206 1187 13223
rect 1613 13206 1619 13223
rect 1181 13203 1619 13206
rect 1731 13223 2169 13226
rect 1731 13206 1737 13223
rect 2163 13206 2169 13223
rect 1731 13203 2169 13206
rect 2281 13223 2719 13226
rect 2281 13206 2287 13223
rect 2713 13206 2719 13223
rect 2281 13203 2719 13206
rect 2831 13223 3269 13226
rect 2831 13206 2837 13223
rect 3263 13206 3269 13223
rect 2831 13203 3269 13206
rect 3381 13223 3819 13226
rect 3381 13206 3387 13223
rect 3813 13206 3819 13223
rect 3381 13203 3819 13206
rect 3931 13223 4369 13226
rect 3931 13206 3937 13223
rect 4363 13206 4369 13223
rect 3931 13203 4369 13206
rect 4481 13223 4919 13226
rect 4481 13206 4487 13223
rect 4913 13206 4919 13223
rect 4481 13203 4919 13206
rect 5031 13223 5469 13226
rect 5031 13206 5037 13223
rect 5463 13206 5469 13223
rect 5031 13203 5469 13206
rect 5581 13223 6019 13226
rect 5581 13206 5587 13223
rect 6013 13206 6019 13223
rect 5581 13203 6019 13206
rect 6131 13223 6569 13226
rect 6131 13206 6137 13223
rect 6563 13206 6569 13223
rect 6131 13203 6569 13206
rect 6681 13223 7119 13226
rect 6681 13206 6687 13223
rect 7113 13206 7119 13223
rect 6681 13203 7119 13206
rect 7231 13223 7669 13226
rect 7231 13206 7237 13223
rect 7663 13206 7669 13223
rect 7231 13203 7669 13206
rect 7781 13223 8219 13226
rect 7781 13206 7787 13223
rect 8213 13206 8219 13223
rect 7781 13203 8219 13206
rect 8331 13223 8769 13226
rect 8331 13206 8337 13223
rect 8763 13206 8769 13223
rect 8331 13203 8769 13206
rect 8881 13223 9319 13226
rect 8881 13206 8887 13223
rect 9313 13206 9319 13223
rect 8881 13203 9319 13206
rect 9431 13223 9869 13226
rect 9431 13206 9437 13223
rect 9863 13206 9869 13223
rect 9431 13203 9869 13206
rect 9981 13223 10419 13226
rect 9981 13206 9987 13223
rect 10413 13206 10419 13223
rect 9981 13203 10419 13206
rect 10531 13223 10969 13226
rect 10531 13206 10537 13223
rect 10963 13206 10969 13223
rect 10531 13203 10969 13206
rect 11081 13223 11519 13226
rect 11081 13206 11087 13223
rect 11513 13206 11519 13223
rect 11081 13203 11519 13206
rect 11631 13223 12069 13226
rect 11631 13206 11637 13223
rect 12063 13206 12069 13223
rect 11631 13203 12069 13206
rect 12181 13223 12619 13226
rect 12181 13206 12187 13223
rect 12613 13206 12619 13223
rect 12181 13203 12619 13206
rect 12731 13223 13169 13226
rect 12731 13206 12737 13223
rect 13163 13206 13169 13223
rect 12731 13203 13169 13206
rect 13281 13223 13719 13226
rect 13281 13206 13287 13223
rect 13713 13206 13719 13223
rect 13281 13203 13719 13206
rect 13975 13219 13987 13925
rect 14263 13219 14275 14213
rect 13975 13200 14275 13219
rect -1025 12669 -1013 13200
rect -737 12669 -725 13200
rect -550 13192 -500 13200
rect -550 13158 -542 13192
rect -508 13158 -500 13192
rect -550 13150 -500 13158
rect 0 13192 50 13200
rect 0 13158 8 13192
rect 42 13158 50 13192
rect 0 13150 50 13158
rect 550 13192 600 13200
rect 550 13158 558 13192
rect 592 13158 600 13192
rect 550 13150 600 13158
rect 1100 13192 1150 13200
rect 1100 13158 1108 13192
rect 1142 13158 1150 13192
rect 1100 13150 1150 13158
rect 1650 13192 1700 13200
rect 1650 13158 1658 13192
rect 1692 13158 1700 13192
rect 1650 13150 1700 13158
rect 2200 13192 2250 13200
rect 2200 13158 2208 13192
rect 2242 13158 2250 13192
rect 2200 13150 2250 13158
rect 2750 13192 2800 13200
rect 2750 13158 2758 13192
rect 2792 13158 2800 13192
rect 2750 13150 2800 13158
rect 3300 13192 3350 13200
rect 3300 13158 3308 13192
rect 3342 13158 3350 13192
rect 3300 13150 3350 13158
rect 3850 13192 3900 13200
rect 3850 13158 3858 13192
rect 3892 13158 3900 13192
rect 3850 13150 3900 13158
rect 4400 13192 4450 13200
rect 4400 13158 4408 13192
rect 4442 13158 4450 13192
rect 4400 13150 4450 13158
rect 4950 13192 5000 13200
rect 4950 13158 4958 13192
rect 4992 13158 5000 13192
rect 4950 13150 5000 13158
rect 5500 13192 5550 13200
rect 5500 13158 5508 13192
rect 5542 13158 5550 13192
rect 5500 13150 5550 13158
rect 6050 13192 6100 13200
rect 6050 13158 6058 13192
rect 6092 13158 6100 13192
rect 6050 13150 6100 13158
rect 6600 13192 6650 13200
rect 6600 13158 6608 13192
rect 6642 13158 6650 13192
rect 6600 13150 6650 13158
rect 7150 13192 7200 13200
rect 7150 13158 7158 13192
rect 7192 13158 7200 13192
rect 7150 13150 7200 13158
rect 7700 13192 7750 13200
rect 7700 13158 7708 13192
rect 7742 13158 7750 13192
rect 7700 13150 7750 13158
rect 8250 13192 8300 13200
rect 8250 13158 8258 13192
rect 8292 13158 8300 13192
rect 8250 13150 8300 13158
rect 8800 13192 8850 13200
rect 8800 13158 8808 13192
rect 8842 13158 8850 13192
rect 8800 13150 8850 13158
rect 9350 13192 9400 13200
rect 9350 13158 9358 13192
rect 9392 13158 9400 13192
rect 9350 13150 9400 13158
rect 9900 13192 9950 13200
rect 9900 13158 9908 13192
rect 9942 13158 9950 13192
rect 9900 13150 9950 13158
rect 10450 13192 10500 13200
rect 10450 13158 10458 13192
rect 10492 13158 10500 13192
rect 10450 13150 10500 13158
rect 11000 13192 11050 13200
rect 11000 13158 11008 13192
rect 11042 13158 11050 13192
rect 11000 13150 11050 13158
rect 11550 13192 11600 13200
rect 11550 13158 11558 13192
rect 11592 13158 11600 13192
rect 11550 13150 11600 13158
rect 12100 13192 12150 13200
rect 12100 13158 12108 13192
rect 12142 13158 12150 13192
rect 12100 13150 12150 13158
rect 12650 13192 12700 13200
rect 12650 13158 12658 13192
rect 12692 13158 12700 13192
rect 12650 13150 12700 13158
rect 13200 13192 13250 13200
rect 13200 13158 13208 13192
rect 13242 13158 13250 13192
rect 13200 13150 13250 13158
rect 13750 13192 13800 13200
rect 13750 13158 13758 13192
rect 13792 13158 13800 13192
rect 13750 13150 13800 13158
rect -469 13144 -31 13147
rect -469 13127 -463 13144
rect -37 13127 -31 13144
rect -469 13124 -31 13127
rect 81 13144 519 13147
rect 81 13127 87 13144
rect 513 13127 519 13144
rect 81 13124 519 13127
rect 631 13144 1069 13147
rect 631 13127 637 13144
rect 1063 13127 1069 13144
rect 631 13124 1069 13127
rect 1181 13144 1619 13147
rect 1181 13127 1187 13144
rect 1613 13127 1619 13144
rect 1181 13124 1619 13127
rect 1731 13144 2169 13147
rect 1731 13127 1737 13144
rect 2163 13127 2169 13144
rect 1731 13124 2169 13127
rect 2281 13144 2719 13147
rect 2281 13127 2287 13144
rect 2713 13127 2719 13144
rect 2281 13124 2719 13127
rect 2831 13144 3269 13147
rect 2831 13127 2837 13144
rect 3263 13127 3269 13144
rect 2831 13124 3269 13127
rect 3381 13144 3819 13147
rect 3381 13127 3387 13144
rect 3813 13127 3819 13144
rect 3381 13124 3819 13127
rect 3931 13144 4369 13147
rect 3931 13127 3937 13144
rect 4363 13127 4369 13144
rect 3931 13124 4369 13127
rect 4481 13144 4919 13147
rect 4481 13127 4487 13144
rect 4913 13127 4919 13144
rect 4481 13124 4919 13127
rect 5031 13144 5469 13147
rect 5031 13127 5037 13144
rect 5463 13127 5469 13144
rect 5031 13124 5469 13127
rect 5581 13144 6019 13147
rect 5581 13127 5587 13144
rect 6013 13127 6019 13144
rect 5581 13124 6019 13127
rect 6131 13144 6569 13147
rect 6131 13127 6137 13144
rect 6563 13127 6569 13144
rect 6131 13124 6569 13127
rect 6681 13144 7119 13147
rect 6681 13127 6687 13144
rect 7113 13127 7119 13144
rect 6681 13124 7119 13127
rect 7231 13144 7669 13147
rect 7231 13127 7237 13144
rect 7663 13127 7669 13144
rect 7231 13124 7669 13127
rect 7781 13144 8219 13147
rect 7781 13127 7787 13144
rect 8213 13127 8219 13144
rect 7781 13124 8219 13127
rect 8331 13144 8769 13147
rect 8331 13127 8337 13144
rect 8763 13127 8769 13144
rect 8331 13124 8769 13127
rect 8881 13144 9319 13147
rect 8881 13127 8887 13144
rect 9313 13127 9319 13144
rect 8881 13124 9319 13127
rect 9431 13144 9869 13147
rect 9431 13127 9437 13144
rect 9863 13127 9869 13144
rect 9431 13124 9869 13127
rect 9981 13144 10419 13147
rect 9981 13127 9987 13144
rect 10413 13127 10419 13144
rect 9981 13124 10419 13127
rect 10531 13144 10969 13147
rect 10531 13127 10537 13144
rect 10963 13127 10969 13144
rect 10531 13124 10969 13127
rect 11081 13144 11519 13147
rect 11081 13127 11087 13144
rect 11513 13127 11519 13144
rect 11081 13124 11519 13127
rect 11631 13144 12069 13147
rect 11631 13127 11637 13144
rect 12063 13127 12069 13144
rect 11631 13124 12069 13127
rect 12181 13144 12619 13147
rect 12181 13127 12187 13144
rect 12613 13127 12619 13144
rect 12181 13124 12619 13127
rect 12731 13144 13169 13147
rect 12731 13127 12737 13144
rect 13163 13127 13169 13144
rect 12731 13124 13169 13127
rect 13281 13144 13719 13147
rect 13281 13127 13287 13144
rect 13713 13127 13719 13144
rect 13281 13124 13719 13127
rect -474 13119 -26 13124
rect 76 13119 524 13124
rect 626 13119 1074 13124
rect 1176 13119 1624 13124
rect 1726 13119 2174 13124
rect 2276 13119 2724 13124
rect 2826 13119 3274 13124
rect 3376 13119 3824 13124
rect 3926 13119 4374 13124
rect 4476 13119 4924 13124
rect 5026 13119 5474 13124
rect 5576 13119 6024 13124
rect 6126 13119 6574 13124
rect 6676 13119 7124 13124
rect 7226 13119 7674 13124
rect 7776 13119 8224 13124
rect 8326 13119 8774 13124
rect 8876 13119 9324 13124
rect 9426 13119 9874 13124
rect 9976 13119 10424 13124
rect 10526 13119 10974 13124
rect 11076 13119 11524 13124
rect 11626 13119 12074 13124
rect 12176 13119 12624 13124
rect 12726 13119 13174 13124
rect 13276 13119 13724 13124
rect -474 13113 -3 13119
rect -474 13065 -23 13113
rect -474 12735 -415 13065
rect -85 12735 -23 13065
rect -474 12687 -23 12735
rect -6 12687 -3 13113
rect -474 12681 -3 12687
rect 53 13113 547 13119
rect 53 12687 56 13113
rect 73 13065 527 13113
rect 73 12735 135 13065
rect 465 12735 527 13065
rect 73 12687 527 12735
rect 544 12687 547 13113
rect 53 12681 547 12687
rect 603 13113 1097 13119
rect 603 12687 606 13113
rect 623 13065 1077 13113
rect 623 12735 685 13065
rect 1015 12735 1077 13065
rect 623 12687 1077 12735
rect 1094 12687 1097 13113
rect 603 12681 1097 12687
rect 1153 13113 1647 13119
rect 1153 12687 1156 13113
rect 1173 13065 1627 13113
rect 1173 12735 1235 13065
rect 1565 12735 1627 13065
rect 1173 12687 1627 12735
rect 1644 12687 1647 13113
rect 1153 12681 1647 12687
rect 1703 13113 2197 13119
rect 1703 12687 1706 13113
rect 1723 13065 2177 13113
rect 1723 12735 1785 13065
rect 2115 12735 2177 13065
rect 1723 12687 2177 12735
rect 2194 12687 2197 13113
rect 1703 12681 2197 12687
rect 2253 13113 2747 13119
rect 2253 12687 2256 13113
rect 2273 13065 2727 13113
rect 2273 12735 2335 13065
rect 2665 12735 2727 13065
rect 2273 12687 2727 12735
rect 2744 12687 2747 13113
rect 2253 12681 2747 12687
rect 2803 13113 3297 13119
rect 2803 12687 2806 13113
rect 2823 13065 3277 13113
rect 2823 12735 2885 13065
rect 3215 12735 3277 13065
rect 2823 12687 3277 12735
rect 3294 12687 3297 13113
rect 2803 12681 3297 12687
rect 3353 13113 3847 13119
rect 3353 12687 3356 13113
rect 3373 13065 3827 13113
rect 3373 12735 3435 13065
rect 3765 12735 3827 13065
rect 3373 12687 3827 12735
rect 3844 12687 3847 13113
rect 3353 12681 3847 12687
rect 3903 13113 4397 13119
rect 3903 12687 3906 13113
rect 3923 13065 4377 13113
rect 3923 12735 3985 13065
rect 4315 12735 4377 13065
rect 3923 12687 4377 12735
rect 4394 12687 4397 13113
rect 3903 12681 4397 12687
rect 4453 13113 4947 13119
rect 4453 12687 4456 13113
rect 4473 13065 4927 13113
rect 4473 12735 4535 13065
rect 4865 12735 4927 13065
rect 4473 12687 4927 12735
rect 4944 12687 4947 13113
rect 4453 12681 4947 12687
rect 5003 13113 5497 13119
rect 5003 12687 5006 13113
rect 5023 13065 5477 13113
rect 5023 12735 5085 13065
rect 5415 12735 5477 13065
rect 5023 12687 5477 12735
rect 5494 12687 5497 13113
rect 5003 12681 5497 12687
rect 5553 13113 6047 13119
rect 5553 12687 5556 13113
rect 5573 13065 6027 13113
rect 5573 12735 5635 13065
rect 5965 12735 6027 13065
rect 5573 12687 6027 12735
rect 6044 12687 6047 13113
rect 5553 12681 6047 12687
rect 6103 13113 6597 13119
rect 6103 12687 6106 13113
rect 6123 13065 6577 13113
rect 6123 12735 6185 13065
rect 6515 12735 6577 13065
rect 6123 12687 6577 12735
rect 6594 12687 6597 13113
rect 6103 12681 6597 12687
rect 6653 13113 7147 13119
rect 6653 12687 6656 13113
rect 6673 13065 7127 13113
rect 6673 12735 6735 13065
rect 7065 12735 7127 13065
rect 6673 12687 7127 12735
rect 7144 12687 7147 13113
rect 6653 12681 7147 12687
rect 7203 13113 7697 13119
rect 7203 12687 7206 13113
rect 7223 13065 7677 13113
rect 7223 12735 7285 13065
rect 7615 12735 7677 13065
rect 7223 12687 7677 12735
rect 7694 12687 7697 13113
rect 7203 12681 7697 12687
rect 7753 13113 8247 13119
rect 7753 12687 7756 13113
rect 7773 13065 8227 13113
rect 7773 12735 7835 13065
rect 8165 12735 8227 13065
rect 7773 12687 8227 12735
rect 8244 12687 8247 13113
rect 7753 12681 8247 12687
rect 8303 13113 8797 13119
rect 8303 12687 8306 13113
rect 8323 13065 8777 13113
rect 8323 12735 8385 13065
rect 8715 12735 8777 13065
rect 8323 12687 8777 12735
rect 8794 12687 8797 13113
rect 8303 12681 8797 12687
rect 8853 13113 9347 13119
rect 8853 12687 8856 13113
rect 8873 13065 9327 13113
rect 8873 12735 8935 13065
rect 9265 12735 9327 13065
rect 8873 12687 9327 12735
rect 9344 12687 9347 13113
rect 8853 12681 9347 12687
rect 9403 13113 9897 13119
rect 9403 12687 9406 13113
rect 9423 13065 9877 13113
rect 9423 12735 9485 13065
rect 9815 12735 9877 13065
rect 9423 12687 9877 12735
rect 9894 12687 9897 13113
rect 9403 12681 9897 12687
rect 9953 13113 10447 13119
rect 9953 12687 9956 13113
rect 9973 13065 10427 13113
rect 9973 12735 10035 13065
rect 10365 12735 10427 13065
rect 9973 12687 10427 12735
rect 10444 12687 10447 13113
rect 9953 12681 10447 12687
rect 10503 13113 10997 13119
rect 10503 12687 10506 13113
rect 10523 13065 10977 13113
rect 10523 12735 10585 13065
rect 10915 12735 10977 13065
rect 10523 12687 10977 12735
rect 10994 12687 10997 13113
rect 10503 12681 10997 12687
rect 11053 13113 11547 13119
rect 11053 12687 11056 13113
rect 11073 13065 11527 13113
rect 11073 12735 11135 13065
rect 11465 12735 11527 13065
rect 11073 12687 11527 12735
rect 11544 12687 11547 13113
rect 11053 12681 11547 12687
rect 11603 13113 12097 13119
rect 11603 12687 11606 13113
rect 11623 13065 12077 13113
rect 11623 12735 11685 13065
rect 12015 12735 12077 13065
rect 11623 12687 12077 12735
rect 12094 12687 12097 13113
rect 11603 12681 12097 12687
rect 12153 13113 12647 13119
rect 12153 12687 12156 13113
rect 12173 13065 12627 13113
rect 12173 12735 12235 13065
rect 12565 12735 12627 13065
rect 12173 12687 12627 12735
rect 12644 12687 12647 13113
rect 12153 12681 12647 12687
rect 12703 13113 13197 13119
rect 12703 12687 12706 13113
rect 12723 13065 13177 13113
rect 12723 12735 12785 13065
rect 13115 12735 13177 13065
rect 12723 12687 13177 12735
rect 13194 12687 13197 13113
rect 12703 12681 13197 12687
rect 13253 13113 13724 13119
rect 13253 12687 13256 13113
rect 13273 13065 13724 13113
rect 13273 12735 13335 13065
rect 13665 12735 13724 13065
rect 13273 12687 13724 12735
rect 13253 12681 13724 12687
rect -474 12676 -26 12681
rect 76 12676 524 12681
rect 626 12676 1074 12681
rect 1176 12676 1624 12681
rect 1726 12676 2174 12681
rect 2276 12676 2724 12681
rect 2826 12676 3274 12681
rect 3376 12676 3824 12681
rect 3926 12676 4374 12681
rect 4476 12676 4924 12681
rect 5026 12676 5474 12681
rect 5576 12676 6024 12681
rect 6126 12676 6574 12681
rect 6676 12676 7124 12681
rect 7226 12676 7674 12681
rect 7776 12676 8224 12681
rect 8326 12676 8774 12681
rect 8876 12676 9324 12681
rect 9426 12676 9874 12681
rect 9976 12676 10424 12681
rect 10526 12676 10974 12681
rect 11076 12676 11524 12681
rect 11626 12676 12074 12681
rect 12176 12676 12624 12681
rect 12726 12676 13174 12681
rect 13276 12676 13724 12681
rect -1025 12650 -725 12669
rect -469 12673 -31 12676
rect -469 12656 -463 12673
rect -37 12656 -31 12673
rect -469 12653 -31 12656
rect 81 12673 519 12676
rect 81 12656 87 12673
rect 513 12656 519 12673
rect 81 12653 519 12656
rect 631 12673 1069 12676
rect 631 12656 637 12673
rect 1063 12656 1069 12673
rect 631 12653 1069 12656
rect 1181 12673 1619 12676
rect 1181 12656 1187 12673
rect 1613 12656 1619 12673
rect 1181 12653 1619 12656
rect 1731 12673 2169 12676
rect 1731 12656 1737 12673
rect 2163 12656 2169 12673
rect 1731 12653 2169 12656
rect 2281 12673 2719 12676
rect 2281 12656 2287 12673
rect 2713 12656 2719 12673
rect 2281 12653 2719 12656
rect 2831 12673 3269 12676
rect 2831 12656 2837 12673
rect 3263 12656 3269 12673
rect 2831 12653 3269 12656
rect 3381 12673 3819 12676
rect 3381 12656 3387 12673
rect 3813 12656 3819 12673
rect 3381 12653 3819 12656
rect 3931 12673 4369 12676
rect 3931 12656 3937 12673
rect 4363 12656 4369 12673
rect 3931 12653 4369 12656
rect 4481 12673 4919 12676
rect 4481 12656 4487 12673
rect 4913 12656 4919 12673
rect 4481 12653 4919 12656
rect 5031 12673 5469 12676
rect 5031 12656 5037 12673
rect 5463 12656 5469 12673
rect 5031 12653 5469 12656
rect 5581 12673 6019 12676
rect 5581 12656 5587 12673
rect 6013 12656 6019 12673
rect 5581 12653 6019 12656
rect 6131 12673 6569 12676
rect 6131 12656 6137 12673
rect 6563 12656 6569 12673
rect 6131 12653 6569 12656
rect 6681 12673 7119 12676
rect 6681 12656 6687 12673
rect 7113 12656 7119 12673
rect 6681 12653 7119 12656
rect 7231 12673 7669 12676
rect 7231 12656 7237 12673
rect 7663 12656 7669 12673
rect 7231 12653 7669 12656
rect 7781 12673 8219 12676
rect 7781 12656 7787 12673
rect 8213 12656 8219 12673
rect 7781 12653 8219 12656
rect 8331 12673 8769 12676
rect 8331 12656 8337 12673
rect 8763 12656 8769 12673
rect 8331 12653 8769 12656
rect 8881 12673 9319 12676
rect 8881 12656 8887 12673
rect 9313 12656 9319 12673
rect 8881 12653 9319 12656
rect 9431 12673 9869 12676
rect 9431 12656 9437 12673
rect 9863 12656 9869 12673
rect 9431 12653 9869 12656
rect 9981 12673 10419 12676
rect 9981 12656 9987 12673
rect 10413 12656 10419 12673
rect 9981 12653 10419 12656
rect 10531 12673 10969 12676
rect 10531 12656 10537 12673
rect 10963 12656 10969 12673
rect 10531 12653 10969 12656
rect 11081 12673 11519 12676
rect 11081 12656 11087 12673
rect 11513 12656 11519 12673
rect 11081 12653 11519 12656
rect 11631 12673 12069 12676
rect 11631 12656 11637 12673
rect 12063 12656 12069 12673
rect 11631 12653 12069 12656
rect 12181 12673 12619 12676
rect 12181 12656 12187 12673
rect 12613 12656 12619 12673
rect 12181 12653 12619 12656
rect 12731 12673 13169 12676
rect 12731 12656 12737 12673
rect 13163 12656 13169 12673
rect 12731 12653 13169 12656
rect 13281 12673 13719 12676
rect 13281 12656 13287 12673
rect 13713 12656 13719 12673
rect 13281 12653 13719 12656
rect 13975 12669 13987 13200
rect 14263 12669 14275 13200
rect 13975 12650 14275 12669
rect -1025 12119 -1013 12650
rect -737 12119 -725 12650
rect -550 12642 -500 12650
rect -550 12608 -542 12642
rect -508 12608 -500 12642
rect -550 12600 -500 12608
rect 0 12642 50 12650
rect 0 12608 8 12642
rect 42 12608 50 12642
rect 0 12600 50 12608
rect 550 12642 600 12650
rect 550 12608 558 12642
rect 592 12608 600 12642
rect 550 12600 600 12608
rect 1100 12642 1150 12650
rect 1100 12608 1108 12642
rect 1142 12608 1150 12642
rect 1100 12600 1150 12608
rect 1650 12642 1700 12650
rect 1650 12608 1658 12642
rect 1692 12608 1700 12642
rect 1650 12600 1700 12608
rect 2200 12642 2250 12650
rect 2200 12608 2208 12642
rect 2242 12608 2250 12642
rect 2200 12600 2250 12608
rect 2750 12642 2800 12650
rect 2750 12608 2758 12642
rect 2792 12608 2800 12642
rect 2750 12600 2800 12608
rect 3300 12642 3350 12650
rect 3300 12608 3308 12642
rect 3342 12608 3350 12642
rect 3300 12600 3350 12608
rect 3850 12642 3900 12650
rect 3850 12608 3858 12642
rect 3892 12608 3900 12642
rect 3850 12600 3900 12608
rect 4400 12642 4450 12650
rect 4400 12608 4408 12642
rect 4442 12608 4450 12642
rect 4400 12600 4450 12608
rect 4950 12642 5000 12650
rect 4950 12608 4958 12642
rect 4992 12608 5000 12642
rect 4950 12600 5000 12608
rect 5500 12642 5550 12650
rect 5500 12608 5508 12642
rect 5542 12608 5550 12642
rect 5500 12600 5550 12608
rect 6050 12642 6100 12650
rect 6050 12608 6058 12642
rect 6092 12608 6100 12642
rect 6050 12600 6100 12608
rect 6600 12642 6650 12650
rect 6600 12608 6608 12642
rect 6642 12608 6650 12642
rect 6600 12600 6650 12608
rect 7150 12642 7200 12650
rect 7150 12608 7158 12642
rect 7192 12608 7200 12642
rect 7150 12600 7200 12608
rect 7700 12642 7750 12650
rect 7700 12608 7708 12642
rect 7742 12608 7750 12642
rect 7700 12600 7750 12608
rect 8250 12642 8300 12650
rect 8250 12608 8258 12642
rect 8292 12608 8300 12642
rect 8250 12600 8300 12608
rect 8800 12642 8850 12650
rect 8800 12608 8808 12642
rect 8842 12608 8850 12642
rect 8800 12600 8850 12608
rect 9350 12642 9400 12650
rect 9350 12608 9358 12642
rect 9392 12608 9400 12642
rect 9350 12600 9400 12608
rect 9900 12642 9950 12650
rect 9900 12608 9908 12642
rect 9942 12608 9950 12642
rect 9900 12600 9950 12608
rect 10450 12642 10500 12650
rect 10450 12608 10458 12642
rect 10492 12608 10500 12642
rect 10450 12600 10500 12608
rect 11000 12642 11050 12650
rect 11000 12608 11008 12642
rect 11042 12608 11050 12642
rect 11000 12600 11050 12608
rect 11550 12642 11600 12650
rect 11550 12608 11558 12642
rect 11592 12608 11600 12642
rect 11550 12600 11600 12608
rect 12100 12642 12150 12650
rect 12100 12608 12108 12642
rect 12142 12608 12150 12642
rect 12100 12600 12150 12608
rect 12650 12642 12700 12650
rect 12650 12608 12658 12642
rect 12692 12608 12700 12642
rect 12650 12600 12700 12608
rect 13200 12642 13250 12650
rect 13200 12608 13208 12642
rect 13242 12608 13250 12642
rect 13200 12600 13250 12608
rect 13750 12642 13800 12650
rect 13750 12608 13758 12642
rect 13792 12608 13800 12642
rect 13750 12600 13800 12608
rect -469 12594 -31 12597
rect -469 12577 -463 12594
rect -37 12577 -31 12594
rect -469 12574 -31 12577
rect 81 12594 519 12597
rect 81 12577 87 12594
rect 513 12577 519 12594
rect 81 12574 519 12577
rect 631 12594 1069 12597
rect 631 12577 637 12594
rect 1063 12577 1069 12594
rect 631 12574 1069 12577
rect 1181 12594 1619 12597
rect 1181 12577 1187 12594
rect 1613 12577 1619 12594
rect 1181 12574 1619 12577
rect 1731 12594 2169 12597
rect 1731 12577 1737 12594
rect 2163 12577 2169 12594
rect 1731 12574 2169 12577
rect 2281 12594 2719 12597
rect 2281 12577 2287 12594
rect 2713 12577 2719 12594
rect 2281 12574 2719 12577
rect 2831 12594 3269 12597
rect 2831 12577 2837 12594
rect 3263 12577 3269 12594
rect 2831 12574 3269 12577
rect 3381 12594 3819 12597
rect 3381 12577 3387 12594
rect 3813 12577 3819 12594
rect 3381 12574 3819 12577
rect 3931 12594 4369 12597
rect 3931 12577 3937 12594
rect 4363 12577 4369 12594
rect 3931 12574 4369 12577
rect 4481 12594 4919 12597
rect 4481 12577 4487 12594
rect 4913 12577 4919 12594
rect 4481 12574 4919 12577
rect 5031 12594 5469 12597
rect 5031 12577 5037 12594
rect 5463 12577 5469 12594
rect 5031 12574 5469 12577
rect 5581 12594 6019 12597
rect 5581 12577 5587 12594
rect 6013 12577 6019 12594
rect 5581 12574 6019 12577
rect 6131 12594 6569 12597
rect 6131 12577 6137 12594
rect 6563 12577 6569 12594
rect 6131 12574 6569 12577
rect 6681 12594 7119 12597
rect 6681 12577 6687 12594
rect 7113 12577 7119 12594
rect 6681 12574 7119 12577
rect 7231 12594 7669 12597
rect 7231 12577 7237 12594
rect 7663 12577 7669 12594
rect 7231 12574 7669 12577
rect 7781 12594 8219 12597
rect 7781 12577 7787 12594
rect 8213 12577 8219 12594
rect 7781 12574 8219 12577
rect 8331 12594 8769 12597
rect 8331 12577 8337 12594
rect 8763 12577 8769 12594
rect 8331 12574 8769 12577
rect 8881 12594 9319 12597
rect 8881 12577 8887 12594
rect 9313 12577 9319 12594
rect 8881 12574 9319 12577
rect 9431 12594 9869 12597
rect 9431 12577 9437 12594
rect 9863 12577 9869 12594
rect 9431 12574 9869 12577
rect 9981 12594 10419 12597
rect 9981 12577 9987 12594
rect 10413 12577 10419 12594
rect 9981 12574 10419 12577
rect 10531 12594 10969 12597
rect 10531 12577 10537 12594
rect 10963 12577 10969 12594
rect 10531 12574 10969 12577
rect 11081 12594 11519 12597
rect 11081 12577 11087 12594
rect 11513 12577 11519 12594
rect 11081 12574 11519 12577
rect 11631 12594 12069 12597
rect 11631 12577 11637 12594
rect 12063 12577 12069 12594
rect 11631 12574 12069 12577
rect 12181 12594 12619 12597
rect 12181 12577 12187 12594
rect 12613 12577 12619 12594
rect 12181 12574 12619 12577
rect 12731 12594 13169 12597
rect 12731 12577 12737 12594
rect 13163 12577 13169 12594
rect 12731 12574 13169 12577
rect 13281 12594 13719 12597
rect 13281 12577 13287 12594
rect 13713 12577 13719 12594
rect 13281 12574 13719 12577
rect -474 12569 -26 12574
rect 76 12569 524 12574
rect 626 12569 1074 12574
rect 1176 12569 1624 12574
rect 1726 12569 2174 12574
rect 2276 12569 2724 12574
rect 2826 12569 3274 12574
rect 3376 12569 3824 12574
rect 3926 12569 4374 12574
rect 4476 12569 4924 12574
rect 5026 12569 5474 12574
rect 5576 12569 6024 12574
rect 6126 12569 6574 12574
rect 6676 12569 7124 12574
rect 7226 12569 7674 12574
rect 7776 12569 8224 12574
rect 8326 12569 8774 12574
rect 8876 12569 9324 12574
rect 9426 12569 9874 12574
rect 9976 12569 10424 12574
rect 10526 12569 10974 12574
rect 11076 12569 11524 12574
rect 11626 12569 12074 12574
rect 12176 12569 12624 12574
rect 12726 12569 13174 12574
rect 13276 12569 13724 12574
rect -474 12563 -3 12569
rect -474 12515 -23 12563
rect -474 12185 -415 12515
rect -85 12185 -23 12515
rect -474 12137 -23 12185
rect -6 12137 -3 12563
rect -474 12131 -3 12137
rect 53 12563 547 12569
rect 53 12137 56 12563
rect 73 12515 527 12563
rect 73 12185 135 12515
rect 465 12185 527 12515
rect 73 12137 527 12185
rect 544 12137 547 12563
rect 53 12131 547 12137
rect 603 12563 1097 12569
rect 603 12137 606 12563
rect 623 12515 1077 12563
rect 623 12185 685 12515
rect 1015 12185 1077 12515
rect 623 12137 1077 12185
rect 1094 12137 1097 12563
rect 603 12131 1097 12137
rect 1153 12563 1647 12569
rect 1153 12137 1156 12563
rect 1173 12515 1627 12563
rect 1173 12185 1235 12515
rect 1565 12185 1627 12515
rect 1173 12137 1627 12185
rect 1644 12137 1647 12563
rect 1153 12131 1647 12137
rect 1703 12563 2197 12569
rect 1703 12137 1706 12563
rect 1723 12515 2177 12563
rect 1723 12185 1785 12515
rect 2115 12185 2177 12515
rect 1723 12137 2177 12185
rect 2194 12137 2197 12563
rect 1703 12131 2197 12137
rect 2253 12563 2747 12569
rect 2253 12137 2256 12563
rect 2273 12515 2727 12563
rect 2273 12185 2335 12515
rect 2665 12185 2727 12515
rect 2273 12137 2727 12185
rect 2744 12137 2747 12563
rect 2253 12131 2747 12137
rect 2803 12563 3297 12569
rect 2803 12137 2806 12563
rect 2823 12515 3277 12563
rect 2823 12185 2885 12515
rect 3215 12185 3277 12515
rect 2823 12137 3277 12185
rect 3294 12137 3297 12563
rect 2803 12131 3297 12137
rect 3353 12563 3847 12569
rect 3353 12137 3356 12563
rect 3373 12515 3827 12563
rect 3373 12185 3435 12515
rect 3765 12185 3827 12515
rect 3373 12137 3827 12185
rect 3844 12137 3847 12563
rect 3353 12131 3847 12137
rect 3903 12563 4397 12569
rect 3903 12137 3906 12563
rect 3923 12515 4377 12563
rect 3923 12185 3985 12515
rect 4315 12185 4377 12515
rect 3923 12137 4377 12185
rect 4394 12137 4397 12563
rect 3903 12131 4397 12137
rect 4453 12563 4947 12569
rect 4453 12137 4456 12563
rect 4473 12515 4927 12563
rect 4473 12185 4535 12515
rect 4865 12185 4927 12515
rect 4473 12137 4927 12185
rect 4944 12137 4947 12563
rect 4453 12131 4947 12137
rect 5003 12563 5497 12569
rect 5003 12137 5006 12563
rect 5023 12515 5477 12563
rect 5023 12185 5085 12515
rect 5415 12185 5477 12515
rect 5023 12137 5477 12185
rect 5494 12137 5497 12563
rect 5003 12131 5497 12137
rect 5553 12563 6047 12569
rect 5553 12137 5556 12563
rect 5573 12515 6027 12563
rect 5573 12185 5635 12515
rect 5965 12185 6027 12515
rect 5573 12137 6027 12185
rect 6044 12137 6047 12563
rect 5553 12131 6047 12137
rect 6103 12563 6597 12569
rect 6103 12137 6106 12563
rect 6123 12515 6577 12563
rect 6123 12185 6185 12515
rect 6515 12185 6577 12515
rect 6123 12137 6577 12185
rect 6594 12137 6597 12563
rect 6103 12131 6597 12137
rect 6653 12563 7147 12569
rect 6653 12137 6656 12563
rect 6673 12515 7127 12563
rect 6673 12185 6735 12515
rect 7065 12185 7127 12515
rect 6673 12137 7127 12185
rect 7144 12137 7147 12563
rect 6653 12131 7147 12137
rect 7203 12563 7697 12569
rect 7203 12137 7206 12563
rect 7223 12515 7677 12563
rect 7223 12185 7285 12515
rect 7615 12185 7677 12515
rect 7223 12137 7677 12185
rect 7694 12137 7697 12563
rect 7203 12131 7697 12137
rect 7753 12563 8247 12569
rect 7753 12137 7756 12563
rect 7773 12515 8227 12563
rect 7773 12185 7835 12515
rect 8165 12185 8227 12515
rect 7773 12137 8227 12185
rect 8244 12137 8247 12563
rect 7753 12131 8247 12137
rect 8303 12563 8797 12569
rect 8303 12137 8306 12563
rect 8323 12515 8777 12563
rect 8323 12185 8385 12515
rect 8715 12185 8777 12515
rect 8323 12137 8777 12185
rect 8794 12137 8797 12563
rect 8303 12131 8797 12137
rect 8853 12563 9347 12569
rect 8853 12137 8856 12563
rect 8873 12515 9327 12563
rect 8873 12185 8935 12515
rect 9265 12185 9327 12515
rect 8873 12137 9327 12185
rect 9344 12137 9347 12563
rect 8853 12131 9347 12137
rect 9403 12563 9897 12569
rect 9403 12137 9406 12563
rect 9423 12515 9877 12563
rect 9423 12185 9485 12515
rect 9815 12185 9877 12515
rect 9423 12137 9877 12185
rect 9894 12137 9897 12563
rect 9403 12131 9897 12137
rect 9953 12563 10447 12569
rect 9953 12137 9956 12563
rect 9973 12515 10427 12563
rect 9973 12185 10035 12515
rect 10365 12185 10427 12515
rect 9973 12137 10427 12185
rect 10444 12137 10447 12563
rect 9953 12131 10447 12137
rect 10503 12563 10997 12569
rect 10503 12137 10506 12563
rect 10523 12515 10977 12563
rect 10523 12185 10585 12515
rect 10915 12185 10977 12515
rect 10523 12137 10977 12185
rect 10994 12137 10997 12563
rect 10503 12131 10997 12137
rect 11053 12563 11547 12569
rect 11053 12137 11056 12563
rect 11073 12515 11527 12563
rect 11073 12185 11135 12515
rect 11465 12185 11527 12515
rect 11073 12137 11527 12185
rect 11544 12137 11547 12563
rect 11053 12131 11547 12137
rect 11603 12563 12097 12569
rect 11603 12137 11606 12563
rect 11623 12515 12077 12563
rect 11623 12185 11685 12515
rect 12015 12185 12077 12515
rect 11623 12137 12077 12185
rect 12094 12137 12097 12563
rect 11603 12131 12097 12137
rect 12153 12563 12647 12569
rect 12153 12137 12156 12563
rect 12173 12515 12627 12563
rect 12173 12185 12235 12515
rect 12565 12185 12627 12515
rect 12173 12137 12627 12185
rect 12644 12137 12647 12563
rect 12153 12131 12647 12137
rect 12703 12563 13197 12569
rect 12703 12137 12706 12563
rect 12723 12515 13177 12563
rect 12723 12185 12785 12515
rect 13115 12185 13177 12515
rect 12723 12137 13177 12185
rect 13194 12137 13197 12563
rect 12703 12131 13197 12137
rect 13253 12563 13724 12569
rect 13253 12137 13256 12563
rect 13273 12515 13724 12563
rect 13273 12185 13335 12515
rect 13665 12185 13724 12515
rect 13273 12137 13724 12185
rect 13253 12131 13724 12137
rect -474 12126 -26 12131
rect 76 12126 524 12131
rect 626 12126 1074 12131
rect 1176 12126 1624 12131
rect 1726 12126 2174 12131
rect 2276 12126 2724 12131
rect 2826 12126 3274 12131
rect 3376 12126 3824 12131
rect 3926 12126 4374 12131
rect 4476 12126 4924 12131
rect 5026 12126 5474 12131
rect 5576 12126 6024 12131
rect 6126 12126 6574 12131
rect 6676 12126 7124 12131
rect 7226 12126 7674 12131
rect 7776 12126 8224 12131
rect 8326 12126 8774 12131
rect 8876 12126 9324 12131
rect 9426 12126 9874 12131
rect 9976 12126 10424 12131
rect 10526 12126 10974 12131
rect 11076 12126 11524 12131
rect 11626 12126 12074 12131
rect 12176 12126 12624 12131
rect 12726 12126 13174 12131
rect 13276 12126 13724 12131
rect -1025 12100 -725 12119
rect -469 12123 -31 12126
rect -469 12106 -463 12123
rect -37 12106 -31 12123
rect -469 12103 -31 12106
rect 81 12123 519 12126
rect 81 12106 87 12123
rect 513 12106 519 12123
rect 81 12103 519 12106
rect 631 12123 1069 12126
rect 631 12106 637 12123
rect 1063 12106 1069 12123
rect 631 12103 1069 12106
rect 1181 12123 1619 12126
rect 1181 12106 1187 12123
rect 1613 12106 1619 12123
rect 1181 12103 1619 12106
rect 1731 12123 2169 12126
rect 1731 12106 1737 12123
rect 2163 12106 2169 12123
rect 1731 12103 2169 12106
rect 2281 12123 2719 12126
rect 2281 12106 2287 12123
rect 2713 12106 2719 12123
rect 2281 12103 2719 12106
rect 2831 12123 3269 12126
rect 2831 12106 2837 12123
rect 3263 12106 3269 12123
rect 2831 12103 3269 12106
rect 3381 12123 3819 12126
rect 3381 12106 3387 12123
rect 3813 12106 3819 12123
rect 3381 12103 3819 12106
rect 3931 12123 4369 12126
rect 3931 12106 3937 12123
rect 4363 12106 4369 12123
rect 3931 12103 4369 12106
rect 4481 12123 4919 12126
rect 4481 12106 4487 12123
rect 4913 12106 4919 12123
rect 4481 12103 4919 12106
rect 5031 12123 5469 12126
rect 5031 12106 5037 12123
rect 5463 12106 5469 12123
rect 5031 12103 5469 12106
rect 5581 12123 6019 12126
rect 5581 12106 5587 12123
rect 6013 12106 6019 12123
rect 5581 12103 6019 12106
rect 6131 12123 6569 12126
rect 6131 12106 6137 12123
rect 6563 12106 6569 12123
rect 6131 12103 6569 12106
rect 6681 12123 7119 12126
rect 6681 12106 6687 12123
rect 7113 12106 7119 12123
rect 6681 12103 7119 12106
rect 7231 12123 7669 12126
rect 7231 12106 7237 12123
rect 7663 12106 7669 12123
rect 7231 12103 7669 12106
rect 7781 12123 8219 12126
rect 7781 12106 7787 12123
rect 8213 12106 8219 12123
rect 7781 12103 8219 12106
rect 8331 12123 8769 12126
rect 8331 12106 8337 12123
rect 8763 12106 8769 12123
rect 8331 12103 8769 12106
rect 8881 12123 9319 12126
rect 8881 12106 8887 12123
rect 9313 12106 9319 12123
rect 8881 12103 9319 12106
rect 9431 12123 9869 12126
rect 9431 12106 9437 12123
rect 9863 12106 9869 12123
rect 9431 12103 9869 12106
rect 9981 12123 10419 12126
rect 9981 12106 9987 12123
rect 10413 12106 10419 12123
rect 9981 12103 10419 12106
rect 10531 12123 10969 12126
rect 10531 12106 10537 12123
rect 10963 12106 10969 12123
rect 10531 12103 10969 12106
rect 11081 12123 11519 12126
rect 11081 12106 11087 12123
rect 11513 12106 11519 12123
rect 11081 12103 11519 12106
rect 11631 12123 12069 12126
rect 11631 12106 11637 12123
rect 12063 12106 12069 12123
rect 11631 12103 12069 12106
rect 12181 12123 12619 12126
rect 12181 12106 12187 12123
rect 12613 12106 12619 12123
rect 12181 12103 12619 12106
rect 12731 12123 13169 12126
rect 12731 12106 12737 12123
rect 13163 12106 13169 12123
rect 12731 12103 13169 12106
rect 13281 12123 13719 12126
rect 13281 12106 13287 12123
rect 13713 12106 13719 12123
rect 13281 12103 13719 12106
rect 13975 12119 13987 12650
rect 14263 12119 14275 12650
rect 13975 12100 14275 12119
rect -1025 11569 -1013 12100
rect -737 11569 -725 12100
rect -550 12092 -500 12100
rect -550 12058 -542 12092
rect -508 12058 -500 12092
rect -550 12050 -500 12058
rect 0 12092 50 12100
rect 0 12058 8 12092
rect 42 12058 50 12092
rect 0 12050 50 12058
rect 550 12092 600 12100
rect 550 12058 558 12092
rect 592 12058 600 12092
rect 550 12050 600 12058
rect 1100 12092 1150 12100
rect 1100 12058 1108 12092
rect 1142 12058 1150 12092
rect 1100 12050 1150 12058
rect 1650 12092 1700 12100
rect 1650 12058 1658 12092
rect 1692 12058 1700 12092
rect 1650 12050 1700 12058
rect 2200 12092 2250 12100
rect 2200 12058 2208 12092
rect 2242 12058 2250 12092
rect 2200 12050 2250 12058
rect 2750 12092 2800 12100
rect 2750 12058 2758 12092
rect 2792 12058 2800 12092
rect 2750 12050 2800 12058
rect 3300 12092 3350 12100
rect 3300 12058 3308 12092
rect 3342 12058 3350 12092
rect 3300 12050 3350 12058
rect 3850 12092 3900 12100
rect 3850 12058 3858 12092
rect 3892 12058 3900 12092
rect 3850 12050 3900 12058
rect 4400 12092 4450 12100
rect 4400 12058 4408 12092
rect 4442 12058 4450 12092
rect 4400 12050 4450 12058
rect 4950 12092 5000 12100
rect 4950 12058 4958 12092
rect 4992 12058 5000 12092
rect 4950 12050 5000 12058
rect 5500 12092 5550 12100
rect 5500 12058 5508 12092
rect 5542 12058 5550 12092
rect 5500 12050 5550 12058
rect 6050 12092 6100 12100
rect 6050 12058 6058 12092
rect 6092 12058 6100 12092
rect 6050 12050 6100 12058
rect 6600 12092 6650 12100
rect 6600 12058 6608 12092
rect 6642 12058 6650 12092
rect 6600 12050 6650 12058
rect 7150 12092 7200 12100
rect 7150 12058 7158 12092
rect 7192 12058 7200 12092
rect 7150 12050 7200 12058
rect 7700 12092 7750 12100
rect 7700 12058 7708 12092
rect 7742 12058 7750 12092
rect 7700 12050 7750 12058
rect 8250 12092 8300 12100
rect 8250 12058 8258 12092
rect 8292 12058 8300 12092
rect 8250 12050 8300 12058
rect 8800 12092 8850 12100
rect 8800 12058 8808 12092
rect 8842 12058 8850 12092
rect 8800 12050 8850 12058
rect 9350 12092 9400 12100
rect 9350 12058 9358 12092
rect 9392 12058 9400 12092
rect 9350 12050 9400 12058
rect 9900 12092 9950 12100
rect 9900 12058 9908 12092
rect 9942 12058 9950 12092
rect 9900 12050 9950 12058
rect 10450 12092 10500 12100
rect 10450 12058 10458 12092
rect 10492 12058 10500 12092
rect 10450 12050 10500 12058
rect 11000 12092 11050 12100
rect 11000 12058 11008 12092
rect 11042 12058 11050 12092
rect 11000 12050 11050 12058
rect 11550 12092 11600 12100
rect 11550 12058 11558 12092
rect 11592 12058 11600 12092
rect 11550 12050 11600 12058
rect 12100 12092 12150 12100
rect 12100 12058 12108 12092
rect 12142 12058 12150 12092
rect 12100 12050 12150 12058
rect 12650 12092 12700 12100
rect 12650 12058 12658 12092
rect 12692 12058 12700 12092
rect 12650 12050 12700 12058
rect 13200 12092 13250 12100
rect 13200 12058 13208 12092
rect 13242 12058 13250 12092
rect 13200 12050 13250 12058
rect 13750 12092 13800 12100
rect 13750 12058 13758 12092
rect 13792 12058 13800 12092
rect 13750 12050 13800 12058
rect -469 12044 -31 12047
rect -469 12027 -463 12044
rect -37 12027 -31 12044
rect -469 12024 -31 12027
rect 81 12044 519 12047
rect 81 12027 87 12044
rect 513 12027 519 12044
rect 81 12024 519 12027
rect 631 12044 1069 12047
rect 631 12027 637 12044
rect 1063 12027 1069 12044
rect 631 12024 1069 12027
rect 1181 12044 1619 12047
rect 1181 12027 1187 12044
rect 1613 12027 1619 12044
rect 1181 12024 1619 12027
rect 1731 12044 2169 12047
rect 1731 12027 1737 12044
rect 2163 12027 2169 12044
rect 1731 12024 2169 12027
rect 2281 12044 2719 12047
rect 2281 12027 2287 12044
rect 2713 12027 2719 12044
rect 2281 12024 2719 12027
rect 2831 12044 3269 12047
rect 2831 12027 2837 12044
rect 3263 12027 3269 12044
rect 2831 12024 3269 12027
rect 3381 12044 3819 12047
rect 3381 12027 3387 12044
rect 3813 12027 3819 12044
rect 3381 12024 3819 12027
rect 3931 12044 4369 12047
rect 3931 12027 3937 12044
rect 4363 12027 4369 12044
rect 3931 12024 4369 12027
rect 4481 12044 4919 12047
rect 4481 12027 4487 12044
rect 4913 12027 4919 12044
rect 4481 12024 4919 12027
rect 5031 12044 5469 12047
rect 5031 12027 5037 12044
rect 5463 12027 5469 12044
rect 5031 12024 5469 12027
rect 5581 12044 6019 12047
rect 5581 12027 5587 12044
rect 6013 12027 6019 12044
rect 5581 12024 6019 12027
rect 6131 12044 6569 12047
rect 6131 12027 6137 12044
rect 6563 12027 6569 12044
rect 6131 12024 6569 12027
rect 6681 12044 7119 12047
rect 6681 12027 6687 12044
rect 7113 12027 7119 12044
rect 6681 12024 7119 12027
rect 7231 12044 7669 12047
rect 7231 12027 7237 12044
rect 7663 12027 7669 12044
rect 7231 12024 7669 12027
rect 7781 12044 8219 12047
rect 7781 12027 7787 12044
rect 8213 12027 8219 12044
rect 7781 12024 8219 12027
rect 8331 12044 8769 12047
rect 8331 12027 8337 12044
rect 8763 12027 8769 12044
rect 8331 12024 8769 12027
rect 8881 12044 9319 12047
rect 8881 12027 8887 12044
rect 9313 12027 9319 12044
rect 8881 12024 9319 12027
rect 9431 12044 9869 12047
rect 9431 12027 9437 12044
rect 9863 12027 9869 12044
rect 9431 12024 9869 12027
rect 9981 12044 10419 12047
rect 9981 12027 9987 12044
rect 10413 12027 10419 12044
rect 9981 12024 10419 12027
rect 10531 12044 10969 12047
rect 10531 12027 10537 12044
rect 10963 12027 10969 12044
rect 10531 12024 10969 12027
rect 11081 12044 11519 12047
rect 11081 12027 11087 12044
rect 11513 12027 11519 12044
rect 11081 12024 11519 12027
rect 11631 12044 12069 12047
rect 11631 12027 11637 12044
rect 12063 12027 12069 12044
rect 11631 12024 12069 12027
rect 12181 12044 12619 12047
rect 12181 12027 12187 12044
rect 12613 12027 12619 12044
rect 12181 12024 12619 12027
rect 12731 12044 13169 12047
rect 12731 12027 12737 12044
rect 13163 12027 13169 12044
rect 12731 12024 13169 12027
rect 13281 12044 13719 12047
rect 13281 12027 13287 12044
rect 13713 12027 13719 12044
rect 13281 12024 13719 12027
rect -474 12019 -26 12024
rect 76 12019 524 12024
rect 626 12019 1074 12024
rect 1176 12019 1624 12024
rect 1726 12019 2174 12024
rect 2276 12019 2724 12024
rect 2826 12019 3274 12024
rect 3376 12019 3824 12024
rect 3926 12019 4374 12024
rect 4476 12019 4924 12024
rect 5026 12019 5474 12024
rect 5576 12019 6024 12024
rect 6126 12019 6574 12024
rect 6676 12019 7124 12024
rect 7226 12019 7674 12024
rect 7776 12019 8224 12024
rect 8326 12019 8774 12024
rect 8876 12019 9324 12024
rect 9426 12019 9874 12024
rect 9976 12019 10424 12024
rect 10526 12019 10974 12024
rect 11076 12019 11524 12024
rect 11626 12019 12074 12024
rect 12176 12019 12624 12024
rect 12726 12019 13174 12024
rect 13276 12019 13724 12024
rect -474 12013 -3 12019
rect -474 11965 -23 12013
rect -474 11635 -415 11965
rect -85 11635 -23 11965
rect -474 11587 -23 11635
rect -6 11587 -3 12013
rect -474 11581 -3 11587
rect 53 12013 547 12019
rect 53 11587 56 12013
rect 73 11965 527 12013
rect 73 11635 135 11965
rect 465 11635 527 11965
rect 73 11587 527 11635
rect 544 11587 547 12013
rect 53 11581 547 11587
rect 603 12013 1097 12019
rect 603 11587 606 12013
rect 623 11965 1077 12013
rect 623 11635 685 11965
rect 1015 11635 1077 11965
rect 623 11587 1077 11635
rect 1094 11587 1097 12013
rect 603 11581 1097 11587
rect 1153 12013 1647 12019
rect 1153 11587 1156 12013
rect 1173 11965 1627 12013
rect 1173 11635 1235 11965
rect 1565 11635 1627 11965
rect 1173 11587 1627 11635
rect 1644 11587 1647 12013
rect 1153 11581 1647 11587
rect 1703 12013 2197 12019
rect 1703 11587 1706 12013
rect 1723 11965 2177 12013
rect 1723 11635 1785 11965
rect 2115 11635 2177 11965
rect 1723 11587 2177 11635
rect 2194 11587 2197 12013
rect 1703 11581 2197 11587
rect 2253 12013 2747 12019
rect 2253 11587 2256 12013
rect 2273 11965 2727 12013
rect 2273 11635 2335 11965
rect 2665 11635 2727 11965
rect 2273 11587 2727 11635
rect 2744 11587 2747 12013
rect 2253 11581 2747 11587
rect 2803 12013 3297 12019
rect 2803 11587 2806 12013
rect 2823 11965 3277 12013
rect 2823 11635 2885 11965
rect 3215 11635 3277 11965
rect 2823 11587 3277 11635
rect 3294 11587 3297 12013
rect 2803 11581 3297 11587
rect 3353 12013 3847 12019
rect 3353 11587 3356 12013
rect 3373 11965 3827 12013
rect 3373 11635 3435 11965
rect 3765 11635 3827 11965
rect 3373 11587 3827 11635
rect 3844 11587 3847 12013
rect 3353 11581 3847 11587
rect 3903 12013 4397 12019
rect 3903 11587 3906 12013
rect 3923 11965 4377 12013
rect 3923 11635 3985 11965
rect 4315 11635 4377 11965
rect 3923 11587 4377 11635
rect 4394 11587 4397 12013
rect 3903 11581 4397 11587
rect 4453 12013 4947 12019
rect 4453 11587 4456 12013
rect 4473 11965 4927 12013
rect 4473 11635 4535 11965
rect 4865 11635 4927 11965
rect 4473 11587 4927 11635
rect 4944 11587 4947 12013
rect 4453 11581 4947 11587
rect 5003 12013 5497 12019
rect 5003 11587 5006 12013
rect 5023 11965 5477 12013
rect 5023 11635 5085 11965
rect 5415 11635 5477 11965
rect 5023 11587 5477 11635
rect 5494 11587 5497 12013
rect 5003 11581 5497 11587
rect 5553 12013 6047 12019
rect 5553 11587 5556 12013
rect 5573 11965 6027 12013
rect 5573 11635 5635 11965
rect 5965 11635 6027 11965
rect 5573 11587 6027 11635
rect 6044 11587 6047 12013
rect 5553 11581 6047 11587
rect 6103 12013 6597 12019
rect 6103 11587 6106 12013
rect 6123 11965 6577 12013
rect 6123 11635 6185 11965
rect 6515 11635 6577 11965
rect 6123 11587 6577 11635
rect 6594 11587 6597 12013
rect 6103 11581 6597 11587
rect 6653 12013 7147 12019
rect 6653 11587 6656 12013
rect 6673 11965 7127 12013
rect 6673 11635 6735 11965
rect 7065 11635 7127 11965
rect 6673 11587 7127 11635
rect 7144 11587 7147 12013
rect 6653 11581 7147 11587
rect 7203 12013 7697 12019
rect 7203 11587 7206 12013
rect 7223 11965 7677 12013
rect 7223 11635 7285 11965
rect 7615 11635 7677 11965
rect 7223 11587 7677 11635
rect 7694 11587 7697 12013
rect 7203 11581 7697 11587
rect 7753 12013 8247 12019
rect 7753 11587 7756 12013
rect 7773 11965 8227 12013
rect 7773 11635 7835 11965
rect 8165 11635 8227 11965
rect 7773 11587 8227 11635
rect 8244 11587 8247 12013
rect 7753 11581 8247 11587
rect 8303 12013 8797 12019
rect 8303 11587 8306 12013
rect 8323 11965 8777 12013
rect 8323 11635 8385 11965
rect 8715 11635 8777 11965
rect 8323 11587 8777 11635
rect 8794 11587 8797 12013
rect 8303 11581 8797 11587
rect 8853 12013 9347 12019
rect 8853 11587 8856 12013
rect 8873 11965 9327 12013
rect 8873 11635 8935 11965
rect 9265 11635 9327 11965
rect 8873 11587 9327 11635
rect 9344 11587 9347 12013
rect 8853 11581 9347 11587
rect 9403 12013 9897 12019
rect 9403 11587 9406 12013
rect 9423 11965 9877 12013
rect 9423 11635 9485 11965
rect 9815 11635 9877 11965
rect 9423 11587 9877 11635
rect 9894 11587 9897 12013
rect 9403 11581 9897 11587
rect 9953 12013 10447 12019
rect 9953 11587 9956 12013
rect 9973 11965 10427 12013
rect 9973 11635 10035 11965
rect 10365 11635 10427 11965
rect 9973 11587 10427 11635
rect 10444 11587 10447 12013
rect 9953 11581 10447 11587
rect 10503 12013 10997 12019
rect 10503 11587 10506 12013
rect 10523 11965 10977 12013
rect 10523 11635 10585 11965
rect 10915 11635 10977 11965
rect 10523 11587 10977 11635
rect 10994 11587 10997 12013
rect 10503 11581 10997 11587
rect 11053 12013 11547 12019
rect 11053 11587 11056 12013
rect 11073 11965 11527 12013
rect 11073 11635 11135 11965
rect 11465 11635 11527 11965
rect 11073 11587 11527 11635
rect 11544 11587 11547 12013
rect 11053 11581 11547 11587
rect 11603 12013 12097 12019
rect 11603 11587 11606 12013
rect 11623 11965 12077 12013
rect 11623 11635 11685 11965
rect 12015 11635 12077 11965
rect 11623 11587 12077 11635
rect 12094 11587 12097 12013
rect 11603 11581 12097 11587
rect 12153 12013 12647 12019
rect 12153 11587 12156 12013
rect 12173 11965 12627 12013
rect 12173 11635 12235 11965
rect 12565 11635 12627 11965
rect 12173 11587 12627 11635
rect 12644 11587 12647 12013
rect 12153 11581 12647 11587
rect 12703 12013 13197 12019
rect 12703 11587 12706 12013
rect 12723 11965 13177 12013
rect 12723 11635 12785 11965
rect 13115 11635 13177 11965
rect 12723 11587 13177 11635
rect 13194 11587 13197 12013
rect 12703 11581 13197 11587
rect 13253 12013 13724 12019
rect 13253 11587 13256 12013
rect 13273 11965 13724 12013
rect 13273 11635 13335 11965
rect 13665 11635 13724 11965
rect 13273 11587 13724 11635
rect 13253 11581 13724 11587
rect -474 11576 -26 11581
rect 76 11576 524 11581
rect 626 11576 1074 11581
rect 1176 11576 1624 11581
rect 1726 11576 2174 11581
rect 2276 11576 2724 11581
rect 2826 11576 3274 11581
rect 3376 11576 3824 11581
rect 3926 11576 4374 11581
rect 4476 11576 4924 11581
rect 5026 11576 5474 11581
rect 5576 11576 6024 11581
rect 6126 11576 6574 11581
rect 6676 11576 7124 11581
rect 7226 11576 7674 11581
rect 7776 11576 8224 11581
rect 8326 11576 8774 11581
rect 8876 11576 9324 11581
rect 9426 11576 9874 11581
rect 9976 11576 10424 11581
rect 10526 11576 10974 11581
rect 11076 11576 11524 11581
rect 11626 11576 12074 11581
rect 12176 11576 12624 11581
rect 12726 11576 13174 11581
rect 13276 11576 13724 11581
rect -1025 11550 -725 11569
rect -469 11573 -31 11576
rect -469 11556 -463 11573
rect -37 11556 -31 11573
rect -469 11553 -31 11556
rect 81 11573 519 11576
rect 81 11556 87 11573
rect 513 11556 519 11573
rect 81 11553 519 11556
rect 631 11573 1069 11576
rect 631 11556 637 11573
rect 1063 11556 1069 11573
rect 631 11553 1069 11556
rect 1181 11573 1619 11576
rect 1181 11556 1187 11573
rect 1613 11556 1619 11573
rect 1181 11553 1619 11556
rect 1731 11573 2169 11576
rect 1731 11556 1737 11573
rect 2163 11556 2169 11573
rect 1731 11553 2169 11556
rect 2281 11573 2719 11576
rect 2281 11556 2287 11573
rect 2713 11556 2719 11573
rect 2281 11553 2719 11556
rect 2831 11573 3269 11576
rect 2831 11556 2837 11573
rect 3263 11556 3269 11573
rect 2831 11553 3269 11556
rect 3381 11573 3819 11576
rect 3381 11556 3387 11573
rect 3813 11556 3819 11573
rect 3381 11553 3819 11556
rect 3931 11573 4369 11576
rect 3931 11556 3937 11573
rect 4363 11556 4369 11573
rect 3931 11553 4369 11556
rect 4481 11573 4919 11576
rect 4481 11556 4487 11573
rect 4913 11556 4919 11573
rect 4481 11553 4919 11556
rect 5031 11573 5469 11576
rect 5031 11556 5037 11573
rect 5463 11556 5469 11573
rect 5031 11553 5469 11556
rect 5581 11573 6019 11576
rect 5581 11556 5587 11573
rect 6013 11556 6019 11573
rect 5581 11553 6019 11556
rect 6131 11573 6569 11576
rect 6131 11556 6137 11573
rect 6563 11556 6569 11573
rect 6131 11553 6569 11556
rect 6681 11573 7119 11576
rect 6681 11556 6687 11573
rect 7113 11556 7119 11573
rect 6681 11553 7119 11556
rect 7231 11573 7669 11576
rect 7231 11556 7237 11573
rect 7663 11556 7669 11573
rect 7231 11553 7669 11556
rect 7781 11573 8219 11576
rect 7781 11556 7787 11573
rect 8213 11556 8219 11573
rect 7781 11553 8219 11556
rect 8331 11573 8769 11576
rect 8331 11556 8337 11573
rect 8763 11556 8769 11573
rect 8331 11553 8769 11556
rect 8881 11573 9319 11576
rect 8881 11556 8887 11573
rect 9313 11556 9319 11573
rect 8881 11553 9319 11556
rect 9431 11573 9869 11576
rect 9431 11556 9437 11573
rect 9863 11556 9869 11573
rect 9431 11553 9869 11556
rect 9981 11573 10419 11576
rect 9981 11556 9987 11573
rect 10413 11556 10419 11573
rect 9981 11553 10419 11556
rect 10531 11573 10969 11576
rect 10531 11556 10537 11573
rect 10963 11556 10969 11573
rect 10531 11553 10969 11556
rect 11081 11573 11519 11576
rect 11081 11556 11087 11573
rect 11513 11556 11519 11573
rect 11081 11553 11519 11556
rect 11631 11573 12069 11576
rect 11631 11556 11637 11573
rect 12063 11556 12069 11573
rect 11631 11553 12069 11556
rect 12181 11573 12619 11576
rect 12181 11556 12187 11573
rect 12613 11556 12619 11573
rect 12181 11553 12619 11556
rect 12731 11573 13169 11576
rect 12731 11556 12737 11573
rect 13163 11556 13169 11573
rect 12731 11553 13169 11556
rect 13281 11573 13719 11576
rect 13281 11556 13287 11573
rect 13713 11556 13719 11573
rect 13281 11553 13719 11556
rect 13975 11569 13987 12100
rect 14263 11569 14275 12100
rect 13975 11550 14275 11569
rect -1025 11019 -1013 11550
rect -737 11019 -725 11550
rect -550 11542 -500 11550
rect -550 11508 -542 11542
rect -508 11508 -500 11542
rect -550 11500 -500 11508
rect 0 11542 50 11550
rect 0 11508 8 11542
rect 42 11508 50 11542
rect 0 11500 50 11508
rect 550 11542 600 11550
rect 550 11508 558 11542
rect 592 11508 600 11542
rect 550 11500 600 11508
rect 1100 11542 1150 11550
rect 1100 11508 1108 11542
rect 1142 11508 1150 11542
rect 1100 11500 1150 11508
rect 1650 11542 1700 11550
rect 1650 11508 1658 11542
rect 1692 11508 1700 11542
rect 1650 11500 1700 11508
rect 2200 11542 2250 11550
rect 2200 11508 2208 11542
rect 2242 11508 2250 11542
rect 2200 11500 2250 11508
rect 2750 11542 2800 11550
rect 2750 11508 2758 11542
rect 2792 11508 2800 11542
rect 2750 11500 2800 11508
rect 3300 11542 3350 11550
rect 3300 11508 3308 11542
rect 3342 11508 3350 11542
rect 3300 11500 3350 11508
rect 3850 11542 3900 11550
rect 3850 11508 3858 11542
rect 3892 11508 3900 11542
rect 3850 11500 3900 11508
rect 4400 11542 4450 11550
rect 4400 11508 4408 11542
rect 4442 11508 4450 11542
rect 4400 11500 4450 11508
rect 4950 11542 5000 11550
rect 4950 11508 4958 11542
rect 4992 11508 5000 11542
rect 4950 11500 5000 11508
rect 5500 11542 5550 11550
rect 5500 11508 5508 11542
rect 5542 11508 5550 11542
rect 5500 11500 5550 11508
rect 6050 11542 6100 11550
rect 6050 11508 6058 11542
rect 6092 11508 6100 11542
rect 6050 11500 6100 11508
rect 6600 11542 6650 11550
rect 6600 11508 6608 11542
rect 6642 11508 6650 11542
rect 6600 11500 6650 11508
rect 7150 11542 7200 11550
rect 7150 11508 7158 11542
rect 7192 11508 7200 11542
rect 7150 11500 7200 11508
rect 7700 11542 7750 11550
rect 7700 11508 7708 11542
rect 7742 11508 7750 11542
rect 7700 11500 7750 11508
rect 8250 11542 8300 11550
rect 8250 11508 8258 11542
rect 8292 11508 8300 11542
rect 8250 11500 8300 11508
rect 8800 11542 8850 11550
rect 8800 11508 8808 11542
rect 8842 11508 8850 11542
rect 8800 11500 8850 11508
rect 9350 11542 9400 11550
rect 9350 11508 9358 11542
rect 9392 11508 9400 11542
rect 9350 11500 9400 11508
rect 9900 11542 9950 11550
rect 9900 11508 9908 11542
rect 9942 11508 9950 11542
rect 9900 11500 9950 11508
rect 10450 11542 10500 11550
rect 10450 11508 10458 11542
rect 10492 11508 10500 11542
rect 10450 11500 10500 11508
rect 11000 11542 11050 11550
rect 11000 11508 11008 11542
rect 11042 11508 11050 11542
rect 11000 11500 11050 11508
rect 11550 11542 11600 11550
rect 11550 11508 11558 11542
rect 11592 11508 11600 11542
rect 11550 11500 11600 11508
rect 12100 11542 12150 11550
rect 12100 11508 12108 11542
rect 12142 11508 12150 11542
rect 12100 11500 12150 11508
rect 12650 11542 12700 11550
rect 12650 11508 12658 11542
rect 12692 11508 12700 11542
rect 12650 11500 12700 11508
rect 13200 11542 13250 11550
rect 13200 11508 13208 11542
rect 13242 11508 13250 11542
rect 13200 11500 13250 11508
rect 13750 11542 13800 11550
rect 13750 11508 13758 11542
rect 13792 11508 13800 11542
rect 13750 11500 13800 11508
rect -469 11494 -31 11497
rect -469 11477 -463 11494
rect -37 11477 -31 11494
rect -469 11474 -31 11477
rect 81 11494 519 11497
rect 81 11477 87 11494
rect 513 11477 519 11494
rect 81 11474 519 11477
rect 631 11494 1069 11497
rect 631 11477 637 11494
rect 1063 11477 1069 11494
rect 631 11474 1069 11477
rect 1181 11494 1619 11497
rect 1181 11477 1187 11494
rect 1613 11477 1619 11494
rect 1181 11474 1619 11477
rect 1731 11494 2169 11497
rect 1731 11477 1737 11494
rect 2163 11477 2169 11494
rect 1731 11474 2169 11477
rect 2281 11494 2719 11497
rect 2281 11477 2287 11494
rect 2713 11477 2719 11494
rect 2281 11474 2719 11477
rect 2831 11494 3269 11497
rect 2831 11477 2837 11494
rect 3263 11477 3269 11494
rect 2831 11474 3269 11477
rect 3381 11494 3819 11497
rect 3381 11477 3387 11494
rect 3813 11477 3819 11494
rect 3381 11474 3819 11477
rect 3931 11494 4369 11497
rect 3931 11477 3937 11494
rect 4363 11477 4369 11494
rect 3931 11474 4369 11477
rect 4481 11494 4919 11497
rect 4481 11477 4487 11494
rect 4913 11477 4919 11494
rect 4481 11474 4919 11477
rect 5031 11494 5469 11497
rect 5031 11477 5037 11494
rect 5463 11477 5469 11494
rect 5031 11474 5469 11477
rect 5581 11494 6019 11497
rect 5581 11477 5587 11494
rect 6013 11477 6019 11494
rect 5581 11474 6019 11477
rect 6131 11494 6569 11497
rect 6131 11477 6137 11494
rect 6563 11477 6569 11494
rect 6131 11474 6569 11477
rect 6681 11494 7119 11497
rect 6681 11477 6687 11494
rect 7113 11477 7119 11494
rect 6681 11474 7119 11477
rect 7231 11494 7669 11497
rect 7231 11477 7237 11494
rect 7663 11477 7669 11494
rect 7231 11474 7669 11477
rect 7781 11494 8219 11497
rect 7781 11477 7787 11494
rect 8213 11477 8219 11494
rect 7781 11474 8219 11477
rect 8331 11494 8769 11497
rect 8331 11477 8337 11494
rect 8763 11477 8769 11494
rect 8331 11474 8769 11477
rect 8881 11494 9319 11497
rect 8881 11477 8887 11494
rect 9313 11477 9319 11494
rect 8881 11474 9319 11477
rect 9431 11494 9869 11497
rect 9431 11477 9437 11494
rect 9863 11477 9869 11494
rect 9431 11474 9869 11477
rect 9981 11494 10419 11497
rect 9981 11477 9987 11494
rect 10413 11477 10419 11494
rect 9981 11474 10419 11477
rect 10531 11494 10969 11497
rect 10531 11477 10537 11494
rect 10963 11477 10969 11494
rect 10531 11474 10969 11477
rect 11081 11494 11519 11497
rect 11081 11477 11087 11494
rect 11513 11477 11519 11494
rect 11081 11474 11519 11477
rect 11631 11494 12069 11497
rect 11631 11477 11637 11494
rect 12063 11477 12069 11494
rect 11631 11474 12069 11477
rect 12181 11494 12619 11497
rect 12181 11477 12187 11494
rect 12613 11477 12619 11494
rect 12181 11474 12619 11477
rect 12731 11494 13169 11497
rect 12731 11477 12737 11494
rect 13163 11477 13169 11494
rect 12731 11474 13169 11477
rect 13281 11494 13719 11497
rect 13281 11477 13287 11494
rect 13713 11477 13719 11494
rect 13281 11474 13719 11477
rect -474 11469 -26 11474
rect 76 11469 524 11474
rect 626 11469 1074 11474
rect 1176 11469 1624 11474
rect 1726 11469 2174 11474
rect 2276 11469 2724 11474
rect 2826 11469 3274 11474
rect 3376 11469 3824 11474
rect 3926 11469 4374 11474
rect 4476 11469 4924 11474
rect 5026 11469 5474 11474
rect 5576 11469 6024 11474
rect 6126 11469 6574 11474
rect 6676 11469 7124 11474
rect 7226 11469 7674 11474
rect 7776 11469 8224 11474
rect 8326 11469 8774 11474
rect 8876 11469 9324 11474
rect 9426 11469 9874 11474
rect 9976 11469 10424 11474
rect 10526 11469 10974 11474
rect 11076 11469 11524 11474
rect 11626 11469 12074 11474
rect 12176 11469 12624 11474
rect 12726 11469 13174 11474
rect 13276 11469 13724 11474
rect -474 11463 -3 11469
rect -474 11415 -23 11463
rect -474 11085 -415 11415
rect -85 11085 -23 11415
rect -474 11037 -23 11085
rect -6 11037 -3 11463
rect -474 11031 -3 11037
rect 53 11463 547 11469
rect 53 11037 56 11463
rect 73 11415 527 11463
rect 73 11085 135 11415
rect 465 11085 527 11415
rect 73 11037 527 11085
rect 544 11037 547 11463
rect 53 11031 547 11037
rect 603 11463 1097 11469
rect 603 11037 606 11463
rect 623 11415 1077 11463
rect 623 11085 685 11415
rect 1015 11085 1077 11415
rect 623 11037 1077 11085
rect 1094 11037 1097 11463
rect 603 11031 1097 11037
rect 1153 11463 1647 11469
rect 1153 11037 1156 11463
rect 1173 11415 1627 11463
rect 1173 11085 1235 11415
rect 1565 11085 1627 11415
rect 1173 11037 1627 11085
rect 1644 11037 1647 11463
rect 1153 11031 1647 11037
rect 1703 11463 2197 11469
rect 1703 11037 1706 11463
rect 1723 11415 2177 11463
rect 1723 11085 1785 11415
rect 2115 11085 2177 11415
rect 1723 11037 2177 11085
rect 2194 11037 2197 11463
rect 1703 11031 2197 11037
rect 2253 11463 2747 11469
rect 2253 11037 2256 11463
rect 2273 11415 2727 11463
rect 2273 11085 2335 11415
rect 2665 11085 2727 11415
rect 2273 11037 2727 11085
rect 2744 11037 2747 11463
rect 2253 11031 2747 11037
rect 2803 11463 3297 11469
rect 2803 11037 2806 11463
rect 2823 11415 3277 11463
rect 2823 11085 2885 11415
rect 3215 11085 3277 11415
rect 2823 11037 3277 11085
rect 3294 11037 3297 11463
rect 2803 11031 3297 11037
rect 3353 11463 3847 11469
rect 3353 11037 3356 11463
rect 3373 11415 3827 11463
rect 3373 11085 3435 11415
rect 3765 11085 3827 11415
rect 3373 11037 3827 11085
rect 3844 11037 3847 11463
rect 3353 11031 3847 11037
rect 3903 11463 4397 11469
rect 3903 11037 3906 11463
rect 3923 11415 4377 11463
rect 3923 11085 3985 11415
rect 4315 11085 4377 11415
rect 3923 11037 4377 11085
rect 4394 11037 4397 11463
rect 3903 11031 4397 11037
rect 4453 11463 4947 11469
rect 4453 11037 4456 11463
rect 4473 11415 4927 11463
rect 4473 11085 4535 11415
rect 4865 11085 4927 11415
rect 4473 11037 4927 11085
rect 4944 11037 4947 11463
rect 4453 11031 4947 11037
rect 5003 11463 5497 11469
rect 5003 11037 5006 11463
rect 5023 11415 5477 11463
rect 5023 11085 5085 11415
rect 5415 11085 5477 11415
rect 5023 11037 5477 11085
rect 5494 11037 5497 11463
rect 5003 11031 5497 11037
rect 5553 11463 6047 11469
rect 5553 11037 5556 11463
rect 5573 11415 6027 11463
rect 5573 11085 5635 11415
rect 5965 11085 6027 11415
rect 5573 11037 6027 11085
rect 6044 11037 6047 11463
rect 5553 11031 6047 11037
rect 6103 11463 6597 11469
rect 6103 11037 6106 11463
rect 6123 11415 6577 11463
rect 6123 11085 6185 11415
rect 6515 11085 6577 11415
rect 6123 11037 6577 11085
rect 6594 11037 6597 11463
rect 6103 11031 6597 11037
rect 6653 11463 7147 11469
rect 6653 11037 6656 11463
rect 6673 11415 7127 11463
rect 6673 11085 6735 11415
rect 7065 11085 7127 11415
rect 6673 11037 7127 11085
rect 7144 11037 7147 11463
rect 6653 11031 7147 11037
rect 7203 11463 7697 11469
rect 7203 11037 7206 11463
rect 7223 11415 7677 11463
rect 7223 11085 7285 11415
rect 7615 11085 7677 11415
rect 7223 11037 7677 11085
rect 7694 11037 7697 11463
rect 7203 11031 7697 11037
rect 7753 11463 8247 11469
rect 7753 11037 7756 11463
rect 7773 11415 8227 11463
rect 7773 11085 7835 11415
rect 8165 11085 8227 11415
rect 7773 11037 8227 11085
rect 8244 11037 8247 11463
rect 7753 11031 8247 11037
rect 8303 11463 8797 11469
rect 8303 11037 8306 11463
rect 8323 11415 8777 11463
rect 8323 11085 8385 11415
rect 8715 11085 8777 11415
rect 8323 11037 8777 11085
rect 8794 11037 8797 11463
rect 8303 11031 8797 11037
rect 8853 11463 9347 11469
rect 8853 11037 8856 11463
rect 8873 11415 9327 11463
rect 8873 11085 8935 11415
rect 9265 11085 9327 11415
rect 8873 11037 9327 11085
rect 9344 11037 9347 11463
rect 8853 11031 9347 11037
rect 9403 11463 9897 11469
rect 9403 11037 9406 11463
rect 9423 11415 9877 11463
rect 9423 11085 9485 11415
rect 9815 11085 9877 11415
rect 9423 11037 9877 11085
rect 9894 11037 9897 11463
rect 9403 11031 9897 11037
rect 9953 11463 10447 11469
rect 9953 11037 9956 11463
rect 9973 11415 10427 11463
rect 9973 11085 10035 11415
rect 10365 11085 10427 11415
rect 9973 11037 10427 11085
rect 10444 11037 10447 11463
rect 9953 11031 10447 11037
rect 10503 11463 10997 11469
rect 10503 11037 10506 11463
rect 10523 11415 10977 11463
rect 10523 11085 10585 11415
rect 10915 11085 10977 11415
rect 10523 11037 10977 11085
rect 10994 11037 10997 11463
rect 10503 11031 10997 11037
rect 11053 11463 11547 11469
rect 11053 11037 11056 11463
rect 11073 11415 11527 11463
rect 11073 11085 11135 11415
rect 11465 11085 11527 11415
rect 11073 11037 11527 11085
rect 11544 11037 11547 11463
rect 11053 11031 11547 11037
rect 11603 11463 12097 11469
rect 11603 11037 11606 11463
rect 11623 11415 12077 11463
rect 11623 11085 11685 11415
rect 12015 11085 12077 11415
rect 11623 11037 12077 11085
rect 12094 11037 12097 11463
rect 11603 11031 12097 11037
rect 12153 11463 12647 11469
rect 12153 11037 12156 11463
rect 12173 11415 12627 11463
rect 12173 11085 12235 11415
rect 12565 11085 12627 11415
rect 12173 11037 12627 11085
rect 12644 11037 12647 11463
rect 12153 11031 12647 11037
rect 12703 11463 13197 11469
rect 12703 11037 12706 11463
rect 12723 11415 13177 11463
rect 12723 11085 12785 11415
rect 13115 11085 13177 11415
rect 12723 11037 13177 11085
rect 13194 11037 13197 11463
rect 12703 11031 13197 11037
rect 13253 11463 13724 11469
rect 13253 11037 13256 11463
rect 13273 11415 13724 11463
rect 13273 11085 13335 11415
rect 13665 11085 13724 11415
rect 13273 11037 13724 11085
rect 13253 11031 13724 11037
rect -474 11026 -26 11031
rect 76 11026 524 11031
rect 626 11026 1074 11031
rect 1176 11026 1624 11031
rect 1726 11026 2174 11031
rect 2276 11026 2724 11031
rect 2826 11026 3274 11031
rect 3376 11026 3824 11031
rect 3926 11026 4374 11031
rect 4476 11026 4924 11031
rect 5026 11026 5474 11031
rect 5576 11026 6024 11031
rect 6126 11026 6574 11031
rect 6676 11026 7124 11031
rect 7226 11026 7674 11031
rect 7776 11026 8224 11031
rect 8326 11026 8774 11031
rect 8876 11026 9324 11031
rect 9426 11026 9874 11031
rect 9976 11026 10424 11031
rect 10526 11026 10974 11031
rect 11076 11026 11524 11031
rect 11626 11026 12074 11031
rect 12176 11026 12624 11031
rect 12726 11026 13174 11031
rect 13276 11026 13724 11031
rect -1025 11000 -725 11019
rect -469 11023 -31 11026
rect -469 11006 -463 11023
rect -37 11006 -31 11023
rect -469 11003 -31 11006
rect 81 11023 519 11026
rect 81 11006 87 11023
rect 513 11006 519 11023
rect 81 11003 519 11006
rect 631 11023 1069 11026
rect 631 11006 637 11023
rect 1063 11006 1069 11023
rect 631 11003 1069 11006
rect 1181 11023 1619 11026
rect 1181 11006 1187 11023
rect 1613 11006 1619 11023
rect 1181 11003 1619 11006
rect 1731 11023 2169 11026
rect 1731 11006 1737 11023
rect 2163 11006 2169 11023
rect 1731 11003 2169 11006
rect 2281 11023 2719 11026
rect 2281 11006 2287 11023
rect 2713 11006 2719 11023
rect 2281 11003 2719 11006
rect 2831 11023 3269 11026
rect 2831 11006 2837 11023
rect 3263 11006 3269 11023
rect 2831 11003 3269 11006
rect 3381 11023 3819 11026
rect 3381 11006 3387 11023
rect 3813 11006 3819 11023
rect 3381 11003 3819 11006
rect 3931 11023 4369 11026
rect 3931 11006 3937 11023
rect 4363 11006 4369 11023
rect 3931 11003 4369 11006
rect 4481 11023 4919 11026
rect 4481 11006 4487 11023
rect 4913 11006 4919 11023
rect 4481 11003 4919 11006
rect 5031 11023 5469 11026
rect 5031 11006 5037 11023
rect 5463 11006 5469 11023
rect 5031 11003 5469 11006
rect 5581 11023 6019 11026
rect 5581 11006 5587 11023
rect 6013 11006 6019 11023
rect 5581 11003 6019 11006
rect 6131 11023 6569 11026
rect 6131 11006 6137 11023
rect 6563 11006 6569 11023
rect 6131 11003 6569 11006
rect 6681 11023 7119 11026
rect 6681 11006 6687 11023
rect 7113 11006 7119 11023
rect 6681 11003 7119 11006
rect 7231 11023 7669 11026
rect 7231 11006 7237 11023
rect 7663 11006 7669 11023
rect 7231 11003 7669 11006
rect 7781 11023 8219 11026
rect 7781 11006 7787 11023
rect 8213 11006 8219 11023
rect 7781 11003 8219 11006
rect 8331 11023 8769 11026
rect 8331 11006 8337 11023
rect 8763 11006 8769 11023
rect 8331 11003 8769 11006
rect 8881 11023 9319 11026
rect 8881 11006 8887 11023
rect 9313 11006 9319 11023
rect 8881 11003 9319 11006
rect 9431 11023 9869 11026
rect 9431 11006 9437 11023
rect 9863 11006 9869 11023
rect 9431 11003 9869 11006
rect 9981 11023 10419 11026
rect 9981 11006 9987 11023
rect 10413 11006 10419 11023
rect 9981 11003 10419 11006
rect 10531 11023 10969 11026
rect 10531 11006 10537 11023
rect 10963 11006 10969 11023
rect 10531 11003 10969 11006
rect 11081 11023 11519 11026
rect 11081 11006 11087 11023
rect 11513 11006 11519 11023
rect 11081 11003 11519 11006
rect 11631 11023 12069 11026
rect 11631 11006 11637 11023
rect 12063 11006 12069 11023
rect 11631 11003 12069 11006
rect 12181 11023 12619 11026
rect 12181 11006 12187 11023
rect 12613 11006 12619 11023
rect 12181 11003 12619 11006
rect 12731 11023 13169 11026
rect 12731 11006 12737 11023
rect 13163 11006 13169 11023
rect 12731 11003 13169 11006
rect 13281 11023 13719 11026
rect 13281 11006 13287 11023
rect 13713 11006 13719 11023
rect 13281 11003 13719 11006
rect 13975 11019 13987 11550
rect 14263 11019 14275 11550
rect 13975 11000 14275 11019
rect -1025 10469 -1013 11000
rect -737 10469 -725 11000
rect -550 10992 -500 11000
rect -550 10958 -542 10992
rect -508 10958 -500 10992
rect -550 10950 -500 10958
rect 0 10992 50 11000
rect 0 10958 8 10992
rect 42 10958 50 10992
rect 0 10950 50 10958
rect 550 10992 600 11000
rect 550 10958 558 10992
rect 592 10958 600 10992
rect 550 10950 600 10958
rect 1100 10992 1150 11000
rect 1100 10958 1108 10992
rect 1142 10958 1150 10992
rect 1100 10950 1150 10958
rect 1650 10992 1700 11000
rect 1650 10958 1658 10992
rect 1692 10958 1700 10992
rect 1650 10950 1700 10958
rect 2200 10992 2250 11000
rect 2200 10958 2208 10992
rect 2242 10958 2250 10992
rect 2200 10950 2250 10958
rect 2750 10992 2800 11000
rect 2750 10958 2758 10992
rect 2792 10958 2800 10992
rect 2750 10950 2800 10958
rect 3300 10992 3350 11000
rect 3300 10958 3308 10992
rect 3342 10958 3350 10992
rect 3300 10950 3350 10958
rect 3850 10992 3900 11000
rect 3850 10958 3858 10992
rect 3892 10958 3900 10992
rect 3850 10950 3900 10958
rect 4400 10992 4450 11000
rect 4400 10958 4408 10992
rect 4442 10958 4450 10992
rect 4400 10950 4450 10958
rect 4950 10992 5000 11000
rect 4950 10958 4958 10992
rect 4992 10958 5000 10992
rect 4950 10950 5000 10958
rect 5500 10992 5550 11000
rect 5500 10958 5508 10992
rect 5542 10958 5550 10992
rect 5500 10950 5550 10958
rect 6050 10992 6100 11000
rect 6050 10958 6058 10992
rect 6092 10958 6100 10992
rect 6050 10950 6100 10958
rect 6600 10992 6650 11000
rect 6600 10958 6608 10992
rect 6642 10958 6650 10992
rect 6600 10950 6650 10958
rect 7150 10992 7200 11000
rect 7150 10958 7158 10992
rect 7192 10958 7200 10992
rect 7150 10950 7200 10958
rect 7700 10992 7750 11000
rect 7700 10958 7708 10992
rect 7742 10958 7750 10992
rect 7700 10950 7750 10958
rect 8250 10992 8300 11000
rect 8250 10958 8258 10992
rect 8292 10958 8300 10992
rect 8250 10950 8300 10958
rect 8800 10992 8850 11000
rect 8800 10958 8808 10992
rect 8842 10958 8850 10992
rect 8800 10950 8850 10958
rect 9350 10992 9400 11000
rect 9350 10958 9358 10992
rect 9392 10958 9400 10992
rect 9350 10950 9400 10958
rect 9900 10992 9950 11000
rect 9900 10958 9908 10992
rect 9942 10958 9950 10992
rect 9900 10950 9950 10958
rect 10450 10992 10500 11000
rect 10450 10958 10458 10992
rect 10492 10958 10500 10992
rect 10450 10950 10500 10958
rect 11000 10992 11050 11000
rect 11000 10958 11008 10992
rect 11042 10958 11050 10992
rect 11000 10950 11050 10958
rect 11550 10992 11600 11000
rect 11550 10958 11558 10992
rect 11592 10958 11600 10992
rect 11550 10950 11600 10958
rect 12100 10992 12150 11000
rect 12100 10958 12108 10992
rect 12142 10958 12150 10992
rect 12100 10950 12150 10958
rect 12650 10992 12700 11000
rect 12650 10958 12658 10992
rect 12692 10958 12700 10992
rect 12650 10950 12700 10958
rect 13200 10992 13250 11000
rect 13200 10958 13208 10992
rect 13242 10958 13250 10992
rect 13200 10950 13250 10958
rect 13750 10992 13800 11000
rect 13750 10958 13758 10992
rect 13792 10958 13800 10992
rect 13750 10950 13800 10958
rect -469 10944 -31 10947
rect -469 10927 -463 10944
rect -37 10927 -31 10944
rect -469 10924 -31 10927
rect 81 10944 519 10947
rect 81 10927 87 10944
rect 513 10927 519 10944
rect 81 10924 519 10927
rect 631 10944 1069 10947
rect 631 10927 637 10944
rect 1063 10927 1069 10944
rect 631 10924 1069 10927
rect 1181 10944 1619 10947
rect 1181 10927 1187 10944
rect 1613 10927 1619 10944
rect 1181 10924 1619 10927
rect 1731 10944 2169 10947
rect 1731 10927 1737 10944
rect 2163 10927 2169 10944
rect 1731 10924 2169 10927
rect 2281 10944 2719 10947
rect 2281 10927 2287 10944
rect 2713 10927 2719 10944
rect 2281 10924 2719 10927
rect 2831 10944 3269 10947
rect 2831 10927 2837 10944
rect 3263 10927 3269 10944
rect 2831 10924 3269 10927
rect 3381 10944 3819 10947
rect 3381 10927 3387 10944
rect 3813 10927 3819 10944
rect 3381 10924 3819 10927
rect 3931 10944 4369 10947
rect 3931 10927 3937 10944
rect 4363 10927 4369 10944
rect 3931 10924 4369 10927
rect 4481 10944 4919 10947
rect 4481 10927 4487 10944
rect 4913 10927 4919 10944
rect 4481 10924 4919 10927
rect 5031 10944 5469 10947
rect 5031 10927 5037 10944
rect 5463 10927 5469 10944
rect 5031 10924 5469 10927
rect 5581 10944 6019 10947
rect 5581 10927 5587 10944
rect 6013 10927 6019 10944
rect 5581 10924 6019 10927
rect 6131 10944 6569 10947
rect 6131 10927 6137 10944
rect 6563 10927 6569 10944
rect 6131 10924 6569 10927
rect 6681 10944 7119 10947
rect 6681 10927 6687 10944
rect 7113 10927 7119 10944
rect 6681 10924 7119 10927
rect 7231 10944 7669 10947
rect 7231 10927 7237 10944
rect 7663 10927 7669 10944
rect 7231 10924 7669 10927
rect 7781 10944 8219 10947
rect 7781 10927 7787 10944
rect 8213 10927 8219 10944
rect 7781 10924 8219 10927
rect 8331 10944 8769 10947
rect 8331 10927 8337 10944
rect 8763 10927 8769 10944
rect 8331 10924 8769 10927
rect 8881 10944 9319 10947
rect 8881 10927 8887 10944
rect 9313 10927 9319 10944
rect 8881 10924 9319 10927
rect 9431 10944 9869 10947
rect 9431 10927 9437 10944
rect 9863 10927 9869 10944
rect 9431 10924 9869 10927
rect 9981 10944 10419 10947
rect 9981 10927 9987 10944
rect 10413 10927 10419 10944
rect 9981 10924 10419 10927
rect 10531 10944 10969 10947
rect 10531 10927 10537 10944
rect 10963 10927 10969 10944
rect 10531 10924 10969 10927
rect 11081 10944 11519 10947
rect 11081 10927 11087 10944
rect 11513 10927 11519 10944
rect 11081 10924 11519 10927
rect 11631 10944 12069 10947
rect 11631 10927 11637 10944
rect 12063 10927 12069 10944
rect 11631 10924 12069 10927
rect 12181 10944 12619 10947
rect 12181 10927 12187 10944
rect 12613 10927 12619 10944
rect 12181 10924 12619 10927
rect 12731 10944 13169 10947
rect 12731 10927 12737 10944
rect 13163 10927 13169 10944
rect 12731 10924 13169 10927
rect 13281 10944 13719 10947
rect 13281 10927 13287 10944
rect 13713 10927 13719 10944
rect 13281 10924 13719 10927
rect -474 10919 -26 10924
rect 76 10919 524 10924
rect 626 10919 1074 10924
rect 1176 10919 1624 10924
rect 1726 10919 2174 10924
rect 2276 10919 2724 10924
rect 2826 10919 3274 10924
rect 3376 10919 3824 10924
rect 3926 10919 4374 10924
rect 4476 10919 4924 10924
rect 5026 10919 5474 10924
rect 5576 10919 6024 10924
rect 6126 10919 6574 10924
rect 6676 10919 7124 10924
rect 7226 10919 7674 10924
rect 7776 10919 8224 10924
rect 8326 10919 8774 10924
rect 8876 10919 9324 10924
rect 9426 10919 9874 10924
rect 9976 10919 10424 10924
rect 10526 10919 10974 10924
rect 11076 10919 11524 10924
rect 11626 10919 12074 10924
rect 12176 10919 12624 10924
rect 12726 10919 13174 10924
rect 13276 10919 13724 10924
rect -474 10913 -3 10919
rect -474 10865 -23 10913
rect -474 10535 -415 10865
rect -85 10535 -23 10865
rect -474 10487 -23 10535
rect -6 10487 -3 10913
rect -474 10481 -3 10487
rect 53 10913 547 10919
rect 53 10487 56 10913
rect 73 10865 527 10913
rect 73 10535 135 10865
rect 465 10535 527 10865
rect 73 10487 527 10535
rect 544 10487 547 10913
rect 53 10481 547 10487
rect 603 10913 1097 10919
rect 603 10487 606 10913
rect 623 10865 1077 10913
rect 623 10535 685 10865
rect 1015 10535 1077 10865
rect 623 10487 1077 10535
rect 1094 10487 1097 10913
rect 603 10481 1097 10487
rect 1153 10913 1647 10919
rect 1153 10487 1156 10913
rect 1173 10865 1627 10913
rect 1173 10535 1235 10865
rect 1565 10535 1627 10865
rect 1173 10487 1627 10535
rect 1644 10487 1647 10913
rect 1153 10481 1647 10487
rect 1703 10913 2197 10919
rect 1703 10487 1706 10913
rect 1723 10865 2177 10913
rect 1723 10535 1785 10865
rect 2115 10535 2177 10865
rect 1723 10487 2177 10535
rect 2194 10487 2197 10913
rect 1703 10481 2197 10487
rect 2253 10913 2747 10919
rect 2253 10487 2256 10913
rect 2273 10865 2727 10913
rect 2273 10535 2335 10865
rect 2665 10535 2727 10865
rect 2273 10487 2727 10535
rect 2744 10487 2747 10913
rect 2253 10481 2747 10487
rect 2803 10913 3297 10919
rect 2803 10487 2806 10913
rect 2823 10865 3277 10913
rect 2823 10535 2885 10865
rect 3215 10535 3277 10865
rect 2823 10487 3277 10535
rect 3294 10487 3297 10913
rect 2803 10481 3297 10487
rect 3353 10913 3847 10919
rect 3353 10487 3356 10913
rect 3373 10865 3827 10913
rect 3373 10535 3435 10865
rect 3765 10535 3827 10865
rect 3373 10487 3827 10535
rect 3844 10487 3847 10913
rect 3353 10481 3847 10487
rect 3903 10913 4397 10919
rect 3903 10487 3906 10913
rect 3923 10865 4377 10913
rect 3923 10535 3985 10865
rect 4315 10535 4377 10865
rect 3923 10487 4377 10535
rect 4394 10487 4397 10913
rect 3903 10481 4397 10487
rect 4453 10913 4947 10919
rect 4453 10487 4456 10913
rect 4473 10865 4927 10913
rect 4473 10535 4535 10865
rect 4865 10535 4927 10865
rect 4473 10487 4927 10535
rect 4944 10487 4947 10913
rect 4453 10481 4947 10487
rect 5003 10913 5497 10919
rect 5003 10487 5006 10913
rect 5023 10865 5477 10913
rect 5023 10535 5085 10865
rect 5415 10535 5477 10865
rect 5023 10487 5477 10535
rect 5494 10487 5497 10913
rect 5003 10481 5497 10487
rect 5553 10913 6047 10919
rect 5553 10487 5556 10913
rect 5573 10865 6027 10913
rect 5573 10535 5635 10865
rect 5965 10535 6027 10865
rect 5573 10487 6027 10535
rect 6044 10487 6047 10913
rect 5553 10481 6047 10487
rect 6103 10913 6597 10919
rect 6103 10487 6106 10913
rect 6123 10865 6577 10913
rect 6123 10535 6185 10865
rect 6515 10535 6577 10865
rect 6123 10487 6577 10535
rect 6594 10487 6597 10913
rect 6103 10481 6597 10487
rect 6653 10913 7147 10919
rect 6653 10487 6656 10913
rect 6673 10865 7127 10913
rect 6673 10535 6735 10865
rect 7065 10535 7127 10865
rect 6673 10487 7127 10535
rect 7144 10487 7147 10913
rect 6653 10481 7147 10487
rect 7203 10913 7697 10919
rect 7203 10487 7206 10913
rect 7223 10865 7677 10913
rect 7223 10535 7285 10865
rect 7615 10535 7677 10865
rect 7223 10487 7677 10535
rect 7694 10487 7697 10913
rect 7203 10481 7697 10487
rect 7753 10913 8247 10919
rect 7753 10487 7756 10913
rect 7773 10865 8227 10913
rect 7773 10535 7835 10865
rect 8165 10535 8227 10865
rect 7773 10487 8227 10535
rect 8244 10487 8247 10913
rect 7753 10481 8247 10487
rect 8303 10913 8797 10919
rect 8303 10487 8306 10913
rect 8323 10865 8777 10913
rect 8323 10535 8385 10865
rect 8715 10535 8777 10865
rect 8323 10487 8777 10535
rect 8794 10487 8797 10913
rect 8303 10481 8797 10487
rect 8853 10913 9347 10919
rect 8853 10487 8856 10913
rect 8873 10865 9327 10913
rect 8873 10535 8935 10865
rect 9265 10535 9327 10865
rect 8873 10487 9327 10535
rect 9344 10487 9347 10913
rect 8853 10481 9347 10487
rect 9403 10913 9897 10919
rect 9403 10487 9406 10913
rect 9423 10865 9877 10913
rect 9423 10535 9485 10865
rect 9815 10535 9877 10865
rect 9423 10487 9877 10535
rect 9894 10487 9897 10913
rect 9403 10481 9897 10487
rect 9953 10913 10447 10919
rect 9953 10487 9956 10913
rect 9973 10865 10427 10913
rect 9973 10535 10035 10865
rect 10365 10535 10427 10865
rect 9973 10487 10427 10535
rect 10444 10487 10447 10913
rect 9953 10481 10447 10487
rect 10503 10913 10997 10919
rect 10503 10487 10506 10913
rect 10523 10865 10977 10913
rect 10523 10535 10585 10865
rect 10915 10535 10977 10865
rect 10523 10487 10977 10535
rect 10994 10487 10997 10913
rect 10503 10481 10997 10487
rect 11053 10913 11547 10919
rect 11053 10487 11056 10913
rect 11073 10865 11527 10913
rect 11073 10535 11135 10865
rect 11465 10535 11527 10865
rect 11073 10487 11527 10535
rect 11544 10487 11547 10913
rect 11053 10481 11547 10487
rect 11603 10913 12097 10919
rect 11603 10487 11606 10913
rect 11623 10865 12077 10913
rect 11623 10535 11685 10865
rect 12015 10535 12077 10865
rect 11623 10487 12077 10535
rect 12094 10487 12097 10913
rect 11603 10481 12097 10487
rect 12153 10913 12647 10919
rect 12153 10487 12156 10913
rect 12173 10865 12627 10913
rect 12173 10535 12235 10865
rect 12565 10535 12627 10865
rect 12173 10487 12627 10535
rect 12644 10487 12647 10913
rect 12153 10481 12647 10487
rect 12703 10913 13197 10919
rect 12703 10487 12706 10913
rect 12723 10865 13177 10913
rect 12723 10535 12785 10865
rect 13115 10535 13177 10865
rect 12723 10487 13177 10535
rect 13194 10487 13197 10913
rect 12703 10481 13197 10487
rect 13253 10913 13724 10919
rect 13253 10487 13256 10913
rect 13273 10865 13724 10913
rect 13273 10535 13335 10865
rect 13665 10535 13724 10865
rect 13273 10487 13724 10535
rect 13253 10481 13724 10487
rect -474 10476 -26 10481
rect 76 10476 524 10481
rect 626 10476 1074 10481
rect 1176 10476 1624 10481
rect 1726 10476 2174 10481
rect 2276 10476 2724 10481
rect 2826 10476 3274 10481
rect 3376 10476 3824 10481
rect 3926 10476 4374 10481
rect 4476 10476 4924 10481
rect 5026 10476 5474 10481
rect 5576 10476 6024 10481
rect 6126 10476 6574 10481
rect 6676 10476 7124 10481
rect 7226 10476 7674 10481
rect 7776 10476 8224 10481
rect 8326 10476 8774 10481
rect 8876 10476 9324 10481
rect 9426 10476 9874 10481
rect 9976 10476 10424 10481
rect 10526 10476 10974 10481
rect 11076 10476 11524 10481
rect 11626 10476 12074 10481
rect 12176 10476 12624 10481
rect 12726 10476 13174 10481
rect 13276 10476 13724 10481
rect -1025 10450 -725 10469
rect -469 10473 -31 10476
rect -469 10456 -463 10473
rect -37 10456 -31 10473
rect -469 10453 -31 10456
rect 81 10473 519 10476
rect 81 10456 87 10473
rect 513 10456 519 10473
rect 81 10453 519 10456
rect 631 10473 1069 10476
rect 631 10456 637 10473
rect 1063 10456 1069 10473
rect 631 10453 1069 10456
rect 1181 10473 1619 10476
rect 1181 10456 1187 10473
rect 1613 10456 1619 10473
rect 1181 10453 1619 10456
rect 1731 10473 2169 10476
rect 1731 10456 1737 10473
rect 2163 10456 2169 10473
rect 1731 10453 2169 10456
rect 2281 10473 2719 10476
rect 2281 10456 2287 10473
rect 2713 10456 2719 10473
rect 2281 10453 2719 10456
rect 2831 10473 3269 10476
rect 2831 10456 2837 10473
rect 3263 10456 3269 10473
rect 2831 10453 3269 10456
rect 3381 10473 3819 10476
rect 3381 10456 3387 10473
rect 3813 10456 3819 10473
rect 3381 10453 3819 10456
rect 3931 10473 4369 10476
rect 3931 10456 3937 10473
rect 4363 10456 4369 10473
rect 3931 10453 4369 10456
rect 4481 10473 4919 10476
rect 4481 10456 4487 10473
rect 4913 10456 4919 10473
rect 4481 10453 4919 10456
rect 5031 10473 5469 10476
rect 5031 10456 5037 10473
rect 5463 10456 5469 10473
rect 5031 10453 5469 10456
rect 5581 10473 6019 10476
rect 5581 10456 5587 10473
rect 6013 10456 6019 10473
rect 5581 10453 6019 10456
rect 6131 10473 6569 10476
rect 6131 10456 6137 10473
rect 6563 10456 6569 10473
rect 6131 10453 6569 10456
rect 6681 10473 7119 10476
rect 6681 10456 6687 10473
rect 7113 10456 7119 10473
rect 6681 10453 7119 10456
rect 7231 10473 7669 10476
rect 7231 10456 7237 10473
rect 7663 10456 7669 10473
rect 7231 10453 7669 10456
rect 7781 10473 8219 10476
rect 7781 10456 7787 10473
rect 8213 10456 8219 10473
rect 7781 10453 8219 10456
rect 8331 10473 8769 10476
rect 8331 10456 8337 10473
rect 8763 10456 8769 10473
rect 8331 10453 8769 10456
rect 8881 10473 9319 10476
rect 8881 10456 8887 10473
rect 9313 10456 9319 10473
rect 8881 10453 9319 10456
rect 9431 10473 9869 10476
rect 9431 10456 9437 10473
rect 9863 10456 9869 10473
rect 9431 10453 9869 10456
rect 9981 10473 10419 10476
rect 9981 10456 9987 10473
rect 10413 10456 10419 10473
rect 9981 10453 10419 10456
rect 10531 10473 10969 10476
rect 10531 10456 10537 10473
rect 10963 10456 10969 10473
rect 10531 10453 10969 10456
rect 11081 10473 11519 10476
rect 11081 10456 11087 10473
rect 11513 10456 11519 10473
rect 11081 10453 11519 10456
rect 11631 10473 12069 10476
rect 11631 10456 11637 10473
rect 12063 10456 12069 10473
rect 11631 10453 12069 10456
rect 12181 10473 12619 10476
rect 12181 10456 12187 10473
rect 12613 10456 12619 10473
rect 12181 10453 12619 10456
rect 12731 10473 13169 10476
rect 12731 10456 12737 10473
rect 13163 10456 13169 10473
rect 12731 10453 13169 10456
rect 13281 10473 13719 10476
rect 13281 10456 13287 10473
rect 13713 10456 13719 10473
rect 13281 10453 13719 10456
rect 13975 10469 13987 11000
rect 14263 10469 14275 11000
rect 13975 10450 14275 10469
rect -1025 9919 -1013 10450
rect -737 9919 -725 10450
rect -550 10442 -500 10450
rect -550 10408 -542 10442
rect -508 10408 -500 10442
rect -550 10400 -500 10408
rect 0 10442 50 10450
rect 0 10408 8 10442
rect 42 10408 50 10442
rect 0 10400 50 10408
rect 550 10442 600 10450
rect 550 10408 558 10442
rect 592 10408 600 10442
rect 550 10400 600 10408
rect 1100 10442 1150 10450
rect 1100 10408 1108 10442
rect 1142 10408 1150 10442
rect 1100 10400 1150 10408
rect 1650 10442 1700 10450
rect 1650 10408 1658 10442
rect 1692 10408 1700 10442
rect 1650 10400 1700 10408
rect 2200 10442 2250 10450
rect 2200 10408 2208 10442
rect 2242 10408 2250 10442
rect 2200 10400 2250 10408
rect 2750 10442 2800 10450
rect 2750 10408 2758 10442
rect 2792 10408 2800 10442
rect 2750 10400 2800 10408
rect 3300 10442 3350 10450
rect 3300 10408 3308 10442
rect 3342 10408 3350 10442
rect 3300 10400 3350 10408
rect 3850 10442 3900 10450
rect 3850 10408 3858 10442
rect 3892 10408 3900 10442
rect 3850 10400 3900 10408
rect 4400 10442 4450 10450
rect 4400 10408 4408 10442
rect 4442 10408 4450 10442
rect 4400 10400 4450 10408
rect 4950 10442 5000 10450
rect 4950 10408 4958 10442
rect 4992 10408 5000 10442
rect 4950 10400 5000 10408
rect 5500 10442 5550 10450
rect 5500 10408 5508 10442
rect 5542 10408 5550 10442
rect 5500 10400 5550 10408
rect 6050 10442 6100 10450
rect 6050 10408 6058 10442
rect 6092 10408 6100 10442
rect 6050 10400 6100 10408
rect 6600 10442 6650 10450
rect 6600 10408 6608 10442
rect 6642 10408 6650 10442
rect 6600 10400 6650 10408
rect 7150 10442 7200 10450
rect 7150 10408 7158 10442
rect 7192 10408 7200 10442
rect 7150 10400 7200 10408
rect 7700 10442 7750 10450
rect 7700 10408 7708 10442
rect 7742 10408 7750 10442
rect 7700 10400 7750 10408
rect 8250 10442 8300 10450
rect 8250 10408 8258 10442
rect 8292 10408 8300 10442
rect 8250 10400 8300 10408
rect 8800 10442 8850 10450
rect 8800 10408 8808 10442
rect 8842 10408 8850 10442
rect 8800 10400 8850 10408
rect 9350 10442 9400 10450
rect 9350 10408 9358 10442
rect 9392 10408 9400 10442
rect 9350 10400 9400 10408
rect 9900 10442 9950 10450
rect 9900 10408 9908 10442
rect 9942 10408 9950 10442
rect 9900 10400 9950 10408
rect 10450 10442 10500 10450
rect 10450 10408 10458 10442
rect 10492 10408 10500 10442
rect 10450 10400 10500 10408
rect 11000 10442 11050 10450
rect 11000 10408 11008 10442
rect 11042 10408 11050 10442
rect 11000 10400 11050 10408
rect 11550 10442 11600 10450
rect 11550 10408 11558 10442
rect 11592 10408 11600 10442
rect 11550 10400 11600 10408
rect 12100 10442 12150 10450
rect 12100 10408 12108 10442
rect 12142 10408 12150 10442
rect 12100 10400 12150 10408
rect 12650 10442 12700 10450
rect 12650 10408 12658 10442
rect 12692 10408 12700 10442
rect 12650 10400 12700 10408
rect 13200 10442 13250 10450
rect 13200 10408 13208 10442
rect 13242 10408 13250 10442
rect 13200 10400 13250 10408
rect 13750 10442 13800 10450
rect 13750 10408 13758 10442
rect 13792 10408 13800 10442
rect 13750 10400 13800 10408
rect -469 10394 -31 10397
rect -469 10377 -463 10394
rect -37 10377 -31 10394
rect -469 10374 -31 10377
rect 81 10394 519 10397
rect 81 10377 87 10394
rect 513 10377 519 10394
rect 81 10374 519 10377
rect 631 10394 1069 10397
rect 631 10377 637 10394
rect 1063 10377 1069 10394
rect 631 10374 1069 10377
rect 1181 10394 1619 10397
rect 1181 10377 1187 10394
rect 1613 10377 1619 10394
rect 1181 10374 1619 10377
rect 1731 10394 2169 10397
rect 1731 10377 1737 10394
rect 2163 10377 2169 10394
rect 1731 10374 2169 10377
rect 2281 10394 2719 10397
rect 2281 10377 2287 10394
rect 2713 10377 2719 10394
rect 2281 10374 2719 10377
rect 2831 10394 3269 10397
rect 2831 10377 2837 10394
rect 3263 10377 3269 10394
rect 2831 10374 3269 10377
rect 3381 10394 3819 10397
rect 3381 10377 3387 10394
rect 3813 10377 3819 10394
rect 3381 10374 3819 10377
rect 3931 10394 4369 10397
rect 3931 10377 3937 10394
rect 4363 10377 4369 10394
rect 3931 10374 4369 10377
rect 4481 10394 4919 10397
rect 4481 10377 4487 10394
rect 4913 10377 4919 10394
rect 4481 10374 4919 10377
rect 5031 10394 5469 10397
rect 5031 10377 5037 10394
rect 5463 10377 5469 10394
rect 5031 10374 5469 10377
rect 5581 10394 6019 10397
rect 5581 10377 5587 10394
rect 6013 10377 6019 10394
rect 5581 10374 6019 10377
rect 6131 10394 6569 10397
rect 6131 10377 6137 10394
rect 6563 10377 6569 10394
rect 6131 10374 6569 10377
rect 6681 10394 7119 10397
rect 6681 10377 6687 10394
rect 7113 10377 7119 10394
rect 6681 10374 7119 10377
rect 7231 10394 7669 10397
rect 7231 10377 7237 10394
rect 7663 10377 7669 10394
rect 7231 10374 7669 10377
rect 7781 10394 8219 10397
rect 7781 10377 7787 10394
rect 8213 10377 8219 10394
rect 7781 10374 8219 10377
rect 8331 10394 8769 10397
rect 8331 10377 8337 10394
rect 8763 10377 8769 10394
rect 8331 10374 8769 10377
rect 8881 10394 9319 10397
rect 8881 10377 8887 10394
rect 9313 10377 9319 10394
rect 8881 10374 9319 10377
rect 9431 10394 9869 10397
rect 9431 10377 9437 10394
rect 9863 10377 9869 10394
rect 9431 10374 9869 10377
rect 9981 10394 10419 10397
rect 9981 10377 9987 10394
rect 10413 10377 10419 10394
rect 9981 10374 10419 10377
rect 10531 10394 10969 10397
rect 10531 10377 10537 10394
rect 10963 10377 10969 10394
rect 10531 10374 10969 10377
rect 11081 10394 11519 10397
rect 11081 10377 11087 10394
rect 11513 10377 11519 10394
rect 11081 10374 11519 10377
rect 11631 10394 12069 10397
rect 11631 10377 11637 10394
rect 12063 10377 12069 10394
rect 11631 10374 12069 10377
rect 12181 10394 12619 10397
rect 12181 10377 12187 10394
rect 12613 10377 12619 10394
rect 12181 10374 12619 10377
rect 12731 10394 13169 10397
rect 12731 10377 12737 10394
rect 13163 10377 13169 10394
rect 12731 10374 13169 10377
rect 13281 10394 13719 10397
rect 13281 10377 13287 10394
rect 13713 10377 13719 10394
rect 13281 10374 13719 10377
rect -474 10369 -26 10374
rect 76 10369 524 10374
rect 626 10369 1074 10374
rect 1176 10369 1624 10374
rect 1726 10369 2174 10374
rect 2276 10369 2724 10374
rect 2826 10369 3274 10374
rect 3376 10369 3824 10374
rect 3926 10369 4374 10374
rect 4476 10369 4924 10374
rect 5026 10369 5474 10374
rect 5576 10369 6024 10374
rect 6126 10369 6574 10374
rect 6676 10369 7124 10374
rect 7226 10369 7674 10374
rect 7776 10369 8224 10374
rect 8326 10369 8774 10374
rect 8876 10369 9324 10374
rect 9426 10369 9874 10374
rect 9976 10369 10424 10374
rect 10526 10369 10974 10374
rect 11076 10369 11524 10374
rect 11626 10369 12074 10374
rect 12176 10369 12624 10374
rect 12726 10369 13174 10374
rect 13276 10369 13724 10374
rect -474 10363 -3 10369
rect -474 10315 -23 10363
rect -474 9985 -415 10315
rect -85 9985 -23 10315
rect -474 9937 -23 9985
rect -6 9937 -3 10363
rect -474 9931 -3 9937
rect 53 10363 547 10369
rect 53 9937 56 10363
rect 73 10315 527 10363
rect 73 9985 135 10315
rect 465 9985 527 10315
rect 73 9937 527 9985
rect 544 9937 547 10363
rect 53 9931 547 9937
rect 603 10363 1097 10369
rect 603 9937 606 10363
rect 623 10315 1077 10363
rect 623 9985 685 10315
rect 1015 9985 1077 10315
rect 623 9937 1077 9985
rect 1094 9937 1097 10363
rect 603 9931 1097 9937
rect 1153 10363 1647 10369
rect 1153 9937 1156 10363
rect 1173 10315 1627 10363
rect 1173 9985 1235 10315
rect 1565 9985 1627 10315
rect 1173 9937 1627 9985
rect 1644 9937 1647 10363
rect 1153 9931 1647 9937
rect 1703 10363 2197 10369
rect 1703 9937 1706 10363
rect 1723 10315 2177 10363
rect 1723 9985 1785 10315
rect 2115 9985 2177 10315
rect 1723 9937 2177 9985
rect 2194 9937 2197 10363
rect 1703 9931 2197 9937
rect 2253 10363 2747 10369
rect 2253 9937 2256 10363
rect 2273 10315 2727 10363
rect 2273 9985 2335 10315
rect 2665 9985 2727 10315
rect 2273 9937 2727 9985
rect 2744 9937 2747 10363
rect 2253 9931 2747 9937
rect 2803 10363 3297 10369
rect 2803 9937 2806 10363
rect 2823 10315 3277 10363
rect 2823 9985 2885 10315
rect 3215 9985 3277 10315
rect 2823 9937 3277 9985
rect 3294 9937 3297 10363
rect 2803 9931 3297 9937
rect 3353 10363 3847 10369
rect 3353 9937 3356 10363
rect 3373 10315 3827 10363
rect 3373 9985 3435 10315
rect 3765 9985 3827 10315
rect 3373 9937 3827 9985
rect 3844 9937 3847 10363
rect 3353 9931 3847 9937
rect 3903 10363 4397 10369
rect 3903 9937 3906 10363
rect 3923 10315 4377 10363
rect 3923 9985 3985 10315
rect 4315 9985 4377 10315
rect 3923 9937 4377 9985
rect 4394 9937 4397 10363
rect 3903 9931 4397 9937
rect 4453 10363 4947 10369
rect 4453 9937 4456 10363
rect 4473 10315 4927 10363
rect 4473 9985 4535 10315
rect 4865 9985 4927 10315
rect 4473 9937 4927 9985
rect 4944 9937 4947 10363
rect 4453 9931 4947 9937
rect 5003 10363 5497 10369
rect 5003 9937 5006 10363
rect 5023 10315 5477 10363
rect 5023 9985 5085 10315
rect 5415 9985 5477 10315
rect 5023 9937 5477 9985
rect 5494 9937 5497 10363
rect 5003 9931 5497 9937
rect 5553 10363 6047 10369
rect 5553 9937 5556 10363
rect 5573 10315 6027 10363
rect 5573 9985 5635 10315
rect 5965 9985 6027 10315
rect 5573 9937 6027 9985
rect 6044 9937 6047 10363
rect 5553 9931 6047 9937
rect 6103 10363 6597 10369
rect 6103 9937 6106 10363
rect 6123 10315 6577 10363
rect 6123 9985 6185 10315
rect 6515 9985 6577 10315
rect 6123 9937 6577 9985
rect 6594 9937 6597 10363
rect 6103 9931 6597 9937
rect 6653 10363 7147 10369
rect 6653 9937 6656 10363
rect 6673 10315 7127 10363
rect 6673 9985 6735 10315
rect 7065 9985 7127 10315
rect 6673 9937 7127 9985
rect 7144 9937 7147 10363
rect 6653 9931 7147 9937
rect 7203 10363 7697 10369
rect 7203 9937 7206 10363
rect 7223 10315 7677 10363
rect 7223 9985 7285 10315
rect 7615 9985 7677 10315
rect 7223 9937 7677 9985
rect 7694 9937 7697 10363
rect 7203 9931 7697 9937
rect 7753 10363 8247 10369
rect 7753 9937 7756 10363
rect 7773 10315 8227 10363
rect 7773 9985 7835 10315
rect 8165 9985 8227 10315
rect 7773 9937 8227 9985
rect 8244 9937 8247 10363
rect 7753 9931 8247 9937
rect 8303 10363 8797 10369
rect 8303 9937 8306 10363
rect 8323 10315 8777 10363
rect 8323 9985 8385 10315
rect 8715 9985 8777 10315
rect 8323 9937 8777 9985
rect 8794 9937 8797 10363
rect 8303 9931 8797 9937
rect 8853 10363 9347 10369
rect 8853 9937 8856 10363
rect 8873 10315 9327 10363
rect 8873 9985 8935 10315
rect 9265 9985 9327 10315
rect 8873 9937 9327 9985
rect 9344 9937 9347 10363
rect 8853 9931 9347 9937
rect 9403 10363 9897 10369
rect 9403 9937 9406 10363
rect 9423 10315 9877 10363
rect 9423 9985 9485 10315
rect 9815 9985 9877 10315
rect 9423 9937 9877 9985
rect 9894 9937 9897 10363
rect 9403 9931 9897 9937
rect 9953 10363 10447 10369
rect 9953 9937 9956 10363
rect 9973 10315 10427 10363
rect 9973 9985 10035 10315
rect 10365 9985 10427 10315
rect 9973 9937 10427 9985
rect 10444 9937 10447 10363
rect 9953 9931 10447 9937
rect 10503 10363 10997 10369
rect 10503 9937 10506 10363
rect 10523 10315 10977 10363
rect 10523 9985 10585 10315
rect 10915 9985 10977 10315
rect 10523 9937 10977 9985
rect 10994 9937 10997 10363
rect 10503 9931 10997 9937
rect 11053 10363 11547 10369
rect 11053 9937 11056 10363
rect 11073 10315 11527 10363
rect 11073 9985 11135 10315
rect 11465 9985 11527 10315
rect 11073 9937 11527 9985
rect 11544 9937 11547 10363
rect 11053 9931 11547 9937
rect 11603 10363 12097 10369
rect 11603 9937 11606 10363
rect 11623 10315 12077 10363
rect 11623 9985 11685 10315
rect 12015 9985 12077 10315
rect 11623 9937 12077 9985
rect 12094 9937 12097 10363
rect 11603 9931 12097 9937
rect 12153 10363 12647 10369
rect 12153 9937 12156 10363
rect 12173 10315 12627 10363
rect 12173 9985 12235 10315
rect 12565 9985 12627 10315
rect 12173 9937 12627 9985
rect 12644 9937 12647 10363
rect 12153 9931 12647 9937
rect 12703 10363 13197 10369
rect 12703 9937 12706 10363
rect 12723 10315 13177 10363
rect 12723 9985 12785 10315
rect 13115 9985 13177 10315
rect 12723 9937 13177 9985
rect 13194 9937 13197 10363
rect 12703 9931 13197 9937
rect 13253 10363 13724 10369
rect 13253 9937 13256 10363
rect 13273 10315 13724 10363
rect 13273 9985 13335 10315
rect 13665 9985 13724 10315
rect 13273 9937 13724 9985
rect 13253 9931 13724 9937
rect -474 9926 -26 9931
rect 76 9926 524 9931
rect 626 9926 1074 9931
rect 1176 9926 1624 9931
rect 1726 9926 2174 9931
rect 2276 9926 2724 9931
rect 2826 9926 3274 9931
rect 3376 9926 3824 9931
rect 3926 9926 4374 9931
rect 4476 9926 4924 9931
rect 5026 9926 5474 9931
rect 5576 9926 6024 9931
rect 6126 9926 6574 9931
rect 6676 9926 7124 9931
rect 7226 9926 7674 9931
rect 7776 9926 8224 9931
rect 8326 9926 8774 9931
rect 8876 9926 9324 9931
rect 9426 9926 9874 9931
rect 9976 9926 10424 9931
rect 10526 9926 10974 9931
rect 11076 9926 11524 9931
rect 11626 9926 12074 9931
rect 12176 9926 12624 9931
rect 12726 9926 13174 9931
rect 13276 9926 13724 9931
rect -1025 9900 -725 9919
rect -469 9923 -31 9926
rect -469 9906 -463 9923
rect -37 9906 -31 9923
rect -469 9903 -31 9906
rect 81 9923 519 9926
rect 81 9906 87 9923
rect 513 9906 519 9923
rect 81 9903 519 9906
rect 631 9923 1069 9926
rect 631 9906 637 9923
rect 1063 9906 1069 9923
rect 631 9903 1069 9906
rect 1181 9923 1619 9926
rect 1181 9906 1187 9923
rect 1613 9906 1619 9923
rect 1181 9903 1619 9906
rect 1731 9923 2169 9926
rect 1731 9906 1737 9923
rect 2163 9906 2169 9923
rect 1731 9903 2169 9906
rect 2281 9923 2719 9926
rect 2281 9906 2287 9923
rect 2713 9906 2719 9923
rect 2281 9903 2719 9906
rect 2831 9923 3269 9926
rect 2831 9906 2837 9923
rect 3263 9906 3269 9923
rect 2831 9903 3269 9906
rect 3381 9923 3819 9926
rect 3381 9906 3387 9923
rect 3813 9906 3819 9923
rect 3381 9903 3819 9906
rect 3931 9923 4369 9926
rect 3931 9906 3937 9923
rect 4363 9906 4369 9923
rect 3931 9903 4369 9906
rect 4481 9923 4919 9926
rect 4481 9906 4487 9923
rect 4913 9906 4919 9923
rect 4481 9903 4919 9906
rect 5031 9923 5469 9926
rect 5031 9906 5037 9923
rect 5463 9906 5469 9923
rect 5031 9903 5469 9906
rect 5581 9923 6019 9926
rect 5581 9906 5587 9923
rect 6013 9906 6019 9923
rect 5581 9903 6019 9906
rect 6131 9923 6569 9926
rect 6131 9906 6137 9923
rect 6563 9906 6569 9923
rect 6131 9903 6569 9906
rect 6681 9923 7119 9926
rect 6681 9906 6687 9923
rect 7113 9906 7119 9923
rect 6681 9903 7119 9906
rect 7231 9923 7669 9926
rect 7231 9906 7237 9923
rect 7663 9906 7669 9923
rect 7231 9903 7669 9906
rect 7781 9923 8219 9926
rect 7781 9906 7787 9923
rect 8213 9906 8219 9923
rect 7781 9903 8219 9906
rect 8331 9923 8769 9926
rect 8331 9906 8337 9923
rect 8763 9906 8769 9923
rect 8331 9903 8769 9906
rect 8881 9923 9319 9926
rect 8881 9906 8887 9923
rect 9313 9906 9319 9923
rect 8881 9903 9319 9906
rect 9431 9923 9869 9926
rect 9431 9906 9437 9923
rect 9863 9906 9869 9923
rect 9431 9903 9869 9906
rect 9981 9923 10419 9926
rect 9981 9906 9987 9923
rect 10413 9906 10419 9923
rect 9981 9903 10419 9906
rect 10531 9923 10969 9926
rect 10531 9906 10537 9923
rect 10963 9906 10969 9923
rect 10531 9903 10969 9906
rect 11081 9923 11519 9926
rect 11081 9906 11087 9923
rect 11513 9906 11519 9923
rect 11081 9903 11519 9906
rect 11631 9923 12069 9926
rect 11631 9906 11637 9923
rect 12063 9906 12069 9923
rect 11631 9903 12069 9906
rect 12181 9923 12619 9926
rect 12181 9906 12187 9923
rect 12613 9906 12619 9923
rect 12181 9903 12619 9906
rect 12731 9923 13169 9926
rect 12731 9906 12737 9923
rect 13163 9906 13169 9923
rect 12731 9903 13169 9906
rect 13281 9923 13719 9926
rect 13281 9906 13287 9923
rect 13713 9906 13719 9923
rect 13281 9903 13719 9906
rect 13975 9919 13987 10450
rect 14263 9919 14275 10450
rect 13975 9900 14275 9919
rect -1025 9369 -1013 9900
rect -737 9369 -725 9900
rect -550 9892 -500 9900
rect -550 9858 -542 9892
rect -508 9858 -500 9892
rect -550 9850 -500 9858
rect 0 9892 50 9900
rect 0 9858 8 9892
rect 42 9858 50 9892
rect 0 9850 50 9858
rect 550 9892 600 9900
rect 550 9858 558 9892
rect 592 9858 600 9892
rect 550 9850 600 9858
rect 1100 9892 1150 9900
rect 1100 9858 1108 9892
rect 1142 9858 1150 9892
rect 1100 9850 1150 9858
rect 1650 9892 1700 9900
rect 1650 9858 1658 9892
rect 1692 9858 1700 9892
rect 1650 9850 1700 9858
rect 2200 9892 2250 9900
rect 2200 9858 2208 9892
rect 2242 9858 2250 9892
rect 2200 9850 2250 9858
rect 2750 9892 2800 9900
rect 2750 9858 2758 9892
rect 2792 9858 2800 9892
rect 2750 9850 2800 9858
rect 3300 9892 3350 9900
rect 3300 9858 3308 9892
rect 3342 9858 3350 9892
rect 3300 9850 3350 9858
rect 3850 9892 3900 9900
rect 3850 9858 3858 9892
rect 3892 9858 3900 9892
rect 3850 9850 3900 9858
rect 4400 9892 4450 9900
rect 4400 9858 4408 9892
rect 4442 9858 4450 9892
rect 4400 9850 4450 9858
rect 4950 9892 5000 9900
rect 4950 9858 4958 9892
rect 4992 9858 5000 9892
rect 4950 9850 5000 9858
rect 5500 9892 5550 9900
rect 5500 9858 5508 9892
rect 5542 9858 5550 9892
rect 5500 9850 5550 9858
rect 6050 9892 6100 9900
rect 6050 9858 6058 9892
rect 6092 9858 6100 9892
rect 6050 9850 6100 9858
rect 6600 9892 6650 9900
rect 6600 9858 6608 9892
rect 6642 9858 6650 9892
rect 6600 9850 6650 9858
rect 7150 9892 7200 9900
rect 7150 9858 7158 9892
rect 7192 9858 7200 9892
rect 7150 9850 7200 9858
rect 7700 9892 7750 9900
rect 7700 9858 7708 9892
rect 7742 9858 7750 9892
rect 7700 9850 7750 9858
rect 8250 9892 8300 9900
rect 8250 9858 8258 9892
rect 8292 9858 8300 9892
rect 8250 9850 8300 9858
rect 8800 9892 8850 9900
rect 8800 9858 8808 9892
rect 8842 9858 8850 9892
rect 8800 9850 8850 9858
rect 9350 9892 9400 9900
rect 9350 9858 9358 9892
rect 9392 9858 9400 9892
rect 9350 9850 9400 9858
rect 9900 9892 9950 9900
rect 9900 9858 9908 9892
rect 9942 9858 9950 9892
rect 9900 9850 9950 9858
rect 10450 9892 10500 9900
rect 10450 9858 10458 9892
rect 10492 9858 10500 9892
rect 10450 9850 10500 9858
rect 11000 9892 11050 9900
rect 11000 9858 11008 9892
rect 11042 9858 11050 9892
rect 11000 9850 11050 9858
rect 11550 9892 11600 9900
rect 11550 9858 11558 9892
rect 11592 9858 11600 9892
rect 11550 9850 11600 9858
rect 12100 9892 12150 9900
rect 12100 9858 12108 9892
rect 12142 9858 12150 9892
rect 12100 9850 12150 9858
rect 12650 9892 12700 9900
rect 12650 9858 12658 9892
rect 12692 9858 12700 9892
rect 12650 9850 12700 9858
rect 13200 9892 13250 9900
rect 13200 9858 13208 9892
rect 13242 9858 13250 9892
rect 13200 9850 13250 9858
rect 13750 9892 13800 9900
rect 13750 9858 13758 9892
rect 13792 9858 13800 9892
rect 13750 9850 13800 9858
rect -469 9844 -31 9847
rect -469 9827 -463 9844
rect -37 9827 -31 9844
rect -469 9824 -31 9827
rect 81 9844 519 9847
rect 81 9827 87 9844
rect 513 9827 519 9844
rect 81 9824 519 9827
rect 631 9844 1069 9847
rect 631 9827 637 9844
rect 1063 9827 1069 9844
rect 631 9824 1069 9827
rect 1181 9844 1619 9847
rect 1181 9827 1187 9844
rect 1613 9827 1619 9844
rect 1181 9824 1619 9827
rect 1731 9844 2169 9847
rect 1731 9827 1737 9844
rect 2163 9827 2169 9844
rect 1731 9824 2169 9827
rect 2281 9844 2719 9847
rect 2281 9827 2287 9844
rect 2713 9827 2719 9844
rect 2281 9824 2719 9827
rect 2831 9844 3269 9847
rect 2831 9827 2837 9844
rect 3263 9827 3269 9844
rect 2831 9824 3269 9827
rect 3381 9844 3819 9847
rect 3381 9827 3387 9844
rect 3813 9827 3819 9844
rect 3381 9824 3819 9827
rect 3931 9844 4369 9847
rect 3931 9827 3937 9844
rect 4363 9827 4369 9844
rect 3931 9824 4369 9827
rect 4481 9844 4919 9847
rect 4481 9827 4487 9844
rect 4913 9827 4919 9844
rect 4481 9824 4919 9827
rect 5031 9844 5469 9847
rect 5031 9827 5037 9844
rect 5463 9827 5469 9844
rect 5031 9824 5469 9827
rect 5581 9844 6019 9847
rect 5581 9827 5587 9844
rect 6013 9827 6019 9844
rect 5581 9824 6019 9827
rect 6131 9844 6569 9847
rect 6131 9827 6137 9844
rect 6563 9827 6569 9844
rect 6131 9824 6569 9827
rect 6681 9844 7119 9847
rect 6681 9827 6687 9844
rect 7113 9827 7119 9844
rect 6681 9824 7119 9827
rect 7231 9844 7669 9847
rect 7231 9827 7237 9844
rect 7663 9827 7669 9844
rect 7231 9824 7669 9827
rect 7781 9844 8219 9847
rect 7781 9827 7787 9844
rect 8213 9827 8219 9844
rect 7781 9824 8219 9827
rect 8331 9844 8769 9847
rect 8331 9827 8337 9844
rect 8763 9827 8769 9844
rect 8331 9824 8769 9827
rect 8881 9844 9319 9847
rect 8881 9827 8887 9844
rect 9313 9827 9319 9844
rect 8881 9824 9319 9827
rect 9431 9844 9869 9847
rect 9431 9827 9437 9844
rect 9863 9827 9869 9844
rect 9431 9824 9869 9827
rect 9981 9844 10419 9847
rect 9981 9827 9987 9844
rect 10413 9827 10419 9844
rect 9981 9824 10419 9827
rect 10531 9844 10969 9847
rect 10531 9827 10537 9844
rect 10963 9827 10969 9844
rect 10531 9824 10969 9827
rect 11081 9844 11519 9847
rect 11081 9827 11087 9844
rect 11513 9827 11519 9844
rect 11081 9824 11519 9827
rect 11631 9844 12069 9847
rect 11631 9827 11637 9844
rect 12063 9827 12069 9844
rect 11631 9824 12069 9827
rect 12181 9844 12619 9847
rect 12181 9827 12187 9844
rect 12613 9827 12619 9844
rect 12181 9824 12619 9827
rect 12731 9844 13169 9847
rect 12731 9827 12737 9844
rect 13163 9827 13169 9844
rect 12731 9824 13169 9827
rect 13281 9844 13719 9847
rect 13281 9827 13287 9844
rect 13713 9827 13719 9844
rect 13281 9824 13719 9827
rect -474 9819 -26 9824
rect 76 9819 524 9824
rect 626 9819 1074 9824
rect 1176 9819 1624 9824
rect 1726 9819 2174 9824
rect 2276 9819 2724 9824
rect 2826 9819 3274 9824
rect 3376 9819 3824 9824
rect 3926 9819 4374 9824
rect 4476 9819 4924 9824
rect 5026 9819 5474 9824
rect 5576 9819 6024 9824
rect 6126 9819 6574 9824
rect 6676 9819 7124 9824
rect 7226 9819 7674 9824
rect 7776 9819 8224 9824
rect 8326 9819 8774 9824
rect 8876 9819 9324 9824
rect 9426 9819 9874 9824
rect 9976 9819 10424 9824
rect 10526 9819 10974 9824
rect 11076 9819 11524 9824
rect 11626 9819 12074 9824
rect 12176 9819 12624 9824
rect 12726 9819 13174 9824
rect 13276 9819 13724 9824
rect -474 9813 -3 9819
rect -474 9765 -23 9813
rect -474 9435 -415 9765
rect -85 9435 -23 9765
rect -474 9387 -23 9435
rect -6 9387 -3 9813
rect -474 9381 -3 9387
rect 53 9813 547 9819
rect 53 9387 56 9813
rect 73 9765 527 9813
rect 73 9435 135 9765
rect 465 9435 527 9765
rect 73 9387 527 9435
rect 544 9387 547 9813
rect 53 9381 547 9387
rect 603 9813 1097 9819
rect 603 9387 606 9813
rect 623 9765 1077 9813
rect 623 9435 685 9765
rect 1015 9435 1077 9765
rect 623 9387 1077 9435
rect 1094 9387 1097 9813
rect 603 9381 1097 9387
rect 1153 9813 1647 9819
rect 1153 9387 1156 9813
rect 1173 9765 1627 9813
rect 1173 9435 1235 9765
rect 1565 9435 1627 9765
rect 1173 9387 1627 9435
rect 1644 9387 1647 9813
rect 1153 9381 1647 9387
rect 1703 9813 2197 9819
rect 1703 9387 1706 9813
rect 1723 9765 2177 9813
rect 1723 9435 1785 9765
rect 2115 9435 2177 9765
rect 1723 9387 2177 9435
rect 2194 9387 2197 9813
rect 1703 9381 2197 9387
rect 2253 9813 2747 9819
rect 2253 9387 2256 9813
rect 2273 9765 2727 9813
rect 2273 9435 2335 9765
rect 2665 9435 2727 9765
rect 2273 9387 2727 9435
rect 2744 9387 2747 9813
rect 2253 9381 2747 9387
rect 2803 9813 3297 9819
rect 2803 9387 2806 9813
rect 2823 9765 3277 9813
rect 2823 9435 2885 9765
rect 3215 9435 3277 9765
rect 2823 9387 3277 9435
rect 3294 9387 3297 9813
rect 2803 9381 3297 9387
rect 3353 9813 3847 9819
rect 3353 9387 3356 9813
rect 3373 9765 3827 9813
rect 3373 9435 3435 9765
rect 3765 9435 3827 9765
rect 3373 9387 3827 9435
rect 3844 9387 3847 9813
rect 3353 9381 3847 9387
rect 3903 9813 4397 9819
rect 3903 9387 3906 9813
rect 3923 9765 4377 9813
rect 3923 9435 3985 9765
rect 4315 9435 4377 9765
rect 3923 9387 4377 9435
rect 4394 9387 4397 9813
rect 3903 9381 4397 9387
rect 4453 9813 4947 9819
rect 4453 9387 4456 9813
rect 4473 9765 4927 9813
rect 4473 9435 4535 9765
rect 4865 9435 4927 9765
rect 4473 9387 4927 9435
rect 4944 9387 4947 9813
rect 4453 9381 4947 9387
rect 5003 9813 5497 9819
rect 5003 9387 5006 9813
rect 5023 9765 5477 9813
rect 5023 9435 5085 9765
rect 5415 9435 5477 9765
rect 5023 9387 5477 9435
rect 5494 9387 5497 9813
rect 5003 9381 5497 9387
rect 5553 9813 6047 9819
rect 5553 9387 5556 9813
rect 5573 9765 6027 9813
rect 5573 9435 5635 9765
rect 5965 9435 6027 9765
rect 5573 9387 6027 9435
rect 6044 9387 6047 9813
rect 5553 9381 6047 9387
rect 6103 9813 6597 9819
rect 6103 9387 6106 9813
rect 6123 9765 6577 9813
rect 6123 9435 6185 9765
rect 6515 9435 6577 9765
rect 6123 9387 6577 9435
rect 6594 9387 6597 9813
rect 6103 9381 6597 9387
rect 6653 9813 7147 9819
rect 6653 9387 6656 9813
rect 6673 9765 7127 9813
rect 6673 9435 6735 9765
rect 7065 9435 7127 9765
rect 6673 9387 7127 9435
rect 7144 9387 7147 9813
rect 6653 9381 7147 9387
rect 7203 9813 7697 9819
rect 7203 9387 7206 9813
rect 7223 9765 7677 9813
rect 7223 9435 7285 9765
rect 7615 9435 7677 9765
rect 7223 9387 7677 9435
rect 7694 9387 7697 9813
rect 7203 9381 7697 9387
rect 7753 9813 8247 9819
rect 7753 9387 7756 9813
rect 7773 9765 8227 9813
rect 7773 9435 7835 9765
rect 8165 9435 8227 9765
rect 7773 9387 8227 9435
rect 8244 9387 8247 9813
rect 7753 9381 8247 9387
rect 8303 9813 8797 9819
rect 8303 9387 8306 9813
rect 8323 9765 8777 9813
rect 8323 9435 8385 9765
rect 8715 9435 8777 9765
rect 8323 9387 8777 9435
rect 8794 9387 8797 9813
rect 8303 9381 8797 9387
rect 8853 9813 9347 9819
rect 8853 9387 8856 9813
rect 8873 9765 9327 9813
rect 8873 9435 8935 9765
rect 9265 9435 9327 9765
rect 8873 9387 9327 9435
rect 9344 9387 9347 9813
rect 8853 9381 9347 9387
rect 9403 9813 9897 9819
rect 9403 9387 9406 9813
rect 9423 9765 9877 9813
rect 9423 9435 9485 9765
rect 9815 9435 9877 9765
rect 9423 9387 9877 9435
rect 9894 9387 9897 9813
rect 9403 9381 9897 9387
rect 9953 9813 10447 9819
rect 9953 9387 9956 9813
rect 9973 9765 10427 9813
rect 9973 9435 10035 9765
rect 10365 9435 10427 9765
rect 9973 9387 10427 9435
rect 10444 9387 10447 9813
rect 9953 9381 10447 9387
rect 10503 9813 10997 9819
rect 10503 9387 10506 9813
rect 10523 9765 10977 9813
rect 10523 9435 10585 9765
rect 10915 9435 10977 9765
rect 10523 9387 10977 9435
rect 10994 9387 10997 9813
rect 10503 9381 10997 9387
rect 11053 9813 11547 9819
rect 11053 9387 11056 9813
rect 11073 9765 11527 9813
rect 11073 9435 11135 9765
rect 11465 9435 11527 9765
rect 11073 9387 11527 9435
rect 11544 9387 11547 9813
rect 11053 9381 11547 9387
rect 11603 9813 12097 9819
rect 11603 9387 11606 9813
rect 11623 9765 12077 9813
rect 11623 9435 11685 9765
rect 12015 9435 12077 9765
rect 11623 9387 12077 9435
rect 12094 9387 12097 9813
rect 11603 9381 12097 9387
rect 12153 9813 12647 9819
rect 12153 9387 12156 9813
rect 12173 9765 12627 9813
rect 12173 9435 12235 9765
rect 12565 9435 12627 9765
rect 12173 9387 12627 9435
rect 12644 9387 12647 9813
rect 12153 9381 12647 9387
rect 12703 9813 13197 9819
rect 12703 9387 12706 9813
rect 12723 9765 13177 9813
rect 12723 9435 12785 9765
rect 13115 9435 13177 9765
rect 12723 9387 13177 9435
rect 13194 9387 13197 9813
rect 12703 9381 13197 9387
rect 13253 9813 13724 9819
rect 13253 9387 13256 9813
rect 13273 9765 13724 9813
rect 13273 9435 13335 9765
rect 13665 9435 13724 9765
rect 13273 9387 13724 9435
rect 13253 9381 13724 9387
rect -474 9376 -26 9381
rect 76 9376 524 9381
rect 626 9376 1074 9381
rect 1176 9376 1624 9381
rect 1726 9376 2174 9381
rect 2276 9376 2724 9381
rect 2826 9376 3274 9381
rect 3376 9376 3824 9381
rect 3926 9376 4374 9381
rect 4476 9376 4924 9381
rect 5026 9376 5474 9381
rect 5576 9376 6024 9381
rect 6126 9376 6574 9381
rect 6676 9376 7124 9381
rect 7226 9376 7674 9381
rect 7776 9376 8224 9381
rect 8326 9376 8774 9381
rect 8876 9376 9324 9381
rect 9426 9376 9874 9381
rect 9976 9376 10424 9381
rect 10526 9376 10974 9381
rect 11076 9376 11524 9381
rect 11626 9376 12074 9381
rect 12176 9376 12624 9381
rect 12726 9376 13174 9381
rect 13276 9376 13724 9381
rect -1025 9350 -725 9369
rect -469 9373 -31 9376
rect -469 9356 -463 9373
rect -37 9356 -31 9373
rect -469 9353 -31 9356
rect 81 9373 519 9376
rect 81 9356 87 9373
rect 513 9356 519 9373
rect 81 9353 519 9356
rect 631 9373 1069 9376
rect 631 9356 637 9373
rect 1063 9356 1069 9373
rect 631 9353 1069 9356
rect 1181 9373 1619 9376
rect 1181 9356 1187 9373
rect 1613 9356 1619 9373
rect 1181 9353 1619 9356
rect 1731 9373 2169 9376
rect 1731 9356 1737 9373
rect 2163 9356 2169 9373
rect 1731 9353 2169 9356
rect 2281 9373 2719 9376
rect 2281 9356 2287 9373
rect 2713 9356 2719 9373
rect 2281 9353 2719 9356
rect 2831 9373 3269 9376
rect 2831 9356 2837 9373
rect 3263 9356 3269 9373
rect 2831 9353 3269 9356
rect 3381 9373 3819 9376
rect 3381 9356 3387 9373
rect 3813 9356 3819 9373
rect 3381 9353 3819 9356
rect 3931 9373 4369 9376
rect 3931 9356 3937 9373
rect 4363 9356 4369 9373
rect 3931 9353 4369 9356
rect 4481 9373 4919 9376
rect 4481 9356 4487 9373
rect 4913 9356 4919 9373
rect 4481 9353 4919 9356
rect 5031 9373 5469 9376
rect 5031 9356 5037 9373
rect 5463 9356 5469 9373
rect 5031 9353 5469 9356
rect 5581 9373 6019 9376
rect 5581 9356 5587 9373
rect 6013 9356 6019 9373
rect 5581 9353 6019 9356
rect 6131 9373 6569 9376
rect 6131 9356 6137 9373
rect 6563 9356 6569 9373
rect 6131 9353 6569 9356
rect 6681 9373 7119 9376
rect 6681 9356 6687 9373
rect 7113 9356 7119 9373
rect 6681 9353 7119 9356
rect 7231 9373 7669 9376
rect 7231 9356 7237 9373
rect 7663 9356 7669 9373
rect 7231 9353 7669 9356
rect 7781 9373 8219 9376
rect 7781 9356 7787 9373
rect 8213 9356 8219 9373
rect 7781 9353 8219 9356
rect 8331 9373 8769 9376
rect 8331 9356 8337 9373
rect 8763 9356 8769 9373
rect 8331 9353 8769 9356
rect 8881 9373 9319 9376
rect 8881 9356 8887 9373
rect 9313 9356 9319 9373
rect 8881 9353 9319 9356
rect 9431 9373 9869 9376
rect 9431 9356 9437 9373
rect 9863 9356 9869 9373
rect 9431 9353 9869 9356
rect 9981 9373 10419 9376
rect 9981 9356 9987 9373
rect 10413 9356 10419 9373
rect 9981 9353 10419 9356
rect 10531 9373 10969 9376
rect 10531 9356 10537 9373
rect 10963 9356 10969 9373
rect 10531 9353 10969 9356
rect 11081 9373 11519 9376
rect 11081 9356 11087 9373
rect 11513 9356 11519 9373
rect 11081 9353 11519 9356
rect 11631 9373 12069 9376
rect 11631 9356 11637 9373
rect 12063 9356 12069 9373
rect 11631 9353 12069 9356
rect 12181 9373 12619 9376
rect 12181 9356 12187 9373
rect 12613 9356 12619 9373
rect 12181 9353 12619 9356
rect 12731 9373 13169 9376
rect 12731 9356 12737 9373
rect 13163 9356 13169 9373
rect 12731 9353 13169 9356
rect 13281 9373 13719 9376
rect 13281 9356 13287 9373
rect 13713 9356 13719 9373
rect 13281 9353 13719 9356
rect 13975 9369 13987 9900
rect 14263 9369 14275 9900
rect 13975 9350 14275 9369
rect -1025 8819 -1013 9350
rect -737 8819 -725 9350
rect -550 9342 -500 9350
rect -550 9308 -542 9342
rect -508 9308 -500 9342
rect -550 9300 -500 9308
rect 0 9342 50 9350
rect 0 9308 8 9342
rect 42 9308 50 9342
rect 0 9300 50 9308
rect 550 9342 600 9350
rect 550 9308 558 9342
rect 592 9308 600 9342
rect 550 9300 600 9308
rect 1100 9342 1150 9350
rect 1100 9308 1108 9342
rect 1142 9308 1150 9342
rect 1100 9300 1150 9308
rect 1650 9342 1700 9350
rect 1650 9308 1658 9342
rect 1692 9308 1700 9342
rect 1650 9300 1700 9308
rect 2200 9342 2250 9350
rect 2200 9308 2208 9342
rect 2242 9308 2250 9342
rect 2200 9300 2250 9308
rect 2750 9342 2800 9350
rect 2750 9308 2758 9342
rect 2792 9308 2800 9342
rect 2750 9300 2800 9308
rect 3300 9342 3350 9350
rect 3300 9308 3308 9342
rect 3342 9308 3350 9342
rect 3300 9300 3350 9308
rect 3850 9342 3900 9350
rect 3850 9308 3858 9342
rect 3892 9308 3900 9342
rect 3850 9300 3900 9308
rect 4400 9342 4450 9350
rect 4400 9308 4408 9342
rect 4442 9308 4450 9342
rect 4400 9300 4450 9308
rect 4950 9342 5000 9350
rect 4950 9308 4958 9342
rect 4992 9308 5000 9342
rect 4950 9300 5000 9308
rect 5500 9342 5550 9350
rect 5500 9308 5508 9342
rect 5542 9308 5550 9342
rect 5500 9300 5550 9308
rect 6050 9342 6100 9350
rect 6050 9308 6058 9342
rect 6092 9308 6100 9342
rect 6050 9300 6100 9308
rect 6600 9342 6650 9350
rect 6600 9308 6608 9342
rect 6642 9308 6650 9342
rect 6600 9300 6650 9308
rect 7150 9342 7200 9350
rect 7150 9308 7158 9342
rect 7192 9308 7200 9342
rect 7150 9300 7200 9308
rect 7700 9342 7750 9350
rect 7700 9308 7708 9342
rect 7742 9308 7750 9342
rect 7700 9300 7750 9308
rect 8250 9342 8300 9350
rect 8250 9308 8258 9342
rect 8292 9308 8300 9342
rect 8250 9300 8300 9308
rect 8800 9342 8850 9350
rect 8800 9308 8808 9342
rect 8842 9308 8850 9342
rect 8800 9300 8850 9308
rect 9350 9342 9400 9350
rect 9350 9308 9358 9342
rect 9392 9308 9400 9342
rect 9350 9300 9400 9308
rect 9900 9342 9950 9350
rect 9900 9308 9908 9342
rect 9942 9308 9950 9342
rect 9900 9300 9950 9308
rect 10450 9342 10500 9350
rect 10450 9308 10458 9342
rect 10492 9308 10500 9342
rect 10450 9300 10500 9308
rect 11000 9342 11050 9350
rect 11000 9308 11008 9342
rect 11042 9308 11050 9342
rect 11000 9300 11050 9308
rect 11550 9342 11600 9350
rect 11550 9308 11558 9342
rect 11592 9308 11600 9342
rect 11550 9300 11600 9308
rect 12100 9342 12150 9350
rect 12100 9308 12108 9342
rect 12142 9308 12150 9342
rect 12100 9300 12150 9308
rect 12650 9342 12700 9350
rect 12650 9308 12658 9342
rect 12692 9308 12700 9342
rect 12650 9300 12700 9308
rect 13200 9342 13250 9350
rect 13200 9308 13208 9342
rect 13242 9308 13250 9342
rect 13200 9300 13250 9308
rect 13750 9342 13800 9350
rect 13750 9308 13758 9342
rect 13792 9308 13800 9342
rect 13750 9300 13800 9308
rect -469 9294 -31 9297
rect -469 9277 -463 9294
rect -37 9277 -31 9294
rect -469 9274 -31 9277
rect 81 9294 519 9297
rect 81 9277 87 9294
rect 513 9277 519 9294
rect 81 9274 519 9277
rect 631 9294 1069 9297
rect 631 9277 637 9294
rect 1063 9277 1069 9294
rect 631 9274 1069 9277
rect 1181 9294 1619 9297
rect 1181 9277 1187 9294
rect 1613 9277 1619 9294
rect 1181 9274 1619 9277
rect 1731 9294 2169 9297
rect 1731 9277 1737 9294
rect 2163 9277 2169 9294
rect 1731 9274 2169 9277
rect 2281 9294 2719 9297
rect 2281 9277 2287 9294
rect 2713 9277 2719 9294
rect 2281 9274 2719 9277
rect 2831 9294 3269 9297
rect 2831 9277 2837 9294
rect 3263 9277 3269 9294
rect 2831 9274 3269 9277
rect 3381 9294 3819 9297
rect 3381 9277 3387 9294
rect 3813 9277 3819 9294
rect 3381 9274 3819 9277
rect 3931 9294 4369 9297
rect 3931 9277 3937 9294
rect 4363 9277 4369 9294
rect 3931 9274 4369 9277
rect 4481 9294 4919 9297
rect 4481 9277 4487 9294
rect 4913 9277 4919 9294
rect 4481 9274 4919 9277
rect 5031 9294 5469 9297
rect 5031 9277 5037 9294
rect 5463 9277 5469 9294
rect 5031 9274 5469 9277
rect 5581 9294 6019 9297
rect 5581 9277 5587 9294
rect 6013 9277 6019 9294
rect 5581 9274 6019 9277
rect 6131 9294 6569 9297
rect 6131 9277 6137 9294
rect 6563 9277 6569 9294
rect 6131 9274 6569 9277
rect 6681 9294 7119 9297
rect 6681 9277 6687 9294
rect 7113 9277 7119 9294
rect 6681 9274 7119 9277
rect 7231 9294 7669 9297
rect 7231 9277 7237 9294
rect 7663 9277 7669 9294
rect 7231 9274 7669 9277
rect 7781 9294 8219 9297
rect 7781 9277 7787 9294
rect 8213 9277 8219 9294
rect 7781 9274 8219 9277
rect 8331 9294 8769 9297
rect 8331 9277 8337 9294
rect 8763 9277 8769 9294
rect 8331 9274 8769 9277
rect 8881 9294 9319 9297
rect 8881 9277 8887 9294
rect 9313 9277 9319 9294
rect 8881 9274 9319 9277
rect 9431 9294 9869 9297
rect 9431 9277 9437 9294
rect 9863 9277 9869 9294
rect 9431 9274 9869 9277
rect 9981 9294 10419 9297
rect 9981 9277 9987 9294
rect 10413 9277 10419 9294
rect 9981 9274 10419 9277
rect 10531 9294 10969 9297
rect 10531 9277 10537 9294
rect 10963 9277 10969 9294
rect 10531 9274 10969 9277
rect 11081 9294 11519 9297
rect 11081 9277 11087 9294
rect 11513 9277 11519 9294
rect 11081 9274 11519 9277
rect 11631 9294 12069 9297
rect 11631 9277 11637 9294
rect 12063 9277 12069 9294
rect 11631 9274 12069 9277
rect 12181 9294 12619 9297
rect 12181 9277 12187 9294
rect 12613 9277 12619 9294
rect 12181 9274 12619 9277
rect 12731 9294 13169 9297
rect 12731 9277 12737 9294
rect 13163 9277 13169 9294
rect 12731 9274 13169 9277
rect 13281 9294 13719 9297
rect 13281 9277 13287 9294
rect 13713 9277 13719 9294
rect 13281 9274 13719 9277
rect -474 9269 -26 9274
rect 76 9269 524 9274
rect 626 9269 1074 9274
rect 1176 9269 1624 9274
rect 1726 9269 2174 9274
rect 2276 9269 2724 9274
rect 2826 9269 3274 9274
rect 3376 9269 3824 9274
rect 3926 9269 4374 9274
rect 4476 9269 4924 9274
rect 5026 9269 5474 9274
rect 5576 9269 6024 9274
rect 6126 9269 6574 9274
rect 6676 9269 7124 9274
rect 7226 9269 7674 9274
rect 7776 9269 8224 9274
rect 8326 9269 8774 9274
rect 8876 9269 9324 9274
rect 9426 9269 9874 9274
rect 9976 9269 10424 9274
rect 10526 9269 10974 9274
rect 11076 9269 11524 9274
rect 11626 9269 12074 9274
rect 12176 9269 12624 9274
rect 12726 9269 13174 9274
rect 13276 9269 13724 9274
rect -474 9263 -3 9269
rect -474 9215 -23 9263
rect -474 8885 -415 9215
rect -85 8885 -23 9215
rect -474 8837 -23 8885
rect -6 8837 -3 9263
rect -474 8831 -3 8837
rect 53 9263 547 9269
rect 53 8837 56 9263
rect 73 9215 527 9263
rect 73 8885 135 9215
rect 465 8885 527 9215
rect 73 8837 527 8885
rect 544 8837 547 9263
rect 53 8831 547 8837
rect 603 9263 1097 9269
rect 603 8837 606 9263
rect 623 9215 1077 9263
rect 623 8885 685 9215
rect 1015 8885 1077 9215
rect 623 8837 1077 8885
rect 1094 8837 1097 9263
rect 603 8831 1097 8837
rect 1153 9263 1647 9269
rect 1153 8837 1156 9263
rect 1173 9215 1627 9263
rect 1173 8885 1235 9215
rect 1565 8885 1627 9215
rect 1173 8837 1627 8885
rect 1644 8837 1647 9263
rect 1153 8831 1647 8837
rect 1703 9263 2197 9269
rect 1703 8837 1706 9263
rect 1723 9215 2177 9263
rect 1723 8885 1785 9215
rect 2115 8885 2177 9215
rect 1723 8837 2177 8885
rect 2194 8837 2197 9263
rect 1703 8831 2197 8837
rect 2253 9263 2747 9269
rect 2253 8837 2256 9263
rect 2273 9215 2727 9263
rect 2273 8885 2335 9215
rect 2665 8885 2727 9215
rect 2273 8837 2727 8885
rect 2744 8837 2747 9263
rect 2253 8831 2747 8837
rect 2803 9263 3297 9269
rect 2803 8837 2806 9263
rect 2823 9215 3277 9263
rect 2823 8885 2885 9215
rect 3215 8885 3277 9215
rect 2823 8837 3277 8885
rect 3294 8837 3297 9263
rect 2803 8831 3297 8837
rect 3353 9263 3847 9269
rect 3353 8837 3356 9263
rect 3373 9215 3827 9263
rect 3373 8885 3435 9215
rect 3765 8885 3827 9215
rect 3373 8837 3827 8885
rect 3844 8837 3847 9263
rect 3353 8831 3847 8837
rect 3903 9263 4397 9269
rect 3903 8837 3906 9263
rect 3923 9215 4377 9263
rect 3923 8885 3985 9215
rect 4315 8885 4377 9215
rect 3923 8837 4377 8885
rect 4394 8837 4397 9263
rect 3903 8831 4397 8837
rect 4453 9263 4947 9269
rect 4453 8837 4456 9263
rect 4473 9215 4927 9263
rect 4473 8885 4535 9215
rect 4865 8885 4927 9215
rect 4473 8837 4927 8885
rect 4944 8837 4947 9263
rect 4453 8831 4947 8837
rect 5003 9263 5497 9269
rect 5003 8837 5006 9263
rect 5023 9215 5477 9263
rect 5023 8885 5085 9215
rect 5415 8885 5477 9215
rect 5023 8837 5477 8885
rect 5494 8837 5497 9263
rect 5003 8831 5497 8837
rect 5553 9263 6047 9269
rect 5553 8837 5556 9263
rect 5573 9215 6027 9263
rect 5573 8885 5635 9215
rect 5965 8885 6027 9215
rect 5573 8837 6027 8885
rect 6044 8837 6047 9263
rect 5553 8831 6047 8837
rect 6103 9263 6597 9269
rect 6103 8837 6106 9263
rect 6123 9215 6577 9263
rect 6123 8885 6185 9215
rect 6515 8885 6577 9215
rect 6123 8837 6577 8885
rect 6594 8837 6597 9263
rect 6103 8831 6597 8837
rect 6653 9263 7147 9269
rect 6653 8837 6656 9263
rect 6673 9215 7127 9263
rect 6673 8885 6735 9215
rect 7065 8885 7127 9215
rect 6673 8837 7127 8885
rect 7144 8837 7147 9263
rect 6653 8831 7147 8837
rect 7203 9263 7697 9269
rect 7203 8837 7206 9263
rect 7223 9215 7677 9263
rect 7223 8885 7285 9215
rect 7615 8885 7677 9215
rect 7223 8837 7677 8885
rect 7694 8837 7697 9263
rect 7203 8831 7697 8837
rect 7753 9263 8247 9269
rect 7753 8837 7756 9263
rect 7773 9215 8227 9263
rect 7773 8885 7835 9215
rect 8165 8885 8227 9215
rect 7773 8837 8227 8885
rect 8244 8837 8247 9263
rect 7753 8831 8247 8837
rect 8303 9263 8797 9269
rect 8303 8837 8306 9263
rect 8323 9215 8777 9263
rect 8323 8885 8385 9215
rect 8715 8885 8777 9215
rect 8323 8837 8777 8885
rect 8794 8837 8797 9263
rect 8303 8831 8797 8837
rect 8853 9263 9347 9269
rect 8853 8837 8856 9263
rect 8873 9215 9327 9263
rect 8873 8885 8935 9215
rect 9265 8885 9327 9215
rect 8873 8837 9327 8885
rect 9344 8837 9347 9263
rect 8853 8831 9347 8837
rect 9403 9263 9897 9269
rect 9403 8837 9406 9263
rect 9423 9215 9877 9263
rect 9423 8885 9485 9215
rect 9815 8885 9877 9215
rect 9423 8837 9877 8885
rect 9894 8837 9897 9263
rect 9403 8831 9897 8837
rect 9953 9263 10447 9269
rect 9953 8837 9956 9263
rect 9973 9215 10427 9263
rect 9973 8885 10035 9215
rect 10365 8885 10427 9215
rect 9973 8837 10427 8885
rect 10444 8837 10447 9263
rect 9953 8831 10447 8837
rect 10503 9263 10997 9269
rect 10503 8837 10506 9263
rect 10523 9215 10977 9263
rect 10523 8885 10585 9215
rect 10915 8885 10977 9215
rect 10523 8837 10977 8885
rect 10994 8837 10997 9263
rect 10503 8831 10997 8837
rect 11053 9263 11547 9269
rect 11053 8837 11056 9263
rect 11073 9215 11527 9263
rect 11073 8885 11135 9215
rect 11465 8885 11527 9215
rect 11073 8837 11527 8885
rect 11544 8837 11547 9263
rect 11053 8831 11547 8837
rect 11603 9263 12097 9269
rect 11603 8837 11606 9263
rect 11623 9215 12077 9263
rect 11623 8885 11685 9215
rect 12015 8885 12077 9215
rect 11623 8837 12077 8885
rect 12094 8837 12097 9263
rect 11603 8831 12097 8837
rect 12153 9263 12647 9269
rect 12153 8837 12156 9263
rect 12173 9215 12627 9263
rect 12173 8885 12235 9215
rect 12565 8885 12627 9215
rect 12173 8837 12627 8885
rect 12644 8837 12647 9263
rect 12153 8831 12647 8837
rect 12703 9263 13197 9269
rect 12703 8837 12706 9263
rect 12723 9215 13177 9263
rect 12723 8885 12785 9215
rect 13115 8885 13177 9215
rect 12723 8837 13177 8885
rect 13194 8837 13197 9263
rect 12703 8831 13197 8837
rect 13253 9263 13724 9269
rect 13253 8837 13256 9263
rect 13273 9215 13724 9263
rect 13273 8885 13335 9215
rect 13665 8885 13724 9215
rect 13273 8837 13724 8885
rect 13253 8831 13724 8837
rect -474 8826 -26 8831
rect 76 8826 524 8831
rect 626 8826 1074 8831
rect 1176 8826 1624 8831
rect 1726 8826 2174 8831
rect 2276 8826 2724 8831
rect 2826 8826 3274 8831
rect 3376 8826 3824 8831
rect 3926 8826 4374 8831
rect 4476 8826 4924 8831
rect 5026 8826 5474 8831
rect 5576 8826 6024 8831
rect 6126 8826 6574 8831
rect 6676 8826 7124 8831
rect 7226 8826 7674 8831
rect 7776 8826 8224 8831
rect 8326 8826 8774 8831
rect 8876 8826 9324 8831
rect 9426 8826 9874 8831
rect 9976 8826 10424 8831
rect 10526 8826 10974 8831
rect 11076 8826 11524 8831
rect 11626 8826 12074 8831
rect 12176 8826 12624 8831
rect 12726 8826 13174 8831
rect 13276 8826 13724 8831
rect -1025 8800 -725 8819
rect -469 8823 -31 8826
rect -469 8806 -463 8823
rect -37 8806 -31 8823
rect -469 8803 -31 8806
rect 81 8823 519 8826
rect 81 8806 87 8823
rect 513 8806 519 8823
rect 81 8803 519 8806
rect 631 8823 1069 8826
rect 631 8806 637 8823
rect 1063 8806 1069 8823
rect 631 8803 1069 8806
rect 1181 8823 1619 8826
rect 1181 8806 1187 8823
rect 1613 8806 1619 8823
rect 1181 8803 1619 8806
rect 1731 8823 2169 8826
rect 1731 8806 1737 8823
rect 2163 8806 2169 8823
rect 1731 8803 2169 8806
rect 2281 8823 2719 8826
rect 2281 8806 2287 8823
rect 2713 8806 2719 8823
rect 2281 8803 2719 8806
rect 2831 8823 3269 8826
rect 2831 8806 2837 8823
rect 3263 8806 3269 8823
rect 2831 8803 3269 8806
rect 3381 8823 3819 8826
rect 3381 8806 3387 8823
rect 3813 8806 3819 8823
rect 3381 8803 3819 8806
rect 3931 8823 4369 8826
rect 3931 8806 3937 8823
rect 4363 8806 4369 8823
rect 3931 8803 4369 8806
rect 4481 8823 4919 8826
rect 4481 8806 4487 8823
rect 4913 8806 4919 8823
rect 4481 8803 4919 8806
rect 5031 8823 5469 8826
rect 5031 8806 5037 8823
rect 5463 8806 5469 8823
rect 5031 8803 5469 8806
rect 5581 8823 6019 8826
rect 5581 8806 5587 8823
rect 6013 8806 6019 8823
rect 5581 8803 6019 8806
rect 6131 8823 6569 8826
rect 6131 8806 6137 8823
rect 6563 8806 6569 8823
rect 6131 8803 6569 8806
rect 6681 8823 7119 8826
rect 6681 8806 6687 8823
rect 7113 8806 7119 8823
rect 6681 8803 7119 8806
rect 7231 8823 7669 8826
rect 7231 8806 7237 8823
rect 7663 8806 7669 8823
rect 7231 8803 7669 8806
rect 7781 8823 8219 8826
rect 7781 8806 7787 8823
rect 8213 8806 8219 8823
rect 7781 8803 8219 8806
rect 8331 8823 8769 8826
rect 8331 8806 8337 8823
rect 8763 8806 8769 8823
rect 8331 8803 8769 8806
rect 8881 8823 9319 8826
rect 8881 8806 8887 8823
rect 9313 8806 9319 8823
rect 8881 8803 9319 8806
rect 9431 8823 9869 8826
rect 9431 8806 9437 8823
rect 9863 8806 9869 8823
rect 9431 8803 9869 8806
rect 9981 8823 10419 8826
rect 9981 8806 9987 8823
rect 10413 8806 10419 8823
rect 9981 8803 10419 8806
rect 10531 8823 10969 8826
rect 10531 8806 10537 8823
rect 10963 8806 10969 8823
rect 10531 8803 10969 8806
rect 11081 8823 11519 8826
rect 11081 8806 11087 8823
rect 11513 8806 11519 8823
rect 11081 8803 11519 8806
rect 11631 8823 12069 8826
rect 11631 8806 11637 8823
rect 12063 8806 12069 8823
rect 11631 8803 12069 8806
rect 12181 8823 12619 8826
rect 12181 8806 12187 8823
rect 12613 8806 12619 8823
rect 12181 8803 12619 8806
rect 12731 8823 13169 8826
rect 12731 8806 12737 8823
rect 13163 8806 13169 8823
rect 12731 8803 13169 8806
rect 13281 8823 13719 8826
rect 13281 8806 13287 8823
rect 13713 8806 13719 8823
rect 13281 8803 13719 8806
rect 13975 8819 13987 9350
rect 14263 8819 14275 9350
rect 13975 8800 14275 8819
rect -1025 8269 -1013 8800
rect -737 8269 -725 8800
rect -550 8792 -500 8800
rect -550 8758 -542 8792
rect -508 8758 -500 8792
rect -550 8750 -500 8758
rect 0 8792 50 8800
rect 0 8758 8 8792
rect 42 8758 50 8792
rect 0 8750 50 8758
rect 550 8792 600 8800
rect 550 8758 558 8792
rect 592 8758 600 8792
rect 550 8750 600 8758
rect 1100 8792 1150 8800
rect 1100 8758 1108 8792
rect 1142 8758 1150 8792
rect 1100 8750 1150 8758
rect 1650 8792 1700 8800
rect 1650 8758 1658 8792
rect 1692 8758 1700 8792
rect 1650 8750 1700 8758
rect 2200 8792 2250 8800
rect 2200 8758 2208 8792
rect 2242 8758 2250 8792
rect 2200 8750 2250 8758
rect 2750 8792 2800 8800
rect 2750 8758 2758 8792
rect 2792 8758 2800 8792
rect 2750 8750 2800 8758
rect 3300 8792 3350 8800
rect 3300 8758 3308 8792
rect 3342 8758 3350 8792
rect 3300 8750 3350 8758
rect 3850 8792 3900 8800
rect 3850 8758 3858 8792
rect 3892 8758 3900 8792
rect 3850 8750 3900 8758
rect 4400 8792 4450 8800
rect 4400 8758 4408 8792
rect 4442 8758 4450 8792
rect 4400 8750 4450 8758
rect 4950 8792 5000 8800
rect 4950 8758 4958 8792
rect 4992 8758 5000 8792
rect 4950 8750 5000 8758
rect 5500 8792 5550 8800
rect 5500 8758 5508 8792
rect 5542 8758 5550 8792
rect 5500 8750 5550 8758
rect 6050 8792 6100 8800
rect 6050 8758 6058 8792
rect 6092 8758 6100 8792
rect 6050 8750 6100 8758
rect 6600 8792 6650 8800
rect 6600 8758 6608 8792
rect 6642 8758 6650 8792
rect 6600 8750 6650 8758
rect 7150 8792 7200 8800
rect 7150 8758 7158 8792
rect 7192 8758 7200 8792
rect 7150 8750 7200 8758
rect 7700 8792 7750 8800
rect 7700 8758 7708 8792
rect 7742 8758 7750 8792
rect 7700 8750 7750 8758
rect 8250 8792 8300 8800
rect 8250 8758 8258 8792
rect 8292 8758 8300 8792
rect 8250 8750 8300 8758
rect 8800 8792 8850 8800
rect 8800 8758 8808 8792
rect 8842 8758 8850 8792
rect 8800 8750 8850 8758
rect 9350 8792 9400 8800
rect 9350 8758 9358 8792
rect 9392 8758 9400 8792
rect 9350 8750 9400 8758
rect 9900 8792 9950 8800
rect 9900 8758 9908 8792
rect 9942 8758 9950 8792
rect 9900 8750 9950 8758
rect 10450 8792 10500 8800
rect 10450 8758 10458 8792
rect 10492 8758 10500 8792
rect 10450 8750 10500 8758
rect 11000 8792 11050 8800
rect 11000 8758 11008 8792
rect 11042 8758 11050 8792
rect 11000 8750 11050 8758
rect 11550 8792 11600 8800
rect 11550 8758 11558 8792
rect 11592 8758 11600 8792
rect 11550 8750 11600 8758
rect 12100 8792 12150 8800
rect 12100 8758 12108 8792
rect 12142 8758 12150 8792
rect 12100 8750 12150 8758
rect 12650 8792 12700 8800
rect 12650 8758 12658 8792
rect 12692 8758 12700 8792
rect 12650 8750 12700 8758
rect 13200 8792 13250 8800
rect 13200 8758 13208 8792
rect 13242 8758 13250 8792
rect 13200 8750 13250 8758
rect 13750 8792 13800 8800
rect 13750 8758 13758 8792
rect 13792 8758 13800 8792
rect 13750 8750 13800 8758
rect -469 8744 -31 8747
rect -469 8727 -463 8744
rect -37 8727 -31 8744
rect -469 8724 -31 8727
rect 81 8744 519 8747
rect 81 8727 87 8744
rect 513 8727 519 8744
rect 81 8724 519 8727
rect 631 8744 1069 8747
rect 631 8727 637 8744
rect 1063 8727 1069 8744
rect 631 8724 1069 8727
rect 1181 8744 1619 8747
rect 1181 8727 1187 8744
rect 1613 8727 1619 8744
rect 1181 8724 1619 8727
rect 1731 8744 2169 8747
rect 1731 8727 1737 8744
rect 2163 8727 2169 8744
rect 1731 8724 2169 8727
rect 2281 8744 2719 8747
rect 2281 8727 2287 8744
rect 2713 8727 2719 8744
rect 2281 8724 2719 8727
rect 2831 8744 3269 8747
rect 2831 8727 2837 8744
rect 3263 8727 3269 8744
rect 2831 8724 3269 8727
rect 3381 8744 3819 8747
rect 3381 8727 3387 8744
rect 3813 8727 3819 8744
rect 3381 8724 3819 8727
rect 3931 8744 4369 8747
rect 3931 8727 3937 8744
rect 4363 8727 4369 8744
rect 3931 8724 4369 8727
rect 4481 8744 4919 8747
rect 4481 8727 4487 8744
rect 4913 8727 4919 8744
rect 4481 8724 4919 8727
rect 5031 8744 5469 8747
rect 5031 8727 5037 8744
rect 5463 8727 5469 8744
rect 5031 8724 5469 8727
rect 5581 8744 6019 8747
rect 5581 8727 5587 8744
rect 6013 8727 6019 8744
rect 5581 8724 6019 8727
rect 6131 8744 6569 8747
rect 6131 8727 6137 8744
rect 6563 8727 6569 8744
rect 6131 8724 6569 8727
rect 6681 8744 7119 8747
rect 6681 8727 6687 8744
rect 7113 8727 7119 8744
rect 6681 8724 7119 8727
rect 7231 8744 7669 8747
rect 7231 8727 7237 8744
rect 7663 8727 7669 8744
rect 7231 8724 7669 8727
rect 7781 8744 8219 8747
rect 7781 8727 7787 8744
rect 8213 8727 8219 8744
rect 7781 8724 8219 8727
rect 8331 8744 8769 8747
rect 8331 8727 8337 8744
rect 8763 8727 8769 8744
rect 8331 8724 8769 8727
rect 8881 8744 9319 8747
rect 8881 8727 8887 8744
rect 9313 8727 9319 8744
rect 8881 8724 9319 8727
rect 9431 8744 9869 8747
rect 9431 8727 9437 8744
rect 9863 8727 9869 8744
rect 9431 8724 9869 8727
rect 9981 8744 10419 8747
rect 9981 8727 9987 8744
rect 10413 8727 10419 8744
rect 9981 8724 10419 8727
rect 10531 8744 10969 8747
rect 10531 8727 10537 8744
rect 10963 8727 10969 8744
rect 10531 8724 10969 8727
rect 11081 8744 11519 8747
rect 11081 8727 11087 8744
rect 11513 8727 11519 8744
rect 11081 8724 11519 8727
rect 11631 8744 12069 8747
rect 11631 8727 11637 8744
rect 12063 8727 12069 8744
rect 11631 8724 12069 8727
rect 12181 8744 12619 8747
rect 12181 8727 12187 8744
rect 12613 8727 12619 8744
rect 12181 8724 12619 8727
rect 12731 8744 13169 8747
rect 12731 8727 12737 8744
rect 13163 8727 13169 8744
rect 12731 8724 13169 8727
rect 13281 8744 13719 8747
rect 13281 8727 13287 8744
rect 13713 8727 13719 8744
rect 13281 8724 13719 8727
rect -474 8719 -26 8724
rect 76 8719 524 8724
rect 626 8719 1074 8724
rect 1176 8719 1624 8724
rect 1726 8719 2174 8724
rect 2276 8719 2724 8724
rect 2826 8719 3274 8724
rect 3376 8719 3824 8724
rect 3926 8719 4374 8724
rect 4476 8719 4924 8724
rect 5026 8719 5474 8724
rect 5576 8719 6024 8724
rect 6126 8719 6574 8724
rect 6676 8719 7124 8724
rect 7226 8719 7674 8724
rect 7776 8719 8224 8724
rect 8326 8719 8774 8724
rect 8876 8719 9324 8724
rect 9426 8719 9874 8724
rect 9976 8719 10424 8724
rect 10526 8719 10974 8724
rect 11076 8719 11524 8724
rect 11626 8719 12074 8724
rect 12176 8719 12624 8724
rect 12726 8719 13174 8724
rect 13276 8719 13724 8724
rect -474 8713 -3 8719
rect -474 8665 -23 8713
rect -474 8335 -415 8665
rect -85 8335 -23 8665
rect -474 8287 -23 8335
rect -6 8287 -3 8713
rect -474 8281 -3 8287
rect 53 8713 547 8719
rect 53 8287 56 8713
rect 73 8665 527 8713
rect 73 8335 135 8665
rect 465 8335 527 8665
rect 73 8287 527 8335
rect 544 8287 547 8713
rect 53 8281 547 8287
rect 603 8713 1097 8719
rect 603 8287 606 8713
rect 623 8665 1077 8713
rect 623 8335 685 8665
rect 1015 8335 1077 8665
rect 623 8287 1077 8335
rect 1094 8287 1097 8713
rect 603 8281 1097 8287
rect 1153 8713 1647 8719
rect 1153 8287 1156 8713
rect 1173 8665 1627 8713
rect 1173 8335 1235 8665
rect 1565 8335 1627 8665
rect 1173 8287 1627 8335
rect 1644 8287 1647 8713
rect 1153 8281 1647 8287
rect 1703 8713 2197 8719
rect 1703 8287 1706 8713
rect 1723 8665 2177 8713
rect 1723 8335 1785 8665
rect 2115 8335 2177 8665
rect 1723 8287 2177 8335
rect 2194 8287 2197 8713
rect 1703 8281 2197 8287
rect 2253 8713 2747 8719
rect 2253 8287 2256 8713
rect 2273 8665 2727 8713
rect 2273 8335 2335 8665
rect 2665 8335 2727 8665
rect 2273 8287 2727 8335
rect 2744 8287 2747 8713
rect 2253 8281 2747 8287
rect 2803 8713 3297 8719
rect 2803 8287 2806 8713
rect 2823 8665 3277 8713
rect 2823 8335 2885 8665
rect 3215 8335 3277 8665
rect 2823 8287 3277 8335
rect 3294 8287 3297 8713
rect 2803 8281 3297 8287
rect 3353 8713 3847 8719
rect 3353 8287 3356 8713
rect 3373 8665 3827 8713
rect 3373 8335 3435 8665
rect 3765 8335 3827 8665
rect 3373 8287 3827 8335
rect 3844 8287 3847 8713
rect 3353 8281 3847 8287
rect 3903 8713 4397 8719
rect 3903 8287 3906 8713
rect 3923 8665 4377 8713
rect 3923 8335 3985 8665
rect 4315 8335 4377 8665
rect 3923 8287 4377 8335
rect 4394 8287 4397 8713
rect 3903 8281 4397 8287
rect 4453 8713 4947 8719
rect 4453 8287 4456 8713
rect 4473 8665 4927 8713
rect 4473 8335 4535 8665
rect 4865 8335 4927 8665
rect 4473 8287 4927 8335
rect 4944 8287 4947 8713
rect 4453 8281 4947 8287
rect 5003 8713 5497 8719
rect 5003 8287 5006 8713
rect 5023 8665 5477 8713
rect 5023 8335 5085 8665
rect 5415 8335 5477 8665
rect 5023 8287 5477 8335
rect 5494 8287 5497 8713
rect 5003 8281 5497 8287
rect 5553 8713 6047 8719
rect 5553 8287 5556 8713
rect 5573 8665 6027 8713
rect 5573 8335 5635 8665
rect 5965 8335 6027 8665
rect 5573 8287 6027 8335
rect 6044 8287 6047 8713
rect 5553 8281 6047 8287
rect 6103 8713 6597 8719
rect 6103 8287 6106 8713
rect 6123 8665 6577 8713
rect 6123 8335 6185 8665
rect 6515 8335 6577 8665
rect 6123 8287 6577 8335
rect 6594 8287 6597 8713
rect 6103 8281 6597 8287
rect 6653 8713 7147 8719
rect 6653 8287 6656 8713
rect 6673 8665 7127 8713
rect 6673 8335 6735 8665
rect 7065 8335 7127 8665
rect 6673 8287 7127 8335
rect 7144 8287 7147 8713
rect 6653 8281 7147 8287
rect 7203 8713 7697 8719
rect 7203 8287 7206 8713
rect 7223 8665 7677 8713
rect 7223 8335 7285 8665
rect 7615 8335 7677 8665
rect 7223 8287 7677 8335
rect 7694 8287 7697 8713
rect 7203 8281 7697 8287
rect 7753 8713 8247 8719
rect 7753 8287 7756 8713
rect 7773 8665 8227 8713
rect 7773 8335 7835 8665
rect 8165 8335 8227 8665
rect 7773 8287 8227 8335
rect 8244 8287 8247 8713
rect 7753 8281 8247 8287
rect 8303 8713 8797 8719
rect 8303 8287 8306 8713
rect 8323 8665 8777 8713
rect 8323 8335 8385 8665
rect 8715 8335 8777 8665
rect 8323 8287 8777 8335
rect 8794 8287 8797 8713
rect 8303 8281 8797 8287
rect 8853 8713 9347 8719
rect 8853 8287 8856 8713
rect 8873 8665 9327 8713
rect 8873 8335 8935 8665
rect 9265 8335 9327 8665
rect 8873 8287 9327 8335
rect 9344 8287 9347 8713
rect 8853 8281 9347 8287
rect 9403 8713 9897 8719
rect 9403 8287 9406 8713
rect 9423 8665 9877 8713
rect 9423 8335 9485 8665
rect 9815 8335 9877 8665
rect 9423 8287 9877 8335
rect 9894 8287 9897 8713
rect 9403 8281 9897 8287
rect 9953 8713 10447 8719
rect 9953 8287 9956 8713
rect 9973 8665 10427 8713
rect 9973 8335 10035 8665
rect 10365 8335 10427 8665
rect 9973 8287 10427 8335
rect 10444 8287 10447 8713
rect 9953 8281 10447 8287
rect 10503 8713 10997 8719
rect 10503 8287 10506 8713
rect 10523 8665 10977 8713
rect 10523 8335 10585 8665
rect 10915 8335 10977 8665
rect 10523 8287 10977 8335
rect 10994 8287 10997 8713
rect 10503 8281 10997 8287
rect 11053 8713 11547 8719
rect 11053 8287 11056 8713
rect 11073 8665 11527 8713
rect 11073 8335 11135 8665
rect 11465 8335 11527 8665
rect 11073 8287 11527 8335
rect 11544 8287 11547 8713
rect 11053 8281 11547 8287
rect 11603 8713 12097 8719
rect 11603 8287 11606 8713
rect 11623 8665 12077 8713
rect 11623 8335 11685 8665
rect 12015 8335 12077 8665
rect 11623 8287 12077 8335
rect 12094 8287 12097 8713
rect 11603 8281 12097 8287
rect 12153 8713 12647 8719
rect 12153 8287 12156 8713
rect 12173 8665 12627 8713
rect 12173 8335 12235 8665
rect 12565 8335 12627 8665
rect 12173 8287 12627 8335
rect 12644 8287 12647 8713
rect 12153 8281 12647 8287
rect 12703 8713 13197 8719
rect 12703 8287 12706 8713
rect 12723 8665 13177 8713
rect 12723 8335 12785 8665
rect 13115 8335 13177 8665
rect 12723 8287 13177 8335
rect 13194 8287 13197 8713
rect 12703 8281 13197 8287
rect 13253 8713 13724 8719
rect 13253 8287 13256 8713
rect 13273 8665 13724 8713
rect 13273 8335 13335 8665
rect 13665 8335 13724 8665
rect 13273 8287 13724 8335
rect 13253 8281 13724 8287
rect -474 8276 -26 8281
rect 76 8276 524 8281
rect 626 8276 1074 8281
rect 1176 8276 1624 8281
rect 1726 8276 2174 8281
rect 2276 8276 2724 8281
rect 2826 8276 3274 8281
rect 3376 8276 3824 8281
rect 3926 8276 4374 8281
rect 4476 8276 4924 8281
rect 5026 8276 5474 8281
rect 5576 8276 6024 8281
rect 6126 8276 6574 8281
rect 6676 8276 7124 8281
rect 7226 8276 7674 8281
rect 7776 8276 8224 8281
rect 8326 8276 8774 8281
rect 8876 8276 9324 8281
rect 9426 8276 9874 8281
rect 9976 8276 10424 8281
rect 10526 8276 10974 8281
rect 11076 8276 11524 8281
rect 11626 8276 12074 8281
rect 12176 8276 12624 8281
rect 12726 8276 13174 8281
rect 13276 8276 13724 8281
rect -1025 8250 -725 8269
rect -469 8273 -31 8276
rect -469 8256 -463 8273
rect -37 8256 -31 8273
rect -469 8253 -31 8256
rect 81 8273 519 8276
rect 81 8256 87 8273
rect 513 8256 519 8273
rect 81 8253 519 8256
rect 631 8273 1069 8276
rect 631 8256 637 8273
rect 1063 8256 1069 8273
rect 631 8253 1069 8256
rect 1181 8273 1619 8276
rect 1181 8256 1187 8273
rect 1613 8256 1619 8273
rect 1181 8253 1619 8256
rect 1731 8273 2169 8276
rect 1731 8256 1737 8273
rect 2163 8256 2169 8273
rect 1731 8253 2169 8256
rect 2281 8273 2719 8276
rect 2281 8256 2287 8273
rect 2713 8256 2719 8273
rect 2281 8253 2719 8256
rect 2831 8273 3269 8276
rect 2831 8256 2837 8273
rect 3263 8256 3269 8273
rect 2831 8253 3269 8256
rect 3381 8273 3819 8276
rect 3381 8256 3387 8273
rect 3813 8256 3819 8273
rect 3381 8253 3819 8256
rect 3931 8273 4369 8276
rect 3931 8256 3937 8273
rect 4363 8256 4369 8273
rect 3931 8253 4369 8256
rect 4481 8273 4919 8276
rect 4481 8256 4487 8273
rect 4913 8256 4919 8273
rect 4481 8253 4919 8256
rect 5031 8273 5469 8276
rect 5031 8256 5037 8273
rect 5463 8256 5469 8273
rect 5031 8253 5469 8256
rect 5581 8273 6019 8276
rect 5581 8256 5587 8273
rect 6013 8256 6019 8273
rect 5581 8253 6019 8256
rect 6131 8273 6569 8276
rect 6131 8256 6137 8273
rect 6563 8256 6569 8273
rect 6131 8253 6569 8256
rect 6681 8273 7119 8276
rect 6681 8256 6687 8273
rect 7113 8256 7119 8273
rect 6681 8253 7119 8256
rect 7231 8273 7669 8276
rect 7231 8256 7237 8273
rect 7663 8256 7669 8273
rect 7231 8253 7669 8256
rect 7781 8273 8219 8276
rect 7781 8256 7787 8273
rect 8213 8256 8219 8273
rect 7781 8253 8219 8256
rect 8331 8273 8769 8276
rect 8331 8256 8337 8273
rect 8763 8256 8769 8273
rect 8331 8253 8769 8256
rect 8881 8273 9319 8276
rect 8881 8256 8887 8273
rect 9313 8256 9319 8273
rect 8881 8253 9319 8256
rect 9431 8273 9869 8276
rect 9431 8256 9437 8273
rect 9863 8256 9869 8273
rect 9431 8253 9869 8256
rect 9981 8273 10419 8276
rect 9981 8256 9987 8273
rect 10413 8256 10419 8273
rect 9981 8253 10419 8256
rect 10531 8273 10969 8276
rect 10531 8256 10537 8273
rect 10963 8256 10969 8273
rect 10531 8253 10969 8256
rect 11081 8273 11519 8276
rect 11081 8256 11087 8273
rect 11513 8256 11519 8273
rect 11081 8253 11519 8256
rect 11631 8273 12069 8276
rect 11631 8256 11637 8273
rect 12063 8256 12069 8273
rect 11631 8253 12069 8256
rect 12181 8273 12619 8276
rect 12181 8256 12187 8273
rect 12613 8256 12619 8273
rect 12181 8253 12619 8256
rect 12731 8273 13169 8276
rect 12731 8256 12737 8273
rect 13163 8256 13169 8273
rect 12731 8253 13169 8256
rect 13281 8273 13719 8276
rect 13281 8256 13287 8273
rect 13713 8256 13719 8273
rect 13281 8253 13719 8256
rect 13975 8269 13987 8800
rect 14263 8269 14275 8800
rect 13975 8250 14275 8269
rect -1025 7719 -1013 8250
rect -737 7719 -725 8250
rect -550 8242 -500 8250
rect -550 8208 -542 8242
rect -508 8208 -500 8242
rect -550 8200 -500 8208
rect 0 8242 50 8250
rect 0 8208 8 8242
rect 42 8208 50 8242
rect 0 8200 50 8208
rect 550 8242 600 8250
rect 550 8208 558 8242
rect 592 8208 600 8242
rect 550 8200 600 8208
rect 1100 8242 1150 8250
rect 1100 8208 1108 8242
rect 1142 8208 1150 8242
rect 1100 8200 1150 8208
rect 1650 8242 1700 8250
rect 1650 8208 1658 8242
rect 1692 8208 1700 8242
rect 1650 8200 1700 8208
rect 2200 8242 2250 8250
rect 2200 8208 2208 8242
rect 2242 8208 2250 8242
rect 2200 8200 2250 8208
rect 2750 8242 2800 8250
rect 2750 8208 2758 8242
rect 2792 8208 2800 8242
rect 2750 8200 2800 8208
rect 3300 8242 3350 8250
rect 3300 8208 3308 8242
rect 3342 8208 3350 8242
rect 3300 8200 3350 8208
rect 3850 8242 3900 8250
rect 3850 8208 3858 8242
rect 3892 8208 3900 8242
rect 3850 8200 3900 8208
rect 4400 8242 4450 8250
rect 4400 8208 4408 8242
rect 4442 8208 4450 8242
rect 4400 8200 4450 8208
rect 4950 8242 5000 8250
rect 4950 8208 4958 8242
rect 4992 8208 5000 8242
rect 4950 8200 5000 8208
rect 5500 8242 5550 8250
rect 5500 8208 5508 8242
rect 5542 8208 5550 8242
rect 5500 8200 5550 8208
rect 6050 8242 6100 8250
rect 6050 8208 6058 8242
rect 6092 8208 6100 8242
rect 6050 8200 6100 8208
rect 6600 8242 6650 8250
rect 6600 8208 6608 8242
rect 6642 8208 6650 8242
rect 6600 8200 6650 8208
rect 7150 8242 7200 8250
rect 7150 8208 7158 8242
rect 7192 8208 7200 8242
rect 7150 8200 7200 8208
rect 7700 8242 7750 8250
rect 7700 8208 7708 8242
rect 7742 8208 7750 8242
rect 7700 8200 7750 8208
rect 8250 8242 8300 8250
rect 8250 8208 8258 8242
rect 8292 8208 8300 8242
rect 8250 8200 8300 8208
rect 8800 8242 8850 8250
rect 8800 8208 8808 8242
rect 8842 8208 8850 8242
rect 8800 8200 8850 8208
rect 9350 8242 9400 8250
rect 9350 8208 9358 8242
rect 9392 8208 9400 8242
rect 9350 8200 9400 8208
rect 9900 8242 9950 8250
rect 9900 8208 9908 8242
rect 9942 8208 9950 8242
rect 9900 8200 9950 8208
rect 10450 8242 10500 8250
rect 10450 8208 10458 8242
rect 10492 8208 10500 8242
rect 10450 8200 10500 8208
rect 11000 8242 11050 8250
rect 11000 8208 11008 8242
rect 11042 8208 11050 8242
rect 11000 8200 11050 8208
rect 11550 8242 11600 8250
rect 11550 8208 11558 8242
rect 11592 8208 11600 8242
rect 11550 8200 11600 8208
rect 12100 8242 12150 8250
rect 12100 8208 12108 8242
rect 12142 8208 12150 8242
rect 12100 8200 12150 8208
rect 12650 8242 12700 8250
rect 12650 8208 12658 8242
rect 12692 8208 12700 8242
rect 12650 8200 12700 8208
rect 13200 8242 13250 8250
rect 13200 8208 13208 8242
rect 13242 8208 13250 8242
rect 13200 8200 13250 8208
rect 13750 8242 13800 8250
rect 13750 8208 13758 8242
rect 13792 8208 13800 8242
rect 13750 8200 13800 8208
rect -469 8194 -31 8197
rect -469 8177 -463 8194
rect -37 8177 -31 8194
rect -469 8174 -31 8177
rect 81 8194 519 8197
rect 81 8177 87 8194
rect 513 8177 519 8194
rect 81 8174 519 8177
rect 631 8194 1069 8197
rect 631 8177 637 8194
rect 1063 8177 1069 8194
rect 631 8174 1069 8177
rect 1181 8194 1619 8197
rect 1181 8177 1187 8194
rect 1613 8177 1619 8194
rect 1181 8174 1619 8177
rect 1731 8194 2169 8197
rect 1731 8177 1737 8194
rect 2163 8177 2169 8194
rect 1731 8174 2169 8177
rect 2281 8194 2719 8197
rect 2281 8177 2287 8194
rect 2713 8177 2719 8194
rect 2281 8174 2719 8177
rect 2831 8194 3269 8197
rect 2831 8177 2837 8194
rect 3263 8177 3269 8194
rect 2831 8174 3269 8177
rect 3381 8194 3819 8197
rect 3381 8177 3387 8194
rect 3813 8177 3819 8194
rect 3381 8174 3819 8177
rect 3931 8194 4369 8197
rect 3931 8177 3937 8194
rect 4363 8177 4369 8194
rect 3931 8174 4369 8177
rect 4481 8194 4919 8197
rect 4481 8177 4487 8194
rect 4913 8177 4919 8194
rect 4481 8174 4919 8177
rect 5031 8194 5469 8197
rect 5031 8177 5037 8194
rect 5463 8177 5469 8194
rect 5031 8174 5469 8177
rect 5581 8194 6019 8197
rect 5581 8177 5587 8194
rect 6013 8177 6019 8194
rect 5581 8174 6019 8177
rect 6131 8194 6569 8197
rect 6131 8177 6137 8194
rect 6563 8177 6569 8194
rect 6131 8174 6569 8177
rect 6681 8194 7119 8197
rect 6681 8177 6687 8194
rect 7113 8177 7119 8194
rect 6681 8174 7119 8177
rect 7231 8194 7669 8197
rect 7231 8177 7237 8194
rect 7663 8177 7669 8194
rect 7231 8174 7669 8177
rect 7781 8194 8219 8197
rect 7781 8177 7787 8194
rect 8213 8177 8219 8194
rect 7781 8174 8219 8177
rect 8331 8194 8769 8197
rect 8331 8177 8337 8194
rect 8763 8177 8769 8194
rect 8331 8174 8769 8177
rect 8881 8194 9319 8197
rect 8881 8177 8887 8194
rect 9313 8177 9319 8194
rect 8881 8174 9319 8177
rect 9431 8194 9869 8197
rect 9431 8177 9437 8194
rect 9863 8177 9869 8194
rect 9431 8174 9869 8177
rect 9981 8194 10419 8197
rect 9981 8177 9987 8194
rect 10413 8177 10419 8194
rect 9981 8174 10419 8177
rect 10531 8194 10969 8197
rect 10531 8177 10537 8194
rect 10963 8177 10969 8194
rect 10531 8174 10969 8177
rect 11081 8194 11519 8197
rect 11081 8177 11087 8194
rect 11513 8177 11519 8194
rect 11081 8174 11519 8177
rect 11631 8194 12069 8197
rect 11631 8177 11637 8194
rect 12063 8177 12069 8194
rect 11631 8174 12069 8177
rect 12181 8194 12619 8197
rect 12181 8177 12187 8194
rect 12613 8177 12619 8194
rect 12181 8174 12619 8177
rect 12731 8194 13169 8197
rect 12731 8177 12737 8194
rect 13163 8177 13169 8194
rect 12731 8174 13169 8177
rect 13281 8194 13719 8197
rect 13281 8177 13287 8194
rect 13713 8177 13719 8194
rect 13281 8174 13719 8177
rect -474 8169 -26 8174
rect 76 8169 524 8174
rect 626 8169 1074 8174
rect 1176 8169 1624 8174
rect 1726 8169 2174 8174
rect 2276 8169 2724 8174
rect 2826 8169 3274 8174
rect 3376 8169 3824 8174
rect 3926 8169 4374 8174
rect 4476 8169 4924 8174
rect 5026 8169 5474 8174
rect 5576 8169 6024 8174
rect 6126 8169 6574 8174
rect 6676 8169 7124 8174
rect 7226 8169 7674 8174
rect 7776 8169 8224 8174
rect 8326 8169 8774 8174
rect 8876 8169 9324 8174
rect 9426 8169 9874 8174
rect 9976 8169 10424 8174
rect 10526 8169 10974 8174
rect 11076 8169 11524 8174
rect 11626 8169 12074 8174
rect 12176 8169 12624 8174
rect 12726 8169 13174 8174
rect 13276 8169 13724 8174
rect -474 8163 -3 8169
rect -474 8115 -23 8163
rect -474 7785 -415 8115
rect -85 7785 -23 8115
rect -474 7737 -23 7785
rect -6 7737 -3 8163
rect -474 7731 -3 7737
rect 53 8163 547 8169
rect 53 7737 56 8163
rect 73 8115 527 8163
rect 73 7785 135 8115
rect 465 7785 527 8115
rect 73 7737 527 7785
rect 544 7737 547 8163
rect 53 7731 547 7737
rect 603 8163 1097 8169
rect 603 7737 606 8163
rect 623 8115 1077 8163
rect 623 7785 685 8115
rect 1015 7785 1077 8115
rect 623 7737 1077 7785
rect 1094 7737 1097 8163
rect 603 7731 1097 7737
rect 1153 8163 1647 8169
rect 1153 7737 1156 8163
rect 1173 8115 1627 8163
rect 1173 7785 1235 8115
rect 1565 7785 1627 8115
rect 1173 7737 1627 7785
rect 1644 7737 1647 8163
rect 1153 7731 1647 7737
rect 1703 8163 2197 8169
rect 1703 7737 1706 8163
rect 1723 8115 2177 8163
rect 1723 7785 1785 8115
rect 2115 7785 2177 8115
rect 1723 7737 2177 7785
rect 2194 7737 2197 8163
rect 1703 7731 2197 7737
rect 2253 8163 2747 8169
rect 2253 7737 2256 8163
rect 2273 8115 2727 8163
rect 2273 7785 2335 8115
rect 2665 7785 2727 8115
rect 2273 7737 2727 7785
rect 2744 7737 2747 8163
rect 2253 7731 2747 7737
rect 2803 8163 3297 8169
rect 2803 7737 2806 8163
rect 2823 8115 3277 8163
rect 2823 7785 2885 8115
rect 3215 7785 3277 8115
rect 2823 7737 3277 7785
rect 3294 7737 3297 8163
rect 2803 7731 3297 7737
rect 3353 8163 3847 8169
rect 3353 7737 3356 8163
rect 3373 8115 3827 8163
rect 3373 7785 3435 8115
rect 3765 7785 3827 8115
rect 3373 7737 3827 7785
rect 3844 7737 3847 8163
rect 3353 7731 3847 7737
rect 3903 8163 4397 8169
rect 3903 7737 3906 8163
rect 3923 8115 4377 8163
rect 3923 7785 3985 8115
rect 4315 7785 4377 8115
rect 3923 7737 4377 7785
rect 4394 7737 4397 8163
rect 3903 7731 4397 7737
rect 4453 8163 4947 8169
rect 4453 7737 4456 8163
rect 4473 8115 4927 8163
rect 4473 7785 4535 8115
rect 4865 7785 4927 8115
rect 4473 7737 4927 7785
rect 4944 7737 4947 8163
rect 4453 7731 4947 7737
rect 5003 8163 5497 8169
rect 5003 7737 5006 8163
rect 5023 8115 5477 8163
rect 5023 7785 5085 8115
rect 5415 7785 5477 8115
rect 5023 7737 5477 7785
rect 5494 7737 5497 8163
rect 5003 7731 5497 7737
rect 5553 8163 6047 8169
rect 5553 7737 5556 8163
rect 5573 8115 6027 8163
rect 5573 7785 5635 8115
rect 5965 7785 6027 8115
rect 5573 7737 6027 7785
rect 6044 7737 6047 8163
rect 5553 7731 6047 7737
rect 6103 8163 6597 8169
rect 6103 7737 6106 8163
rect 6123 8115 6577 8163
rect 6123 7785 6185 8115
rect 6515 7785 6577 8115
rect 6123 7737 6577 7785
rect 6594 7737 6597 8163
rect 6103 7731 6597 7737
rect 6653 8163 7147 8169
rect 6653 7737 6656 8163
rect 6673 8115 7127 8163
rect 6673 7785 6735 8115
rect 7065 7785 7127 8115
rect 6673 7737 7127 7785
rect 7144 7737 7147 8163
rect 6653 7731 7147 7737
rect 7203 8163 7697 8169
rect 7203 7737 7206 8163
rect 7223 8115 7677 8163
rect 7223 7785 7285 8115
rect 7615 7785 7677 8115
rect 7223 7737 7677 7785
rect 7694 7737 7697 8163
rect 7203 7731 7697 7737
rect 7753 8163 8247 8169
rect 7753 7737 7756 8163
rect 7773 8115 8227 8163
rect 7773 7785 7835 8115
rect 8165 7785 8227 8115
rect 7773 7737 8227 7785
rect 8244 7737 8247 8163
rect 7753 7731 8247 7737
rect 8303 8163 8797 8169
rect 8303 7737 8306 8163
rect 8323 8115 8777 8163
rect 8323 7785 8385 8115
rect 8715 7785 8777 8115
rect 8323 7737 8777 7785
rect 8794 7737 8797 8163
rect 8303 7731 8797 7737
rect 8853 8163 9347 8169
rect 8853 7737 8856 8163
rect 8873 8115 9327 8163
rect 8873 7785 8935 8115
rect 9265 7785 9327 8115
rect 8873 7737 9327 7785
rect 9344 7737 9347 8163
rect 8853 7731 9347 7737
rect 9403 8163 9897 8169
rect 9403 7737 9406 8163
rect 9423 8115 9877 8163
rect 9423 7785 9485 8115
rect 9815 7785 9877 8115
rect 9423 7737 9877 7785
rect 9894 7737 9897 8163
rect 9403 7731 9897 7737
rect 9953 8163 10447 8169
rect 9953 7737 9956 8163
rect 9973 8115 10427 8163
rect 9973 7785 10035 8115
rect 10365 7785 10427 8115
rect 9973 7737 10427 7785
rect 10444 7737 10447 8163
rect 9953 7731 10447 7737
rect 10503 8163 10997 8169
rect 10503 7737 10506 8163
rect 10523 8115 10977 8163
rect 10523 7785 10585 8115
rect 10915 7785 10977 8115
rect 10523 7737 10977 7785
rect 10994 7737 10997 8163
rect 10503 7731 10997 7737
rect 11053 8163 11547 8169
rect 11053 7737 11056 8163
rect 11073 8115 11527 8163
rect 11073 7785 11135 8115
rect 11465 7785 11527 8115
rect 11073 7737 11527 7785
rect 11544 7737 11547 8163
rect 11053 7731 11547 7737
rect 11603 8163 12097 8169
rect 11603 7737 11606 8163
rect 11623 8115 12077 8163
rect 11623 7785 11685 8115
rect 12015 7785 12077 8115
rect 11623 7737 12077 7785
rect 12094 7737 12097 8163
rect 11603 7731 12097 7737
rect 12153 8163 12647 8169
rect 12153 7737 12156 8163
rect 12173 8115 12627 8163
rect 12173 7785 12235 8115
rect 12565 7785 12627 8115
rect 12173 7737 12627 7785
rect 12644 7737 12647 8163
rect 12153 7731 12647 7737
rect 12703 8163 13197 8169
rect 12703 7737 12706 8163
rect 12723 8115 13177 8163
rect 12723 7785 12785 8115
rect 13115 7785 13177 8115
rect 12723 7737 13177 7785
rect 13194 7737 13197 8163
rect 12703 7731 13197 7737
rect 13253 8163 13724 8169
rect 13253 7737 13256 8163
rect 13273 8115 13724 8163
rect 13273 7785 13335 8115
rect 13665 7785 13724 8115
rect 13273 7737 13724 7785
rect 13253 7731 13724 7737
rect -474 7726 -26 7731
rect 76 7726 524 7731
rect 626 7726 1074 7731
rect 1176 7726 1624 7731
rect 1726 7726 2174 7731
rect 2276 7726 2724 7731
rect 2826 7726 3274 7731
rect 3376 7726 3824 7731
rect 3926 7726 4374 7731
rect 4476 7726 4924 7731
rect 5026 7726 5474 7731
rect 5576 7726 6024 7731
rect 6126 7726 6574 7731
rect 6676 7726 7124 7731
rect 7226 7726 7674 7731
rect 7776 7726 8224 7731
rect 8326 7726 8774 7731
rect 8876 7726 9324 7731
rect 9426 7726 9874 7731
rect 9976 7726 10424 7731
rect 10526 7726 10974 7731
rect 11076 7726 11524 7731
rect 11626 7726 12074 7731
rect 12176 7726 12624 7731
rect 12726 7726 13174 7731
rect 13276 7726 13724 7731
rect -1025 7700 -725 7719
rect -469 7723 -31 7726
rect -469 7706 -463 7723
rect -37 7706 -31 7723
rect -469 7703 -31 7706
rect 81 7723 519 7726
rect 81 7706 87 7723
rect 513 7706 519 7723
rect 81 7703 519 7706
rect 631 7723 1069 7726
rect 631 7706 637 7723
rect 1063 7706 1069 7723
rect 631 7703 1069 7706
rect 1181 7723 1619 7726
rect 1181 7706 1187 7723
rect 1613 7706 1619 7723
rect 1181 7703 1619 7706
rect 1731 7723 2169 7726
rect 1731 7706 1737 7723
rect 2163 7706 2169 7723
rect 1731 7703 2169 7706
rect 2281 7723 2719 7726
rect 2281 7706 2287 7723
rect 2713 7706 2719 7723
rect 2281 7703 2719 7706
rect 2831 7723 3269 7726
rect 2831 7706 2837 7723
rect 3263 7706 3269 7723
rect 2831 7703 3269 7706
rect 3381 7723 3819 7726
rect 3381 7706 3387 7723
rect 3813 7706 3819 7723
rect 3381 7703 3819 7706
rect 3931 7723 4369 7726
rect 3931 7706 3937 7723
rect 4363 7706 4369 7723
rect 3931 7703 4369 7706
rect 4481 7723 4919 7726
rect 4481 7706 4487 7723
rect 4913 7706 4919 7723
rect 4481 7703 4919 7706
rect 5031 7723 5469 7726
rect 5031 7706 5037 7723
rect 5463 7706 5469 7723
rect 5031 7703 5469 7706
rect 5581 7723 6019 7726
rect 5581 7706 5587 7723
rect 6013 7706 6019 7723
rect 5581 7703 6019 7706
rect 6131 7723 6569 7726
rect 6131 7706 6137 7723
rect 6563 7706 6569 7723
rect 6131 7703 6569 7706
rect 6681 7723 7119 7726
rect 6681 7706 6687 7723
rect 7113 7706 7119 7723
rect 6681 7703 7119 7706
rect 7231 7723 7669 7726
rect 7231 7706 7237 7723
rect 7663 7706 7669 7723
rect 7231 7703 7669 7706
rect 7781 7723 8219 7726
rect 7781 7706 7787 7723
rect 8213 7706 8219 7723
rect 7781 7703 8219 7706
rect 8331 7723 8769 7726
rect 8331 7706 8337 7723
rect 8763 7706 8769 7723
rect 8331 7703 8769 7706
rect 8881 7723 9319 7726
rect 8881 7706 8887 7723
rect 9313 7706 9319 7723
rect 8881 7703 9319 7706
rect 9431 7723 9869 7726
rect 9431 7706 9437 7723
rect 9863 7706 9869 7723
rect 9431 7703 9869 7706
rect 9981 7723 10419 7726
rect 9981 7706 9987 7723
rect 10413 7706 10419 7723
rect 9981 7703 10419 7706
rect 10531 7723 10969 7726
rect 10531 7706 10537 7723
rect 10963 7706 10969 7723
rect 10531 7703 10969 7706
rect 11081 7723 11519 7726
rect 11081 7706 11087 7723
rect 11513 7706 11519 7723
rect 11081 7703 11519 7706
rect 11631 7723 12069 7726
rect 11631 7706 11637 7723
rect 12063 7706 12069 7723
rect 11631 7703 12069 7706
rect 12181 7723 12619 7726
rect 12181 7706 12187 7723
rect 12613 7706 12619 7723
rect 12181 7703 12619 7706
rect 12731 7723 13169 7726
rect 12731 7706 12737 7723
rect 13163 7706 13169 7723
rect 12731 7703 13169 7706
rect 13281 7723 13719 7726
rect 13281 7706 13287 7723
rect 13713 7706 13719 7723
rect 13281 7703 13719 7706
rect 13975 7719 13987 8250
rect 14263 7719 14275 8250
rect 13975 7700 14275 7719
rect -1025 7169 -1013 7700
rect -737 7169 -725 7700
rect -550 7692 -500 7700
rect -550 7658 -542 7692
rect -508 7658 -500 7692
rect -550 7650 -500 7658
rect 0 7692 50 7700
rect 0 7658 8 7692
rect 42 7658 50 7692
rect 0 7650 50 7658
rect 550 7692 600 7700
rect 550 7658 558 7692
rect 592 7658 600 7692
rect 550 7650 600 7658
rect 1100 7692 1150 7700
rect 1100 7658 1108 7692
rect 1142 7658 1150 7692
rect 1100 7650 1150 7658
rect 1650 7692 1700 7700
rect 1650 7658 1658 7692
rect 1692 7658 1700 7692
rect 1650 7650 1700 7658
rect 2200 7692 2250 7700
rect 2200 7658 2208 7692
rect 2242 7658 2250 7692
rect 2200 7650 2250 7658
rect 2750 7692 2800 7700
rect 2750 7658 2758 7692
rect 2792 7658 2800 7692
rect 2750 7650 2800 7658
rect 3300 7692 3350 7700
rect 3300 7658 3308 7692
rect 3342 7658 3350 7692
rect 3300 7650 3350 7658
rect 3850 7692 3900 7700
rect 3850 7658 3858 7692
rect 3892 7658 3900 7692
rect 3850 7650 3900 7658
rect 4400 7692 4450 7700
rect 4400 7658 4408 7692
rect 4442 7658 4450 7692
rect 4400 7650 4450 7658
rect 4950 7692 5000 7700
rect 4950 7658 4958 7692
rect 4992 7658 5000 7692
rect 4950 7650 5000 7658
rect 5500 7692 5550 7700
rect 5500 7658 5508 7692
rect 5542 7658 5550 7692
rect 5500 7650 5550 7658
rect 6050 7692 6100 7700
rect 6050 7658 6058 7692
rect 6092 7658 6100 7692
rect 6050 7650 6100 7658
rect 6600 7692 6650 7700
rect 6600 7658 6608 7692
rect 6642 7658 6650 7692
rect 6600 7650 6650 7658
rect 7150 7692 7200 7700
rect 7150 7658 7158 7692
rect 7192 7658 7200 7692
rect 7150 7650 7200 7658
rect 7700 7692 7750 7700
rect 7700 7658 7708 7692
rect 7742 7658 7750 7692
rect 7700 7650 7750 7658
rect 8250 7692 8300 7700
rect 8250 7658 8258 7692
rect 8292 7658 8300 7692
rect 8250 7650 8300 7658
rect 8800 7692 8850 7700
rect 8800 7658 8808 7692
rect 8842 7658 8850 7692
rect 8800 7650 8850 7658
rect 9350 7692 9400 7700
rect 9350 7658 9358 7692
rect 9392 7658 9400 7692
rect 9350 7650 9400 7658
rect 9900 7692 9950 7700
rect 9900 7658 9908 7692
rect 9942 7658 9950 7692
rect 9900 7650 9950 7658
rect 10450 7692 10500 7700
rect 10450 7658 10458 7692
rect 10492 7658 10500 7692
rect 10450 7650 10500 7658
rect 11000 7692 11050 7700
rect 11000 7658 11008 7692
rect 11042 7658 11050 7692
rect 11000 7650 11050 7658
rect 11550 7692 11600 7700
rect 11550 7658 11558 7692
rect 11592 7658 11600 7692
rect 11550 7650 11600 7658
rect 12100 7692 12150 7700
rect 12100 7658 12108 7692
rect 12142 7658 12150 7692
rect 12100 7650 12150 7658
rect 12650 7692 12700 7700
rect 12650 7658 12658 7692
rect 12692 7658 12700 7692
rect 12650 7650 12700 7658
rect 13200 7692 13250 7700
rect 13200 7658 13208 7692
rect 13242 7658 13250 7692
rect 13200 7650 13250 7658
rect 13750 7692 13800 7700
rect 13750 7658 13758 7692
rect 13792 7658 13800 7692
rect 13750 7650 13800 7658
rect -469 7644 -31 7647
rect -469 7627 -463 7644
rect -37 7627 -31 7644
rect -469 7624 -31 7627
rect 81 7644 519 7647
rect 81 7627 87 7644
rect 513 7627 519 7644
rect 81 7624 519 7627
rect 631 7644 1069 7647
rect 631 7627 637 7644
rect 1063 7627 1069 7644
rect 631 7624 1069 7627
rect 1181 7644 1619 7647
rect 1181 7627 1187 7644
rect 1613 7627 1619 7644
rect 1181 7624 1619 7627
rect 1731 7644 2169 7647
rect 1731 7627 1737 7644
rect 2163 7627 2169 7644
rect 1731 7624 2169 7627
rect 2281 7644 2719 7647
rect 2281 7627 2287 7644
rect 2713 7627 2719 7644
rect 2281 7624 2719 7627
rect 2831 7644 3269 7647
rect 2831 7627 2837 7644
rect 3263 7627 3269 7644
rect 2831 7624 3269 7627
rect 3381 7644 3819 7647
rect 3381 7627 3387 7644
rect 3813 7627 3819 7644
rect 3381 7624 3819 7627
rect 3931 7644 4369 7647
rect 3931 7627 3937 7644
rect 4363 7627 4369 7644
rect 3931 7624 4369 7627
rect 4481 7644 4919 7647
rect 4481 7627 4487 7644
rect 4913 7627 4919 7644
rect 4481 7624 4919 7627
rect 5031 7644 5469 7647
rect 5031 7627 5037 7644
rect 5463 7627 5469 7644
rect 5031 7624 5469 7627
rect 5581 7644 6019 7647
rect 5581 7627 5587 7644
rect 6013 7627 6019 7644
rect 5581 7624 6019 7627
rect 6131 7644 6569 7647
rect 6131 7627 6137 7644
rect 6563 7627 6569 7644
rect 6131 7624 6569 7627
rect 6681 7644 7119 7647
rect 6681 7627 6687 7644
rect 7113 7627 7119 7644
rect 6681 7624 7119 7627
rect 7231 7644 7669 7647
rect 7231 7627 7237 7644
rect 7663 7627 7669 7644
rect 7231 7624 7669 7627
rect 7781 7644 8219 7647
rect 7781 7627 7787 7644
rect 8213 7627 8219 7644
rect 7781 7624 8219 7627
rect 8331 7644 8769 7647
rect 8331 7627 8337 7644
rect 8763 7627 8769 7644
rect 8331 7624 8769 7627
rect 8881 7644 9319 7647
rect 8881 7627 8887 7644
rect 9313 7627 9319 7644
rect 8881 7624 9319 7627
rect 9431 7644 9869 7647
rect 9431 7627 9437 7644
rect 9863 7627 9869 7644
rect 9431 7624 9869 7627
rect 9981 7644 10419 7647
rect 9981 7627 9987 7644
rect 10413 7627 10419 7644
rect 9981 7624 10419 7627
rect 10531 7644 10969 7647
rect 10531 7627 10537 7644
rect 10963 7627 10969 7644
rect 10531 7624 10969 7627
rect 11081 7644 11519 7647
rect 11081 7627 11087 7644
rect 11513 7627 11519 7644
rect 11081 7624 11519 7627
rect 11631 7644 12069 7647
rect 11631 7627 11637 7644
rect 12063 7627 12069 7644
rect 11631 7624 12069 7627
rect 12181 7644 12619 7647
rect 12181 7627 12187 7644
rect 12613 7627 12619 7644
rect 12181 7624 12619 7627
rect 12731 7644 13169 7647
rect 12731 7627 12737 7644
rect 13163 7627 13169 7644
rect 12731 7624 13169 7627
rect 13281 7644 13719 7647
rect 13281 7627 13287 7644
rect 13713 7627 13719 7644
rect 13281 7624 13719 7627
rect -474 7619 -26 7624
rect 76 7619 524 7624
rect 626 7619 1074 7624
rect 1176 7619 1624 7624
rect 1726 7619 2174 7624
rect 2276 7619 2724 7624
rect 2826 7619 3274 7624
rect 3376 7619 3824 7624
rect 3926 7619 4374 7624
rect 4476 7619 4924 7624
rect 5026 7619 5474 7624
rect 5576 7619 6024 7624
rect 6126 7619 6574 7624
rect 6676 7619 7124 7624
rect 7226 7619 7674 7624
rect 7776 7619 8224 7624
rect 8326 7619 8774 7624
rect 8876 7619 9324 7624
rect 9426 7619 9874 7624
rect 9976 7619 10424 7624
rect 10526 7619 10974 7624
rect 11076 7619 11524 7624
rect 11626 7619 12074 7624
rect 12176 7619 12624 7624
rect 12726 7619 13174 7624
rect 13276 7619 13724 7624
rect -474 7613 -3 7619
rect -474 7565 -23 7613
rect -474 7235 -415 7565
rect -85 7235 -23 7565
rect -474 7187 -23 7235
rect -6 7187 -3 7613
rect -474 7181 -3 7187
rect 53 7613 547 7619
rect 53 7187 56 7613
rect 73 7565 527 7613
rect 73 7235 135 7565
rect 465 7235 527 7565
rect 73 7187 527 7235
rect 544 7187 547 7613
rect 53 7181 547 7187
rect 603 7613 1097 7619
rect 603 7187 606 7613
rect 623 7565 1077 7613
rect 623 7235 685 7565
rect 1015 7235 1077 7565
rect 623 7187 1077 7235
rect 1094 7187 1097 7613
rect 603 7181 1097 7187
rect 1153 7613 1647 7619
rect 1153 7187 1156 7613
rect 1173 7565 1627 7613
rect 1173 7235 1235 7565
rect 1565 7235 1627 7565
rect 1173 7187 1627 7235
rect 1644 7187 1647 7613
rect 1153 7181 1647 7187
rect 1703 7613 2197 7619
rect 1703 7187 1706 7613
rect 1723 7565 2177 7613
rect 1723 7235 1785 7565
rect 2115 7235 2177 7565
rect 1723 7187 2177 7235
rect 2194 7187 2197 7613
rect 1703 7181 2197 7187
rect 2253 7613 2747 7619
rect 2253 7187 2256 7613
rect 2273 7565 2727 7613
rect 2273 7235 2335 7565
rect 2665 7235 2727 7565
rect 2273 7187 2727 7235
rect 2744 7187 2747 7613
rect 2253 7181 2747 7187
rect 2803 7613 3297 7619
rect 2803 7187 2806 7613
rect 2823 7565 3277 7613
rect 2823 7235 2885 7565
rect 3215 7235 3277 7565
rect 2823 7187 3277 7235
rect 3294 7187 3297 7613
rect 2803 7181 3297 7187
rect 3353 7613 3847 7619
rect 3353 7187 3356 7613
rect 3373 7565 3827 7613
rect 3373 7235 3435 7565
rect 3765 7235 3827 7565
rect 3373 7187 3827 7235
rect 3844 7187 3847 7613
rect 3353 7181 3847 7187
rect 3903 7613 4397 7619
rect 3903 7187 3906 7613
rect 3923 7565 4377 7613
rect 3923 7235 3985 7565
rect 4315 7235 4377 7565
rect 3923 7187 4377 7235
rect 4394 7187 4397 7613
rect 3903 7181 4397 7187
rect 4453 7613 4947 7619
rect 4453 7187 4456 7613
rect 4473 7565 4927 7613
rect 4473 7235 4535 7565
rect 4865 7235 4927 7565
rect 4473 7187 4927 7235
rect 4944 7187 4947 7613
rect 4453 7181 4947 7187
rect 5003 7613 5497 7619
rect 5003 7187 5006 7613
rect 5023 7565 5477 7613
rect 5023 7235 5085 7565
rect 5415 7235 5477 7565
rect 5023 7187 5477 7235
rect 5494 7187 5497 7613
rect 5003 7181 5497 7187
rect 5553 7613 6047 7619
rect 5553 7187 5556 7613
rect 5573 7565 6027 7613
rect 5573 7235 5635 7565
rect 5965 7235 6027 7565
rect 5573 7187 6027 7235
rect 6044 7187 6047 7613
rect 5553 7181 6047 7187
rect 6103 7613 6597 7619
rect 6103 7187 6106 7613
rect 6123 7565 6577 7613
rect 6123 7235 6185 7565
rect 6515 7235 6577 7565
rect 6123 7187 6577 7235
rect 6594 7187 6597 7613
rect 6103 7181 6597 7187
rect 6653 7613 7147 7619
rect 6653 7187 6656 7613
rect 6673 7565 7127 7613
rect 6673 7235 6735 7565
rect 7065 7235 7127 7565
rect 6673 7187 7127 7235
rect 7144 7187 7147 7613
rect 6653 7181 7147 7187
rect 7203 7613 7697 7619
rect 7203 7187 7206 7613
rect 7223 7565 7677 7613
rect 7223 7235 7285 7565
rect 7615 7235 7677 7565
rect 7223 7187 7677 7235
rect 7694 7187 7697 7613
rect 7203 7181 7697 7187
rect 7753 7613 8247 7619
rect 7753 7187 7756 7613
rect 7773 7565 8227 7613
rect 7773 7235 7835 7565
rect 8165 7235 8227 7565
rect 7773 7187 8227 7235
rect 8244 7187 8247 7613
rect 7753 7181 8247 7187
rect 8303 7613 8797 7619
rect 8303 7187 8306 7613
rect 8323 7565 8777 7613
rect 8323 7235 8385 7565
rect 8715 7235 8777 7565
rect 8323 7187 8777 7235
rect 8794 7187 8797 7613
rect 8303 7181 8797 7187
rect 8853 7613 9347 7619
rect 8853 7187 8856 7613
rect 8873 7565 9327 7613
rect 8873 7235 8935 7565
rect 9265 7235 9327 7565
rect 8873 7187 9327 7235
rect 9344 7187 9347 7613
rect 8853 7181 9347 7187
rect 9403 7613 9897 7619
rect 9403 7187 9406 7613
rect 9423 7565 9877 7613
rect 9423 7235 9485 7565
rect 9815 7235 9877 7565
rect 9423 7187 9877 7235
rect 9894 7187 9897 7613
rect 9403 7181 9897 7187
rect 9953 7613 10447 7619
rect 9953 7187 9956 7613
rect 9973 7565 10427 7613
rect 9973 7235 10035 7565
rect 10365 7235 10427 7565
rect 9973 7187 10427 7235
rect 10444 7187 10447 7613
rect 9953 7181 10447 7187
rect 10503 7613 10997 7619
rect 10503 7187 10506 7613
rect 10523 7565 10977 7613
rect 10523 7235 10585 7565
rect 10915 7235 10977 7565
rect 10523 7187 10977 7235
rect 10994 7187 10997 7613
rect 10503 7181 10997 7187
rect 11053 7613 11547 7619
rect 11053 7187 11056 7613
rect 11073 7565 11527 7613
rect 11073 7235 11135 7565
rect 11465 7235 11527 7565
rect 11073 7187 11527 7235
rect 11544 7187 11547 7613
rect 11053 7181 11547 7187
rect 11603 7613 12097 7619
rect 11603 7187 11606 7613
rect 11623 7565 12077 7613
rect 11623 7235 11685 7565
rect 12015 7235 12077 7565
rect 11623 7187 12077 7235
rect 12094 7187 12097 7613
rect 11603 7181 12097 7187
rect 12153 7613 12647 7619
rect 12153 7187 12156 7613
rect 12173 7565 12627 7613
rect 12173 7235 12235 7565
rect 12565 7235 12627 7565
rect 12173 7187 12627 7235
rect 12644 7187 12647 7613
rect 12153 7181 12647 7187
rect 12703 7613 13197 7619
rect 12703 7187 12706 7613
rect 12723 7565 13177 7613
rect 12723 7235 12785 7565
rect 13115 7235 13177 7565
rect 12723 7187 13177 7235
rect 13194 7187 13197 7613
rect 12703 7181 13197 7187
rect 13253 7613 13724 7619
rect 13253 7187 13256 7613
rect 13273 7565 13724 7613
rect 13273 7235 13335 7565
rect 13665 7235 13724 7565
rect 13273 7187 13724 7235
rect 13253 7181 13724 7187
rect -474 7176 -26 7181
rect 76 7176 524 7181
rect 626 7176 1074 7181
rect 1176 7176 1624 7181
rect 1726 7176 2174 7181
rect 2276 7176 2724 7181
rect 2826 7176 3274 7181
rect 3376 7176 3824 7181
rect 3926 7176 4374 7181
rect 4476 7176 4924 7181
rect 5026 7176 5474 7181
rect 5576 7176 6024 7181
rect 6126 7176 6574 7181
rect 6676 7176 7124 7181
rect 7226 7176 7674 7181
rect 7776 7176 8224 7181
rect 8326 7176 8774 7181
rect 8876 7176 9324 7181
rect 9426 7176 9874 7181
rect 9976 7176 10424 7181
rect 10526 7176 10974 7181
rect 11076 7176 11524 7181
rect 11626 7176 12074 7181
rect 12176 7176 12624 7181
rect 12726 7176 13174 7181
rect 13276 7176 13724 7181
rect -1025 7150 -725 7169
rect -469 7173 -31 7176
rect -469 7156 -463 7173
rect -37 7156 -31 7173
rect -469 7153 -31 7156
rect 81 7173 519 7176
rect 81 7156 87 7173
rect 513 7156 519 7173
rect 81 7153 519 7156
rect 631 7173 1069 7176
rect 631 7156 637 7173
rect 1063 7156 1069 7173
rect 631 7153 1069 7156
rect 1181 7173 1619 7176
rect 1181 7156 1187 7173
rect 1613 7156 1619 7173
rect 1181 7153 1619 7156
rect 1731 7173 2169 7176
rect 1731 7156 1737 7173
rect 2163 7156 2169 7173
rect 1731 7153 2169 7156
rect 2281 7173 2719 7176
rect 2281 7156 2287 7173
rect 2713 7156 2719 7173
rect 2281 7153 2719 7156
rect 2831 7173 3269 7176
rect 2831 7156 2837 7173
rect 3263 7156 3269 7173
rect 2831 7153 3269 7156
rect 3381 7173 3819 7176
rect 3381 7156 3387 7173
rect 3813 7156 3819 7173
rect 3381 7153 3819 7156
rect 3931 7173 4369 7176
rect 3931 7156 3937 7173
rect 4363 7156 4369 7173
rect 3931 7153 4369 7156
rect 4481 7173 4919 7176
rect 4481 7156 4487 7173
rect 4913 7156 4919 7173
rect 4481 7153 4919 7156
rect 5031 7173 5469 7176
rect 5031 7156 5037 7173
rect 5463 7156 5469 7173
rect 5031 7153 5469 7156
rect 5581 7173 6019 7176
rect 5581 7156 5587 7173
rect 6013 7156 6019 7173
rect 5581 7153 6019 7156
rect 6131 7173 6569 7176
rect 6131 7156 6137 7173
rect 6563 7156 6569 7173
rect 6131 7153 6569 7156
rect 6681 7173 7119 7176
rect 6681 7156 6687 7173
rect 7113 7156 7119 7173
rect 6681 7153 7119 7156
rect 7231 7173 7669 7176
rect 7231 7156 7237 7173
rect 7663 7156 7669 7173
rect 7231 7153 7669 7156
rect 7781 7173 8219 7176
rect 7781 7156 7787 7173
rect 8213 7156 8219 7173
rect 7781 7153 8219 7156
rect 8331 7173 8769 7176
rect 8331 7156 8337 7173
rect 8763 7156 8769 7173
rect 8331 7153 8769 7156
rect 8881 7173 9319 7176
rect 8881 7156 8887 7173
rect 9313 7156 9319 7173
rect 8881 7153 9319 7156
rect 9431 7173 9869 7176
rect 9431 7156 9437 7173
rect 9863 7156 9869 7173
rect 9431 7153 9869 7156
rect 9981 7173 10419 7176
rect 9981 7156 9987 7173
rect 10413 7156 10419 7173
rect 9981 7153 10419 7156
rect 10531 7173 10969 7176
rect 10531 7156 10537 7173
rect 10963 7156 10969 7173
rect 10531 7153 10969 7156
rect 11081 7173 11519 7176
rect 11081 7156 11087 7173
rect 11513 7156 11519 7173
rect 11081 7153 11519 7156
rect 11631 7173 12069 7176
rect 11631 7156 11637 7173
rect 12063 7156 12069 7173
rect 11631 7153 12069 7156
rect 12181 7173 12619 7176
rect 12181 7156 12187 7173
rect 12613 7156 12619 7173
rect 12181 7153 12619 7156
rect 12731 7173 13169 7176
rect 12731 7156 12737 7173
rect 13163 7156 13169 7173
rect 12731 7153 13169 7156
rect 13281 7173 13719 7176
rect 13281 7156 13287 7173
rect 13713 7156 13719 7173
rect 13281 7153 13719 7156
rect 13975 7169 13987 7700
rect 14263 7169 14275 7700
rect 13975 7150 14275 7169
rect -1025 6619 -1013 7150
rect -737 6619 -725 7150
rect -550 7142 -500 7150
rect -550 7108 -542 7142
rect -508 7108 -500 7142
rect -550 7100 -500 7108
rect 0 7142 50 7150
rect 0 7108 8 7142
rect 42 7108 50 7142
rect 0 7100 50 7108
rect 550 7142 600 7150
rect 550 7108 558 7142
rect 592 7108 600 7142
rect 550 7100 600 7108
rect 1100 7142 1150 7150
rect 1100 7108 1108 7142
rect 1142 7108 1150 7142
rect 1100 7100 1150 7108
rect 1650 7142 1700 7150
rect 1650 7108 1658 7142
rect 1692 7108 1700 7142
rect 1650 7100 1700 7108
rect 2200 7142 2250 7150
rect 2200 7108 2208 7142
rect 2242 7108 2250 7142
rect 2200 7100 2250 7108
rect 2750 7142 2800 7150
rect 2750 7108 2758 7142
rect 2792 7108 2800 7142
rect 2750 7100 2800 7108
rect 3300 7142 3350 7150
rect 3300 7108 3308 7142
rect 3342 7108 3350 7142
rect 3300 7100 3350 7108
rect 3850 7142 3900 7150
rect 3850 7108 3858 7142
rect 3892 7108 3900 7142
rect 3850 7100 3900 7108
rect 4400 7142 4450 7150
rect 4400 7108 4408 7142
rect 4442 7108 4450 7142
rect 4400 7100 4450 7108
rect 4950 7142 5000 7150
rect 4950 7108 4958 7142
rect 4992 7108 5000 7142
rect 4950 7100 5000 7108
rect 5500 7142 5550 7150
rect 5500 7108 5508 7142
rect 5542 7108 5550 7142
rect 5500 7100 5550 7108
rect 6050 7142 6100 7150
rect 6050 7108 6058 7142
rect 6092 7108 6100 7142
rect 6050 7100 6100 7108
rect 6600 7142 6650 7150
rect 6600 7108 6608 7142
rect 6642 7108 6650 7142
rect 6600 7100 6650 7108
rect 7150 7142 7200 7150
rect 7150 7108 7158 7142
rect 7192 7108 7200 7142
rect 7150 7100 7200 7108
rect 7700 7142 7750 7150
rect 7700 7108 7708 7142
rect 7742 7108 7750 7142
rect 7700 7100 7750 7108
rect 8250 7142 8300 7150
rect 8250 7108 8258 7142
rect 8292 7108 8300 7142
rect 8250 7100 8300 7108
rect 8800 7142 8850 7150
rect 8800 7108 8808 7142
rect 8842 7108 8850 7142
rect 8800 7100 8850 7108
rect 9350 7142 9400 7150
rect 9350 7108 9358 7142
rect 9392 7108 9400 7142
rect 9350 7100 9400 7108
rect 9900 7142 9950 7150
rect 9900 7108 9908 7142
rect 9942 7108 9950 7142
rect 9900 7100 9950 7108
rect 10450 7142 10500 7150
rect 10450 7108 10458 7142
rect 10492 7108 10500 7142
rect 10450 7100 10500 7108
rect 11000 7142 11050 7150
rect 11000 7108 11008 7142
rect 11042 7108 11050 7142
rect 11000 7100 11050 7108
rect 11550 7142 11600 7150
rect 11550 7108 11558 7142
rect 11592 7108 11600 7142
rect 11550 7100 11600 7108
rect 12100 7142 12150 7150
rect 12100 7108 12108 7142
rect 12142 7108 12150 7142
rect 12100 7100 12150 7108
rect 12650 7142 12700 7150
rect 12650 7108 12658 7142
rect 12692 7108 12700 7142
rect 12650 7100 12700 7108
rect 13200 7142 13250 7150
rect 13200 7108 13208 7142
rect 13242 7108 13250 7142
rect 13200 7100 13250 7108
rect 13750 7142 13800 7150
rect 13750 7108 13758 7142
rect 13792 7108 13800 7142
rect 13750 7100 13800 7108
rect -469 7094 -31 7097
rect -469 7077 -463 7094
rect -37 7077 -31 7094
rect -469 7074 -31 7077
rect 81 7094 519 7097
rect 81 7077 87 7094
rect 513 7077 519 7094
rect 81 7074 519 7077
rect 631 7094 1069 7097
rect 631 7077 637 7094
rect 1063 7077 1069 7094
rect 631 7074 1069 7077
rect 1181 7094 1619 7097
rect 1181 7077 1187 7094
rect 1613 7077 1619 7094
rect 1181 7074 1619 7077
rect 1731 7094 2169 7097
rect 1731 7077 1737 7094
rect 2163 7077 2169 7094
rect 1731 7074 2169 7077
rect 2281 7094 2719 7097
rect 2281 7077 2287 7094
rect 2713 7077 2719 7094
rect 2281 7074 2719 7077
rect 2831 7094 3269 7097
rect 2831 7077 2837 7094
rect 3263 7077 3269 7094
rect 2831 7074 3269 7077
rect 3381 7094 3819 7097
rect 3381 7077 3387 7094
rect 3813 7077 3819 7094
rect 3381 7074 3819 7077
rect 3931 7094 4369 7097
rect 3931 7077 3937 7094
rect 4363 7077 4369 7094
rect 3931 7074 4369 7077
rect 4481 7094 4919 7097
rect 4481 7077 4487 7094
rect 4913 7077 4919 7094
rect 4481 7074 4919 7077
rect 5031 7094 5469 7097
rect 5031 7077 5037 7094
rect 5463 7077 5469 7094
rect 5031 7074 5469 7077
rect 5581 7094 6019 7097
rect 5581 7077 5587 7094
rect 6013 7077 6019 7094
rect 5581 7074 6019 7077
rect 6131 7094 6569 7097
rect 6131 7077 6137 7094
rect 6563 7077 6569 7094
rect 6131 7074 6569 7077
rect 6681 7094 7119 7097
rect 6681 7077 6687 7094
rect 7113 7077 7119 7094
rect 6681 7074 7119 7077
rect 7231 7094 7669 7097
rect 7231 7077 7237 7094
rect 7663 7077 7669 7094
rect 7231 7074 7669 7077
rect 7781 7094 8219 7097
rect 7781 7077 7787 7094
rect 8213 7077 8219 7094
rect 7781 7074 8219 7077
rect 8331 7094 8769 7097
rect 8331 7077 8337 7094
rect 8763 7077 8769 7094
rect 8331 7074 8769 7077
rect 8881 7094 9319 7097
rect 8881 7077 8887 7094
rect 9313 7077 9319 7094
rect 8881 7074 9319 7077
rect 9431 7094 9869 7097
rect 9431 7077 9437 7094
rect 9863 7077 9869 7094
rect 9431 7074 9869 7077
rect 9981 7094 10419 7097
rect 9981 7077 9987 7094
rect 10413 7077 10419 7094
rect 9981 7074 10419 7077
rect 10531 7094 10969 7097
rect 10531 7077 10537 7094
rect 10963 7077 10969 7094
rect 10531 7074 10969 7077
rect 11081 7094 11519 7097
rect 11081 7077 11087 7094
rect 11513 7077 11519 7094
rect 11081 7074 11519 7077
rect 11631 7094 12069 7097
rect 11631 7077 11637 7094
rect 12063 7077 12069 7094
rect 11631 7074 12069 7077
rect 12181 7094 12619 7097
rect 12181 7077 12187 7094
rect 12613 7077 12619 7094
rect 12181 7074 12619 7077
rect 12731 7094 13169 7097
rect 12731 7077 12737 7094
rect 13163 7077 13169 7094
rect 12731 7074 13169 7077
rect 13281 7094 13719 7097
rect 13281 7077 13287 7094
rect 13713 7077 13719 7094
rect 13281 7074 13719 7077
rect -474 7069 -26 7074
rect 76 7069 524 7074
rect 626 7069 1074 7074
rect 1176 7069 1624 7074
rect 1726 7069 2174 7074
rect 2276 7069 2724 7074
rect 2826 7069 3274 7074
rect 3376 7069 3824 7074
rect 3926 7069 4374 7074
rect 4476 7069 4924 7074
rect 5026 7069 5474 7074
rect 5576 7069 6024 7074
rect 6126 7069 6574 7074
rect 6676 7069 7124 7074
rect 7226 7069 7674 7074
rect 7776 7069 8224 7074
rect 8326 7069 8774 7074
rect 8876 7069 9324 7074
rect 9426 7069 9874 7074
rect 9976 7069 10424 7074
rect 10526 7069 10974 7074
rect 11076 7069 11524 7074
rect 11626 7069 12074 7074
rect 12176 7069 12624 7074
rect 12726 7069 13174 7074
rect 13276 7069 13724 7074
rect -474 7063 -3 7069
rect -474 7015 -23 7063
rect -474 6685 -415 7015
rect -85 6685 -23 7015
rect -474 6637 -23 6685
rect -6 6637 -3 7063
rect -474 6631 -3 6637
rect 53 7063 547 7069
rect 53 6637 56 7063
rect 73 7015 527 7063
rect 73 6685 135 7015
rect 465 6685 527 7015
rect 73 6637 527 6685
rect 544 6637 547 7063
rect 53 6631 547 6637
rect 603 7063 1097 7069
rect 603 6637 606 7063
rect 623 7015 1077 7063
rect 623 6685 685 7015
rect 1015 6685 1077 7015
rect 623 6637 1077 6685
rect 1094 6637 1097 7063
rect 603 6631 1097 6637
rect 1153 7063 1647 7069
rect 1153 6637 1156 7063
rect 1173 7015 1627 7063
rect 1173 6685 1235 7015
rect 1565 6685 1627 7015
rect 1173 6637 1627 6685
rect 1644 6637 1647 7063
rect 1153 6631 1647 6637
rect 1703 7063 2197 7069
rect 1703 6637 1706 7063
rect 1723 7015 2177 7063
rect 1723 6685 1785 7015
rect 2115 6685 2177 7015
rect 1723 6637 2177 6685
rect 2194 6637 2197 7063
rect 1703 6631 2197 6637
rect 2253 7063 2747 7069
rect 2253 6637 2256 7063
rect 2273 7015 2727 7063
rect 2273 6685 2335 7015
rect 2665 6685 2727 7015
rect 2273 6637 2727 6685
rect 2744 6637 2747 7063
rect 2253 6631 2747 6637
rect 2803 7063 3297 7069
rect 2803 6637 2806 7063
rect 2823 7015 3277 7063
rect 2823 6685 2885 7015
rect 3215 6685 3277 7015
rect 2823 6637 3277 6685
rect 3294 6637 3297 7063
rect 2803 6631 3297 6637
rect 3353 7063 3847 7069
rect 3353 6637 3356 7063
rect 3373 7015 3827 7063
rect 3373 6685 3435 7015
rect 3765 6685 3827 7015
rect 3373 6637 3827 6685
rect 3844 6637 3847 7063
rect 3353 6631 3847 6637
rect 3903 7063 4397 7069
rect 3903 6637 3906 7063
rect 3923 7015 4377 7063
rect 3923 6685 3985 7015
rect 4315 6685 4377 7015
rect 3923 6637 4377 6685
rect 4394 6637 4397 7063
rect 3903 6631 4397 6637
rect 4453 7063 4947 7069
rect 4453 6637 4456 7063
rect 4473 7015 4927 7063
rect 4473 6685 4535 7015
rect 4865 6685 4927 7015
rect 4473 6637 4927 6685
rect 4944 6637 4947 7063
rect 4453 6631 4947 6637
rect 5003 7063 5497 7069
rect 5003 6637 5006 7063
rect 5023 7015 5477 7063
rect 5023 6685 5085 7015
rect 5415 6685 5477 7015
rect 5023 6637 5477 6685
rect 5494 6637 5497 7063
rect 5003 6631 5497 6637
rect 5553 7063 6047 7069
rect 5553 6637 5556 7063
rect 5573 7015 6027 7063
rect 5573 6685 5635 7015
rect 5965 6685 6027 7015
rect 5573 6637 6027 6685
rect 6044 6637 6047 7063
rect 5553 6631 6047 6637
rect 6103 7063 6597 7069
rect 6103 6637 6106 7063
rect 6123 7015 6577 7063
rect 6123 6685 6185 7015
rect 6515 6685 6577 7015
rect 6123 6637 6577 6685
rect 6594 6637 6597 7063
rect 6103 6631 6597 6637
rect 6653 7063 7147 7069
rect 6653 6637 6656 7063
rect 6673 7015 7127 7063
rect 6673 6685 6735 7015
rect 7065 6685 7127 7015
rect 6673 6637 7127 6685
rect 7144 6637 7147 7063
rect 6653 6631 7147 6637
rect 7203 7063 7697 7069
rect 7203 6637 7206 7063
rect 7223 7015 7677 7063
rect 7223 6685 7285 7015
rect 7615 6685 7677 7015
rect 7223 6637 7677 6685
rect 7694 6637 7697 7063
rect 7203 6631 7697 6637
rect 7753 7063 8247 7069
rect 7753 6637 7756 7063
rect 7773 7015 8227 7063
rect 7773 6685 7835 7015
rect 8165 6685 8227 7015
rect 7773 6637 8227 6685
rect 8244 6637 8247 7063
rect 7753 6631 8247 6637
rect 8303 7063 8797 7069
rect 8303 6637 8306 7063
rect 8323 7015 8777 7063
rect 8323 6685 8385 7015
rect 8715 6685 8777 7015
rect 8323 6637 8777 6685
rect 8794 6637 8797 7063
rect 8303 6631 8797 6637
rect 8853 7063 9347 7069
rect 8853 6637 8856 7063
rect 8873 7015 9327 7063
rect 8873 6685 8935 7015
rect 9265 6685 9327 7015
rect 8873 6637 9327 6685
rect 9344 6637 9347 7063
rect 8853 6631 9347 6637
rect 9403 7063 9897 7069
rect 9403 6637 9406 7063
rect 9423 7015 9877 7063
rect 9423 6685 9485 7015
rect 9815 6685 9877 7015
rect 9423 6637 9877 6685
rect 9894 6637 9897 7063
rect 9403 6631 9897 6637
rect 9953 7063 10447 7069
rect 9953 6637 9956 7063
rect 9973 7015 10427 7063
rect 9973 6685 10035 7015
rect 10365 6685 10427 7015
rect 9973 6637 10427 6685
rect 10444 6637 10447 7063
rect 9953 6631 10447 6637
rect 10503 7063 10997 7069
rect 10503 6637 10506 7063
rect 10523 7015 10977 7063
rect 10523 6685 10585 7015
rect 10915 6685 10977 7015
rect 10523 6637 10977 6685
rect 10994 6637 10997 7063
rect 10503 6631 10997 6637
rect 11053 7063 11547 7069
rect 11053 6637 11056 7063
rect 11073 7015 11527 7063
rect 11073 6685 11135 7015
rect 11465 6685 11527 7015
rect 11073 6637 11527 6685
rect 11544 6637 11547 7063
rect 11053 6631 11547 6637
rect 11603 7063 12097 7069
rect 11603 6637 11606 7063
rect 11623 7015 12077 7063
rect 11623 6685 11685 7015
rect 12015 6685 12077 7015
rect 11623 6637 12077 6685
rect 12094 6637 12097 7063
rect 11603 6631 12097 6637
rect 12153 7063 12647 7069
rect 12153 6637 12156 7063
rect 12173 7015 12627 7063
rect 12173 6685 12235 7015
rect 12565 6685 12627 7015
rect 12173 6637 12627 6685
rect 12644 6637 12647 7063
rect 12153 6631 12647 6637
rect 12703 7063 13197 7069
rect 12703 6637 12706 7063
rect 12723 7015 13177 7063
rect 12723 6685 12785 7015
rect 13115 6685 13177 7015
rect 12723 6637 13177 6685
rect 13194 6637 13197 7063
rect 12703 6631 13197 6637
rect 13253 7063 13724 7069
rect 13253 6637 13256 7063
rect 13273 7015 13724 7063
rect 13273 6685 13335 7015
rect 13665 6685 13724 7015
rect 13273 6637 13724 6685
rect 13253 6631 13724 6637
rect -474 6626 -26 6631
rect 76 6626 524 6631
rect 626 6626 1074 6631
rect 1176 6626 1624 6631
rect 1726 6626 2174 6631
rect 2276 6626 2724 6631
rect 2826 6626 3274 6631
rect 3376 6626 3824 6631
rect 3926 6626 4374 6631
rect 4476 6626 4924 6631
rect 5026 6626 5474 6631
rect 5576 6626 6024 6631
rect 6126 6626 6574 6631
rect 6676 6626 7124 6631
rect 7226 6626 7674 6631
rect 7776 6626 8224 6631
rect 8326 6626 8774 6631
rect 8876 6626 9324 6631
rect 9426 6626 9874 6631
rect 9976 6626 10424 6631
rect 10526 6626 10974 6631
rect 11076 6626 11524 6631
rect 11626 6626 12074 6631
rect 12176 6626 12624 6631
rect 12726 6626 13174 6631
rect 13276 6626 13724 6631
rect -1025 6600 -725 6619
rect -469 6623 -31 6626
rect -469 6606 -463 6623
rect -37 6606 -31 6623
rect -469 6603 -31 6606
rect 81 6623 519 6626
rect 81 6606 87 6623
rect 513 6606 519 6623
rect 81 6603 519 6606
rect 631 6623 1069 6626
rect 631 6606 637 6623
rect 1063 6606 1069 6623
rect 631 6603 1069 6606
rect 1181 6623 1619 6626
rect 1181 6606 1187 6623
rect 1613 6606 1619 6623
rect 1181 6603 1619 6606
rect 1731 6623 2169 6626
rect 1731 6606 1737 6623
rect 2163 6606 2169 6623
rect 1731 6603 2169 6606
rect 2281 6623 2719 6626
rect 2281 6606 2287 6623
rect 2713 6606 2719 6623
rect 2281 6603 2719 6606
rect 2831 6623 3269 6626
rect 2831 6606 2837 6623
rect 3263 6606 3269 6623
rect 2831 6603 3269 6606
rect 3381 6623 3819 6626
rect 3381 6606 3387 6623
rect 3813 6606 3819 6623
rect 3381 6603 3819 6606
rect 3931 6623 4369 6626
rect 3931 6606 3937 6623
rect 4363 6606 4369 6623
rect 3931 6603 4369 6606
rect 4481 6623 4919 6626
rect 4481 6606 4487 6623
rect 4913 6606 4919 6623
rect 4481 6603 4919 6606
rect 5031 6623 5469 6626
rect 5031 6606 5037 6623
rect 5463 6606 5469 6623
rect 5031 6603 5469 6606
rect 5581 6623 6019 6626
rect 5581 6606 5587 6623
rect 6013 6606 6019 6623
rect 5581 6603 6019 6606
rect 6131 6623 6569 6626
rect 6131 6606 6137 6623
rect 6563 6606 6569 6623
rect 6131 6603 6569 6606
rect 6681 6623 7119 6626
rect 6681 6606 6687 6623
rect 7113 6606 7119 6623
rect 6681 6603 7119 6606
rect 7231 6623 7669 6626
rect 7231 6606 7237 6623
rect 7663 6606 7669 6623
rect 7231 6603 7669 6606
rect 7781 6623 8219 6626
rect 7781 6606 7787 6623
rect 8213 6606 8219 6623
rect 7781 6603 8219 6606
rect 8331 6623 8769 6626
rect 8331 6606 8337 6623
rect 8763 6606 8769 6623
rect 8331 6603 8769 6606
rect 8881 6623 9319 6626
rect 8881 6606 8887 6623
rect 9313 6606 9319 6623
rect 8881 6603 9319 6606
rect 9431 6623 9869 6626
rect 9431 6606 9437 6623
rect 9863 6606 9869 6623
rect 9431 6603 9869 6606
rect 9981 6623 10419 6626
rect 9981 6606 9987 6623
rect 10413 6606 10419 6623
rect 9981 6603 10419 6606
rect 10531 6623 10969 6626
rect 10531 6606 10537 6623
rect 10963 6606 10969 6623
rect 10531 6603 10969 6606
rect 11081 6623 11519 6626
rect 11081 6606 11087 6623
rect 11513 6606 11519 6623
rect 11081 6603 11519 6606
rect 11631 6623 12069 6626
rect 11631 6606 11637 6623
rect 12063 6606 12069 6623
rect 11631 6603 12069 6606
rect 12181 6623 12619 6626
rect 12181 6606 12187 6623
rect 12613 6606 12619 6623
rect 12181 6603 12619 6606
rect 12731 6623 13169 6626
rect 12731 6606 12737 6623
rect 13163 6606 13169 6623
rect 12731 6603 13169 6606
rect 13281 6623 13719 6626
rect 13281 6606 13287 6623
rect 13713 6606 13719 6623
rect 13281 6603 13719 6606
rect 13975 6619 13987 7150
rect 14263 6619 14275 7150
rect 13975 6600 14275 6619
rect -1025 6069 -1013 6600
rect -737 6069 -725 6600
rect -550 6592 -500 6600
rect -550 6558 -542 6592
rect -508 6558 -500 6592
rect -550 6550 -500 6558
rect 0 6592 50 6600
rect 0 6558 8 6592
rect 42 6558 50 6592
rect 0 6550 50 6558
rect 550 6592 600 6600
rect 550 6558 558 6592
rect 592 6558 600 6592
rect 550 6550 600 6558
rect 1100 6592 1150 6600
rect 1100 6558 1108 6592
rect 1142 6558 1150 6592
rect 1100 6550 1150 6558
rect 1650 6592 1700 6600
rect 1650 6558 1658 6592
rect 1692 6558 1700 6592
rect 1650 6550 1700 6558
rect 2200 6592 2250 6600
rect 2200 6558 2208 6592
rect 2242 6558 2250 6592
rect 2200 6550 2250 6558
rect 2750 6592 2800 6600
rect 2750 6558 2758 6592
rect 2792 6558 2800 6592
rect 2750 6550 2800 6558
rect 3300 6592 3350 6600
rect 3300 6558 3308 6592
rect 3342 6558 3350 6592
rect 3300 6550 3350 6558
rect 3850 6592 3900 6600
rect 3850 6558 3858 6592
rect 3892 6558 3900 6592
rect 3850 6550 3900 6558
rect 4400 6592 4450 6600
rect 4400 6558 4408 6592
rect 4442 6558 4450 6592
rect 4400 6550 4450 6558
rect 4950 6592 5000 6600
rect 4950 6558 4958 6592
rect 4992 6558 5000 6592
rect 4950 6550 5000 6558
rect 5500 6592 5550 6600
rect 5500 6558 5508 6592
rect 5542 6558 5550 6592
rect 5500 6550 5550 6558
rect 6050 6592 6100 6600
rect 6050 6558 6058 6592
rect 6092 6558 6100 6592
rect 6050 6550 6100 6558
rect 6600 6592 6650 6600
rect 6600 6558 6608 6592
rect 6642 6558 6650 6592
rect 6600 6550 6650 6558
rect 7150 6592 7200 6600
rect 7150 6558 7158 6592
rect 7192 6558 7200 6592
rect 7150 6550 7200 6558
rect 7700 6592 7750 6600
rect 7700 6558 7708 6592
rect 7742 6558 7750 6592
rect 7700 6550 7750 6558
rect 8250 6592 8300 6600
rect 8250 6558 8258 6592
rect 8292 6558 8300 6592
rect 8250 6550 8300 6558
rect 8800 6592 8850 6600
rect 8800 6558 8808 6592
rect 8842 6558 8850 6592
rect 8800 6550 8850 6558
rect 9350 6592 9400 6600
rect 9350 6558 9358 6592
rect 9392 6558 9400 6592
rect 9350 6550 9400 6558
rect 9900 6592 9950 6600
rect 9900 6558 9908 6592
rect 9942 6558 9950 6592
rect 9900 6550 9950 6558
rect 10450 6592 10500 6600
rect 10450 6558 10458 6592
rect 10492 6558 10500 6592
rect 10450 6550 10500 6558
rect 11000 6592 11050 6600
rect 11000 6558 11008 6592
rect 11042 6558 11050 6592
rect 11000 6550 11050 6558
rect 11550 6592 11600 6600
rect 11550 6558 11558 6592
rect 11592 6558 11600 6592
rect 11550 6550 11600 6558
rect 12100 6592 12150 6600
rect 12100 6558 12108 6592
rect 12142 6558 12150 6592
rect 12100 6550 12150 6558
rect 12650 6592 12700 6600
rect 12650 6558 12658 6592
rect 12692 6558 12700 6592
rect 12650 6550 12700 6558
rect 13200 6592 13250 6600
rect 13200 6558 13208 6592
rect 13242 6558 13250 6592
rect 13200 6550 13250 6558
rect 13750 6592 13800 6600
rect 13750 6558 13758 6592
rect 13792 6558 13800 6592
rect 13750 6550 13800 6558
rect -469 6544 -31 6547
rect -469 6527 -463 6544
rect -37 6527 -31 6544
rect -469 6524 -31 6527
rect 81 6544 519 6547
rect 81 6527 87 6544
rect 513 6527 519 6544
rect 81 6524 519 6527
rect 631 6544 1069 6547
rect 631 6527 637 6544
rect 1063 6527 1069 6544
rect 631 6524 1069 6527
rect 1181 6544 1619 6547
rect 1181 6527 1187 6544
rect 1613 6527 1619 6544
rect 1181 6524 1619 6527
rect 1731 6544 2169 6547
rect 1731 6527 1737 6544
rect 2163 6527 2169 6544
rect 1731 6524 2169 6527
rect 2281 6544 2719 6547
rect 2281 6527 2287 6544
rect 2713 6527 2719 6544
rect 2281 6524 2719 6527
rect 2831 6544 3269 6547
rect 2831 6527 2837 6544
rect 3263 6527 3269 6544
rect 2831 6524 3269 6527
rect 3381 6544 3819 6547
rect 3381 6527 3387 6544
rect 3813 6527 3819 6544
rect 3381 6524 3819 6527
rect 3931 6544 4369 6547
rect 3931 6527 3937 6544
rect 4363 6527 4369 6544
rect 3931 6524 4369 6527
rect 4481 6544 4919 6547
rect 4481 6527 4487 6544
rect 4913 6527 4919 6544
rect 4481 6524 4919 6527
rect 5031 6544 5469 6547
rect 5031 6527 5037 6544
rect 5463 6527 5469 6544
rect 5031 6524 5469 6527
rect 5581 6544 6019 6547
rect 5581 6527 5587 6544
rect 6013 6527 6019 6544
rect 5581 6524 6019 6527
rect 6131 6544 6569 6547
rect 6131 6527 6137 6544
rect 6563 6527 6569 6544
rect 6131 6524 6569 6527
rect 6681 6544 7119 6547
rect 6681 6527 6687 6544
rect 7113 6527 7119 6544
rect 6681 6524 7119 6527
rect 7231 6544 7669 6547
rect 7231 6527 7237 6544
rect 7663 6527 7669 6544
rect 7231 6524 7669 6527
rect 7781 6544 8219 6547
rect 7781 6527 7787 6544
rect 8213 6527 8219 6544
rect 7781 6524 8219 6527
rect 8331 6544 8769 6547
rect 8331 6527 8337 6544
rect 8763 6527 8769 6544
rect 8331 6524 8769 6527
rect 8881 6544 9319 6547
rect 8881 6527 8887 6544
rect 9313 6527 9319 6544
rect 8881 6524 9319 6527
rect 9431 6544 9869 6547
rect 9431 6527 9437 6544
rect 9863 6527 9869 6544
rect 9431 6524 9869 6527
rect 9981 6544 10419 6547
rect 9981 6527 9987 6544
rect 10413 6527 10419 6544
rect 9981 6524 10419 6527
rect 10531 6544 10969 6547
rect 10531 6527 10537 6544
rect 10963 6527 10969 6544
rect 10531 6524 10969 6527
rect 11081 6544 11519 6547
rect 11081 6527 11087 6544
rect 11513 6527 11519 6544
rect 11081 6524 11519 6527
rect 11631 6544 12069 6547
rect 11631 6527 11637 6544
rect 12063 6527 12069 6544
rect 11631 6524 12069 6527
rect 12181 6544 12619 6547
rect 12181 6527 12187 6544
rect 12613 6527 12619 6544
rect 12181 6524 12619 6527
rect 12731 6544 13169 6547
rect 12731 6527 12737 6544
rect 13163 6527 13169 6544
rect 12731 6524 13169 6527
rect 13281 6544 13719 6547
rect 13281 6527 13287 6544
rect 13713 6527 13719 6544
rect 13281 6524 13719 6527
rect -474 6519 -26 6524
rect 76 6519 524 6524
rect 626 6519 1074 6524
rect 1176 6519 1624 6524
rect 1726 6519 2174 6524
rect 2276 6519 2724 6524
rect 2826 6519 3274 6524
rect 3376 6519 3824 6524
rect 3926 6519 4374 6524
rect 4476 6519 4924 6524
rect 5026 6519 5474 6524
rect 5576 6519 6024 6524
rect 6126 6519 6574 6524
rect 6676 6519 7124 6524
rect 7226 6519 7674 6524
rect 7776 6519 8224 6524
rect 8326 6519 8774 6524
rect 8876 6519 9324 6524
rect 9426 6519 9874 6524
rect 9976 6519 10424 6524
rect 10526 6519 10974 6524
rect 11076 6519 11524 6524
rect 11626 6519 12074 6524
rect 12176 6519 12624 6524
rect 12726 6519 13174 6524
rect 13276 6519 13724 6524
rect -474 6513 -3 6519
rect -474 6465 -23 6513
rect -474 6135 -415 6465
rect -85 6135 -23 6465
rect -474 6087 -23 6135
rect -6 6087 -3 6513
rect -474 6081 -3 6087
rect 53 6513 547 6519
rect 53 6087 56 6513
rect 73 6465 527 6513
rect 73 6135 135 6465
rect 465 6135 527 6465
rect 73 6087 527 6135
rect 544 6087 547 6513
rect 53 6081 547 6087
rect 603 6513 1097 6519
rect 603 6087 606 6513
rect 623 6465 1077 6513
rect 623 6135 685 6465
rect 1015 6135 1077 6465
rect 623 6087 1077 6135
rect 1094 6087 1097 6513
rect 603 6081 1097 6087
rect 1153 6513 1647 6519
rect 1153 6087 1156 6513
rect 1173 6465 1627 6513
rect 1173 6135 1235 6465
rect 1565 6135 1627 6465
rect 1173 6087 1627 6135
rect 1644 6087 1647 6513
rect 1153 6081 1647 6087
rect 1703 6513 2197 6519
rect 1703 6087 1706 6513
rect 1723 6465 2177 6513
rect 1723 6135 1785 6465
rect 2115 6135 2177 6465
rect 1723 6087 2177 6135
rect 2194 6087 2197 6513
rect 1703 6081 2197 6087
rect 2253 6513 2747 6519
rect 2253 6087 2256 6513
rect 2273 6465 2727 6513
rect 2273 6135 2335 6465
rect 2665 6135 2727 6465
rect 2273 6087 2727 6135
rect 2744 6087 2747 6513
rect 2253 6081 2747 6087
rect 2803 6513 3297 6519
rect 2803 6087 2806 6513
rect 2823 6465 3277 6513
rect 2823 6135 2885 6465
rect 3215 6135 3277 6465
rect 2823 6087 3277 6135
rect 3294 6087 3297 6513
rect 2803 6081 3297 6087
rect 3353 6513 3847 6519
rect 3353 6087 3356 6513
rect 3373 6465 3827 6513
rect 3373 6135 3435 6465
rect 3765 6135 3827 6465
rect 3373 6087 3827 6135
rect 3844 6087 3847 6513
rect 3353 6081 3847 6087
rect 3903 6513 4397 6519
rect 3903 6087 3906 6513
rect 3923 6465 4377 6513
rect 3923 6135 3985 6465
rect 4315 6135 4377 6465
rect 3923 6087 4377 6135
rect 4394 6087 4397 6513
rect 3903 6081 4397 6087
rect 4453 6513 4947 6519
rect 4453 6087 4456 6513
rect 4473 6465 4927 6513
rect 4473 6135 4535 6465
rect 4865 6135 4927 6465
rect 4473 6087 4927 6135
rect 4944 6087 4947 6513
rect 4453 6081 4947 6087
rect 5003 6513 5497 6519
rect 5003 6087 5006 6513
rect 5023 6465 5477 6513
rect 5023 6135 5085 6465
rect 5415 6135 5477 6465
rect 5023 6087 5477 6135
rect 5494 6087 5497 6513
rect 5003 6081 5497 6087
rect 5553 6513 6047 6519
rect 5553 6087 5556 6513
rect 5573 6465 6027 6513
rect 5573 6135 5635 6465
rect 5965 6135 6027 6465
rect 5573 6087 6027 6135
rect 6044 6087 6047 6513
rect 5553 6081 6047 6087
rect 6103 6513 6597 6519
rect 6103 6087 6106 6513
rect 6123 6465 6577 6513
rect 6123 6135 6185 6465
rect 6515 6135 6577 6465
rect 6123 6087 6577 6135
rect 6594 6087 6597 6513
rect 6103 6081 6597 6087
rect 6653 6513 7147 6519
rect 6653 6087 6656 6513
rect 6673 6465 7127 6513
rect 6673 6135 6735 6465
rect 7065 6135 7127 6465
rect 6673 6087 7127 6135
rect 7144 6087 7147 6513
rect 6653 6081 7147 6087
rect 7203 6513 7697 6519
rect 7203 6087 7206 6513
rect 7223 6465 7677 6513
rect 7223 6135 7285 6465
rect 7615 6135 7677 6465
rect 7223 6087 7677 6135
rect 7694 6087 7697 6513
rect 7203 6081 7697 6087
rect 7753 6513 8247 6519
rect 7753 6087 7756 6513
rect 7773 6465 8227 6513
rect 7773 6135 7835 6465
rect 8165 6135 8227 6465
rect 7773 6087 8227 6135
rect 8244 6087 8247 6513
rect 7753 6081 8247 6087
rect 8303 6513 8797 6519
rect 8303 6087 8306 6513
rect 8323 6465 8777 6513
rect 8323 6135 8385 6465
rect 8715 6135 8777 6465
rect 8323 6087 8777 6135
rect 8794 6087 8797 6513
rect 8303 6081 8797 6087
rect 8853 6513 9347 6519
rect 8853 6087 8856 6513
rect 8873 6465 9327 6513
rect 8873 6135 8935 6465
rect 9265 6135 9327 6465
rect 8873 6087 9327 6135
rect 9344 6087 9347 6513
rect 8853 6081 9347 6087
rect 9403 6513 9897 6519
rect 9403 6087 9406 6513
rect 9423 6465 9877 6513
rect 9423 6135 9485 6465
rect 9815 6135 9877 6465
rect 9423 6087 9877 6135
rect 9894 6087 9897 6513
rect 9403 6081 9897 6087
rect 9953 6513 10447 6519
rect 9953 6087 9956 6513
rect 9973 6465 10427 6513
rect 9973 6135 10035 6465
rect 10365 6135 10427 6465
rect 9973 6087 10427 6135
rect 10444 6087 10447 6513
rect 9953 6081 10447 6087
rect 10503 6513 10997 6519
rect 10503 6087 10506 6513
rect 10523 6465 10977 6513
rect 10523 6135 10585 6465
rect 10915 6135 10977 6465
rect 10523 6087 10977 6135
rect 10994 6087 10997 6513
rect 10503 6081 10997 6087
rect 11053 6513 11547 6519
rect 11053 6087 11056 6513
rect 11073 6465 11527 6513
rect 11073 6135 11135 6465
rect 11465 6135 11527 6465
rect 11073 6087 11527 6135
rect 11544 6087 11547 6513
rect 11053 6081 11547 6087
rect 11603 6513 12097 6519
rect 11603 6087 11606 6513
rect 11623 6465 12077 6513
rect 11623 6135 11685 6465
rect 12015 6135 12077 6465
rect 11623 6087 12077 6135
rect 12094 6087 12097 6513
rect 11603 6081 12097 6087
rect 12153 6513 12647 6519
rect 12153 6087 12156 6513
rect 12173 6465 12627 6513
rect 12173 6135 12235 6465
rect 12565 6135 12627 6465
rect 12173 6087 12627 6135
rect 12644 6087 12647 6513
rect 12153 6081 12647 6087
rect 12703 6513 13197 6519
rect 12703 6087 12706 6513
rect 12723 6465 13177 6513
rect 12723 6135 12785 6465
rect 13115 6135 13177 6465
rect 12723 6087 13177 6135
rect 13194 6087 13197 6513
rect 12703 6081 13197 6087
rect 13253 6513 13724 6519
rect 13253 6087 13256 6513
rect 13273 6465 13724 6513
rect 13273 6135 13335 6465
rect 13665 6135 13724 6465
rect 13273 6087 13724 6135
rect 13253 6081 13724 6087
rect -474 6076 -26 6081
rect 76 6076 524 6081
rect 626 6076 1074 6081
rect 1176 6076 1624 6081
rect 1726 6076 2174 6081
rect 2276 6076 2724 6081
rect 2826 6076 3274 6081
rect 3376 6076 3824 6081
rect 3926 6076 4374 6081
rect 4476 6076 4924 6081
rect 5026 6076 5474 6081
rect 5576 6076 6024 6081
rect 6126 6076 6574 6081
rect 6676 6076 7124 6081
rect 7226 6076 7674 6081
rect 7776 6076 8224 6081
rect 8326 6076 8774 6081
rect 8876 6076 9324 6081
rect 9426 6076 9874 6081
rect 9976 6076 10424 6081
rect 10526 6076 10974 6081
rect 11076 6076 11524 6081
rect 11626 6076 12074 6081
rect 12176 6076 12624 6081
rect 12726 6076 13174 6081
rect 13276 6076 13724 6081
rect -1025 6050 -725 6069
rect -469 6073 -31 6076
rect -469 6056 -463 6073
rect -37 6056 -31 6073
rect -469 6053 -31 6056
rect 81 6073 519 6076
rect 81 6056 87 6073
rect 513 6056 519 6073
rect 81 6053 519 6056
rect 631 6073 1069 6076
rect 631 6056 637 6073
rect 1063 6056 1069 6073
rect 631 6053 1069 6056
rect 1181 6073 1619 6076
rect 1181 6056 1187 6073
rect 1613 6056 1619 6073
rect 1181 6053 1619 6056
rect 1731 6073 2169 6076
rect 1731 6056 1737 6073
rect 2163 6056 2169 6073
rect 1731 6053 2169 6056
rect 2281 6073 2719 6076
rect 2281 6056 2287 6073
rect 2713 6056 2719 6073
rect 2281 6053 2719 6056
rect 2831 6073 3269 6076
rect 2831 6056 2837 6073
rect 3263 6056 3269 6073
rect 2831 6053 3269 6056
rect 3381 6073 3819 6076
rect 3381 6056 3387 6073
rect 3813 6056 3819 6073
rect 3381 6053 3819 6056
rect 3931 6073 4369 6076
rect 3931 6056 3937 6073
rect 4363 6056 4369 6073
rect 3931 6053 4369 6056
rect 4481 6073 4919 6076
rect 4481 6056 4487 6073
rect 4913 6056 4919 6073
rect 4481 6053 4919 6056
rect 5031 6073 5469 6076
rect 5031 6056 5037 6073
rect 5463 6056 5469 6073
rect 5031 6053 5469 6056
rect 5581 6073 6019 6076
rect 5581 6056 5587 6073
rect 6013 6056 6019 6073
rect 5581 6053 6019 6056
rect 6131 6073 6569 6076
rect 6131 6056 6137 6073
rect 6563 6056 6569 6073
rect 6131 6053 6569 6056
rect 6681 6073 7119 6076
rect 6681 6056 6687 6073
rect 7113 6056 7119 6073
rect 6681 6053 7119 6056
rect 7231 6073 7669 6076
rect 7231 6056 7237 6073
rect 7663 6056 7669 6073
rect 7231 6053 7669 6056
rect 7781 6073 8219 6076
rect 7781 6056 7787 6073
rect 8213 6056 8219 6073
rect 7781 6053 8219 6056
rect 8331 6073 8769 6076
rect 8331 6056 8337 6073
rect 8763 6056 8769 6073
rect 8331 6053 8769 6056
rect 8881 6073 9319 6076
rect 8881 6056 8887 6073
rect 9313 6056 9319 6073
rect 8881 6053 9319 6056
rect 9431 6073 9869 6076
rect 9431 6056 9437 6073
rect 9863 6056 9869 6073
rect 9431 6053 9869 6056
rect 9981 6073 10419 6076
rect 9981 6056 9987 6073
rect 10413 6056 10419 6073
rect 9981 6053 10419 6056
rect 10531 6073 10969 6076
rect 10531 6056 10537 6073
rect 10963 6056 10969 6073
rect 10531 6053 10969 6056
rect 11081 6073 11519 6076
rect 11081 6056 11087 6073
rect 11513 6056 11519 6073
rect 11081 6053 11519 6056
rect 11631 6073 12069 6076
rect 11631 6056 11637 6073
rect 12063 6056 12069 6073
rect 11631 6053 12069 6056
rect 12181 6073 12619 6076
rect 12181 6056 12187 6073
rect 12613 6056 12619 6073
rect 12181 6053 12619 6056
rect 12731 6073 13169 6076
rect 12731 6056 12737 6073
rect 13163 6056 13169 6073
rect 12731 6053 13169 6056
rect 13281 6073 13719 6076
rect 13281 6056 13287 6073
rect 13713 6056 13719 6073
rect 13281 6053 13719 6056
rect 13975 6069 13987 6600
rect 14263 6069 14275 6600
rect 13975 6050 14275 6069
rect -1025 5519 -1013 6050
rect -737 5519 -725 6050
rect -550 6042 -500 6050
rect -550 6008 -542 6042
rect -508 6008 -500 6042
rect -550 6000 -500 6008
rect 0 6042 50 6050
rect 0 6008 8 6042
rect 42 6008 50 6042
rect 0 6000 50 6008
rect 550 6042 600 6050
rect 550 6008 558 6042
rect 592 6008 600 6042
rect 550 6000 600 6008
rect 1100 6042 1150 6050
rect 1100 6008 1108 6042
rect 1142 6008 1150 6042
rect 1100 6000 1150 6008
rect 1650 6042 1700 6050
rect 1650 6008 1658 6042
rect 1692 6008 1700 6042
rect 1650 6000 1700 6008
rect 2200 6042 2250 6050
rect 2200 6008 2208 6042
rect 2242 6008 2250 6042
rect 2200 6000 2250 6008
rect 2750 6042 2800 6050
rect 2750 6008 2758 6042
rect 2792 6008 2800 6042
rect 2750 6000 2800 6008
rect 3300 6042 3350 6050
rect 3300 6008 3308 6042
rect 3342 6008 3350 6042
rect 3300 6000 3350 6008
rect 3850 6042 3900 6050
rect 3850 6008 3858 6042
rect 3892 6008 3900 6042
rect 3850 6000 3900 6008
rect 4400 6042 4450 6050
rect 4400 6008 4408 6042
rect 4442 6008 4450 6042
rect 4400 6000 4450 6008
rect 4950 6042 5000 6050
rect 4950 6008 4958 6042
rect 4992 6008 5000 6042
rect 4950 6000 5000 6008
rect 5500 6042 5550 6050
rect 5500 6008 5508 6042
rect 5542 6008 5550 6042
rect 5500 6000 5550 6008
rect 6050 6042 6100 6050
rect 6050 6008 6058 6042
rect 6092 6008 6100 6042
rect 6050 6000 6100 6008
rect 6600 6042 6650 6050
rect 6600 6008 6608 6042
rect 6642 6008 6650 6042
rect 6600 6000 6650 6008
rect 7150 6042 7200 6050
rect 7150 6008 7158 6042
rect 7192 6008 7200 6042
rect 7150 6000 7200 6008
rect 7700 6042 7750 6050
rect 7700 6008 7708 6042
rect 7742 6008 7750 6042
rect 7700 6000 7750 6008
rect 8250 6042 8300 6050
rect 8250 6008 8258 6042
rect 8292 6008 8300 6042
rect 8250 6000 8300 6008
rect 8800 6042 8850 6050
rect 8800 6008 8808 6042
rect 8842 6008 8850 6042
rect 8800 6000 8850 6008
rect 9350 6042 9400 6050
rect 9350 6008 9358 6042
rect 9392 6008 9400 6042
rect 9350 6000 9400 6008
rect 9900 6042 9950 6050
rect 9900 6008 9908 6042
rect 9942 6008 9950 6042
rect 9900 6000 9950 6008
rect 10450 6042 10500 6050
rect 10450 6008 10458 6042
rect 10492 6008 10500 6042
rect 10450 6000 10500 6008
rect 11000 6042 11050 6050
rect 11000 6008 11008 6042
rect 11042 6008 11050 6042
rect 11000 6000 11050 6008
rect 11550 6042 11600 6050
rect 11550 6008 11558 6042
rect 11592 6008 11600 6042
rect 11550 6000 11600 6008
rect 12100 6042 12150 6050
rect 12100 6008 12108 6042
rect 12142 6008 12150 6042
rect 12100 6000 12150 6008
rect 12650 6042 12700 6050
rect 12650 6008 12658 6042
rect 12692 6008 12700 6042
rect 12650 6000 12700 6008
rect 13200 6042 13250 6050
rect 13200 6008 13208 6042
rect 13242 6008 13250 6042
rect 13200 6000 13250 6008
rect 13750 6042 13800 6050
rect 13750 6008 13758 6042
rect 13792 6008 13800 6042
rect 13750 6000 13800 6008
rect -469 5994 -31 5997
rect -469 5977 -463 5994
rect -37 5977 -31 5994
rect -469 5974 -31 5977
rect 81 5994 519 5997
rect 81 5977 87 5994
rect 513 5977 519 5994
rect 81 5974 519 5977
rect 631 5994 1069 5997
rect 631 5977 637 5994
rect 1063 5977 1069 5994
rect 631 5974 1069 5977
rect 1181 5994 1619 5997
rect 1181 5977 1187 5994
rect 1613 5977 1619 5994
rect 1181 5974 1619 5977
rect 1731 5994 2169 5997
rect 1731 5977 1737 5994
rect 2163 5977 2169 5994
rect 1731 5974 2169 5977
rect 2281 5994 2719 5997
rect 2281 5977 2287 5994
rect 2713 5977 2719 5994
rect 2281 5974 2719 5977
rect 2831 5994 3269 5997
rect 2831 5977 2837 5994
rect 3263 5977 3269 5994
rect 2831 5974 3269 5977
rect 3381 5994 3819 5997
rect 3381 5977 3387 5994
rect 3813 5977 3819 5994
rect 3381 5974 3819 5977
rect 3931 5994 4369 5997
rect 3931 5977 3937 5994
rect 4363 5977 4369 5994
rect 3931 5974 4369 5977
rect 4481 5994 4919 5997
rect 4481 5977 4487 5994
rect 4913 5977 4919 5994
rect 4481 5974 4919 5977
rect 5031 5994 5469 5997
rect 5031 5977 5037 5994
rect 5463 5977 5469 5994
rect 5031 5974 5469 5977
rect 5581 5994 6019 5997
rect 5581 5977 5587 5994
rect 6013 5977 6019 5994
rect 5581 5974 6019 5977
rect 6131 5994 6569 5997
rect 6131 5977 6137 5994
rect 6563 5977 6569 5994
rect 6131 5974 6569 5977
rect 6681 5994 7119 5997
rect 6681 5977 6687 5994
rect 7113 5977 7119 5994
rect 6681 5974 7119 5977
rect 7231 5994 7669 5997
rect 7231 5977 7237 5994
rect 7663 5977 7669 5994
rect 7231 5974 7669 5977
rect 7781 5994 8219 5997
rect 7781 5977 7787 5994
rect 8213 5977 8219 5994
rect 7781 5974 8219 5977
rect 8331 5994 8769 5997
rect 8331 5977 8337 5994
rect 8763 5977 8769 5994
rect 8331 5974 8769 5977
rect 8881 5994 9319 5997
rect 8881 5977 8887 5994
rect 9313 5977 9319 5994
rect 8881 5974 9319 5977
rect 9431 5994 9869 5997
rect 9431 5977 9437 5994
rect 9863 5977 9869 5994
rect 9431 5974 9869 5977
rect 9981 5994 10419 5997
rect 9981 5977 9987 5994
rect 10413 5977 10419 5994
rect 9981 5974 10419 5977
rect 10531 5994 10969 5997
rect 10531 5977 10537 5994
rect 10963 5977 10969 5994
rect 10531 5974 10969 5977
rect 11081 5994 11519 5997
rect 11081 5977 11087 5994
rect 11513 5977 11519 5994
rect 11081 5974 11519 5977
rect 11631 5994 12069 5997
rect 11631 5977 11637 5994
rect 12063 5977 12069 5994
rect 11631 5974 12069 5977
rect 12181 5994 12619 5997
rect 12181 5977 12187 5994
rect 12613 5977 12619 5994
rect 12181 5974 12619 5977
rect 12731 5994 13169 5997
rect 12731 5977 12737 5994
rect 13163 5977 13169 5994
rect 12731 5974 13169 5977
rect 13281 5994 13719 5997
rect 13281 5977 13287 5994
rect 13713 5977 13719 5994
rect 13281 5974 13719 5977
rect -474 5969 -26 5974
rect 76 5969 524 5974
rect 626 5969 1074 5974
rect 1176 5969 1624 5974
rect 1726 5969 2174 5974
rect 2276 5969 2724 5974
rect 2826 5969 3274 5974
rect 3376 5969 3824 5974
rect 3926 5969 4374 5974
rect 4476 5969 4924 5974
rect 5026 5969 5474 5974
rect 5576 5969 6024 5974
rect 6126 5969 6574 5974
rect 6676 5969 7124 5974
rect 7226 5969 7674 5974
rect 7776 5969 8224 5974
rect 8326 5969 8774 5974
rect 8876 5969 9324 5974
rect 9426 5969 9874 5974
rect 9976 5969 10424 5974
rect 10526 5969 10974 5974
rect 11076 5969 11524 5974
rect 11626 5969 12074 5974
rect 12176 5969 12624 5974
rect 12726 5969 13174 5974
rect 13276 5969 13724 5974
rect -474 5963 -3 5969
rect -474 5915 -23 5963
rect -474 5585 -415 5915
rect -85 5585 -23 5915
rect -474 5537 -23 5585
rect -6 5537 -3 5963
rect -474 5531 -3 5537
rect 53 5963 547 5969
rect 53 5537 56 5963
rect 73 5915 527 5963
rect 73 5585 135 5915
rect 465 5585 527 5915
rect 73 5537 527 5585
rect 544 5537 547 5963
rect 53 5531 547 5537
rect 603 5963 1097 5969
rect 603 5537 606 5963
rect 623 5915 1077 5963
rect 623 5585 685 5915
rect 1015 5585 1077 5915
rect 623 5537 1077 5585
rect 1094 5537 1097 5963
rect 603 5531 1097 5537
rect 1153 5963 1647 5969
rect 1153 5537 1156 5963
rect 1173 5915 1627 5963
rect 1173 5585 1235 5915
rect 1565 5585 1627 5915
rect 1173 5537 1627 5585
rect 1644 5537 1647 5963
rect 1153 5531 1647 5537
rect 1703 5963 2197 5969
rect 1703 5537 1706 5963
rect 1723 5915 2177 5963
rect 1723 5585 1785 5915
rect 2115 5585 2177 5915
rect 1723 5537 2177 5585
rect 2194 5537 2197 5963
rect 1703 5531 2197 5537
rect 2253 5963 2747 5969
rect 2253 5537 2256 5963
rect 2273 5915 2727 5963
rect 2273 5585 2335 5915
rect 2665 5585 2727 5915
rect 2273 5537 2727 5585
rect 2744 5537 2747 5963
rect 2253 5531 2747 5537
rect 2803 5963 3297 5969
rect 2803 5537 2806 5963
rect 2823 5915 3277 5963
rect 2823 5585 2885 5915
rect 3215 5585 3277 5915
rect 2823 5537 3277 5585
rect 3294 5537 3297 5963
rect 2803 5531 3297 5537
rect 3353 5963 3847 5969
rect 3353 5537 3356 5963
rect 3373 5915 3827 5963
rect 3373 5585 3435 5915
rect 3765 5585 3827 5915
rect 3373 5537 3827 5585
rect 3844 5537 3847 5963
rect 3353 5531 3847 5537
rect 3903 5963 4397 5969
rect 3903 5537 3906 5963
rect 3923 5915 4377 5963
rect 3923 5585 3985 5915
rect 4315 5585 4377 5915
rect 3923 5537 4377 5585
rect 4394 5537 4397 5963
rect 3903 5531 4397 5537
rect 4453 5963 4947 5969
rect 4453 5537 4456 5963
rect 4473 5915 4927 5963
rect 4473 5585 4535 5915
rect 4865 5585 4927 5915
rect 4473 5537 4927 5585
rect 4944 5537 4947 5963
rect 4453 5531 4947 5537
rect 5003 5963 5497 5969
rect 5003 5537 5006 5963
rect 5023 5915 5477 5963
rect 5023 5585 5085 5915
rect 5415 5585 5477 5915
rect 5023 5537 5477 5585
rect 5494 5537 5497 5963
rect 5003 5531 5497 5537
rect 5553 5963 6047 5969
rect 5553 5537 5556 5963
rect 5573 5915 6027 5963
rect 5573 5585 5635 5915
rect 5965 5585 6027 5915
rect 5573 5537 6027 5585
rect 6044 5537 6047 5963
rect 5553 5531 6047 5537
rect 6103 5963 6597 5969
rect 6103 5537 6106 5963
rect 6123 5915 6577 5963
rect 6123 5585 6185 5915
rect 6515 5585 6577 5915
rect 6123 5537 6577 5585
rect 6594 5537 6597 5963
rect 6103 5531 6597 5537
rect 6653 5963 7147 5969
rect 6653 5537 6656 5963
rect 6673 5915 7127 5963
rect 6673 5585 6735 5915
rect 7065 5585 7127 5915
rect 6673 5537 7127 5585
rect 7144 5537 7147 5963
rect 6653 5531 7147 5537
rect 7203 5963 7697 5969
rect 7203 5537 7206 5963
rect 7223 5915 7677 5963
rect 7223 5585 7285 5915
rect 7615 5585 7677 5915
rect 7223 5537 7677 5585
rect 7694 5537 7697 5963
rect 7203 5531 7697 5537
rect 7753 5963 8247 5969
rect 7753 5537 7756 5963
rect 7773 5915 8227 5963
rect 7773 5585 7835 5915
rect 8165 5585 8227 5915
rect 7773 5537 8227 5585
rect 8244 5537 8247 5963
rect 7753 5531 8247 5537
rect 8303 5963 8797 5969
rect 8303 5537 8306 5963
rect 8323 5915 8777 5963
rect 8323 5585 8385 5915
rect 8715 5585 8777 5915
rect 8323 5537 8777 5585
rect 8794 5537 8797 5963
rect 8303 5531 8797 5537
rect 8853 5963 9347 5969
rect 8853 5537 8856 5963
rect 8873 5915 9327 5963
rect 8873 5585 8935 5915
rect 9265 5585 9327 5915
rect 8873 5537 9327 5585
rect 9344 5537 9347 5963
rect 8853 5531 9347 5537
rect 9403 5963 9897 5969
rect 9403 5537 9406 5963
rect 9423 5915 9877 5963
rect 9423 5585 9485 5915
rect 9815 5585 9877 5915
rect 9423 5537 9877 5585
rect 9894 5537 9897 5963
rect 9403 5531 9897 5537
rect 9953 5963 10447 5969
rect 9953 5537 9956 5963
rect 9973 5915 10427 5963
rect 9973 5585 10035 5915
rect 10365 5585 10427 5915
rect 9973 5537 10427 5585
rect 10444 5537 10447 5963
rect 9953 5531 10447 5537
rect 10503 5963 10997 5969
rect 10503 5537 10506 5963
rect 10523 5915 10977 5963
rect 10523 5585 10585 5915
rect 10915 5585 10977 5915
rect 10523 5537 10977 5585
rect 10994 5537 10997 5963
rect 10503 5531 10997 5537
rect 11053 5963 11547 5969
rect 11053 5537 11056 5963
rect 11073 5915 11527 5963
rect 11073 5585 11135 5915
rect 11465 5585 11527 5915
rect 11073 5537 11527 5585
rect 11544 5537 11547 5963
rect 11053 5531 11547 5537
rect 11603 5963 12097 5969
rect 11603 5537 11606 5963
rect 11623 5915 12077 5963
rect 11623 5585 11685 5915
rect 12015 5585 12077 5915
rect 11623 5537 12077 5585
rect 12094 5537 12097 5963
rect 11603 5531 12097 5537
rect 12153 5963 12647 5969
rect 12153 5537 12156 5963
rect 12173 5915 12627 5963
rect 12173 5585 12235 5915
rect 12565 5585 12627 5915
rect 12173 5537 12627 5585
rect 12644 5537 12647 5963
rect 12153 5531 12647 5537
rect 12703 5963 13197 5969
rect 12703 5537 12706 5963
rect 12723 5915 13177 5963
rect 12723 5585 12785 5915
rect 13115 5585 13177 5915
rect 12723 5537 13177 5585
rect 13194 5537 13197 5963
rect 12703 5531 13197 5537
rect 13253 5963 13724 5969
rect 13253 5537 13256 5963
rect 13273 5915 13724 5963
rect 13273 5585 13335 5915
rect 13665 5585 13724 5915
rect 13273 5537 13724 5585
rect 13253 5531 13724 5537
rect -474 5526 -26 5531
rect 76 5526 524 5531
rect 626 5526 1074 5531
rect 1176 5526 1624 5531
rect 1726 5526 2174 5531
rect 2276 5526 2724 5531
rect 2826 5526 3274 5531
rect 3376 5526 3824 5531
rect 3926 5526 4374 5531
rect 4476 5526 4924 5531
rect 5026 5526 5474 5531
rect 5576 5526 6024 5531
rect 6126 5526 6574 5531
rect 6676 5526 7124 5531
rect 7226 5526 7674 5531
rect 7776 5526 8224 5531
rect 8326 5526 8774 5531
rect 8876 5526 9324 5531
rect 9426 5526 9874 5531
rect 9976 5526 10424 5531
rect 10526 5526 10974 5531
rect 11076 5526 11524 5531
rect 11626 5526 12074 5531
rect 12176 5526 12624 5531
rect 12726 5526 13174 5531
rect 13276 5526 13724 5531
rect -1025 5500 -725 5519
rect -469 5523 -31 5526
rect -469 5506 -463 5523
rect -37 5506 -31 5523
rect -469 5503 -31 5506
rect 81 5523 519 5526
rect 81 5506 87 5523
rect 513 5506 519 5523
rect 81 5503 519 5506
rect 631 5523 1069 5526
rect 631 5506 637 5523
rect 1063 5506 1069 5523
rect 631 5503 1069 5506
rect 1181 5523 1619 5526
rect 1181 5506 1187 5523
rect 1613 5506 1619 5523
rect 1181 5503 1619 5506
rect 1731 5523 2169 5526
rect 1731 5506 1737 5523
rect 2163 5506 2169 5523
rect 1731 5503 2169 5506
rect 2281 5523 2719 5526
rect 2281 5506 2287 5523
rect 2713 5506 2719 5523
rect 2281 5503 2719 5506
rect 2831 5523 3269 5526
rect 2831 5506 2837 5523
rect 3263 5506 3269 5523
rect 2831 5503 3269 5506
rect 3381 5523 3819 5526
rect 3381 5506 3387 5523
rect 3813 5506 3819 5523
rect 3381 5503 3819 5506
rect 3931 5523 4369 5526
rect 3931 5506 3937 5523
rect 4363 5506 4369 5523
rect 3931 5503 4369 5506
rect 4481 5523 4919 5526
rect 4481 5506 4487 5523
rect 4913 5506 4919 5523
rect 4481 5503 4919 5506
rect 5031 5523 5469 5526
rect 5031 5506 5037 5523
rect 5463 5506 5469 5523
rect 5031 5503 5469 5506
rect 5581 5523 6019 5526
rect 5581 5506 5587 5523
rect 6013 5506 6019 5523
rect 5581 5503 6019 5506
rect 6131 5523 6569 5526
rect 6131 5506 6137 5523
rect 6563 5506 6569 5523
rect 6131 5503 6569 5506
rect 6681 5523 7119 5526
rect 6681 5506 6687 5523
rect 7113 5506 7119 5523
rect 6681 5503 7119 5506
rect 7231 5523 7669 5526
rect 7231 5506 7237 5523
rect 7663 5506 7669 5523
rect 7231 5503 7669 5506
rect 7781 5523 8219 5526
rect 7781 5506 7787 5523
rect 8213 5506 8219 5523
rect 7781 5503 8219 5506
rect 8331 5523 8769 5526
rect 8331 5506 8337 5523
rect 8763 5506 8769 5523
rect 8331 5503 8769 5506
rect 8881 5523 9319 5526
rect 8881 5506 8887 5523
rect 9313 5506 9319 5523
rect 8881 5503 9319 5506
rect 9431 5523 9869 5526
rect 9431 5506 9437 5523
rect 9863 5506 9869 5523
rect 9431 5503 9869 5506
rect 9981 5523 10419 5526
rect 9981 5506 9987 5523
rect 10413 5506 10419 5523
rect 9981 5503 10419 5506
rect 10531 5523 10969 5526
rect 10531 5506 10537 5523
rect 10963 5506 10969 5523
rect 10531 5503 10969 5506
rect 11081 5523 11519 5526
rect 11081 5506 11087 5523
rect 11513 5506 11519 5523
rect 11081 5503 11519 5506
rect 11631 5523 12069 5526
rect 11631 5506 11637 5523
rect 12063 5506 12069 5523
rect 11631 5503 12069 5506
rect 12181 5523 12619 5526
rect 12181 5506 12187 5523
rect 12613 5506 12619 5523
rect 12181 5503 12619 5506
rect 12731 5523 13169 5526
rect 12731 5506 12737 5523
rect 13163 5506 13169 5523
rect 12731 5503 13169 5506
rect 13281 5523 13719 5526
rect 13281 5506 13287 5523
rect 13713 5506 13719 5523
rect 13281 5503 13719 5506
rect 13975 5519 13987 6050
rect 14263 5519 14275 6050
rect 13975 5500 14275 5519
rect -1025 4969 -1013 5500
rect -737 4969 -725 5500
rect -550 5492 -500 5500
rect -550 5458 -542 5492
rect -508 5458 -500 5492
rect -550 5450 -500 5458
rect 0 5492 50 5500
rect 0 5458 8 5492
rect 42 5458 50 5492
rect 0 5450 50 5458
rect 550 5492 600 5500
rect 550 5458 558 5492
rect 592 5458 600 5492
rect 550 5450 600 5458
rect 1100 5492 1150 5500
rect 1100 5458 1108 5492
rect 1142 5458 1150 5492
rect 1100 5450 1150 5458
rect 1650 5492 1700 5500
rect 1650 5458 1658 5492
rect 1692 5458 1700 5492
rect 1650 5450 1700 5458
rect 2200 5492 2250 5500
rect 2200 5458 2208 5492
rect 2242 5458 2250 5492
rect 2200 5450 2250 5458
rect 2750 5492 2800 5500
rect 2750 5458 2758 5492
rect 2792 5458 2800 5492
rect 2750 5450 2800 5458
rect 3300 5492 3350 5500
rect 3300 5458 3308 5492
rect 3342 5458 3350 5492
rect 3300 5450 3350 5458
rect 3850 5492 3900 5500
rect 3850 5458 3858 5492
rect 3892 5458 3900 5492
rect 3850 5450 3900 5458
rect 4400 5492 4450 5500
rect 4400 5458 4408 5492
rect 4442 5458 4450 5492
rect 4400 5450 4450 5458
rect 4950 5492 5000 5500
rect 4950 5458 4958 5492
rect 4992 5458 5000 5492
rect 4950 5450 5000 5458
rect 5500 5492 5550 5500
rect 5500 5458 5508 5492
rect 5542 5458 5550 5492
rect 5500 5450 5550 5458
rect 6050 5492 6100 5500
rect 6050 5458 6058 5492
rect 6092 5458 6100 5492
rect 6050 5450 6100 5458
rect 6600 5492 6650 5500
rect 6600 5458 6608 5492
rect 6642 5458 6650 5492
rect 6600 5450 6650 5458
rect 7150 5492 7200 5500
rect 7150 5458 7158 5492
rect 7192 5458 7200 5492
rect 7150 5450 7200 5458
rect 7700 5492 7750 5500
rect 7700 5458 7708 5492
rect 7742 5458 7750 5492
rect 7700 5450 7750 5458
rect 8250 5492 8300 5500
rect 8250 5458 8258 5492
rect 8292 5458 8300 5492
rect 8250 5450 8300 5458
rect 8800 5492 8850 5500
rect 8800 5458 8808 5492
rect 8842 5458 8850 5492
rect 8800 5450 8850 5458
rect 9350 5492 9400 5500
rect 9350 5458 9358 5492
rect 9392 5458 9400 5492
rect 9350 5450 9400 5458
rect 9900 5492 9950 5500
rect 9900 5458 9908 5492
rect 9942 5458 9950 5492
rect 9900 5450 9950 5458
rect 10450 5492 10500 5500
rect 10450 5458 10458 5492
rect 10492 5458 10500 5492
rect 10450 5450 10500 5458
rect 11000 5492 11050 5500
rect 11000 5458 11008 5492
rect 11042 5458 11050 5492
rect 11000 5450 11050 5458
rect 11550 5492 11600 5500
rect 11550 5458 11558 5492
rect 11592 5458 11600 5492
rect 11550 5450 11600 5458
rect 12100 5492 12150 5500
rect 12100 5458 12108 5492
rect 12142 5458 12150 5492
rect 12100 5450 12150 5458
rect 12650 5492 12700 5500
rect 12650 5458 12658 5492
rect 12692 5458 12700 5492
rect 12650 5450 12700 5458
rect 13200 5492 13250 5500
rect 13200 5458 13208 5492
rect 13242 5458 13250 5492
rect 13200 5450 13250 5458
rect 13750 5492 13800 5500
rect 13750 5458 13758 5492
rect 13792 5458 13800 5492
rect 13750 5450 13800 5458
rect -469 5444 -31 5447
rect -469 5427 -463 5444
rect -37 5427 -31 5444
rect -469 5424 -31 5427
rect 81 5444 519 5447
rect 81 5427 87 5444
rect 513 5427 519 5444
rect 81 5424 519 5427
rect 631 5444 1069 5447
rect 631 5427 637 5444
rect 1063 5427 1069 5444
rect 631 5424 1069 5427
rect 1181 5444 1619 5447
rect 1181 5427 1187 5444
rect 1613 5427 1619 5444
rect 1181 5424 1619 5427
rect 1731 5444 2169 5447
rect 1731 5427 1737 5444
rect 2163 5427 2169 5444
rect 1731 5424 2169 5427
rect 2281 5444 2719 5447
rect 2281 5427 2287 5444
rect 2713 5427 2719 5444
rect 2281 5424 2719 5427
rect 2831 5444 3269 5447
rect 2831 5427 2837 5444
rect 3263 5427 3269 5444
rect 2831 5424 3269 5427
rect 3381 5444 3819 5447
rect 3381 5427 3387 5444
rect 3813 5427 3819 5444
rect 3381 5424 3819 5427
rect 3931 5444 4369 5447
rect 3931 5427 3937 5444
rect 4363 5427 4369 5444
rect 3931 5424 4369 5427
rect 4481 5444 4919 5447
rect 4481 5427 4487 5444
rect 4913 5427 4919 5444
rect 4481 5424 4919 5427
rect 5031 5444 5469 5447
rect 5031 5427 5037 5444
rect 5463 5427 5469 5444
rect 5031 5424 5469 5427
rect 5581 5444 6019 5447
rect 5581 5427 5587 5444
rect 6013 5427 6019 5444
rect 5581 5424 6019 5427
rect 6131 5444 6569 5447
rect 6131 5427 6137 5444
rect 6563 5427 6569 5444
rect 6131 5424 6569 5427
rect 6681 5444 7119 5447
rect 6681 5427 6687 5444
rect 7113 5427 7119 5444
rect 6681 5424 7119 5427
rect 7231 5444 7669 5447
rect 7231 5427 7237 5444
rect 7663 5427 7669 5444
rect 7231 5424 7669 5427
rect 7781 5444 8219 5447
rect 7781 5427 7787 5444
rect 8213 5427 8219 5444
rect 7781 5424 8219 5427
rect 8331 5444 8769 5447
rect 8331 5427 8337 5444
rect 8763 5427 8769 5444
rect 8331 5424 8769 5427
rect 8881 5444 9319 5447
rect 8881 5427 8887 5444
rect 9313 5427 9319 5444
rect 8881 5424 9319 5427
rect 9431 5444 9869 5447
rect 9431 5427 9437 5444
rect 9863 5427 9869 5444
rect 9431 5424 9869 5427
rect 9981 5444 10419 5447
rect 9981 5427 9987 5444
rect 10413 5427 10419 5444
rect 9981 5424 10419 5427
rect 10531 5444 10969 5447
rect 10531 5427 10537 5444
rect 10963 5427 10969 5444
rect 10531 5424 10969 5427
rect 11081 5444 11519 5447
rect 11081 5427 11087 5444
rect 11513 5427 11519 5444
rect 11081 5424 11519 5427
rect 11631 5444 12069 5447
rect 11631 5427 11637 5444
rect 12063 5427 12069 5444
rect 11631 5424 12069 5427
rect 12181 5444 12619 5447
rect 12181 5427 12187 5444
rect 12613 5427 12619 5444
rect 12181 5424 12619 5427
rect 12731 5444 13169 5447
rect 12731 5427 12737 5444
rect 13163 5427 13169 5444
rect 12731 5424 13169 5427
rect 13281 5444 13719 5447
rect 13281 5427 13287 5444
rect 13713 5427 13719 5444
rect 13281 5424 13719 5427
rect -474 5419 -26 5424
rect 76 5419 524 5424
rect 626 5419 1074 5424
rect 1176 5419 1624 5424
rect 1726 5419 2174 5424
rect 2276 5419 2724 5424
rect 2826 5419 3274 5424
rect 3376 5419 3824 5424
rect 3926 5419 4374 5424
rect 4476 5419 4924 5424
rect 5026 5419 5474 5424
rect 5576 5419 6024 5424
rect 6126 5419 6574 5424
rect 6676 5419 7124 5424
rect 7226 5419 7674 5424
rect 7776 5419 8224 5424
rect 8326 5419 8774 5424
rect 8876 5419 9324 5424
rect 9426 5419 9874 5424
rect 9976 5419 10424 5424
rect 10526 5419 10974 5424
rect 11076 5419 11524 5424
rect 11626 5419 12074 5424
rect 12176 5419 12624 5424
rect 12726 5419 13174 5424
rect 13276 5419 13724 5424
rect -474 5413 -3 5419
rect -474 5365 -23 5413
rect -474 5035 -415 5365
rect -85 5035 -23 5365
rect -474 4987 -23 5035
rect -6 4987 -3 5413
rect -474 4981 -3 4987
rect 53 5413 547 5419
rect 53 4987 56 5413
rect 73 5365 527 5413
rect 73 5035 135 5365
rect 465 5035 527 5365
rect 73 4987 527 5035
rect 544 4987 547 5413
rect 53 4981 547 4987
rect 603 5413 1097 5419
rect 603 4987 606 5413
rect 623 5365 1077 5413
rect 623 5035 685 5365
rect 1015 5035 1077 5365
rect 623 4987 1077 5035
rect 1094 4987 1097 5413
rect 603 4981 1097 4987
rect 1153 5413 1647 5419
rect 1153 4987 1156 5413
rect 1173 5365 1627 5413
rect 1173 5035 1235 5365
rect 1565 5035 1627 5365
rect 1173 4987 1627 5035
rect 1644 4987 1647 5413
rect 1153 4981 1647 4987
rect 1703 5413 2197 5419
rect 1703 4987 1706 5413
rect 1723 5365 2177 5413
rect 1723 5035 1785 5365
rect 2115 5035 2177 5365
rect 1723 4987 2177 5035
rect 2194 4987 2197 5413
rect 1703 4981 2197 4987
rect 2253 5413 2747 5419
rect 2253 4987 2256 5413
rect 2273 5365 2727 5413
rect 2273 5035 2335 5365
rect 2665 5035 2727 5365
rect 2273 4987 2727 5035
rect 2744 4987 2747 5413
rect 2253 4981 2747 4987
rect 2803 5413 3297 5419
rect 2803 4987 2806 5413
rect 2823 5365 3277 5413
rect 2823 5035 2885 5365
rect 3215 5035 3277 5365
rect 2823 4987 3277 5035
rect 3294 4987 3297 5413
rect 2803 4981 3297 4987
rect 3353 5413 3847 5419
rect 3353 4987 3356 5413
rect 3373 5365 3827 5413
rect 3373 5035 3435 5365
rect 3765 5035 3827 5365
rect 3373 4987 3827 5035
rect 3844 4987 3847 5413
rect 3353 4981 3847 4987
rect 3903 5413 4397 5419
rect 3903 4987 3906 5413
rect 3923 5365 4377 5413
rect 3923 5035 3985 5365
rect 4315 5035 4377 5365
rect 3923 4987 4377 5035
rect 4394 4987 4397 5413
rect 3903 4981 4397 4987
rect 4453 5413 4947 5419
rect 4453 4987 4456 5413
rect 4473 5365 4927 5413
rect 4473 5035 4535 5365
rect 4865 5035 4927 5365
rect 4473 4987 4927 5035
rect 4944 4987 4947 5413
rect 4453 4981 4947 4987
rect 5003 5413 5497 5419
rect 5003 4987 5006 5413
rect 5023 5365 5477 5413
rect 5023 5035 5085 5365
rect 5415 5035 5477 5365
rect 5023 4987 5477 5035
rect 5494 4987 5497 5413
rect 5003 4981 5497 4987
rect 5553 5413 6047 5419
rect 5553 4987 5556 5413
rect 5573 5365 6027 5413
rect 5573 5035 5635 5365
rect 5965 5035 6027 5365
rect 5573 4987 6027 5035
rect 6044 4987 6047 5413
rect 5553 4981 6047 4987
rect 6103 5413 6597 5419
rect 6103 4987 6106 5413
rect 6123 5365 6577 5413
rect 6123 5035 6185 5365
rect 6515 5035 6577 5365
rect 6123 4987 6577 5035
rect 6594 4987 6597 5413
rect 6103 4981 6597 4987
rect 6653 5413 7147 5419
rect 6653 4987 6656 5413
rect 6673 5365 7127 5413
rect 6673 5035 6735 5365
rect 7065 5035 7127 5365
rect 6673 4987 7127 5035
rect 7144 4987 7147 5413
rect 6653 4981 7147 4987
rect 7203 5413 7697 5419
rect 7203 4987 7206 5413
rect 7223 5365 7677 5413
rect 7223 5035 7285 5365
rect 7615 5035 7677 5365
rect 7223 4987 7677 5035
rect 7694 4987 7697 5413
rect 7203 4981 7697 4987
rect 7753 5413 8247 5419
rect 7753 4987 7756 5413
rect 7773 5365 8227 5413
rect 7773 5035 7835 5365
rect 8165 5035 8227 5365
rect 7773 4987 8227 5035
rect 8244 4987 8247 5413
rect 7753 4981 8247 4987
rect 8303 5413 8797 5419
rect 8303 4987 8306 5413
rect 8323 5365 8777 5413
rect 8323 5035 8385 5365
rect 8715 5035 8777 5365
rect 8323 4987 8777 5035
rect 8794 4987 8797 5413
rect 8303 4981 8797 4987
rect 8853 5413 9347 5419
rect 8853 4987 8856 5413
rect 8873 5365 9327 5413
rect 8873 5035 8935 5365
rect 9265 5035 9327 5365
rect 8873 4987 9327 5035
rect 9344 4987 9347 5413
rect 8853 4981 9347 4987
rect 9403 5413 9897 5419
rect 9403 4987 9406 5413
rect 9423 5365 9877 5413
rect 9423 5035 9485 5365
rect 9815 5035 9877 5365
rect 9423 4987 9877 5035
rect 9894 4987 9897 5413
rect 9403 4981 9897 4987
rect 9953 5413 10447 5419
rect 9953 4987 9956 5413
rect 9973 5365 10427 5413
rect 9973 5035 10035 5365
rect 10365 5035 10427 5365
rect 9973 4987 10427 5035
rect 10444 4987 10447 5413
rect 9953 4981 10447 4987
rect 10503 5413 10997 5419
rect 10503 4987 10506 5413
rect 10523 5365 10977 5413
rect 10523 5035 10585 5365
rect 10915 5035 10977 5365
rect 10523 4987 10977 5035
rect 10994 4987 10997 5413
rect 10503 4981 10997 4987
rect 11053 5413 11547 5419
rect 11053 4987 11056 5413
rect 11073 5365 11527 5413
rect 11073 5035 11135 5365
rect 11465 5035 11527 5365
rect 11073 4987 11527 5035
rect 11544 4987 11547 5413
rect 11053 4981 11547 4987
rect 11603 5413 12097 5419
rect 11603 4987 11606 5413
rect 11623 5365 12077 5413
rect 11623 5035 11685 5365
rect 12015 5035 12077 5365
rect 11623 4987 12077 5035
rect 12094 4987 12097 5413
rect 11603 4981 12097 4987
rect 12153 5413 12647 5419
rect 12153 4987 12156 5413
rect 12173 5365 12627 5413
rect 12173 5035 12235 5365
rect 12565 5035 12627 5365
rect 12173 4987 12627 5035
rect 12644 4987 12647 5413
rect 12153 4981 12647 4987
rect 12703 5413 13197 5419
rect 12703 4987 12706 5413
rect 12723 5365 13177 5413
rect 12723 5035 12785 5365
rect 13115 5035 13177 5365
rect 12723 4987 13177 5035
rect 13194 4987 13197 5413
rect 12703 4981 13197 4987
rect 13253 5413 13724 5419
rect 13253 4987 13256 5413
rect 13273 5365 13724 5413
rect 13273 5035 13335 5365
rect 13665 5035 13724 5365
rect 13273 4987 13724 5035
rect 13253 4981 13724 4987
rect -474 4976 -26 4981
rect 76 4976 524 4981
rect 626 4976 1074 4981
rect 1176 4976 1624 4981
rect 1726 4976 2174 4981
rect 2276 4976 2724 4981
rect 2826 4976 3274 4981
rect 3376 4976 3824 4981
rect 3926 4976 4374 4981
rect 4476 4976 4924 4981
rect 5026 4976 5474 4981
rect 5576 4976 6024 4981
rect 6126 4976 6574 4981
rect 6676 4976 7124 4981
rect 7226 4976 7674 4981
rect 7776 4976 8224 4981
rect 8326 4976 8774 4981
rect 8876 4976 9324 4981
rect 9426 4976 9874 4981
rect 9976 4976 10424 4981
rect 10526 4976 10974 4981
rect 11076 4976 11524 4981
rect 11626 4976 12074 4981
rect 12176 4976 12624 4981
rect 12726 4976 13174 4981
rect 13276 4976 13724 4981
rect -1025 4950 -725 4969
rect -469 4973 -31 4976
rect -469 4956 -463 4973
rect -37 4956 -31 4973
rect -469 4953 -31 4956
rect 81 4973 519 4976
rect 81 4956 87 4973
rect 513 4956 519 4973
rect 81 4953 519 4956
rect 631 4973 1069 4976
rect 631 4956 637 4973
rect 1063 4956 1069 4973
rect 631 4953 1069 4956
rect 1181 4973 1619 4976
rect 1181 4956 1187 4973
rect 1613 4956 1619 4973
rect 1181 4953 1619 4956
rect 1731 4973 2169 4976
rect 1731 4956 1737 4973
rect 2163 4956 2169 4973
rect 1731 4953 2169 4956
rect 2281 4973 2719 4976
rect 2281 4956 2287 4973
rect 2713 4956 2719 4973
rect 2281 4953 2719 4956
rect 2831 4973 3269 4976
rect 2831 4956 2837 4973
rect 3263 4956 3269 4973
rect 2831 4953 3269 4956
rect 3381 4973 3819 4976
rect 3381 4956 3387 4973
rect 3813 4956 3819 4973
rect 3381 4953 3819 4956
rect 3931 4973 4369 4976
rect 3931 4956 3937 4973
rect 4363 4956 4369 4973
rect 3931 4953 4369 4956
rect 4481 4973 4919 4976
rect 4481 4956 4487 4973
rect 4913 4956 4919 4973
rect 4481 4953 4919 4956
rect 5031 4973 5469 4976
rect 5031 4956 5037 4973
rect 5463 4956 5469 4973
rect 5031 4953 5469 4956
rect 5581 4973 6019 4976
rect 5581 4956 5587 4973
rect 6013 4956 6019 4973
rect 5581 4953 6019 4956
rect 6131 4973 6569 4976
rect 6131 4956 6137 4973
rect 6563 4956 6569 4973
rect 6131 4953 6569 4956
rect 6681 4973 7119 4976
rect 6681 4956 6687 4973
rect 7113 4956 7119 4973
rect 6681 4953 7119 4956
rect 7231 4973 7669 4976
rect 7231 4956 7237 4973
rect 7663 4956 7669 4973
rect 7231 4953 7669 4956
rect 7781 4973 8219 4976
rect 7781 4956 7787 4973
rect 8213 4956 8219 4973
rect 7781 4953 8219 4956
rect 8331 4973 8769 4976
rect 8331 4956 8337 4973
rect 8763 4956 8769 4973
rect 8331 4953 8769 4956
rect 8881 4973 9319 4976
rect 8881 4956 8887 4973
rect 9313 4956 9319 4973
rect 8881 4953 9319 4956
rect 9431 4973 9869 4976
rect 9431 4956 9437 4973
rect 9863 4956 9869 4973
rect 9431 4953 9869 4956
rect 9981 4973 10419 4976
rect 9981 4956 9987 4973
rect 10413 4956 10419 4973
rect 9981 4953 10419 4956
rect 10531 4973 10969 4976
rect 10531 4956 10537 4973
rect 10963 4956 10969 4973
rect 10531 4953 10969 4956
rect 11081 4973 11519 4976
rect 11081 4956 11087 4973
rect 11513 4956 11519 4973
rect 11081 4953 11519 4956
rect 11631 4973 12069 4976
rect 11631 4956 11637 4973
rect 12063 4956 12069 4973
rect 11631 4953 12069 4956
rect 12181 4973 12619 4976
rect 12181 4956 12187 4973
rect 12613 4956 12619 4973
rect 12181 4953 12619 4956
rect 12731 4973 13169 4976
rect 12731 4956 12737 4973
rect 13163 4956 13169 4973
rect 12731 4953 13169 4956
rect 13281 4973 13719 4976
rect 13281 4956 13287 4973
rect 13713 4956 13719 4973
rect 13281 4953 13719 4956
rect 13975 4969 13987 5500
rect 14263 4969 14275 5500
rect 13975 4950 14275 4969
rect -1025 4419 -1013 4950
rect -737 4419 -725 4950
rect -550 4942 -500 4950
rect -550 4908 -542 4942
rect -508 4908 -500 4942
rect -550 4900 -500 4908
rect 0 4942 50 4950
rect 0 4908 8 4942
rect 42 4908 50 4942
rect 0 4900 50 4908
rect 550 4942 600 4950
rect 550 4908 558 4942
rect 592 4908 600 4942
rect 550 4900 600 4908
rect 1100 4942 1150 4950
rect 1100 4908 1108 4942
rect 1142 4908 1150 4942
rect 1100 4900 1150 4908
rect 1650 4942 1700 4950
rect 1650 4908 1658 4942
rect 1692 4908 1700 4942
rect 1650 4900 1700 4908
rect 2200 4942 2250 4950
rect 2200 4908 2208 4942
rect 2242 4908 2250 4942
rect 2200 4900 2250 4908
rect 2750 4942 2800 4950
rect 2750 4908 2758 4942
rect 2792 4908 2800 4942
rect 2750 4900 2800 4908
rect 3300 4942 3350 4950
rect 3300 4908 3308 4942
rect 3342 4908 3350 4942
rect 3300 4900 3350 4908
rect 3850 4942 3900 4950
rect 3850 4908 3858 4942
rect 3892 4908 3900 4942
rect 3850 4900 3900 4908
rect 4400 4942 4450 4950
rect 4400 4908 4408 4942
rect 4442 4908 4450 4942
rect 4400 4900 4450 4908
rect 4950 4942 5000 4950
rect 4950 4908 4958 4942
rect 4992 4908 5000 4942
rect 4950 4900 5000 4908
rect 5500 4942 5550 4950
rect 5500 4908 5508 4942
rect 5542 4908 5550 4942
rect 5500 4900 5550 4908
rect 6050 4942 6100 4950
rect 6050 4908 6058 4942
rect 6092 4908 6100 4942
rect 6050 4900 6100 4908
rect 6600 4942 6650 4950
rect 6600 4908 6608 4942
rect 6642 4908 6650 4942
rect 6600 4900 6650 4908
rect 7150 4942 7200 4950
rect 7150 4908 7158 4942
rect 7192 4908 7200 4942
rect 7150 4900 7200 4908
rect 7700 4942 7750 4950
rect 7700 4908 7708 4942
rect 7742 4908 7750 4942
rect 7700 4900 7750 4908
rect 8250 4942 8300 4950
rect 8250 4908 8258 4942
rect 8292 4908 8300 4942
rect 8250 4900 8300 4908
rect 8800 4942 8850 4950
rect 8800 4908 8808 4942
rect 8842 4908 8850 4942
rect 8800 4900 8850 4908
rect 9350 4942 9400 4950
rect 9350 4908 9358 4942
rect 9392 4908 9400 4942
rect 9350 4900 9400 4908
rect 9900 4942 9950 4950
rect 9900 4908 9908 4942
rect 9942 4908 9950 4942
rect 9900 4900 9950 4908
rect 10450 4942 10500 4950
rect 10450 4908 10458 4942
rect 10492 4908 10500 4942
rect 10450 4900 10500 4908
rect 11000 4942 11050 4950
rect 11000 4908 11008 4942
rect 11042 4908 11050 4942
rect 11000 4900 11050 4908
rect 11550 4942 11600 4950
rect 11550 4908 11558 4942
rect 11592 4908 11600 4942
rect 11550 4900 11600 4908
rect 12100 4942 12150 4950
rect 12100 4908 12108 4942
rect 12142 4908 12150 4942
rect 12100 4900 12150 4908
rect 12650 4942 12700 4950
rect 12650 4908 12658 4942
rect 12692 4908 12700 4942
rect 12650 4900 12700 4908
rect 13200 4942 13250 4950
rect 13200 4908 13208 4942
rect 13242 4908 13250 4942
rect 13200 4900 13250 4908
rect 13750 4942 13800 4950
rect 13750 4908 13758 4942
rect 13792 4908 13800 4942
rect 13750 4900 13800 4908
rect -469 4894 -31 4897
rect -469 4877 -463 4894
rect -37 4877 -31 4894
rect -469 4874 -31 4877
rect 81 4894 519 4897
rect 81 4877 87 4894
rect 513 4877 519 4894
rect 81 4874 519 4877
rect 631 4894 1069 4897
rect 631 4877 637 4894
rect 1063 4877 1069 4894
rect 631 4874 1069 4877
rect 1181 4894 1619 4897
rect 1181 4877 1187 4894
rect 1613 4877 1619 4894
rect 1181 4874 1619 4877
rect 1731 4894 2169 4897
rect 1731 4877 1737 4894
rect 2163 4877 2169 4894
rect 1731 4874 2169 4877
rect 2281 4894 2719 4897
rect 2281 4877 2287 4894
rect 2713 4877 2719 4894
rect 2281 4874 2719 4877
rect 2831 4894 3269 4897
rect 2831 4877 2837 4894
rect 3263 4877 3269 4894
rect 2831 4874 3269 4877
rect 3381 4894 3819 4897
rect 3381 4877 3387 4894
rect 3813 4877 3819 4894
rect 3381 4874 3819 4877
rect 3931 4894 4369 4897
rect 3931 4877 3937 4894
rect 4363 4877 4369 4894
rect 3931 4874 4369 4877
rect 4481 4894 4919 4897
rect 4481 4877 4487 4894
rect 4913 4877 4919 4894
rect 4481 4874 4919 4877
rect 5031 4894 5469 4897
rect 5031 4877 5037 4894
rect 5463 4877 5469 4894
rect 5031 4874 5469 4877
rect 5581 4894 6019 4897
rect 5581 4877 5587 4894
rect 6013 4877 6019 4894
rect 5581 4874 6019 4877
rect 6131 4894 6569 4897
rect 6131 4877 6137 4894
rect 6563 4877 6569 4894
rect 6131 4874 6569 4877
rect 6681 4894 7119 4897
rect 6681 4877 6687 4894
rect 7113 4877 7119 4894
rect 6681 4874 7119 4877
rect 7231 4894 7669 4897
rect 7231 4877 7237 4894
rect 7663 4877 7669 4894
rect 7231 4874 7669 4877
rect 7781 4894 8219 4897
rect 7781 4877 7787 4894
rect 8213 4877 8219 4894
rect 7781 4874 8219 4877
rect 8331 4894 8769 4897
rect 8331 4877 8337 4894
rect 8763 4877 8769 4894
rect 8331 4874 8769 4877
rect 8881 4894 9319 4897
rect 8881 4877 8887 4894
rect 9313 4877 9319 4894
rect 8881 4874 9319 4877
rect 9431 4894 9869 4897
rect 9431 4877 9437 4894
rect 9863 4877 9869 4894
rect 9431 4874 9869 4877
rect 9981 4894 10419 4897
rect 9981 4877 9987 4894
rect 10413 4877 10419 4894
rect 9981 4874 10419 4877
rect 10531 4894 10969 4897
rect 10531 4877 10537 4894
rect 10963 4877 10969 4894
rect 10531 4874 10969 4877
rect 11081 4894 11519 4897
rect 11081 4877 11087 4894
rect 11513 4877 11519 4894
rect 11081 4874 11519 4877
rect 11631 4894 12069 4897
rect 11631 4877 11637 4894
rect 12063 4877 12069 4894
rect 11631 4874 12069 4877
rect 12181 4894 12619 4897
rect 12181 4877 12187 4894
rect 12613 4877 12619 4894
rect 12181 4874 12619 4877
rect 12731 4894 13169 4897
rect 12731 4877 12737 4894
rect 13163 4877 13169 4894
rect 12731 4874 13169 4877
rect 13281 4894 13719 4897
rect 13281 4877 13287 4894
rect 13713 4877 13719 4894
rect 13281 4874 13719 4877
rect -474 4869 -26 4874
rect 76 4869 524 4874
rect 626 4869 1074 4874
rect 1176 4869 1624 4874
rect 1726 4869 2174 4874
rect 2276 4869 2724 4874
rect 2826 4869 3274 4874
rect 3376 4869 3824 4874
rect 3926 4869 4374 4874
rect 4476 4869 4924 4874
rect 5026 4869 5474 4874
rect 5576 4869 6024 4874
rect 6126 4869 6574 4874
rect 6676 4869 7124 4874
rect 7226 4869 7674 4874
rect 7776 4869 8224 4874
rect 8326 4869 8774 4874
rect 8876 4869 9324 4874
rect 9426 4869 9874 4874
rect 9976 4869 10424 4874
rect 10526 4869 10974 4874
rect 11076 4869 11524 4874
rect 11626 4869 12074 4874
rect 12176 4869 12624 4874
rect 12726 4869 13174 4874
rect 13276 4869 13724 4874
rect -474 4863 -3 4869
rect -474 4815 -23 4863
rect -474 4485 -415 4815
rect -85 4485 -23 4815
rect -474 4437 -23 4485
rect -6 4437 -3 4863
rect -474 4431 -3 4437
rect 53 4863 547 4869
rect 53 4437 56 4863
rect 73 4815 527 4863
rect 73 4485 135 4815
rect 465 4485 527 4815
rect 73 4437 527 4485
rect 544 4437 547 4863
rect 53 4431 547 4437
rect 603 4863 1097 4869
rect 603 4437 606 4863
rect 623 4815 1077 4863
rect 623 4485 685 4815
rect 1015 4485 1077 4815
rect 623 4437 1077 4485
rect 1094 4437 1097 4863
rect 603 4431 1097 4437
rect 1153 4863 1647 4869
rect 1153 4437 1156 4863
rect 1173 4815 1627 4863
rect 1173 4485 1235 4815
rect 1565 4485 1627 4815
rect 1173 4437 1627 4485
rect 1644 4437 1647 4863
rect 1153 4431 1647 4437
rect 1703 4863 2197 4869
rect 1703 4437 1706 4863
rect 1723 4815 2177 4863
rect 1723 4485 1785 4815
rect 2115 4485 2177 4815
rect 1723 4437 2177 4485
rect 2194 4437 2197 4863
rect 1703 4431 2197 4437
rect 2253 4863 2747 4869
rect 2253 4437 2256 4863
rect 2273 4815 2727 4863
rect 2273 4485 2335 4815
rect 2665 4485 2727 4815
rect 2273 4437 2727 4485
rect 2744 4437 2747 4863
rect 2253 4431 2747 4437
rect 2803 4863 3297 4869
rect 2803 4437 2806 4863
rect 2823 4815 3277 4863
rect 2823 4485 2885 4815
rect 3215 4485 3277 4815
rect 2823 4437 3277 4485
rect 3294 4437 3297 4863
rect 2803 4431 3297 4437
rect 3353 4863 3847 4869
rect 3353 4437 3356 4863
rect 3373 4815 3827 4863
rect 3373 4485 3435 4815
rect 3765 4485 3827 4815
rect 3373 4437 3827 4485
rect 3844 4437 3847 4863
rect 3353 4431 3847 4437
rect 3903 4863 4397 4869
rect 3903 4437 3906 4863
rect 3923 4815 4377 4863
rect 3923 4485 3985 4815
rect 4315 4485 4377 4815
rect 3923 4437 4377 4485
rect 4394 4437 4397 4863
rect 3903 4431 4397 4437
rect 4453 4863 4947 4869
rect 4453 4437 4456 4863
rect 4473 4815 4927 4863
rect 4473 4485 4535 4815
rect 4865 4485 4927 4815
rect 4473 4437 4927 4485
rect 4944 4437 4947 4863
rect 4453 4431 4947 4437
rect 5003 4863 5497 4869
rect 5003 4437 5006 4863
rect 5023 4815 5477 4863
rect 5023 4485 5085 4815
rect 5415 4485 5477 4815
rect 5023 4437 5477 4485
rect 5494 4437 5497 4863
rect 5003 4431 5497 4437
rect 5553 4863 6047 4869
rect 5553 4437 5556 4863
rect 5573 4815 6027 4863
rect 5573 4485 5635 4815
rect 5965 4485 6027 4815
rect 5573 4437 6027 4485
rect 6044 4437 6047 4863
rect 5553 4431 6047 4437
rect 6103 4863 6597 4869
rect 6103 4437 6106 4863
rect 6123 4815 6577 4863
rect 6123 4485 6185 4815
rect 6515 4485 6577 4815
rect 6123 4437 6577 4485
rect 6594 4437 6597 4863
rect 6103 4431 6597 4437
rect 6653 4863 7147 4869
rect 6653 4437 6656 4863
rect 6673 4815 7127 4863
rect 6673 4485 6735 4815
rect 7065 4485 7127 4815
rect 6673 4437 7127 4485
rect 7144 4437 7147 4863
rect 6653 4431 7147 4437
rect 7203 4863 7697 4869
rect 7203 4437 7206 4863
rect 7223 4815 7677 4863
rect 7223 4485 7285 4815
rect 7615 4485 7677 4815
rect 7223 4437 7677 4485
rect 7694 4437 7697 4863
rect 7203 4431 7697 4437
rect 7753 4863 8247 4869
rect 7753 4437 7756 4863
rect 7773 4815 8227 4863
rect 7773 4485 7835 4815
rect 8165 4485 8227 4815
rect 7773 4437 8227 4485
rect 8244 4437 8247 4863
rect 7753 4431 8247 4437
rect 8303 4863 8797 4869
rect 8303 4437 8306 4863
rect 8323 4815 8777 4863
rect 8323 4485 8385 4815
rect 8715 4485 8777 4815
rect 8323 4437 8777 4485
rect 8794 4437 8797 4863
rect 8303 4431 8797 4437
rect 8853 4863 9347 4869
rect 8853 4437 8856 4863
rect 8873 4815 9327 4863
rect 8873 4485 8935 4815
rect 9265 4485 9327 4815
rect 8873 4437 9327 4485
rect 9344 4437 9347 4863
rect 8853 4431 9347 4437
rect 9403 4863 9897 4869
rect 9403 4437 9406 4863
rect 9423 4815 9877 4863
rect 9423 4485 9485 4815
rect 9815 4485 9877 4815
rect 9423 4437 9877 4485
rect 9894 4437 9897 4863
rect 9403 4431 9897 4437
rect 9953 4863 10447 4869
rect 9953 4437 9956 4863
rect 9973 4815 10427 4863
rect 9973 4485 10035 4815
rect 10365 4485 10427 4815
rect 9973 4437 10427 4485
rect 10444 4437 10447 4863
rect 9953 4431 10447 4437
rect 10503 4863 10997 4869
rect 10503 4437 10506 4863
rect 10523 4815 10977 4863
rect 10523 4485 10585 4815
rect 10915 4485 10977 4815
rect 10523 4437 10977 4485
rect 10994 4437 10997 4863
rect 10503 4431 10997 4437
rect 11053 4863 11547 4869
rect 11053 4437 11056 4863
rect 11073 4815 11527 4863
rect 11073 4485 11135 4815
rect 11465 4485 11527 4815
rect 11073 4437 11527 4485
rect 11544 4437 11547 4863
rect 11053 4431 11547 4437
rect 11603 4863 12097 4869
rect 11603 4437 11606 4863
rect 11623 4815 12077 4863
rect 11623 4485 11685 4815
rect 12015 4485 12077 4815
rect 11623 4437 12077 4485
rect 12094 4437 12097 4863
rect 11603 4431 12097 4437
rect 12153 4863 12647 4869
rect 12153 4437 12156 4863
rect 12173 4815 12627 4863
rect 12173 4485 12235 4815
rect 12565 4485 12627 4815
rect 12173 4437 12627 4485
rect 12644 4437 12647 4863
rect 12153 4431 12647 4437
rect 12703 4863 13197 4869
rect 12703 4437 12706 4863
rect 12723 4815 13177 4863
rect 12723 4485 12785 4815
rect 13115 4485 13177 4815
rect 12723 4437 13177 4485
rect 13194 4437 13197 4863
rect 12703 4431 13197 4437
rect 13253 4863 13724 4869
rect 13253 4437 13256 4863
rect 13273 4815 13724 4863
rect 13273 4485 13335 4815
rect 13665 4485 13724 4815
rect 13273 4437 13724 4485
rect 13253 4431 13724 4437
rect -474 4426 -26 4431
rect 76 4426 524 4431
rect 626 4426 1074 4431
rect 1176 4426 1624 4431
rect 1726 4426 2174 4431
rect 2276 4426 2724 4431
rect 2826 4426 3274 4431
rect 3376 4426 3824 4431
rect 3926 4426 4374 4431
rect 4476 4426 4924 4431
rect 5026 4426 5474 4431
rect 5576 4426 6024 4431
rect 6126 4426 6574 4431
rect 6676 4426 7124 4431
rect 7226 4426 7674 4431
rect 7776 4426 8224 4431
rect 8326 4426 8774 4431
rect 8876 4426 9324 4431
rect 9426 4426 9874 4431
rect 9976 4426 10424 4431
rect 10526 4426 10974 4431
rect 11076 4426 11524 4431
rect 11626 4426 12074 4431
rect 12176 4426 12624 4431
rect 12726 4426 13174 4431
rect 13276 4426 13724 4431
rect -1025 4400 -725 4419
rect -469 4423 -31 4426
rect -469 4406 -463 4423
rect -37 4406 -31 4423
rect -469 4403 -31 4406
rect 81 4423 519 4426
rect 81 4406 87 4423
rect 513 4406 519 4423
rect 81 4403 519 4406
rect 631 4423 1069 4426
rect 631 4406 637 4423
rect 1063 4406 1069 4423
rect 631 4403 1069 4406
rect 1181 4423 1619 4426
rect 1181 4406 1187 4423
rect 1613 4406 1619 4423
rect 1181 4403 1619 4406
rect 1731 4423 2169 4426
rect 1731 4406 1737 4423
rect 2163 4406 2169 4423
rect 1731 4403 2169 4406
rect 2281 4423 2719 4426
rect 2281 4406 2287 4423
rect 2713 4406 2719 4423
rect 2281 4403 2719 4406
rect 2831 4423 3269 4426
rect 2831 4406 2837 4423
rect 3263 4406 3269 4423
rect 2831 4403 3269 4406
rect 3381 4423 3819 4426
rect 3381 4406 3387 4423
rect 3813 4406 3819 4423
rect 3381 4403 3819 4406
rect 3931 4423 4369 4426
rect 3931 4406 3937 4423
rect 4363 4406 4369 4423
rect 3931 4403 4369 4406
rect 4481 4423 4919 4426
rect 4481 4406 4487 4423
rect 4913 4406 4919 4423
rect 4481 4403 4919 4406
rect 5031 4423 5469 4426
rect 5031 4406 5037 4423
rect 5463 4406 5469 4423
rect 5031 4403 5469 4406
rect 5581 4423 6019 4426
rect 5581 4406 5587 4423
rect 6013 4406 6019 4423
rect 5581 4403 6019 4406
rect 6131 4423 6569 4426
rect 6131 4406 6137 4423
rect 6563 4406 6569 4423
rect 6131 4403 6569 4406
rect 6681 4423 7119 4426
rect 6681 4406 6687 4423
rect 7113 4406 7119 4423
rect 6681 4403 7119 4406
rect 7231 4423 7669 4426
rect 7231 4406 7237 4423
rect 7663 4406 7669 4423
rect 7231 4403 7669 4406
rect 7781 4423 8219 4426
rect 7781 4406 7787 4423
rect 8213 4406 8219 4423
rect 7781 4403 8219 4406
rect 8331 4423 8769 4426
rect 8331 4406 8337 4423
rect 8763 4406 8769 4423
rect 8331 4403 8769 4406
rect 8881 4423 9319 4426
rect 8881 4406 8887 4423
rect 9313 4406 9319 4423
rect 8881 4403 9319 4406
rect 9431 4423 9869 4426
rect 9431 4406 9437 4423
rect 9863 4406 9869 4423
rect 9431 4403 9869 4406
rect 9981 4423 10419 4426
rect 9981 4406 9987 4423
rect 10413 4406 10419 4423
rect 9981 4403 10419 4406
rect 10531 4423 10969 4426
rect 10531 4406 10537 4423
rect 10963 4406 10969 4423
rect 10531 4403 10969 4406
rect 11081 4423 11519 4426
rect 11081 4406 11087 4423
rect 11513 4406 11519 4423
rect 11081 4403 11519 4406
rect 11631 4423 12069 4426
rect 11631 4406 11637 4423
rect 12063 4406 12069 4423
rect 11631 4403 12069 4406
rect 12181 4423 12619 4426
rect 12181 4406 12187 4423
rect 12613 4406 12619 4423
rect 12181 4403 12619 4406
rect 12731 4423 13169 4426
rect 12731 4406 12737 4423
rect 13163 4406 13169 4423
rect 12731 4403 13169 4406
rect 13281 4423 13719 4426
rect 13281 4406 13287 4423
rect 13713 4406 13719 4423
rect 13281 4403 13719 4406
rect 13975 4419 13987 4950
rect 14263 4419 14275 4950
rect 13975 4400 14275 4419
rect -1025 3869 -1013 4400
rect -737 3869 -725 4400
rect -550 4392 -500 4400
rect -550 4358 -542 4392
rect -508 4358 -500 4392
rect -550 4350 -500 4358
rect 0 4392 50 4400
rect 0 4358 8 4392
rect 42 4358 50 4392
rect 0 4350 50 4358
rect 550 4392 600 4400
rect 550 4358 558 4392
rect 592 4358 600 4392
rect 550 4350 600 4358
rect 1100 4392 1150 4400
rect 1100 4358 1108 4392
rect 1142 4358 1150 4392
rect 1100 4350 1150 4358
rect 1650 4392 1700 4400
rect 1650 4358 1658 4392
rect 1692 4358 1700 4392
rect 1650 4350 1700 4358
rect 2200 4392 2250 4400
rect 2200 4358 2208 4392
rect 2242 4358 2250 4392
rect 2200 4350 2250 4358
rect 2750 4392 2800 4400
rect 2750 4358 2758 4392
rect 2792 4358 2800 4392
rect 2750 4350 2800 4358
rect 3300 4392 3350 4400
rect 3300 4358 3308 4392
rect 3342 4358 3350 4392
rect 3300 4350 3350 4358
rect 3850 4392 3900 4400
rect 3850 4358 3858 4392
rect 3892 4358 3900 4392
rect 3850 4350 3900 4358
rect 4400 4392 4450 4400
rect 4400 4358 4408 4392
rect 4442 4358 4450 4392
rect 4400 4350 4450 4358
rect 4950 4392 5000 4400
rect 4950 4358 4958 4392
rect 4992 4358 5000 4392
rect 4950 4350 5000 4358
rect 5500 4392 5550 4400
rect 5500 4358 5508 4392
rect 5542 4358 5550 4392
rect 5500 4350 5550 4358
rect 6050 4392 6100 4400
rect 6050 4358 6058 4392
rect 6092 4358 6100 4392
rect 6050 4350 6100 4358
rect 6600 4392 6650 4400
rect 6600 4358 6608 4392
rect 6642 4358 6650 4392
rect 6600 4350 6650 4358
rect 7150 4392 7200 4400
rect 7150 4358 7158 4392
rect 7192 4358 7200 4392
rect 7150 4350 7200 4358
rect 7700 4392 7750 4400
rect 7700 4358 7708 4392
rect 7742 4358 7750 4392
rect 7700 4350 7750 4358
rect 8250 4392 8300 4400
rect 8250 4358 8258 4392
rect 8292 4358 8300 4392
rect 8250 4350 8300 4358
rect 8800 4392 8850 4400
rect 8800 4358 8808 4392
rect 8842 4358 8850 4392
rect 8800 4350 8850 4358
rect 9350 4392 9400 4400
rect 9350 4358 9358 4392
rect 9392 4358 9400 4392
rect 9350 4350 9400 4358
rect 9900 4392 9950 4400
rect 9900 4358 9908 4392
rect 9942 4358 9950 4392
rect 9900 4350 9950 4358
rect 10450 4392 10500 4400
rect 10450 4358 10458 4392
rect 10492 4358 10500 4392
rect 10450 4350 10500 4358
rect 11000 4392 11050 4400
rect 11000 4358 11008 4392
rect 11042 4358 11050 4392
rect 11000 4350 11050 4358
rect 11550 4392 11600 4400
rect 11550 4358 11558 4392
rect 11592 4358 11600 4392
rect 11550 4350 11600 4358
rect 12100 4392 12150 4400
rect 12100 4358 12108 4392
rect 12142 4358 12150 4392
rect 12100 4350 12150 4358
rect 12650 4392 12700 4400
rect 12650 4358 12658 4392
rect 12692 4358 12700 4392
rect 12650 4350 12700 4358
rect 13200 4392 13250 4400
rect 13200 4358 13208 4392
rect 13242 4358 13250 4392
rect 13200 4350 13250 4358
rect 13750 4392 13800 4400
rect 13750 4358 13758 4392
rect 13792 4358 13800 4392
rect 13750 4350 13800 4358
rect -469 4344 -31 4347
rect -469 4327 -463 4344
rect -37 4327 -31 4344
rect -469 4324 -31 4327
rect 81 4344 519 4347
rect 81 4327 87 4344
rect 513 4327 519 4344
rect 81 4324 519 4327
rect 631 4344 1069 4347
rect 631 4327 637 4344
rect 1063 4327 1069 4344
rect 631 4324 1069 4327
rect 1181 4344 1619 4347
rect 1181 4327 1187 4344
rect 1613 4327 1619 4344
rect 1181 4324 1619 4327
rect 1731 4344 2169 4347
rect 1731 4327 1737 4344
rect 2163 4327 2169 4344
rect 1731 4324 2169 4327
rect 2281 4344 2719 4347
rect 2281 4327 2287 4344
rect 2713 4327 2719 4344
rect 2281 4324 2719 4327
rect 2831 4344 3269 4347
rect 2831 4327 2837 4344
rect 3263 4327 3269 4344
rect 2831 4324 3269 4327
rect 3381 4344 3819 4347
rect 3381 4327 3387 4344
rect 3813 4327 3819 4344
rect 3381 4324 3819 4327
rect 3931 4344 4369 4347
rect 3931 4327 3937 4344
rect 4363 4327 4369 4344
rect 3931 4324 4369 4327
rect 4481 4344 4919 4347
rect 4481 4327 4487 4344
rect 4913 4327 4919 4344
rect 4481 4324 4919 4327
rect 5031 4344 5469 4347
rect 5031 4327 5037 4344
rect 5463 4327 5469 4344
rect 5031 4324 5469 4327
rect 5581 4344 6019 4347
rect 5581 4327 5587 4344
rect 6013 4327 6019 4344
rect 5581 4324 6019 4327
rect 6131 4344 6569 4347
rect 6131 4327 6137 4344
rect 6563 4327 6569 4344
rect 6131 4324 6569 4327
rect 6681 4344 7119 4347
rect 6681 4327 6687 4344
rect 7113 4327 7119 4344
rect 6681 4324 7119 4327
rect 7231 4344 7669 4347
rect 7231 4327 7237 4344
rect 7663 4327 7669 4344
rect 7231 4324 7669 4327
rect 7781 4344 8219 4347
rect 7781 4327 7787 4344
rect 8213 4327 8219 4344
rect 7781 4324 8219 4327
rect 8331 4344 8769 4347
rect 8331 4327 8337 4344
rect 8763 4327 8769 4344
rect 8331 4324 8769 4327
rect 8881 4344 9319 4347
rect 8881 4327 8887 4344
rect 9313 4327 9319 4344
rect 8881 4324 9319 4327
rect 9431 4344 9869 4347
rect 9431 4327 9437 4344
rect 9863 4327 9869 4344
rect 9431 4324 9869 4327
rect 9981 4344 10419 4347
rect 9981 4327 9987 4344
rect 10413 4327 10419 4344
rect 9981 4324 10419 4327
rect 10531 4344 10969 4347
rect 10531 4327 10537 4344
rect 10963 4327 10969 4344
rect 10531 4324 10969 4327
rect 11081 4344 11519 4347
rect 11081 4327 11087 4344
rect 11513 4327 11519 4344
rect 11081 4324 11519 4327
rect 11631 4344 12069 4347
rect 11631 4327 11637 4344
rect 12063 4327 12069 4344
rect 11631 4324 12069 4327
rect 12181 4344 12619 4347
rect 12181 4327 12187 4344
rect 12613 4327 12619 4344
rect 12181 4324 12619 4327
rect 12731 4344 13169 4347
rect 12731 4327 12737 4344
rect 13163 4327 13169 4344
rect 12731 4324 13169 4327
rect 13281 4344 13719 4347
rect 13281 4327 13287 4344
rect 13713 4327 13719 4344
rect 13281 4324 13719 4327
rect -474 4319 -26 4324
rect 76 4319 524 4324
rect 626 4319 1074 4324
rect 1176 4319 1624 4324
rect 1726 4319 2174 4324
rect 2276 4319 2724 4324
rect 2826 4319 3274 4324
rect 3376 4319 3824 4324
rect 3926 4319 4374 4324
rect 4476 4319 4924 4324
rect 5026 4319 5474 4324
rect 5576 4319 6024 4324
rect 6126 4319 6574 4324
rect 6676 4319 7124 4324
rect 7226 4319 7674 4324
rect 7776 4319 8224 4324
rect 8326 4319 8774 4324
rect 8876 4319 9324 4324
rect 9426 4319 9874 4324
rect 9976 4319 10424 4324
rect 10526 4319 10974 4324
rect 11076 4319 11524 4324
rect 11626 4319 12074 4324
rect 12176 4319 12624 4324
rect 12726 4319 13174 4324
rect 13276 4319 13724 4324
rect -474 4313 -3 4319
rect -474 4265 -23 4313
rect -474 3935 -415 4265
rect -85 3935 -23 4265
rect -474 3887 -23 3935
rect -6 3887 -3 4313
rect -474 3881 -3 3887
rect 53 4313 547 4319
rect 53 3887 56 4313
rect 73 4265 527 4313
rect 73 3935 135 4265
rect 465 3935 527 4265
rect 73 3887 527 3935
rect 544 3887 547 4313
rect 53 3881 547 3887
rect 603 4313 1097 4319
rect 603 3887 606 4313
rect 623 4265 1077 4313
rect 623 3935 685 4265
rect 1015 3935 1077 4265
rect 623 3887 1077 3935
rect 1094 3887 1097 4313
rect 603 3881 1097 3887
rect 1153 4313 1647 4319
rect 1153 3887 1156 4313
rect 1173 4265 1627 4313
rect 1173 3935 1235 4265
rect 1565 3935 1627 4265
rect 1173 3887 1627 3935
rect 1644 3887 1647 4313
rect 1153 3881 1647 3887
rect 1703 4313 2197 4319
rect 1703 3887 1706 4313
rect 1723 4265 2177 4313
rect 1723 3935 1785 4265
rect 2115 3935 2177 4265
rect 1723 3887 2177 3935
rect 2194 3887 2197 4313
rect 1703 3881 2197 3887
rect 2253 4313 2747 4319
rect 2253 3887 2256 4313
rect 2273 4265 2727 4313
rect 2273 3935 2335 4265
rect 2665 3935 2727 4265
rect 2273 3887 2727 3935
rect 2744 3887 2747 4313
rect 2253 3881 2747 3887
rect 2803 4313 3297 4319
rect 2803 3887 2806 4313
rect 2823 4265 3277 4313
rect 2823 3935 2885 4265
rect 3215 3935 3277 4265
rect 2823 3887 3277 3935
rect 3294 3887 3297 4313
rect 2803 3881 3297 3887
rect 3353 4313 3847 4319
rect 3353 3887 3356 4313
rect 3373 4265 3827 4313
rect 3373 3935 3435 4265
rect 3765 3935 3827 4265
rect 3373 3887 3827 3935
rect 3844 3887 3847 4313
rect 3353 3881 3847 3887
rect 3903 4313 4397 4319
rect 3903 3887 3906 4313
rect 3923 4265 4377 4313
rect 3923 3935 3985 4265
rect 4315 3935 4377 4265
rect 3923 3887 4377 3935
rect 4394 3887 4397 4313
rect 3903 3881 4397 3887
rect 4453 4313 4947 4319
rect 4453 3887 4456 4313
rect 4473 4265 4927 4313
rect 4473 3935 4535 4265
rect 4865 3935 4927 4265
rect 4473 3887 4927 3935
rect 4944 3887 4947 4313
rect 4453 3881 4947 3887
rect 5003 4313 5497 4319
rect 5003 3887 5006 4313
rect 5023 4265 5477 4313
rect 5023 3935 5085 4265
rect 5415 3935 5477 4265
rect 5023 3887 5477 3935
rect 5494 3887 5497 4313
rect 5003 3881 5497 3887
rect 5553 4313 6047 4319
rect 5553 3887 5556 4313
rect 5573 4265 6027 4313
rect 5573 3935 5635 4265
rect 5965 3935 6027 4265
rect 5573 3887 6027 3935
rect 6044 3887 6047 4313
rect 5553 3881 6047 3887
rect 6103 4313 6597 4319
rect 6103 3887 6106 4313
rect 6123 4265 6577 4313
rect 6123 3935 6185 4265
rect 6515 3935 6577 4265
rect 6123 3887 6577 3935
rect 6594 3887 6597 4313
rect 6103 3881 6597 3887
rect 6653 4313 7147 4319
rect 6653 3887 6656 4313
rect 6673 4265 7127 4313
rect 6673 3935 6735 4265
rect 7065 3935 7127 4265
rect 6673 3887 7127 3935
rect 7144 3887 7147 4313
rect 6653 3881 7147 3887
rect 7203 4313 7697 4319
rect 7203 3887 7206 4313
rect 7223 4265 7677 4313
rect 7223 3935 7285 4265
rect 7615 3935 7677 4265
rect 7223 3887 7677 3935
rect 7694 3887 7697 4313
rect 7203 3881 7697 3887
rect 7753 4313 8247 4319
rect 7753 3887 7756 4313
rect 7773 4265 8227 4313
rect 7773 3935 7835 4265
rect 8165 3935 8227 4265
rect 7773 3887 8227 3935
rect 8244 3887 8247 4313
rect 7753 3881 8247 3887
rect 8303 4313 8797 4319
rect 8303 3887 8306 4313
rect 8323 4265 8777 4313
rect 8323 3935 8385 4265
rect 8715 3935 8777 4265
rect 8323 3887 8777 3935
rect 8794 3887 8797 4313
rect 8303 3881 8797 3887
rect 8853 4313 9347 4319
rect 8853 3887 8856 4313
rect 8873 4265 9327 4313
rect 8873 3935 8935 4265
rect 9265 3935 9327 4265
rect 8873 3887 9327 3935
rect 9344 3887 9347 4313
rect 8853 3881 9347 3887
rect 9403 4313 9897 4319
rect 9403 3887 9406 4313
rect 9423 4265 9877 4313
rect 9423 3935 9485 4265
rect 9815 3935 9877 4265
rect 9423 3887 9877 3935
rect 9894 3887 9897 4313
rect 9403 3881 9897 3887
rect 9953 4313 10447 4319
rect 9953 3887 9956 4313
rect 9973 4265 10427 4313
rect 9973 3935 10035 4265
rect 10365 3935 10427 4265
rect 9973 3887 10427 3935
rect 10444 3887 10447 4313
rect 9953 3881 10447 3887
rect 10503 4313 10997 4319
rect 10503 3887 10506 4313
rect 10523 4265 10977 4313
rect 10523 3935 10585 4265
rect 10915 3935 10977 4265
rect 10523 3887 10977 3935
rect 10994 3887 10997 4313
rect 10503 3881 10997 3887
rect 11053 4313 11547 4319
rect 11053 3887 11056 4313
rect 11073 4265 11527 4313
rect 11073 3935 11135 4265
rect 11465 3935 11527 4265
rect 11073 3887 11527 3935
rect 11544 3887 11547 4313
rect 11053 3881 11547 3887
rect 11603 4313 12097 4319
rect 11603 3887 11606 4313
rect 11623 4265 12077 4313
rect 11623 3935 11685 4265
rect 12015 3935 12077 4265
rect 11623 3887 12077 3935
rect 12094 3887 12097 4313
rect 11603 3881 12097 3887
rect 12153 4313 12647 4319
rect 12153 3887 12156 4313
rect 12173 4265 12627 4313
rect 12173 3935 12235 4265
rect 12565 3935 12627 4265
rect 12173 3887 12627 3935
rect 12644 3887 12647 4313
rect 12153 3881 12647 3887
rect 12703 4313 13197 4319
rect 12703 3887 12706 4313
rect 12723 4265 13177 4313
rect 12723 3935 12785 4265
rect 13115 3935 13177 4265
rect 12723 3887 13177 3935
rect 13194 3887 13197 4313
rect 12703 3881 13197 3887
rect 13253 4313 13724 4319
rect 13253 3887 13256 4313
rect 13273 4265 13724 4313
rect 13273 3935 13335 4265
rect 13665 3935 13724 4265
rect 13273 3887 13724 3935
rect 13253 3881 13724 3887
rect -474 3876 -26 3881
rect 76 3876 524 3881
rect 626 3876 1074 3881
rect 1176 3876 1624 3881
rect 1726 3876 2174 3881
rect 2276 3876 2724 3881
rect 2826 3876 3274 3881
rect 3376 3876 3824 3881
rect 3926 3876 4374 3881
rect 4476 3876 4924 3881
rect 5026 3876 5474 3881
rect 5576 3876 6024 3881
rect 6126 3876 6574 3881
rect 6676 3876 7124 3881
rect 7226 3876 7674 3881
rect 7776 3876 8224 3881
rect 8326 3876 8774 3881
rect 8876 3876 9324 3881
rect 9426 3876 9874 3881
rect 9976 3876 10424 3881
rect 10526 3876 10974 3881
rect 11076 3876 11524 3881
rect 11626 3876 12074 3881
rect 12176 3876 12624 3881
rect 12726 3876 13174 3881
rect 13276 3876 13724 3881
rect -1025 3850 -725 3869
rect -469 3873 -31 3876
rect -469 3856 -463 3873
rect -37 3856 -31 3873
rect -469 3853 -31 3856
rect 81 3873 519 3876
rect 81 3856 87 3873
rect 513 3856 519 3873
rect 81 3853 519 3856
rect 631 3873 1069 3876
rect 631 3856 637 3873
rect 1063 3856 1069 3873
rect 631 3853 1069 3856
rect 1181 3873 1619 3876
rect 1181 3856 1187 3873
rect 1613 3856 1619 3873
rect 1181 3853 1619 3856
rect 1731 3873 2169 3876
rect 1731 3856 1737 3873
rect 2163 3856 2169 3873
rect 1731 3853 2169 3856
rect 2281 3873 2719 3876
rect 2281 3856 2287 3873
rect 2713 3856 2719 3873
rect 2281 3853 2719 3856
rect 2831 3873 3269 3876
rect 2831 3856 2837 3873
rect 3263 3856 3269 3873
rect 2831 3853 3269 3856
rect 3381 3873 3819 3876
rect 3381 3856 3387 3873
rect 3813 3856 3819 3873
rect 3381 3853 3819 3856
rect 3931 3873 4369 3876
rect 3931 3856 3937 3873
rect 4363 3856 4369 3873
rect 3931 3853 4369 3856
rect 4481 3873 4919 3876
rect 4481 3856 4487 3873
rect 4913 3856 4919 3873
rect 4481 3853 4919 3856
rect 5031 3873 5469 3876
rect 5031 3856 5037 3873
rect 5463 3856 5469 3873
rect 5031 3853 5469 3856
rect 5581 3873 6019 3876
rect 5581 3856 5587 3873
rect 6013 3856 6019 3873
rect 5581 3853 6019 3856
rect 6131 3873 6569 3876
rect 6131 3856 6137 3873
rect 6563 3856 6569 3873
rect 6131 3853 6569 3856
rect 6681 3873 7119 3876
rect 6681 3856 6687 3873
rect 7113 3856 7119 3873
rect 6681 3853 7119 3856
rect 7231 3873 7669 3876
rect 7231 3856 7237 3873
rect 7663 3856 7669 3873
rect 7231 3853 7669 3856
rect 7781 3873 8219 3876
rect 7781 3856 7787 3873
rect 8213 3856 8219 3873
rect 7781 3853 8219 3856
rect 8331 3873 8769 3876
rect 8331 3856 8337 3873
rect 8763 3856 8769 3873
rect 8331 3853 8769 3856
rect 8881 3873 9319 3876
rect 8881 3856 8887 3873
rect 9313 3856 9319 3873
rect 8881 3853 9319 3856
rect 9431 3873 9869 3876
rect 9431 3856 9437 3873
rect 9863 3856 9869 3873
rect 9431 3853 9869 3856
rect 9981 3873 10419 3876
rect 9981 3856 9987 3873
rect 10413 3856 10419 3873
rect 9981 3853 10419 3856
rect 10531 3873 10969 3876
rect 10531 3856 10537 3873
rect 10963 3856 10969 3873
rect 10531 3853 10969 3856
rect 11081 3873 11519 3876
rect 11081 3856 11087 3873
rect 11513 3856 11519 3873
rect 11081 3853 11519 3856
rect 11631 3873 12069 3876
rect 11631 3856 11637 3873
rect 12063 3856 12069 3873
rect 11631 3853 12069 3856
rect 12181 3873 12619 3876
rect 12181 3856 12187 3873
rect 12613 3856 12619 3873
rect 12181 3853 12619 3856
rect 12731 3873 13169 3876
rect 12731 3856 12737 3873
rect 13163 3856 13169 3873
rect 12731 3853 13169 3856
rect 13281 3873 13719 3876
rect 13281 3856 13287 3873
rect 13713 3856 13719 3873
rect 13281 3853 13719 3856
rect 13975 3869 13987 4400
rect 14263 3869 14275 4400
rect 13975 3850 14275 3869
rect -1025 3319 -1013 3850
rect -737 3319 -725 3850
rect -550 3842 -500 3850
rect -550 3808 -542 3842
rect -508 3808 -500 3842
rect -550 3800 -500 3808
rect 0 3842 50 3850
rect 0 3808 8 3842
rect 42 3808 50 3842
rect 0 3800 50 3808
rect 550 3842 600 3850
rect 550 3808 558 3842
rect 592 3808 600 3842
rect 550 3800 600 3808
rect 1100 3842 1150 3850
rect 1100 3808 1108 3842
rect 1142 3808 1150 3842
rect 1100 3800 1150 3808
rect 1650 3842 1700 3850
rect 1650 3808 1658 3842
rect 1692 3808 1700 3842
rect 1650 3800 1700 3808
rect 2200 3842 2250 3850
rect 2200 3808 2208 3842
rect 2242 3808 2250 3842
rect 2200 3800 2250 3808
rect 2750 3842 2800 3850
rect 2750 3808 2758 3842
rect 2792 3808 2800 3842
rect 2750 3800 2800 3808
rect 3300 3842 3350 3850
rect 3300 3808 3308 3842
rect 3342 3808 3350 3842
rect 3300 3800 3350 3808
rect 3850 3842 3900 3850
rect 3850 3808 3858 3842
rect 3892 3808 3900 3842
rect 3850 3800 3900 3808
rect 4400 3842 4450 3850
rect 4400 3808 4408 3842
rect 4442 3808 4450 3842
rect 4400 3800 4450 3808
rect 4950 3842 5000 3850
rect 4950 3808 4958 3842
rect 4992 3808 5000 3842
rect 4950 3800 5000 3808
rect 5500 3842 5550 3850
rect 5500 3808 5508 3842
rect 5542 3808 5550 3842
rect 5500 3800 5550 3808
rect 6050 3842 6100 3850
rect 6050 3808 6058 3842
rect 6092 3808 6100 3842
rect 6050 3800 6100 3808
rect 6600 3842 6650 3850
rect 6600 3808 6608 3842
rect 6642 3808 6650 3842
rect 6600 3800 6650 3808
rect 7150 3842 7200 3850
rect 7150 3808 7158 3842
rect 7192 3808 7200 3842
rect 7150 3800 7200 3808
rect 7700 3842 7750 3850
rect 7700 3808 7708 3842
rect 7742 3808 7750 3842
rect 7700 3800 7750 3808
rect 8250 3842 8300 3850
rect 8250 3808 8258 3842
rect 8292 3808 8300 3842
rect 8250 3800 8300 3808
rect 8800 3842 8850 3850
rect 8800 3808 8808 3842
rect 8842 3808 8850 3842
rect 8800 3800 8850 3808
rect 9350 3842 9400 3850
rect 9350 3808 9358 3842
rect 9392 3808 9400 3842
rect 9350 3800 9400 3808
rect 9900 3842 9950 3850
rect 9900 3808 9908 3842
rect 9942 3808 9950 3842
rect 9900 3800 9950 3808
rect 10450 3842 10500 3850
rect 10450 3808 10458 3842
rect 10492 3808 10500 3842
rect 10450 3800 10500 3808
rect 11000 3842 11050 3850
rect 11000 3808 11008 3842
rect 11042 3808 11050 3842
rect 11000 3800 11050 3808
rect 11550 3842 11600 3850
rect 11550 3808 11558 3842
rect 11592 3808 11600 3842
rect 11550 3800 11600 3808
rect 12100 3842 12150 3850
rect 12100 3808 12108 3842
rect 12142 3808 12150 3842
rect 12100 3800 12150 3808
rect 12650 3842 12700 3850
rect 12650 3808 12658 3842
rect 12692 3808 12700 3842
rect 12650 3800 12700 3808
rect 13200 3842 13250 3850
rect 13200 3808 13208 3842
rect 13242 3808 13250 3842
rect 13200 3800 13250 3808
rect 13750 3842 13800 3850
rect 13750 3808 13758 3842
rect 13792 3808 13800 3842
rect 13750 3800 13800 3808
rect -469 3794 -31 3797
rect -469 3777 -463 3794
rect -37 3777 -31 3794
rect -469 3774 -31 3777
rect 81 3794 519 3797
rect 81 3777 87 3794
rect 513 3777 519 3794
rect 81 3774 519 3777
rect 631 3794 1069 3797
rect 631 3777 637 3794
rect 1063 3777 1069 3794
rect 631 3774 1069 3777
rect 1181 3794 1619 3797
rect 1181 3777 1187 3794
rect 1613 3777 1619 3794
rect 1181 3774 1619 3777
rect 1731 3794 2169 3797
rect 1731 3777 1737 3794
rect 2163 3777 2169 3794
rect 1731 3774 2169 3777
rect 2281 3794 2719 3797
rect 2281 3777 2287 3794
rect 2713 3777 2719 3794
rect 2281 3774 2719 3777
rect 2831 3794 3269 3797
rect 2831 3777 2837 3794
rect 3263 3777 3269 3794
rect 2831 3774 3269 3777
rect 3381 3794 3819 3797
rect 3381 3777 3387 3794
rect 3813 3777 3819 3794
rect 3381 3774 3819 3777
rect 3931 3794 4369 3797
rect 3931 3777 3937 3794
rect 4363 3777 4369 3794
rect 3931 3774 4369 3777
rect 4481 3794 4919 3797
rect 4481 3777 4487 3794
rect 4913 3777 4919 3794
rect 4481 3774 4919 3777
rect 5031 3794 5469 3797
rect 5031 3777 5037 3794
rect 5463 3777 5469 3794
rect 5031 3774 5469 3777
rect 5581 3794 6019 3797
rect 5581 3777 5587 3794
rect 6013 3777 6019 3794
rect 5581 3774 6019 3777
rect 6131 3794 6569 3797
rect 6131 3777 6137 3794
rect 6563 3777 6569 3794
rect 6131 3774 6569 3777
rect 6681 3794 7119 3797
rect 6681 3777 6687 3794
rect 7113 3777 7119 3794
rect 6681 3774 7119 3777
rect 7231 3794 7669 3797
rect 7231 3777 7237 3794
rect 7663 3777 7669 3794
rect 7231 3774 7669 3777
rect 7781 3794 8219 3797
rect 7781 3777 7787 3794
rect 8213 3777 8219 3794
rect 7781 3774 8219 3777
rect 8331 3794 8769 3797
rect 8331 3777 8337 3794
rect 8763 3777 8769 3794
rect 8331 3774 8769 3777
rect 8881 3794 9319 3797
rect 8881 3777 8887 3794
rect 9313 3777 9319 3794
rect 8881 3774 9319 3777
rect 9431 3794 9869 3797
rect 9431 3777 9437 3794
rect 9863 3777 9869 3794
rect 9431 3774 9869 3777
rect 9981 3794 10419 3797
rect 9981 3777 9987 3794
rect 10413 3777 10419 3794
rect 9981 3774 10419 3777
rect 10531 3794 10969 3797
rect 10531 3777 10537 3794
rect 10963 3777 10969 3794
rect 10531 3774 10969 3777
rect 11081 3794 11519 3797
rect 11081 3777 11087 3794
rect 11513 3777 11519 3794
rect 11081 3774 11519 3777
rect 11631 3794 12069 3797
rect 11631 3777 11637 3794
rect 12063 3777 12069 3794
rect 11631 3774 12069 3777
rect 12181 3794 12619 3797
rect 12181 3777 12187 3794
rect 12613 3777 12619 3794
rect 12181 3774 12619 3777
rect 12731 3794 13169 3797
rect 12731 3777 12737 3794
rect 13163 3777 13169 3794
rect 12731 3774 13169 3777
rect 13281 3794 13719 3797
rect 13281 3777 13287 3794
rect 13713 3777 13719 3794
rect 13281 3774 13719 3777
rect -474 3769 -26 3774
rect 76 3769 524 3774
rect 626 3769 1074 3774
rect 1176 3769 1624 3774
rect 1726 3769 2174 3774
rect 2276 3769 2724 3774
rect 2826 3769 3274 3774
rect 3376 3769 3824 3774
rect 3926 3769 4374 3774
rect 4476 3769 4924 3774
rect 5026 3769 5474 3774
rect 5576 3769 6024 3774
rect 6126 3769 6574 3774
rect 6676 3769 7124 3774
rect 7226 3769 7674 3774
rect 7776 3769 8224 3774
rect 8326 3769 8774 3774
rect 8876 3769 9324 3774
rect 9426 3769 9874 3774
rect 9976 3769 10424 3774
rect 10526 3769 10974 3774
rect 11076 3769 11524 3774
rect 11626 3769 12074 3774
rect 12176 3769 12624 3774
rect 12726 3769 13174 3774
rect 13276 3769 13724 3774
rect -474 3763 -3 3769
rect -474 3715 -23 3763
rect -474 3385 -415 3715
rect -85 3385 -23 3715
rect -474 3337 -23 3385
rect -6 3337 -3 3763
rect -474 3331 -3 3337
rect 53 3763 547 3769
rect 53 3337 56 3763
rect 73 3715 527 3763
rect 73 3385 135 3715
rect 465 3385 527 3715
rect 73 3337 527 3385
rect 544 3337 547 3763
rect 53 3331 547 3337
rect 603 3763 1097 3769
rect 603 3337 606 3763
rect 623 3715 1077 3763
rect 623 3385 685 3715
rect 1015 3385 1077 3715
rect 623 3337 1077 3385
rect 1094 3337 1097 3763
rect 603 3331 1097 3337
rect 1153 3763 1647 3769
rect 1153 3337 1156 3763
rect 1173 3715 1627 3763
rect 1173 3385 1235 3715
rect 1565 3385 1627 3715
rect 1173 3337 1627 3385
rect 1644 3337 1647 3763
rect 1153 3331 1647 3337
rect 1703 3763 2197 3769
rect 1703 3337 1706 3763
rect 1723 3715 2177 3763
rect 1723 3385 1785 3715
rect 2115 3385 2177 3715
rect 1723 3337 2177 3385
rect 2194 3337 2197 3763
rect 1703 3331 2197 3337
rect 2253 3763 2747 3769
rect 2253 3337 2256 3763
rect 2273 3715 2727 3763
rect 2273 3385 2335 3715
rect 2665 3385 2727 3715
rect 2273 3337 2727 3385
rect 2744 3337 2747 3763
rect 2253 3331 2747 3337
rect 2803 3763 3297 3769
rect 2803 3337 2806 3763
rect 2823 3715 3277 3763
rect 2823 3385 2885 3715
rect 3215 3385 3277 3715
rect 2823 3337 3277 3385
rect 3294 3337 3297 3763
rect 2803 3331 3297 3337
rect 3353 3763 3847 3769
rect 3353 3337 3356 3763
rect 3373 3715 3827 3763
rect 3373 3385 3435 3715
rect 3765 3385 3827 3715
rect 3373 3337 3827 3385
rect 3844 3337 3847 3763
rect 3353 3331 3847 3337
rect 3903 3763 4397 3769
rect 3903 3337 3906 3763
rect 3923 3715 4377 3763
rect 3923 3385 3985 3715
rect 4315 3385 4377 3715
rect 3923 3337 4377 3385
rect 4394 3337 4397 3763
rect 3903 3331 4397 3337
rect 4453 3763 4947 3769
rect 4453 3337 4456 3763
rect 4473 3715 4927 3763
rect 4473 3385 4535 3715
rect 4865 3385 4927 3715
rect 4473 3337 4927 3385
rect 4944 3337 4947 3763
rect 4453 3331 4947 3337
rect 5003 3763 5497 3769
rect 5003 3337 5006 3763
rect 5023 3715 5477 3763
rect 5023 3385 5085 3715
rect 5415 3385 5477 3715
rect 5023 3337 5477 3385
rect 5494 3337 5497 3763
rect 5003 3331 5497 3337
rect 5553 3763 6047 3769
rect 5553 3337 5556 3763
rect 5573 3715 6027 3763
rect 5573 3385 5635 3715
rect 5965 3385 6027 3715
rect 5573 3337 6027 3385
rect 6044 3337 6047 3763
rect 5553 3331 6047 3337
rect 6103 3763 6597 3769
rect 6103 3337 6106 3763
rect 6123 3715 6577 3763
rect 6123 3385 6185 3715
rect 6515 3385 6577 3715
rect 6123 3337 6577 3385
rect 6594 3337 6597 3763
rect 6103 3331 6597 3337
rect 6653 3763 7147 3769
rect 6653 3337 6656 3763
rect 6673 3715 7127 3763
rect 6673 3385 6735 3715
rect 7065 3385 7127 3715
rect 6673 3337 7127 3385
rect 7144 3337 7147 3763
rect 6653 3331 7147 3337
rect 7203 3763 7697 3769
rect 7203 3337 7206 3763
rect 7223 3715 7677 3763
rect 7223 3385 7285 3715
rect 7615 3385 7677 3715
rect 7223 3337 7677 3385
rect 7694 3337 7697 3763
rect 7203 3331 7697 3337
rect 7753 3763 8247 3769
rect 7753 3337 7756 3763
rect 7773 3715 8227 3763
rect 7773 3385 7835 3715
rect 8165 3385 8227 3715
rect 7773 3337 8227 3385
rect 8244 3337 8247 3763
rect 7753 3331 8247 3337
rect 8303 3763 8797 3769
rect 8303 3337 8306 3763
rect 8323 3715 8777 3763
rect 8323 3385 8385 3715
rect 8715 3385 8777 3715
rect 8323 3337 8777 3385
rect 8794 3337 8797 3763
rect 8303 3331 8797 3337
rect 8853 3763 9347 3769
rect 8853 3337 8856 3763
rect 8873 3715 9327 3763
rect 8873 3385 8935 3715
rect 9265 3385 9327 3715
rect 8873 3337 9327 3385
rect 9344 3337 9347 3763
rect 8853 3331 9347 3337
rect 9403 3763 9897 3769
rect 9403 3337 9406 3763
rect 9423 3715 9877 3763
rect 9423 3385 9485 3715
rect 9815 3385 9877 3715
rect 9423 3337 9877 3385
rect 9894 3337 9897 3763
rect 9403 3331 9897 3337
rect 9953 3763 10447 3769
rect 9953 3337 9956 3763
rect 9973 3715 10427 3763
rect 9973 3385 10035 3715
rect 10365 3385 10427 3715
rect 9973 3337 10427 3385
rect 10444 3337 10447 3763
rect 9953 3331 10447 3337
rect 10503 3763 10997 3769
rect 10503 3337 10506 3763
rect 10523 3715 10977 3763
rect 10523 3385 10585 3715
rect 10915 3385 10977 3715
rect 10523 3337 10977 3385
rect 10994 3337 10997 3763
rect 10503 3331 10997 3337
rect 11053 3763 11547 3769
rect 11053 3337 11056 3763
rect 11073 3715 11527 3763
rect 11073 3385 11135 3715
rect 11465 3385 11527 3715
rect 11073 3337 11527 3385
rect 11544 3337 11547 3763
rect 11053 3331 11547 3337
rect 11603 3763 12097 3769
rect 11603 3337 11606 3763
rect 11623 3715 12077 3763
rect 11623 3385 11685 3715
rect 12015 3385 12077 3715
rect 11623 3337 12077 3385
rect 12094 3337 12097 3763
rect 11603 3331 12097 3337
rect 12153 3763 12647 3769
rect 12153 3337 12156 3763
rect 12173 3715 12627 3763
rect 12173 3385 12235 3715
rect 12565 3385 12627 3715
rect 12173 3337 12627 3385
rect 12644 3337 12647 3763
rect 12153 3331 12647 3337
rect 12703 3763 13197 3769
rect 12703 3337 12706 3763
rect 12723 3715 13177 3763
rect 12723 3385 12785 3715
rect 13115 3385 13177 3715
rect 12723 3337 13177 3385
rect 13194 3337 13197 3763
rect 12703 3331 13197 3337
rect 13253 3763 13724 3769
rect 13253 3337 13256 3763
rect 13273 3715 13724 3763
rect 13273 3385 13335 3715
rect 13665 3385 13724 3715
rect 13273 3337 13724 3385
rect 13253 3331 13724 3337
rect -474 3326 -26 3331
rect 76 3326 524 3331
rect 626 3326 1074 3331
rect 1176 3326 1624 3331
rect 1726 3326 2174 3331
rect 2276 3326 2724 3331
rect 2826 3326 3274 3331
rect 3376 3326 3824 3331
rect 3926 3326 4374 3331
rect 4476 3326 4924 3331
rect 5026 3326 5474 3331
rect 5576 3326 6024 3331
rect 6126 3326 6574 3331
rect 6676 3326 7124 3331
rect 7226 3326 7674 3331
rect 7776 3326 8224 3331
rect 8326 3326 8774 3331
rect 8876 3326 9324 3331
rect 9426 3326 9874 3331
rect 9976 3326 10424 3331
rect 10526 3326 10974 3331
rect 11076 3326 11524 3331
rect 11626 3326 12074 3331
rect 12176 3326 12624 3331
rect 12726 3326 13174 3331
rect 13276 3326 13724 3331
rect -1025 3300 -725 3319
rect -469 3323 -31 3326
rect -469 3306 -463 3323
rect -37 3306 -31 3323
rect -469 3303 -31 3306
rect 81 3323 519 3326
rect 81 3306 87 3323
rect 513 3306 519 3323
rect 81 3303 519 3306
rect 631 3323 1069 3326
rect 631 3306 637 3323
rect 1063 3306 1069 3323
rect 631 3303 1069 3306
rect 1181 3323 1619 3326
rect 1181 3306 1187 3323
rect 1613 3306 1619 3323
rect 1181 3303 1619 3306
rect 1731 3323 2169 3326
rect 1731 3306 1737 3323
rect 2163 3306 2169 3323
rect 1731 3303 2169 3306
rect 2281 3323 2719 3326
rect 2281 3306 2287 3323
rect 2713 3306 2719 3323
rect 2281 3303 2719 3306
rect 2831 3323 3269 3326
rect 2831 3306 2837 3323
rect 3263 3306 3269 3323
rect 2831 3303 3269 3306
rect 3381 3323 3819 3326
rect 3381 3306 3387 3323
rect 3813 3306 3819 3323
rect 3381 3303 3819 3306
rect 3931 3323 4369 3326
rect 3931 3306 3937 3323
rect 4363 3306 4369 3323
rect 3931 3303 4369 3306
rect 4481 3323 4919 3326
rect 4481 3306 4487 3323
rect 4913 3306 4919 3323
rect 4481 3303 4919 3306
rect 5031 3323 5469 3326
rect 5031 3306 5037 3323
rect 5463 3306 5469 3323
rect 5031 3303 5469 3306
rect 5581 3323 6019 3326
rect 5581 3306 5587 3323
rect 6013 3306 6019 3323
rect 5581 3303 6019 3306
rect 6131 3323 6569 3326
rect 6131 3306 6137 3323
rect 6563 3306 6569 3323
rect 6131 3303 6569 3306
rect 6681 3323 7119 3326
rect 6681 3306 6687 3323
rect 7113 3306 7119 3323
rect 6681 3303 7119 3306
rect 7231 3323 7669 3326
rect 7231 3306 7237 3323
rect 7663 3306 7669 3323
rect 7231 3303 7669 3306
rect 7781 3323 8219 3326
rect 7781 3306 7787 3323
rect 8213 3306 8219 3323
rect 7781 3303 8219 3306
rect 8331 3323 8769 3326
rect 8331 3306 8337 3323
rect 8763 3306 8769 3323
rect 8331 3303 8769 3306
rect 8881 3323 9319 3326
rect 8881 3306 8887 3323
rect 9313 3306 9319 3323
rect 8881 3303 9319 3306
rect 9431 3323 9869 3326
rect 9431 3306 9437 3323
rect 9863 3306 9869 3323
rect 9431 3303 9869 3306
rect 9981 3323 10419 3326
rect 9981 3306 9987 3323
rect 10413 3306 10419 3323
rect 9981 3303 10419 3306
rect 10531 3323 10969 3326
rect 10531 3306 10537 3323
rect 10963 3306 10969 3323
rect 10531 3303 10969 3306
rect 11081 3323 11519 3326
rect 11081 3306 11087 3323
rect 11513 3306 11519 3323
rect 11081 3303 11519 3306
rect 11631 3323 12069 3326
rect 11631 3306 11637 3323
rect 12063 3306 12069 3323
rect 11631 3303 12069 3306
rect 12181 3323 12619 3326
rect 12181 3306 12187 3323
rect 12613 3306 12619 3323
rect 12181 3303 12619 3306
rect 12731 3323 13169 3326
rect 12731 3306 12737 3323
rect 13163 3306 13169 3323
rect 12731 3303 13169 3306
rect 13281 3323 13719 3326
rect 13281 3306 13287 3323
rect 13713 3306 13719 3323
rect 13281 3303 13719 3306
rect 13975 3319 13987 3850
rect 14263 3319 14275 3850
rect 13975 3300 14275 3319
rect -1025 2769 -1013 3300
rect -737 2769 -725 3300
rect -550 3292 -500 3300
rect -550 3258 -542 3292
rect -508 3258 -500 3292
rect -550 3250 -500 3258
rect 0 3292 50 3300
rect 0 3258 8 3292
rect 42 3258 50 3292
rect 0 3250 50 3258
rect 550 3292 600 3300
rect 550 3258 558 3292
rect 592 3258 600 3292
rect 550 3250 600 3258
rect 1100 3292 1150 3300
rect 1100 3258 1108 3292
rect 1142 3258 1150 3292
rect 1100 3250 1150 3258
rect 1650 3292 1700 3300
rect 1650 3258 1658 3292
rect 1692 3258 1700 3292
rect 1650 3250 1700 3258
rect 2200 3292 2250 3300
rect 2200 3258 2208 3292
rect 2242 3258 2250 3292
rect 2200 3250 2250 3258
rect 2750 3292 2800 3300
rect 2750 3258 2758 3292
rect 2792 3258 2800 3292
rect 2750 3250 2800 3258
rect 3300 3292 3350 3300
rect 3300 3258 3308 3292
rect 3342 3258 3350 3292
rect 3300 3250 3350 3258
rect 3850 3292 3900 3300
rect 3850 3258 3858 3292
rect 3892 3258 3900 3292
rect 3850 3250 3900 3258
rect 4400 3292 4450 3300
rect 4400 3258 4408 3292
rect 4442 3258 4450 3292
rect 4400 3250 4450 3258
rect 4950 3292 5000 3300
rect 4950 3258 4958 3292
rect 4992 3258 5000 3292
rect 4950 3250 5000 3258
rect 5500 3292 5550 3300
rect 5500 3258 5508 3292
rect 5542 3258 5550 3292
rect 5500 3250 5550 3258
rect 6050 3292 6100 3300
rect 6050 3258 6058 3292
rect 6092 3258 6100 3292
rect 6050 3250 6100 3258
rect 6600 3292 6650 3300
rect 6600 3258 6608 3292
rect 6642 3258 6650 3292
rect 6600 3250 6650 3258
rect 7150 3292 7200 3300
rect 7150 3258 7158 3292
rect 7192 3258 7200 3292
rect 7150 3250 7200 3258
rect 7700 3292 7750 3300
rect 7700 3258 7708 3292
rect 7742 3258 7750 3292
rect 7700 3250 7750 3258
rect 8250 3292 8300 3300
rect 8250 3258 8258 3292
rect 8292 3258 8300 3292
rect 8250 3250 8300 3258
rect 8800 3292 8850 3300
rect 8800 3258 8808 3292
rect 8842 3258 8850 3292
rect 8800 3250 8850 3258
rect 9350 3292 9400 3300
rect 9350 3258 9358 3292
rect 9392 3258 9400 3292
rect 9350 3250 9400 3258
rect 9900 3292 9950 3300
rect 9900 3258 9908 3292
rect 9942 3258 9950 3292
rect 9900 3250 9950 3258
rect 10450 3292 10500 3300
rect 10450 3258 10458 3292
rect 10492 3258 10500 3292
rect 10450 3250 10500 3258
rect 11000 3292 11050 3300
rect 11000 3258 11008 3292
rect 11042 3258 11050 3292
rect 11000 3250 11050 3258
rect 11550 3292 11600 3300
rect 11550 3258 11558 3292
rect 11592 3258 11600 3292
rect 11550 3250 11600 3258
rect 12100 3292 12150 3300
rect 12100 3258 12108 3292
rect 12142 3258 12150 3292
rect 12100 3250 12150 3258
rect 12650 3292 12700 3300
rect 12650 3258 12658 3292
rect 12692 3258 12700 3292
rect 12650 3250 12700 3258
rect 13200 3292 13250 3300
rect 13200 3258 13208 3292
rect 13242 3258 13250 3292
rect 13200 3250 13250 3258
rect 13750 3292 13800 3300
rect 13750 3258 13758 3292
rect 13792 3258 13800 3292
rect 13750 3250 13800 3258
rect -469 3244 -31 3247
rect -469 3227 -463 3244
rect -37 3227 -31 3244
rect -469 3224 -31 3227
rect 81 3244 519 3247
rect 81 3227 87 3244
rect 513 3227 519 3244
rect 81 3224 519 3227
rect 631 3244 1069 3247
rect 631 3227 637 3244
rect 1063 3227 1069 3244
rect 631 3224 1069 3227
rect 1181 3244 1619 3247
rect 1181 3227 1187 3244
rect 1613 3227 1619 3244
rect 1181 3224 1619 3227
rect 1731 3244 2169 3247
rect 1731 3227 1737 3244
rect 2163 3227 2169 3244
rect 1731 3224 2169 3227
rect 2281 3244 2719 3247
rect 2281 3227 2287 3244
rect 2713 3227 2719 3244
rect 2281 3224 2719 3227
rect 2831 3244 3269 3247
rect 2831 3227 2837 3244
rect 3263 3227 3269 3244
rect 2831 3224 3269 3227
rect 3381 3244 3819 3247
rect 3381 3227 3387 3244
rect 3813 3227 3819 3244
rect 3381 3224 3819 3227
rect 3931 3244 4369 3247
rect 3931 3227 3937 3244
rect 4363 3227 4369 3244
rect 3931 3224 4369 3227
rect 4481 3244 4919 3247
rect 4481 3227 4487 3244
rect 4913 3227 4919 3244
rect 4481 3224 4919 3227
rect 5031 3244 5469 3247
rect 5031 3227 5037 3244
rect 5463 3227 5469 3244
rect 5031 3224 5469 3227
rect 5581 3244 6019 3247
rect 5581 3227 5587 3244
rect 6013 3227 6019 3244
rect 5581 3224 6019 3227
rect 6131 3244 6569 3247
rect 6131 3227 6137 3244
rect 6563 3227 6569 3244
rect 6131 3224 6569 3227
rect 6681 3244 7119 3247
rect 6681 3227 6687 3244
rect 7113 3227 7119 3244
rect 6681 3224 7119 3227
rect 7231 3244 7669 3247
rect 7231 3227 7237 3244
rect 7663 3227 7669 3244
rect 7231 3224 7669 3227
rect 7781 3244 8219 3247
rect 7781 3227 7787 3244
rect 8213 3227 8219 3244
rect 7781 3224 8219 3227
rect 8331 3244 8769 3247
rect 8331 3227 8337 3244
rect 8763 3227 8769 3244
rect 8331 3224 8769 3227
rect 8881 3244 9319 3247
rect 8881 3227 8887 3244
rect 9313 3227 9319 3244
rect 8881 3224 9319 3227
rect 9431 3244 9869 3247
rect 9431 3227 9437 3244
rect 9863 3227 9869 3244
rect 9431 3224 9869 3227
rect 9981 3244 10419 3247
rect 9981 3227 9987 3244
rect 10413 3227 10419 3244
rect 9981 3224 10419 3227
rect 10531 3244 10969 3247
rect 10531 3227 10537 3244
rect 10963 3227 10969 3244
rect 10531 3224 10969 3227
rect 11081 3244 11519 3247
rect 11081 3227 11087 3244
rect 11513 3227 11519 3244
rect 11081 3224 11519 3227
rect 11631 3244 12069 3247
rect 11631 3227 11637 3244
rect 12063 3227 12069 3244
rect 11631 3224 12069 3227
rect 12181 3244 12619 3247
rect 12181 3227 12187 3244
rect 12613 3227 12619 3244
rect 12181 3224 12619 3227
rect 12731 3244 13169 3247
rect 12731 3227 12737 3244
rect 13163 3227 13169 3244
rect 12731 3224 13169 3227
rect 13281 3244 13719 3247
rect 13281 3227 13287 3244
rect 13713 3227 13719 3244
rect 13281 3224 13719 3227
rect -474 3219 -26 3224
rect 76 3219 524 3224
rect 626 3219 1074 3224
rect 1176 3219 1624 3224
rect 1726 3219 2174 3224
rect 2276 3219 2724 3224
rect 2826 3219 3274 3224
rect 3376 3219 3824 3224
rect 3926 3219 4374 3224
rect 4476 3219 4924 3224
rect 5026 3219 5474 3224
rect 5576 3219 6024 3224
rect 6126 3219 6574 3224
rect 6676 3219 7124 3224
rect 7226 3219 7674 3224
rect 7776 3219 8224 3224
rect 8326 3219 8774 3224
rect 8876 3219 9324 3224
rect 9426 3219 9874 3224
rect 9976 3219 10424 3224
rect 10526 3219 10974 3224
rect 11076 3219 11524 3224
rect 11626 3219 12074 3224
rect 12176 3219 12624 3224
rect 12726 3219 13174 3224
rect 13276 3219 13724 3224
rect -474 3213 -3 3219
rect -474 3165 -23 3213
rect -474 2835 -415 3165
rect -85 2835 -23 3165
rect -474 2787 -23 2835
rect -6 2787 -3 3213
rect -474 2781 -3 2787
rect 53 3213 547 3219
rect 53 2787 56 3213
rect 73 3165 527 3213
rect 73 2835 135 3165
rect 465 2835 527 3165
rect 73 2787 527 2835
rect 544 2787 547 3213
rect 53 2781 547 2787
rect 603 3213 1097 3219
rect 603 2787 606 3213
rect 623 3165 1077 3213
rect 623 2835 685 3165
rect 1015 2835 1077 3165
rect 623 2787 1077 2835
rect 1094 2787 1097 3213
rect 603 2781 1097 2787
rect 1153 3213 1647 3219
rect 1153 2787 1156 3213
rect 1173 3165 1627 3213
rect 1173 2835 1235 3165
rect 1565 2835 1627 3165
rect 1173 2787 1627 2835
rect 1644 2787 1647 3213
rect 1153 2781 1647 2787
rect 1703 3213 2197 3219
rect 1703 2787 1706 3213
rect 1723 3165 2177 3213
rect 1723 2835 1785 3165
rect 2115 2835 2177 3165
rect 1723 2787 2177 2835
rect 2194 2787 2197 3213
rect 1703 2781 2197 2787
rect 2253 3213 2747 3219
rect 2253 2787 2256 3213
rect 2273 3165 2727 3213
rect 2273 2835 2335 3165
rect 2665 2835 2727 3165
rect 2273 2787 2727 2835
rect 2744 2787 2747 3213
rect 2253 2781 2747 2787
rect 2803 3213 3297 3219
rect 2803 2787 2806 3213
rect 2823 3165 3277 3213
rect 2823 2835 2885 3165
rect 3215 2835 3277 3165
rect 2823 2787 3277 2835
rect 3294 2787 3297 3213
rect 2803 2781 3297 2787
rect 3353 3213 3847 3219
rect 3353 2787 3356 3213
rect 3373 3165 3827 3213
rect 3373 2835 3435 3165
rect 3765 2835 3827 3165
rect 3373 2787 3827 2835
rect 3844 2787 3847 3213
rect 3353 2781 3847 2787
rect 3903 3213 4397 3219
rect 3903 2787 3906 3213
rect 3923 3165 4377 3213
rect 3923 2835 3985 3165
rect 4315 2835 4377 3165
rect 3923 2787 4377 2835
rect 4394 2787 4397 3213
rect 3903 2781 4397 2787
rect 4453 3213 4947 3219
rect 4453 2787 4456 3213
rect 4473 3165 4927 3213
rect 4473 2835 4535 3165
rect 4865 2835 4927 3165
rect 4473 2787 4927 2835
rect 4944 2787 4947 3213
rect 4453 2781 4947 2787
rect 5003 3213 5497 3219
rect 5003 2787 5006 3213
rect 5023 3165 5477 3213
rect 5023 2835 5085 3165
rect 5415 2835 5477 3165
rect 5023 2787 5477 2835
rect 5494 2787 5497 3213
rect 5003 2781 5497 2787
rect 5553 3213 6047 3219
rect 5553 2787 5556 3213
rect 5573 3165 6027 3213
rect 5573 2835 5635 3165
rect 5965 2835 6027 3165
rect 5573 2787 6027 2835
rect 6044 2787 6047 3213
rect 5553 2781 6047 2787
rect 6103 3213 6597 3219
rect 6103 2787 6106 3213
rect 6123 3165 6577 3213
rect 6123 2835 6185 3165
rect 6515 2835 6577 3165
rect 6123 2787 6577 2835
rect 6594 2787 6597 3213
rect 6103 2781 6597 2787
rect 6653 3213 7147 3219
rect 6653 2787 6656 3213
rect 6673 3165 7127 3213
rect 6673 2835 6735 3165
rect 7065 2835 7127 3165
rect 6673 2787 7127 2835
rect 7144 2787 7147 3213
rect 6653 2781 7147 2787
rect 7203 3213 7697 3219
rect 7203 2787 7206 3213
rect 7223 3165 7677 3213
rect 7223 2835 7285 3165
rect 7615 2835 7677 3165
rect 7223 2787 7677 2835
rect 7694 2787 7697 3213
rect 7203 2781 7697 2787
rect 7753 3213 8247 3219
rect 7753 2787 7756 3213
rect 7773 3165 8227 3213
rect 7773 2835 7835 3165
rect 8165 2835 8227 3165
rect 7773 2787 8227 2835
rect 8244 2787 8247 3213
rect 7753 2781 8247 2787
rect 8303 3213 8797 3219
rect 8303 2787 8306 3213
rect 8323 3165 8777 3213
rect 8323 2835 8385 3165
rect 8715 2835 8777 3165
rect 8323 2787 8777 2835
rect 8794 2787 8797 3213
rect 8303 2781 8797 2787
rect 8853 3213 9347 3219
rect 8853 2787 8856 3213
rect 8873 3165 9327 3213
rect 8873 2835 8935 3165
rect 9265 2835 9327 3165
rect 8873 2787 9327 2835
rect 9344 2787 9347 3213
rect 8853 2781 9347 2787
rect 9403 3213 9897 3219
rect 9403 2787 9406 3213
rect 9423 3165 9877 3213
rect 9423 2835 9485 3165
rect 9815 2835 9877 3165
rect 9423 2787 9877 2835
rect 9894 2787 9897 3213
rect 9403 2781 9897 2787
rect 9953 3213 10447 3219
rect 9953 2787 9956 3213
rect 9973 3165 10427 3213
rect 9973 2835 10035 3165
rect 10365 2835 10427 3165
rect 9973 2787 10427 2835
rect 10444 2787 10447 3213
rect 9953 2781 10447 2787
rect 10503 3213 10997 3219
rect 10503 2787 10506 3213
rect 10523 3165 10977 3213
rect 10523 2835 10585 3165
rect 10915 2835 10977 3165
rect 10523 2787 10977 2835
rect 10994 2787 10997 3213
rect 10503 2781 10997 2787
rect 11053 3213 11547 3219
rect 11053 2787 11056 3213
rect 11073 3165 11527 3213
rect 11073 2835 11135 3165
rect 11465 2835 11527 3165
rect 11073 2787 11527 2835
rect 11544 2787 11547 3213
rect 11053 2781 11547 2787
rect 11603 3213 12097 3219
rect 11603 2787 11606 3213
rect 11623 3165 12077 3213
rect 11623 2835 11685 3165
rect 12015 2835 12077 3165
rect 11623 2787 12077 2835
rect 12094 2787 12097 3213
rect 11603 2781 12097 2787
rect 12153 3213 12647 3219
rect 12153 2787 12156 3213
rect 12173 3165 12627 3213
rect 12173 2835 12235 3165
rect 12565 2835 12627 3165
rect 12173 2787 12627 2835
rect 12644 2787 12647 3213
rect 12153 2781 12647 2787
rect 12703 3213 13197 3219
rect 12703 2787 12706 3213
rect 12723 3165 13177 3213
rect 12723 2835 12785 3165
rect 13115 2835 13177 3165
rect 12723 2787 13177 2835
rect 13194 2787 13197 3213
rect 12703 2781 13197 2787
rect 13253 3213 13724 3219
rect 13253 2787 13256 3213
rect 13273 3165 13724 3213
rect 13273 2835 13335 3165
rect 13665 2835 13724 3165
rect 13273 2787 13724 2835
rect 13253 2781 13724 2787
rect -474 2776 -26 2781
rect 76 2776 524 2781
rect 626 2776 1074 2781
rect 1176 2776 1624 2781
rect 1726 2776 2174 2781
rect 2276 2776 2724 2781
rect 2826 2776 3274 2781
rect 3376 2776 3824 2781
rect 3926 2776 4374 2781
rect 4476 2776 4924 2781
rect 5026 2776 5474 2781
rect 5576 2776 6024 2781
rect 6126 2776 6574 2781
rect 6676 2776 7124 2781
rect 7226 2776 7674 2781
rect 7776 2776 8224 2781
rect 8326 2776 8774 2781
rect 8876 2776 9324 2781
rect 9426 2776 9874 2781
rect 9976 2776 10424 2781
rect 10526 2776 10974 2781
rect 11076 2776 11524 2781
rect 11626 2776 12074 2781
rect 12176 2776 12624 2781
rect 12726 2776 13174 2781
rect 13276 2776 13724 2781
rect -1025 2750 -725 2769
rect -469 2773 -31 2776
rect -469 2756 -463 2773
rect -37 2756 -31 2773
rect -469 2753 -31 2756
rect 81 2773 519 2776
rect 81 2756 87 2773
rect 513 2756 519 2773
rect 81 2753 519 2756
rect 631 2773 1069 2776
rect 631 2756 637 2773
rect 1063 2756 1069 2773
rect 631 2753 1069 2756
rect 1181 2773 1619 2776
rect 1181 2756 1187 2773
rect 1613 2756 1619 2773
rect 1181 2753 1619 2756
rect 1731 2773 2169 2776
rect 1731 2756 1737 2773
rect 2163 2756 2169 2773
rect 1731 2753 2169 2756
rect 2281 2773 2719 2776
rect 2281 2756 2287 2773
rect 2713 2756 2719 2773
rect 2281 2753 2719 2756
rect 2831 2773 3269 2776
rect 2831 2756 2837 2773
rect 3263 2756 3269 2773
rect 2831 2753 3269 2756
rect 3381 2773 3819 2776
rect 3381 2756 3387 2773
rect 3813 2756 3819 2773
rect 3381 2753 3819 2756
rect 3931 2773 4369 2776
rect 3931 2756 3937 2773
rect 4363 2756 4369 2773
rect 3931 2753 4369 2756
rect 4481 2773 4919 2776
rect 4481 2756 4487 2773
rect 4913 2756 4919 2773
rect 4481 2753 4919 2756
rect 5031 2773 5469 2776
rect 5031 2756 5037 2773
rect 5463 2756 5469 2773
rect 5031 2753 5469 2756
rect 5581 2773 6019 2776
rect 5581 2756 5587 2773
rect 6013 2756 6019 2773
rect 5581 2753 6019 2756
rect 6131 2773 6569 2776
rect 6131 2756 6137 2773
rect 6563 2756 6569 2773
rect 6131 2753 6569 2756
rect 6681 2773 7119 2776
rect 6681 2756 6687 2773
rect 7113 2756 7119 2773
rect 6681 2753 7119 2756
rect 7231 2773 7669 2776
rect 7231 2756 7237 2773
rect 7663 2756 7669 2773
rect 7231 2753 7669 2756
rect 7781 2773 8219 2776
rect 7781 2756 7787 2773
rect 8213 2756 8219 2773
rect 7781 2753 8219 2756
rect 8331 2773 8769 2776
rect 8331 2756 8337 2773
rect 8763 2756 8769 2773
rect 8331 2753 8769 2756
rect 8881 2773 9319 2776
rect 8881 2756 8887 2773
rect 9313 2756 9319 2773
rect 8881 2753 9319 2756
rect 9431 2773 9869 2776
rect 9431 2756 9437 2773
rect 9863 2756 9869 2773
rect 9431 2753 9869 2756
rect 9981 2773 10419 2776
rect 9981 2756 9987 2773
rect 10413 2756 10419 2773
rect 9981 2753 10419 2756
rect 10531 2773 10969 2776
rect 10531 2756 10537 2773
rect 10963 2756 10969 2773
rect 10531 2753 10969 2756
rect 11081 2773 11519 2776
rect 11081 2756 11087 2773
rect 11513 2756 11519 2773
rect 11081 2753 11519 2756
rect 11631 2773 12069 2776
rect 11631 2756 11637 2773
rect 12063 2756 12069 2773
rect 11631 2753 12069 2756
rect 12181 2773 12619 2776
rect 12181 2756 12187 2773
rect 12613 2756 12619 2773
rect 12181 2753 12619 2756
rect 12731 2773 13169 2776
rect 12731 2756 12737 2773
rect 13163 2756 13169 2773
rect 12731 2753 13169 2756
rect 13281 2773 13719 2776
rect 13281 2756 13287 2773
rect 13713 2756 13719 2773
rect 13281 2753 13719 2756
rect 13975 2769 13987 3300
rect 14263 2769 14275 3300
rect 13975 2750 14275 2769
rect -1025 2219 -1013 2750
rect -737 2219 -725 2750
rect -550 2742 -500 2750
rect -550 2708 -542 2742
rect -508 2708 -500 2742
rect -550 2700 -500 2708
rect 0 2742 50 2750
rect 0 2708 8 2742
rect 42 2708 50 2742
rect 0 2700 50 2708
rect 550 2742 600 2750
rect 550 2708 558 2742
rect 592 2708 600 2742
rect 550 2700 600 2708
rect 1100 2742 1150 2750
rect 1100 2708 1108 2742
rect 1142 2708 1150 2742
rect 1100 2700 1150 2708
rect 1650 2742 1700 2750
rect 1650 2708 1658 2742
rect 1692 2708 1700 2742
rect 1650 2700 1700 2708
rect 2200 2742 2250 2750
rect 2200 2708 2208 2742
rect 2242 2708 2250 2742
rect 2200 2700 2250 2708
rect 2750 2742 2800 2750
rect 2750 2708 2758 2742
rect 2792 2708 2800 2742
rect 2750 2700 2800 2708
rect 3300 2742 3350 2750
rect 3300 2708 3308 2742
rect 3342 2708 3350 2742
rect 3300 2700 3350 2708
rect 3850 2742 3900 2750
rect 3850 2708 3858 2742
rect 3892 2708 3900 2742
rect 3850 2700 3900 2708
rect 4400 2742 4450 2750
rect 4400 2708 4408 2742
rect 4442 2708 4450 2742
rect 4400 2700 4450 2708
rect 4950 2742 5000 2750
rect 4950 2708 4958 2742
rect 4992 2708 5000 2742
rect 4950 2700 5000 2708
rect 5500 2742 5550 2750
rect 5500 2708 5508 2742
rect 5542 2708 5550 2742
rect 5500 2700 5550 2708
rect 6050 2742 6100 2750
rect 6050 2708 6058 2742
rect 6092 2708 6100 2742
rect 6050 2700 6100 2708
rect 6600 2742 6650 2750
rect 6600 2708 6608 2742
rect 6642 2708 6650 2742
rect 6600 2700 6650 2708
rect 7150 2742 7200 2750
rect 7150 2708 7158 2742
rect 7192 2708 7200 2742
rect 7150 2700 7200 2708
rect 7700 2742 7750 2750
rect 7700 2708 7708 2742
rect 7742 2708 7750 2742
rect 7700 2700 7750 2708
rect 8250 2742 8300 2750
rect 8250 2708 8258 2742
rect 8292 2708 8300 2742
rect 8250 2700 8300 2708
rect 8800 2742 8850 2750
rect 8800 2708 8808 2742
rect 8842 2708 8850 2742
rect 8800 2700 8850 2708
rect 9350 2742 9400 2750
rect 9350 2708 9358 2742
rect 9392 2708 9400 2742
rect 9350 2700 9400 2708
rect 9900 2742 9950 2750
rect 9900 2708 9908 2742
rect 9942 2708 9950 2742
rect 9900 2700 9950 2708
rect 10450 2742 10500 2750
rect 10450 2708 10458 2742
rect 10492 2708 10500 2742
rect 10450 2700 10500 2708
rect 11000 2742 11050 2750
rect 11000 2708 11008 2742
rect 11042 2708 11050 2742
rect 11000 2700 11050 2708
rect 11550 2742 11600 2750
rect 11550 2708 11558 2742
rect 11592 2708 11600 2742
rect 11550 2700 11600 2708
rect 12100 2742 12150 2750
rect 12100 2708 12108 2742
rect 12142 2708 12150 2742
rect 12100 2700 12150 2708
rect 12650 2742 12700 2750
rect 12650 2708 12658 2742
rect 12692 2708 12700 2742
rect 12650 2700 12700 2708
rect 13200 2742 13250 2750
rect 13200 2708 13208 2742
rect 13242 2708 13250 2742
rect 13200 2700 13250 2708
rect 13750 2742 13800 2750
rect 13750 2708 13758 2742
rect 13792 2708 13800 2742
rect 13750 2700 13800 2708
rect -469 2694 -31 2697
rect -469 2677 -463 2694
rect -37 2677 -31 2694
rect -469 2674 -31 2677
rect 81 2694 519 2697
rect 81 2677 87 2694
rect 513 2677 519 2694
rect 81 2674 519 2677
rect 631 2694 1069 2697
rect 631 2677 637 2694
rect 1063 2677 1069 2694
rect 631 2674 1069 2677
rect 1181 2694 1619 2697
rect 1181 2677 1187 2694
rect 1613 2677 1619 2694
rect 1181 2674 1619 2677
rect 1731 2694 2169 2697
rect 1731 2677 1737 2694
rect 2163 2677 2169 2694
rect 1731 2674 2169 2677
rect 2281 2694 2719 2697
rect 2281 2677 2287 2694
rect 2713 2677 2719 2694
rect 2281 2674 2719 2677
rect 2831 2694 3269 2697
rect 2831 2677 2837 2694
rect 3263 2677 3269 2694
rect 2831 2674 3269 2677
rect 3381 2694 3819 2697
rect 3381 2677 3387 2694
rect 3813 2677 3819 2694
rect 3381 2674 3819 2677
rect 3931 2694 4369 2697
rect 3931 2677 3937 2694
rect 4363 2677 4369 2694
rect 3931 2674 4369 2677
rect 4481 2694 4919 2697
rect 4481 2677 4487 2694
rect 4913 2677 4919 2694
rect 4481 2674 4919 2677
rect 5031 2694 5469 2697
rect 5031 2677 5037 2694
rect 5463 2677 5469 2694
rect 5031 2674 5469 2677
rect 5581 2694 6019 2697
rect 5581 2677 5587 2694
rect 6013 2677 6019 2694
rect 5581 2674 6019 2677
rect 6131 2694 6569 2697
rect 6131 2677 6137 2694
rect 6563 2677 6569 2694
rect 6131 2674 6569 2677
rect 6681 2694 7119 2697
rect 6681 2677 6687 2694
rect 7113 2677 7119 2694
rect 6681 2674 7119 2677
rect 7231 2694 7669 2697
rect 7231 2677 7237 2694
rect 7663 2677 7669 2694
rect 7231 2674 7669 2677
rect 7781 2694 8219 2697
rect 7781 2677 7787 2694
rect 8213 2677 8219 2694
rect 7781 2674 8219 2677
rect 8331 2694 8769 2697
rect 8331 2677 8337 2694
rect 8763 2677 8769 2694
rect 8331 2674 8769 2677
rect 8881 2694 9319 2697
rect 8881 2677 8887 2694
rect 9313 2677 9319 2694
rect 8881 2674 9319 2677
rect 9431 2694 9869 2697
rect 9431 2677 9437 2694
rect 9863 2677 9869 2694
rect 9431 2674 9869 2677
rect 9981 2694 10419 2697
rect 9981 2677 9987 2694
rect 10413 2677 10419 2694
rect 9981 2674 10419 2677
rect 10531 2694 10969 2697
rect 10531 2677 10537 2694
rect 10963 2677 10969 2694
rect 10531 2674 10969 2677
rect 11081 2694 11519 2697
rect 11081 2677 11087 2694
rect 11513 2677 11519 2694
rect 11081 2674 11519 2677
rect 11631 2694 12069 2697
rect 11631 2677 11637 2694
rect 12063 2677 12069 2694
rect 11631 2674 12069 2677
rect 12181 2694 12619 2697
rect 12181 2677 12187 2694
rect 12613 2677 12619 2694
rect 12181 2674 12619 2677
rect 12731 2694 13169 2697
rect 12731 2677 12737 2694
rect 13163 2677 13169 2694
rect 12731 2674 13169 2677
rect 13281 2694 13719 2697
rect 13281 2677 13287 2694
rect 13713 2677 13719 2694
rect 13281 2674 13719 2677
rect -474 2669 -26 2674
rect 76 2669 524 2674
rect 626 2669 1074 2674
rect 1176 2669 1624 2674
rect 1726 2669 2174 2674
rect 2276 2669 2724 2674
rect 2826 2669 3274 2674
rect 3376 2669 3824 2674
rect 3926 2669 4374 2674
rect 4476 2669 4924 2674
rect 5026 2669 5474 2674
rect 5576 2669 6024 2674
rect 6126 2669 6574 2674
rect 6676 2669 7124 2674
rect 7226 2669 7674 2674
rect 7776 2669 8224 2674
rect 8326 2669 8774 2674
rect 8876 2669 9324 2674
rect 9426 2669 9874 2674
rect 9976 2669 10424 2674
rect 10526 2669 10974 2674
rect 11076 2669 11524 2674
rect 11626 2669 12074 2674
rect 12176 2669 12624 2674
rect 12726 2669 13174 2674
rect 13276 2669 13724 2674
rect -474 2663 -3 2669
rect -474 2615 -23 2663
rect -474 2285 -415 2615
rect -85 2285 -23 2615
rect -474 2237 -23 2285
rect -6 2237 -3 2663
rect -474 2231 -3 2237
rect 53 2663 547 2669
rect 53 2237 56 2663
rect 73 2615 527 2663
rect 73 2285 135 2615
rect 465 2285 527 2615
rect 73 2237 527 2285
rect 544 2237 547 2663
rect 53 2231 547 2237
rect 603 2663 1097 2669
rect 603 2237 606 2663
rect 623 2615 1077 2663
rect 623 2285 685 2615
rect 1015 2285 1077 2615
rect 623 2237 1077 2285
rect 1094 2237 1097 2663
rect 603 2231 1097 2237
rect 1153 2663 1647 2669
rect 1153 2237 1156 2663
rect 1173 2615 1627 2663
rect 1173 2285 1235 2615
rect 1565 2285 1627 2615
rect 1173 2237 1627 2285
rect 1644 2237 1647 2663
rect 1153 2231 1647 2237
rect 1703 2663 2197 2669
rect 1703 2237 1706 2663
rect 1723 2615 2177 2663
rect 1723 2285 1785 2615
rect 2115 2285 2177 2615
rect 1723 2237 2177 2285
rect 2194 2237 2197 2663
rect 1703 2231 2197 2237
rect 2253 2663 2747 2669
rect 2253 2237 2256 2663
rect 2273 2615 2727 2663
rect 2273 2285 2335 2615
rect 2665 2285 2727 2615
rect 2273 2237 2727 2285
rect 2744 2237 2747 2663
rect 2253 2231 2747 2237
rect 2803 2663 3297 2669
rect 2803 2237 2806 2663
rect 2823 2615 3277 2663
rect 2823 2285 2885 2615
rect 3215 2285 3277 2615
rect 2823 2237 3277 2285
rect 3294 2237 3297 2663
rect 2803 2231 3297 2237
rect 3353 2663 3847 2669
rect 3353 2237 3356 2663
rect 3373 2615 3827 2663
rect 3373 2285 3435 2615
rect 3765 2285 3827 2615
rect 3373 2237 3827 2285
rect 3844 2237 3847 2663
rect 3353 2231 3847 2237
rect 3903 2663 4397 2669
rect 3903 2237 3906 2663
rect 3923 2615 4377 2663
rect 3923 2285 3985 2615
rect 4315 2285 4377 2615
rect 3923 2237 4377 2285
rect 4394 2237 4397 2663
rect 3903 2231 4397 2237
rect 4453 2663 4947 2669
rect 4453 2237 4456 2663
rect 4473 2615 4927 2663
rect 4473 2285 4535 2615
rect 4865 2285 4927 2615
rect 4473 2237 4927 2285
rect 4944 2237 4947 2663
rect 4453 2231 4947 2237
rect 5003 2663 5497 2669
rect 5003 2237 5006 2663
rect 5023 2615 5477 2663
rect 5023 2285 5085 2615
rect 5415 2285 5477 2615
rect 5023 2237 5477 2285
rect 5494 2237 5497 2663
rect 5003 2231 5497 2237
rect 5553 2663 6047 2669
rect 5553 2237 5556 2663
rect 5573 2615 6027 2663
rect 5573 2285 5635 2615
rect 5965 2285 6027 2615
rect 5573 2237 6027 2285
rect 6044 2237 6047 2663
rect 5553 2231 6047 2237
rect 6103 2663 6597 2669
rect 6103 2237 6106 2663
rect 6123 2615 6577 2663
rect 6123 2285 6185 2615
rect 6515 2285 6577 2615
rect 6123 2237 6577 2285
rect 6594 2237 6597 2663
rect 6103 2231 6597 2237
rect 6653 2663 7147 2669
rect 6653 2237 6656 2663
rect 6673 2615 7127 2663
rect 6673 2285 6735 2615
rect 7065 2285 7127 2615
rect 6673 2237 7127 2285
rect 7144 2237 7147 2663
rect 6653 2231 7147 2237
rect 7203 2663 7697 2669
rect 7203 2237 7206 2663
rect 7223 2615 7677 2663
rect 7223 2285 7285 2615
rect 7615 2285 7677 2615
rect 7223 2237 7677 2285
rect 7694 2237 7697 2663
rect 7203 2231 7697 2237
rect 7753 2663 8247 2669
rect 7753 2237 7756 2663
rect 7773 2615 8227 2663
rect 7773 2285 7835 2615
rect 8165 2285 8227 2615
rect 7773 2237 8227 2285
rect 8244 2237 8247 2663
rect 7753 2231 8247 2237
rect 8303 2663 8797 2669
rect 8303 2237 8306 2663
rect 8323 2615 8777 2663
rect 8323 2285 8385 2615
rect 8715 2285 8777 2615
rect 8323 2237 8777 2285
rect 8794 2237 8797 2663
rect 8303 2231 8797 2237
rect 8853 2663 9347 2669
rect 8853 2237 8856 2663
rect 8873 2615 9327 2663
rect 8873 2285 8935 2615
rect 9265 2285 9327 2615
rect 8873 2237 9327 2285
rect 9344 2237 9347 2663
rect 8853 2231 9347 2237
rect 9403 2663 9897 2669
rect 9403 2237 9406 2663
rect 9423 2615 9877 2663
rect 9423 2285 9485 2615
rect 9815 2285 9877 2615
rect 9423 2237 9877 2285
rect 9894 2237 9897 2663
rect 9403 2231 9897 2237
rect 9953 2663 10447 2669
rect 9953 2237 9956 2663
rect 9973 2615 10427 2663
rect 9973 2285 10035 2615
rect 10365 2285 10427 2615
rect 9973 2237 10427 2285
rect 10444 2237 10447 2663
rect 9953 2231 10447 2237
rect 10503 2663 10997 2669
rect 10503 2237 10506 2663
rect 10523 2615 10977 2663
rect 10523 2285 10585 2615
rect 10915 2285 10977 2615
rect 10523 2237 10977 2285
rect 10994 2237 10997 2663
rect 10503 2231 10997 2237
rect 11053 2663 11547 2669
rect 11053 2237 11056 2663
rect 11073 2615 11527 2663
rect 11073 2285 11135 2615
rect 11465 2285 11527 2615
rect 11073 2237 11527 2285
rect 11544 2237 11547 2663
rect 11053 2231 11547 2237
rect 11603 2663 12097 2669
rect 11603 2237 11606 2663
rect 11623 2615 12077 2663
rect 11623 2285 11685 2615
rect 12015 2285 12077 2615
rect 11623 2237 12077 2285
rect 12094 2237 12097 2663
rect 11603 2231 12097 2237
rect 12153 2663 12647 2669
rect 12153 2237 12156 2663
rect 12173 2615 12627 2663
rect 12173 2285 12235 2615
rect 12565 2285 12627 2615
rect 12173 2237 12627 2285
rect 12644 2237 12647 2663
rect 12153 2231 12647 2237
rect 12703 2663 13197 2669
rect 12703 2237 12706 2663
rect 12723 2615 13177 2663
rect 12723 2285 12785 2615
rect 13115 2285 13177 2615
rect 12723 2237 13177 2285
rect 13194 2237 13197 2663
rect 12703 2231 13197 2237
rect 13253 2663 13724 2669
rect 13253 2237 13256 2663
rect 13273 2615 13724 2663
rect 13273 2285 13335 2615
rect 13665 2285 13724 2615
rect 13273 2237 13724 2285
rect 13253 2231 13724 2237
rect -474 2226 -26 2231
rect 76 2226 524 2231
rect 626 2226 1074 2231
rect 1176 2226 1624 2231
rect 1726 2226 2174 2231
rect 2276 2226 2724 2231
rect 2826 2226 3274 2231
rect 3376 2226 3824 2231
rect 3926 2226 4374 2231
rect 4476 2226 4924 2231
rect 5026 2226 5474 2231
rect 5576 2226 6024 2231
rect 6126 2226 6574 2231
rect 6676 2226 7124 2231
rect 7226 2226 7674 2231
rect 7776 2226 8224 2231
rect 8326 2226 8774 2231
rect 8876 2226 9324 2231
rect 9426 2226 9874 2231
rect 9976 2226 10424 2231
rect 10526 2226 10974 2231
rect 11076 2226 11524 2231
rect 11626 2226 12074 2231
rect 12176 2226 12624 2231
rect 12726 2226 13174 2231
rect 13276 2226 13724 2231
rect -1025 2200 -725 2219
rect -469 2223 -31 2226
rect -469 2206 -463 2223
rect -37 2206 -31 2223
rect -469 2203 -31 2206
rect 81 2223 519 2226
rect 81 2206 87 2223
rect 513 2206 519 2223
rect 81 2203 519 2206
rect 631 2223 1069 2226
rect 631 2206 637 2223
rect 1063 2206 1069 2223
rect 631 2203 1069 2206
rect 1181 2223 1619 2226
rect 1181 2206 1187 2223
rect 1613 2206 1619 2223
rect 1181 2203 1619 2206
rect 1731 2223 2169 2226
rect 1731 2206 1737 2223
rect 2163 2206 2169 2223
rect 1731 2203 2169 2206
rect 2281 2223 2719 2226
rect 2281 2206 2287 2223
rect 2713 2206 2719 2223
rect 2281 2203 2719 2206
rect 2831 2223 3269 2226
rect 2831 2206 2837 2223
rect 3263 2206 3269 2223
rect 2831 2203 3269 2206
rect 3381 2223 3819 2226
rect 3381 2206 3387 2223
rect 3813 2206 3819 2223
rect 3381 2203 3819 2206
rect 3931 2223 4369 2226
rect 3931 2206 3937 2223
rect 4363 2206 4369 2223
rect 3931 2203 4369 2206
rect 4481 2223 4919 2226
rect 4481 2206 4487 2223
rect 4913 2206 4919 2223
rect 4481 2203 4919 2206
rect 5031 2223 5469 2226
rect 5031 2206 5037 2223
rect 5463 2206 5469 2223
rect 5031 2203 5469 2206
rect 5581 2223 6019 2226
rect 5581 2206 5587 2223
rect 6013 2206 6019 2223
rect 5581 2203 6019 2206
rect 6131 2223 6569 2226
rect 6131 2206 6137 2223
rect 6563 2206 6569 2223
rect 6131 2203 6569 2206
rect 6681 2223 7119 2226
rect 6681 2206 6687 2223
rect 7113 2206 7119 2223
rect 6681 2203 7119 2206
rect 7231 2223 7669 2226
rect 7231 2206 7237 2223
rect 7663 2206 7669 2223
rect 7231 2203 7669 2206
rect 7781 2223 8219 2226
rect 7781 2206 7787 2223
rect 8213 2206 8219 2223
rect 7781 2203 8219 2206
rect 8331 2223 8769 2226
rect 8331 2206 8337 2223
rect 8763 2206 8769 2223
rect 8331 2203 8769 2206
rect 8881 2223 9319 2226
rect 8881 2206 8887 2223
rect 9313 2206 9319 2223
rect 8881 2203 9319 2206
rect 9431 2223 9869 2226
rect 9431 2206 9437 2223
rect 9863 2206 9869 2223
rect 9431 2203 9869 2206
rect 9981 2223 10419 2226
rect 9981 2206 9987 2223
rect 10413 2206 10419 2223
rect 9981 2203 10419 2206
rect 10531 2223 10969 2226
rect 10531 2206 10537 2223
rect 10963 2206 10969 2223
rect 10531 2203 10969 2206
rect 11081 2223 11519 2226
rect 11081 2206 11087 2223
rect 11513 2206 11519 2223
rect 11081 2203 11519 2206
rect 11631 2223 12069 2226
rect 11631 2206 11637 2223
rect 12063 2206 12069 2223
rect 11631 2203 12069 2206
rect 12181 2223 12619 2226
rect 12181 2206 12187 2223
rect 12613 2206 12619 2223
rect 12181 2203 12619 2206
rect 12731 2223 13169 2226
rect 12731 2206 12737 2223
rect 13163 2206 13169 2223
rect 12731 2203 13169 2206
rect 13281 2223 13719 2226
rect 13281 2206 13287 2223
rect 13713 2206 13719 2223
rect 13281 2203 13719 2206
rect 13975 2219 13987 2750
rect 14263 2219 14275 2750
rect 13975 2200 14275 2219
rect -1025 1669 -1013 2200
rect -737 1669 -725 2200
rect -550 2192 -500 2200
rect -550 2158 -542 2192
rect -508 2158 -500 2192
rect -550 2150 -500 2158
rect 0 2192 50 2200
rect 0 2158 8 2192
rect 42 2158 50 2192
rect 0 2150 50 2158
rect 550 2192 600 2200
rect 550 2158 558 2192
rect 592 2158 600 2192
rect 550 2150 600 2158
rect 1100 2192 1150 2200
rect 1100 2158 1108 2192
rect 1142 2158 1150 2192
rect 1100 2150 1150 2158
rect 1650 2192 1700 2200
rect 1650 2158 1658 2192
rect 1692 2158 1700 2192
rect 1650 2150 1700 2158
rect 2200 2192 2250 2200
rect 2200 2158 2208 2192
rect 2242 2158 2250 2192
rect 2200 2150 2250 2158
rect 2750 2192 2800 2200
rect 2750 2158 2758 2192
rect 2792 2158 2800 2192
rect 2750 2150 2800 2158
rect 3300 2192 3350 2200
rect 3300 2158 3308 2192
rect 3342 2158 3350 2192
rect 3300 2150 3350 2158
rect 3850 2192 3900 2200
rect 3850 2158 3858 2192
rect 3892 2158 3900 2192
rect 3850 2150 3900 2158
rect 4400 2192 4450 2200
rect 4400 2158 4408 2192
rect 4442 2158 4450 2192
rect 4400 2150 4450 2158
rect 4950 2192 5000 2200
rect 4950 2158 4958 2192
rect 4992 2158 5000 2192
rect 4950 2150 5000 2158
rect 5500 2192 5550 2200
rect 5500 2158 5508 2192
rect 5542 2158 5550 2192
rect 5500 2150 5550 2158
rect 6050 2192 6100 2200
rect 6050 2158 6058 2192
rect 6092 2158 6100 2192
rect 6050 2150 6100 2158
rect 6600 2192 6650 2200
rect 6600 2158 6608 2192
rect 6642 2158 6650 2192
rect 6600 2150 6650 2158
rect 7150 2192 7200 2200
rect 7150 2158 7158 2192
rect 7192 2158 7200 2192
rect 7150 2150 7200 2158
rect 7700 2192 7750 2200
rect 7700 2158 7708 2192
rect 7742 2158 7750 2192
rect 7700 2150 7750 2158
rect 8250 2192 8300 2200
rect 8250 2158 8258 2192
rect 8292 2158 8300 2192
rect 8250 2150 8300 2158
rect 8800 2192 8850 2200
rect 8800 2158 8808 2192
rect 8842 2158 8850 2192
rect 8800 2150 8850 2158
rect 9350 2192 9400 2200
rect 9350 2158 9358 2192
rect 9392 2158 9400 2192
rect 9350 2150 9400 2158
rect 9900 2192 9950 2200
rect 9900 2158 9908 2192
rect 9942 2158 9950 2192
rect 9900 2150 9950 2158
rect 10450 2192 10500 2200
rect 10450 2158 10458 2192
rect 10492 2158 10500 2192
rect 10450 2150 10500 2158
rect 11000 2192 11050 2200
rect 11000 2158 11008 2192
rect 11042 2158 11050 2192
rect 11000 2150 11050 2158
rect 11550 2192 11600 2200
rect 11550 2158 11558 2192
rect 11592 2158 11600 2192
rect 11550 2150 11600 2158
rect 12100 2192 12150 2200
rect 12100 2158 12108 2192
rect 12142 2158 12150 2192
rect 12100 2150 12150 2158
rect 12650 2192 12700 2200
rect 12650 2158 12658 2192
rect 12692 2158 12700 2192
rect 12650 2150 12700 2158
rect 13200 2192 13250 2200
rect 13200 2158 13208 2192
rect 13242 2158 13250 2192
rect 13200 2150 13250 2158
rect 13750 2192 13800 2200
rect 13750 2158 13758 2192
rect 13792 2158 13800 2192
rect 13750 2150 13800 2158
rect -469 2144 -31 2147
rect -469 2127 -463 2144
rect -37 2127 -31 2144
rect -469 2124 -31 2127
rect 81 2144 519 2147
rect 81 2127 87 2144
rect 513 2127 519 2144
rect 81 2124 519 2127
rect 631 2144 1069 2147
rect 631 2127 637 2144
rect 1063 2127 1069 2144
rect 631 2124 1069 2127
rect 1181 2144 1619 2147
rect 1181 2127 1187 2144
rect 1613 2127 1619 2144
rect 1181 2124 1619 2127
rect 1731 2144 2169 2147
rect 1731 2127 1737 2144
rect 2163 2127 2169 2144
rect 1731 2124 2169 2127
rect 2281 2144 2719 2147
rect 2281 2127 2287 2144
rect 2713 2127 2719 2144
rect 2281 2124 2719 2127
rect 2831 2144 3269 2147
rect 2831 2127 2837 2144
rect 3263 2127 3269 2144
rect 2831 2124 3269 2127
rect 3381 2144 3819 2147
rect 3381 2127 3387 2144
rect 3813 2127 3819 2144
rect 3381 2124 3819 2127
rect 3931 2144 4369 2147
rect 3931 2127 3937 2144
rect 4363 2127 4369 2144
rect 3931 2124 4369 2127
rect 4481 2144 4919 2147
rect 4481 2127 4487 2144
rect 4913 2127 4919 2144
rect 4481 2124 4919 2127
rect 5031 2144 5469 2147
rect 5031 2127 5037 2144
rect 5463 2127 5469 2144
rect 5031 2124 5469 2127
rect 5581 2144 6019 2147
rect 5581 2127 5587 2144
rect 6013 2127 6019 2144
rect 5581 2124 6019 2127
rect 6131 2144 6569 2147
rect 6131 2127 6137 2144
rect 6563 2127 6569 2144
rect 6131 2124 6569 2127
rect 6681 2144 7119 2147
rect 6681 2127 6687 2144
rect 7113 2127 7119 2144
rect 6681 2124 7119 2127
rect 7231 2144 7669 2147
rect 7231 2127 7237 2144
rect 7663 2127 7669 2144
rect 7231 2124 7669 2127
rect 7781 2144 8219 2147
rect 7781 2127 7787 2144
rect 8213 2127 8219 2144
rect 7781 2124 8219 2127
rect 8331 2144 8769 2147
rect 8331 2127 8337 2144
rect 8763 2127 8769 2144
rect 8331 2124 8769 2127
rect 8881 2144 9319 2147
rect 8881 2127 8887 2144
rect 9313 2127 9319 2144
rect 8881 2124 9319 2127
rect 9431 2144 9869 2147
rect 9431 2127 9437 2144
rect 9863 2127 9869 2144
rect 9431 2124 9869 2127
rect 9981 2144 10419 2147
rect 9981 2127 9987 2144
rect 10413 2127 10419 2144
rect 9981 2124 10419 2127
rect 10531 2144 10969 2147
rect 10531 2127 10537 2144
rect 10963 2127 10969 2144
rect 10531 2124 10969 2127
rect 11081 2144 11519 2147
rect 11081 2127 11087 2144
rect 11513 2127 11519 2144
rect 11081 2124 11519 2127
rect 11631 2144 12069 2147
rect 11631 2127 11637 2144
rect 12063 2127 12069 2144
rect 11631 2124 12069 2127
rect 12181 2144 12619 2147
rect 12181 2127 12187 2144
rect 12613 2127 12619 2144
rect 12181 2124 12619 2127
rect 12731 2144 13169 2147
rect 12731 2127 12737 2144
rect 13163 2127 13169 2144
rect 12731 2124 13169 2127
rect 13281 2144 13719 2147
rect 13281 2127 13287 2144
rect 13713 2127 13719 2144
rect 13281 2124 13719 2127
rect -474 2119 -26 2124
rect 76 2119 524 2124
rect 626 2119 1074 2124
rect 1176 2119 1624 2124
rect 1726 2119 2174 2124
rect 2276 2119 2724 2124
rect 2826 2119 3274 2124
rect 3376 2119 3824 2124
rect 3926 2119 4374 2124
rect 4476 2119 4924 2124
rect 5026 2119 5474 2124
rect 5576 2119 6024 2124
rect 6126 2119 6574 2124
rect 6676 2119 7124 2124
rect 7226 2119 7674 2124
rect 7776 2119 8224 2124
rect 8326 2119 8774 2124
rect 8876 2119 9324 2124
rect 9426 2119 9874 2124
rect 9976 2119 10424 2124
rect 10526 2119 10974 2124
rect 11076 2119 11524 2124
rect 11626 2119 12074 2124
rect 12176 2119 12624 2124
rect 12726 2119 13174 2124
rect 13276 2119 13724 2124
rect -474 2113 -3 2119
rect -474 2065 -23 2113
rect -474 1735 -415 2065
rect -85 1735 -23 2065
rect -474 1687 -23 1735
rect -6 1687 -3 2113
rect -474 1681 -3 1687
rect 53 2113 547 2119
rect 53 1687 56 2113
rect 73 2065 527 2113
rect 73 1735 135 2065
rect 465 1735 527 2065
rect 73 1687 527 1735
rect 544 1687 547 2113
rect 53 1681 547 1687
rect 603 2113 1097 2119
rect 603 1687 606 2113
rect 623 2065 1077 2113
rect 623 1735 685 2065
rect 1015 1735 1077 2065
rect 623 1687 1077 1735
rect 1094 1687 1097 2113
rect 603 1681 1097 1687
rect 1153 2113 1647 2119
rect 1153 1687 1156 2113
rect 1173 2065 1627 2113
rect 1173 1735 1235 2065
rect 1565 1735 1627 2065
rect 1173 1687 1627 1735
rect 1644 1687 1647 2113
rect 1153 1681 1647 1687
rect 1703 2113 2197 2119
rect 1703 1687 1706 2113
rect 1723 2065 2177 2113
rect 1723 1735 1785 2065
rect 2115 1735 2177 2065
rect 1723 1687 2177 1735
rect 2194 1687 2197 2113
rect 1703 1681 2197 1687
rect 2253 2113 2747 2119
rect 2253 1687 2256 2113
rect 2273 2065 2727 2113
rect 2273 1735 2335 2065
rect 2665 1735 2727 2065
rect 2273 1687 2727 1735
rect 2744 1687 2747 2113
rect 2253 1681 2747 1687
rect 2803 2113 3297 2119
rect 2803 1687 2806 2113
rect 2823 2065 3277 2113
rect 2823 1735 2885 2065
rect 3215 1735 3277 2065
rect 2823 1687 3277 1735
rect 3294 1687 3297 2113
rect 2803 1681 3297 1687
rect 3353 2113 3847 2119
rect 3353 1687 3356 2113
rect 3373 2065 3827 2113
rect 3373 1735 3435 2065
rect 3765 1735 3827 2065
rect 3373 1687 3827 1735
rect 3844 1687 3847 2113
rect 3353 1681 3847 1687
rect 3903 2113 4397 2119
rect 3903 1687 3906 2113
rect 3923 2065 4377 2113
rect 3923 1735 3985 2065
rect 4315 1735 4377 2065
rect 3923 1687 4377 1735
rect 4394 1687 4397 2113
rect 3903 1681 4397 1687
rect 4453 2113 4947 2119
rect 4453 1687 4456 2113
rect 4473 2065 4927 2113
rect 4473 1735 4535 2065
rect 4865 1735 4927 2065
rect 4473 1687 4927 1735
rect 4944 1687 4947 2113
rect 4453 1681 4947 1687
rect 5003 2113 5497 2119
rect 5003 1687 5006 2113
rect 5023 2065 5477 2113
rect 5023 1735 5085 2065
rect 5415 1735 5477 2065
rect 5023 1687 5477 1735
rect 5494 1687 5497 2113
rect 5003 1681 5497 1687
rect 5553 2113 6047 2119
rect 5553 1687 5556 2113
rect 5573 2065 6027 2113
rect 5573 1735 5635 2065
rect 5965 1735 6027 2065
rect 5573 1687 6027 1735
rect 6044 1687 6047 2113
rect 5553 1681 6047 1687
rect 6103 2113 6597 2119
rect 6103 1687 6106 2113
rect 6123 2065 6577 2113
rect 6123 1735 6185 2065
rect 6515 1735 6577 2065
rect 6123 1687 6577 1735
rect 6594 1687 6597 2113
rect 6103 1681 6597 1687
rect 6653 2113 7147 2119
rect 6653 1687 6656 2113
rect 6673 2065 7127 2113
rect 6673 1735 6735 2065
rect 7065 1735 7127 2065
rect 6673 1687 7127 1735
rect 7144 1687 7147 2113
rect 6653 1681 7147 1687
rect 7203 2113 7697 2119
rect 7203 1687 7206 2113
rect 7223 2065 7677 2113
rect 7223 1735 7285 2065
rect 7615 1735 7677 2065
rect 7223 1687 7677 1735
rect 7694 1687 7697 2113
rect 7203 1681 7697 1687
rect 7753 2113 8247 2119
rect 7753 1687 7756 2113
rect 7773 2065 8227 2113
rect 7773 1735 7835 2065
rect 8165 1735 8227 2065
rect 7773 1687 8227 1735
rect 8244 1687 8247 2113
rect 7753 1681 8247 1687
rect 8303 2113 8797 2119
rect 8303 1687 8306 2113
rect 8323 2065 8777 2113
rect 8323 1735 8385 2065
rect 8715 1735 8777 2065
rect 8323 1687 8777 1735
rect 8794 1687 8797 2113
rect 8303 1681 8797 1687
rect 8853 2113 9347 2119
rect 8853 1687 8856 2113
rect 8873 2065 9327 2113
rect 8873 1735 8935 2065
rect 9265 1735 9327 2065
rect 8873 1687 9327 1735
rect 9344 1687 9347 2113
rect 8853 1681 9347 1687
rect 9403 2113 9897 2119
rect 9403 1687 9406 2113
rect 9423 2065 9877 2113
rect 9423 1735 9485 2065
rect 9815 1735 9877 2065
rect 9423 1687 9877 1735
rect 9894 1687 9897 2113
rect 9403 1681 9897 1687
rect 9953 2113 10447 2119
rect 9953 1687 9956 2113
rect 9973 2065 10427 2113
rect 9973 1735 10035 2065
rect 10365 1735 10427 2065
rect 9973 1687 10427 1735
rect 10444 1687 10447 2113
rect 9953 1681 10447 1687
rect 10503 2113 10997 2119
rect 10503 1687 10506 2113
rect 10523 2065 10977 2113
rect 10523 1735 10585 2065
rect 10915 1735 10977 2065
rect 10523 1687 10977 1735
rect 10994 1687 10997 2113
rect 10503 1681 10997 1687
rect 11053 2113 11547 2119
rect 11053 1687 11056 2113
rect 11073 2065 11527 2113
rect 11073 1735 11135 2065
rect 11465 1735 11527 2065
rect 11073 1687 11527 1735
rect 11544 1687 11547 2113
rect 11053 1681 11547 1687
rect 11603 2113 12097 2119
rect 11603 1687 11606 2113
rect 11623 2065 12077 2113
rect 11623 1735 11685 2065
rect 12015 1735 12077 2065
rect 11623 1687 12077 1735
rect 12094 1687 12097 2113
rect 11603 1681 12097 1687
rect 12153 2113 12647 2119
rect 12153 1687 12156 2113
rect 12173 2065 12627 2113
rect 12173 1735 12235 2065
rect 12565 1735 12627 2065
rect 12173 1687 12627 1735
rect 12644 1687 12647 2113
rect 12153 1681 12647 1687
rect 12703 2113 13197 2119
rect 12703 1687 12706 2113
rect 12723 2065 13177 2113
rect 12723 1735 12785 2065
rect 13115 1735 13177 2065
rect 12723 1687 13177 1735
rect 13194 1687 13197 2113
rect 12703 1681 13197 1687
rect 13253 2113 13724 2119
rect 13253 1687 13256 2113
rect 13273 2065 13724 2113
rect 13273 1735 13335 2065
rect 13665 1735 13724 2065
rect 13273 1687 13724 1735
rect 13253 1681 13724 1687
rect -474 1676 -26 1681
rect 76 1676 524 1681
rect 626 1676 1074 1681
rect 1176 1676 1624 1681
rect 1726 1676 2174 1681
rect 2276 1676 2724 1681
rect 2826 1676 3274 1681
rect 3376 1676 3824 1681
rect 3926 1676 4374 1681
rect 4476 1676 4924 1681
rect 5026 1676 5474 1681
rect 5576 1676 6024 1681
rect 6126 1676 6574 1681
rect 6676 1676 7124 1681
rect 7226 1676 7674 1681
rect 7776 1676 8224 1681
rect 8326 1676 8774 1681
rect 8876 1676 9324 1681
rect 9426 1676 9874 1681
rect 9976 1676 10424 1681
rect 10526 1676 10974 1681
rect 11076 1676 11524 1681
rect 11626 1676 12074 1681
rect 12176 1676 12624 1681
rect 12726 1676 13174 1681
rect 13276 1676 13724 1681
rect -1025 1650 -725 1669
rect -469 1673 -31 1676
rect -469 1656 -463 1673
rect -37 1656 -31 1673
rect -469 1653 -31 1656
rect 81 1673 519 1676
rect 81 1656 87 1673
rect 513 1656 519 1673
rect 81 1653 519 1656
rect 631 1673 1069 1676
rect 631 1656 637 1673
rect 1063 1656 1069 1673
rect 631 1653 1069 1656
rect 1181 1673 1619 1676
rect 1181 1656 1187 1673
rect 1613 1656 1619 1673
rect 1181 1653 1619 1656
rect 1731 1673 2169 1676
rect 1731 1656 1737 1673
rect 2163 1656 2169 1673
rect 1731 1653 2169 1656
rect 2281 1673 2719 1676
rect 2281 1656 2287 1673
rect 2713 1656 2719 1673
rect 2281 1653 2719 1656
rect 2831 1673 3269 1676
rect 2831 1656 2837 1673
rect 3263 1656 3269 1673
rect 2831 1653 3269 1656
rect 3381 1673 3819 1676
rect 3381 1656 3387 1673
rect 3813 1656 3819 1673
rect 3381 1653 3819 1656
rect 3931 1673 4369 1676
rect 3931 1656 3937 1673
rect 4363 1656 4369 1673
rect 3931 1653 4369 1656
rect 4481 1673 4919 1676
rect 4481 1656 4487 1673
rect 4913 1656 4919 1673
rect 4481 1653 4919 1656
rect 5031 1673 5469 1676
rect 5031 1656 5037 1673
rect 5463 1656 5469 1673
rect 5031 1653 5469 1656
rect 5581 1673 6019 1676
rect 5581 1656 5587 1673
rect 6013 1656 6019 1673
rect 5581 1653 6019 1656
rect 6131 1673 6569 1676
rect 6131 1656 6137 1673
rect 6563 1656 6569 1673
rect 6131 1653 6569 1656
rect 6681 1673 7119 1676
rect 6681 1656 6687 1673
rect 7113 1656 7119 1673
rect 6681 1653 7119 1656
rect 7231 1673 7669 1676
rect 7231 1656 7237 1673
rect 7663 1656 7669 1673
rect 7231 1653 7669 1656
rect 7781 1673 8219 1676
rect 7781 1656 7787 1673
rect 8213 1656 8219 1673
rect 7781 1653 8219 1656
rect 8331 1673 8769 1676
rect 8331 1656 8337 1673
rect 8763 1656 8769 1673
rect 8331 1653 8769 1656
rect 8881 1673 9319 1676
rect 8881 1656 8887 1673
rect 9313 1656 9319 1673
rect 8881 1653 9319 1656
rect 9431 1673 9869 1676
rect 9431 1656 9437 1673
rect 9863 1656 9869 1673
rect 9431 1653 9869 1656
rect 9981 1673 10419 1676
rect 9981 1656 9987 1673
rect 10413 1656 10419 1673
rect 9981 1653 10419 1656
rect 10531 1673 10969 1676
rect 10531 1656 10537 1673
rect 10963 1656 10969 1673
rect 10531 1653 10969 1656
rect 11081 1673 11519 1676
rect 11081 1656 11087 1673
rect 11513 1656 11519 1673
rect 11081 1653 11519 1656
rect 11631 1673 12069 1676
rect 11631 1656 11637 1673
rect 12063 1656 12069 1673
rect 11631 1653 12069 1656
rect 12181 1673 12619 1676
rect 12181 1656 12187 1673
rect 12613 1656 12619 1673
rect 12181 1653 12619 1656
rect 12731 1673 13169 1676
rect 12731 1656 12737 1673
rect 13163 1656 13169 1673
rect 12731 1653 13169 1656
rect 13281 1673 13719 1676
rect 13281 1656 13287 1673
rect 13713 1656 13719 1673
rect 13281 1653 13719 1656
rect 13975 1669 13987 2200
rect 14263 1669 14275 2200
rect 13975 1650 14275 1669
rect -1025 1119 -1013 1650
rect -737 1119 -725 1650
rect -550 1642 -500 1650
rect -550 1608 -542 1642
rect -508 1608 -500 1642
rect -550 1600 -500 1608
rect 0 1642 50 1650
rect 0 1608 8 1642
rect 42 1608 50 1642
rect 0 1600 50 1608
rect 550 1642 600 1650
rect 550 1608 558 1642
rect 592 1608 600 1642
rect 550 1600 600 1608
rect 1100 1642 1150 1650
rect 1100 1608 1108 1642
rect 1142 1608 1150 1642
rect 1100 1600 1150 1608
rect 1650 1642 1700 1650
rect 1650 1608 1658 1642
rect 1692 1608 1700 1642
rect 1650 1600 1700 1608
rect 2200 1642 2250 1650
rect 2200 1608 2208 1642
rect 2242 1608 2250 1642
rect 2200 1600 2250 1608
rect 2750 1642 2800 1650
rect 2750 1608 2758 1642
rect 2792 1608 2800 1642
rect 2750 1600 2800 1608
rect 3300 1642 3350 1650
rect 3300 1608 3308 1642
rect 3342 1608 3350 1642
rect 3300 1600 3350 1608
rect 3850 1642 3900 1650
rect 3850 1608 3858 1642
rect 3892 1608 3900 1642
rect 3850 1600 3900 1608
rect 4400 1642 4450 1650
rect 4400 1608 4408 1642
rect 4442 1608 4450 1642
rect 4400 1600 4450 1608
rect 4950 1642 5000 1650
rect 4950 1608 4958 1642
rect 4992 1608 5000 1642
rect 4950 1600 5000 1608
rect 5500 1642 5550 1650
rect 5500 1608 5508 1642
rect 5542 1608 5550 1642
rect 5500 1600 5550 1608
rect 6050 1642 6100 1650
rect 6050 1608 6058 1642
rect 6092 1608 6100 1642
rect 6050 1600 6100 1608
rect 6600 1642 6650 1650
rect 6600 1608 6608 1642
rect 6642 1608 6650 1642
rect 6600 1600 6650 1608
rect 7150 1642 7200 1650
rect 7150 1608 7158 1642
rect 7192 1608 7200 1642
rect 7150 1600 7200 1608
rect 7700 1642 7750 1650
rect 7700 1608 7708 1642
rect 7742 1608 7750 1642
rect 7700 1600 7750 1608
rect 8250 1642 8300 1650
rect 8250 1608 8258 1642
rect 8292 1608 8300 1642
rect 8250 1600 8300 1608
rect 8800 1642 8850 1650
rect 8800 1608 8808 1642
rect 8842 1608 8850 1642
rect 8800 1600 8850 1608
rect 9350 1642 9400 1650
rect 9350 1608 9358 1642
rect 9392 1608 9400 1642
rect 9350 1600 9400 1608
rect 9900 1642 9950 1650
rect 9900 1608 9908 1642
rect 9942 1608 9950 1642
rect 9900 1600 9950 1608
rect 10450 1642 10500 1650
rect 10450 1608 10458 1642
rect 10492 1608 10500 1642
rect 10450 1600 10500 1608
rect 11000 1642 11050 1650
rect 11000 1608 11008 1642
rect 11042 1608 11050 1642
rect 11000 1600 11050 1608
rect 11550 1642 11600 1650
rect 11550 1608 11558 1642
rect 11592 1608 11600 1642
rect 11550 1600 11600 1608
rect 12100 1642 12150 1650
rect 12100 1608 12108 1642
rect 12142 1608 12150 1642
rect 12100 1600 12150 1608
rect 12650 1642 12700 1650
rect 12650 1608 12658 1642
rect 12692 1608 12700 1642
rect 12650 1600 12700 1608
rect 13200 1642 13250 1650
rect 13200 1608 13208 1642
rect 13242 1608 13250 1642
rect 13200 1600 13250 1608
rect 13750 1642 13800 1650
rect 13750 1608 13758 1642
rect 13792 1608 13800 1642
rect 13750 1600 13800 1608
rect -469 1594 -31 1597
rect -469 1577 -463 1594
rect -37 1577 -31 1594
rect -469 1574 -31 1577
rect 81 1594 519 1597
rect 81 1577 87 1594
rect 513 1577 519 1594
rect 81 1574 519 1577
rect 631 1594 1069 1597
rect 631 1577 637 1594
rect 1063 1577 1069 1594
rect 631 1574 1069 1577
rect 1181 1594 1619 1597
rect 1181 1577 1187 1594
rect 1613 1577 1619 1594
rect 1181 1574 1619 1577
rect 1731 1594 2169 1597
rect 1731 1577 1737 1594
rect 2163 1577 2169 1594
rect 1731 1574 2169 1577
rect 2281 1594 2719 1597
rect 2281 1577 2287 1594
rect 2713 1577 2719 1594
rect 2281 1574 2719 1577
rect 2831 1594 3269 1597
rect 2831 1577 2837 1594
rect 3263 1577 3269 1594
rect 2831 1574 3269 1577
rect 3381 1594 3819 1597
rect 3381 1577 3387 1594
rect 3813 1577 3819 1594
rect 3381 1574 3819 1577
rect 3931 1594 4369 1597
rect 3931 1577 3937 1594
rect 4363 1577 4369 1594
rect 3931 1574 4369 1577
rect 4481 1594 4919 1597
rect 4481 1577 4487 1594
rect 4913 1577 4919 1594
rect 4481 1574 4919 1577
rect 5031 1594 5469 1597
rect 5031 1577 5037 1594
rect 5463 1577 5469 1594
rect 5031 1574 5469 1577
rect 5581 1594 6019 1597
rect 5581 1577 5587 1594
rect 6013 1577 6019 1594
rect 5581 1574 6019 1577
rect 6131 1594 6569 1597
rect 6131 1577 6137 1594
rect 6563 1577 6569 1594
rect 6131 1574 6569 1577
rect 6681 1594 7119 1597
rect 6681 1577 6687 1594
rect 7113 1577 7119 1594
rect 6681 1574 7119 1577
rect 7231 1594 7669 1597
rect 7231 1577 7237 1594
rect 7663 1577 7669 1594
rect 7231 1574 7669 1577
rect 7781 1594 8219 1597
rect 7781 1577 7787 1594
rect 8213 1577 8219 1594
rect 7781 1574 8219 1577
rect 8331 1594 8769 1597
rect 8331 1577 8337 1594
rect 8763 1577 8769 1594
rect 8331 1574 8769 1577
rect 8881 1594 9319 1597
rect 8881 1577 8887 1594
rect 9313 1577 9319 1594
rect 8881 1574 9319 1577
rect 9431 1594 9869 1597
rect 9431 1577 9437 1594
rect 9863 1577 9869 1594
rect 9431 1574 9869 1577
rect 9981 1594 10419 1597
rect 9981 1577 9987 1594
rect 10413 1577 10419 1594
rect 9981 1574 10419 1577
rect 10531 1594 10969 1597
rect 10531 1577 10537 1594
rect 10963 1577 10969 1594
rect 10531 1574 10969 1577
rect 11081 1594 11519 1597
rect 11081 1577 11087 1594
rect 11513 1577 11519 1594
rect 11081 1574 11519 1577
rect 11631 1594 12069 1597
rect 11631 1577 11637 1594
rect 12063 1577 12069 1594
rect 11631 1574 12069 1577
rect 12181 1594 12619 1597
rect 12181 1577 12187 1594
rect 12613 1577 12619 1594
rect 12181 1574 12619 1577
rect 12731 1594 13169 1597
rect 12731 1577 12737 1594
rect 13163 1577 13169 1594
rect 12731 1574 13169 1577
rect 13281 1594 13719 1597
rect 13281 1577 13287 1594
rect 13713 1577 13719 1594
rect 13281 1574 13719 1577
rect -474 1569 -26 1574
rect 76 1569 524 1574
rect 626 1569 1074 1574
rect 1176 1569 1624 1574
rect 1726 1569 2174 1574
rect 2276 1569 2724 1574
rect 2826 1569 3274 1574
rect 3376 1569 3824 1574
rect 3926 1569 4374 1574
rect 4476 1569 4924 1574
rect 5026 1569 5474 1574
rect 5576 1569 6024 1574
rect 6126 1569 6574 1574
rect 6676 1569 7124 1574
rect 7226 1569 7674 1574
rect 7776 1569 8224 1574
rect 8326 1569 8774 1574
rect 8876 1569 9324 1574
rect 9426 1569 9874 1574
rect 9976 1569 10424 1574
rect 10526 1569 10974 1574
rect 11076 1569 11524 1574
rect 11626 1569 12074 1574
rect 12176 1569 12624 1574
rect 12726 1569 13174 1574
rect 13276 1569 13724 1574
rect -474 1563 -3 1569
rect -474 1515 -23 1563
rect -474 1185 -415 1515
rect -85 1185 -23 1515
rect -474 1137 -23 1185
rect -6 1137 -3 1563
rect -474 1131 -3 1137
rect 53 1563 547 1569
rect 53 1137 56 1563
rect 73 1515 527 1563
rect 73 1185 135 1515
rect 465 1185 527 1515
rect 73 1137 527 1185
rect 544 1137 547 1563
rect 53 1131 547 1137
rect 603 1563 1097 1569
rect 603 1137 606 1563
rect 623 1515 1077 1563
rect 623 1185 685 1515
rect 1015 1185 1077 1515
rect 623 1137 1077 1185
rect 1094 1137 1097 1563
rect 603 1131 1097 1137
rect 1153 1563 1647 1569
rect 1153 1137 1156 1563
rect 1173 1515 1627 1563
rect 1173 1185 1235 1515
rect 1565 1185 1627 1515
rect 1173 1137 1627 1185
rect 1644 1137 1647 1563
rect 1153 1131 1647 1137
rect 1703 1563 2197 1569
rect 1703 1137 1706 1563
rect 1723 1515 2177 1563
rect 1723 1185 1785 1515
rect 2115 1185 2177 1515
rect 1723 1137 2177 1185
rect 2194 1137 2197 1563
rect 1703 1131 2197 1137
rect 2253 1563 2747 1569
rect 2253 1137 2256 1563
rect 2273 1515 2727 1563
rect 2273 1185 2335 1515
rect 2665 1185 2727 1515
rect 2273 1137 2727 1185
rect 2744 1137 2747 1563
rect 2253 1131 2747 1137
rect 2803 1563 3297 1569
rect 2803 1137 2806 1563
rect 2823 1515 3277 1563
rect 2823 1185 2885 1515
rect 3215 1185 3277 1515
rect 2823 1137 3277 1185
rect 3294 1137 3297 1563
rect 2803 1131 3297 1137
rect 3353 1563 3847 1569
rect 3353 1137 3356 1563
rect 3373 1515 3827 1563
rect 3373 1185 3435 1515
rect 3765 1185 3827 1515
rect 3373 1137 3827 1185
rect 3844 1137 3847 1563
rect 3353 1131 3847 1137
rect 3903 1563 4397 1569
rect 3903 1137 3906 1563
rect 3923 1515 4377 1563
rect 3923 1185 3985 1515
rect 4315 1185 4377 1515
rect 3923 1137 4377 1185
rect 4394 1137 4397 1563
rect 3903 1131 4397 1137
rect 4453 1563 4947 1569
rect 4453 1137 4456 1563
rect 4473 1515 4927 1563
rect 4473 1185 4535 1515
rect 4865 1185 4927 1515
rect 4473 1137 4927 1185
rect 4944 1137 4947 1563
rect 4453 1131 4947 1137
rect 5003 1563 5497 1569
rect 5003 1137 5006 1563
rect 5023 1515 5477 1563
rect 5023 1185 5085 1515
rect 5415 1185 5477 1515
rect 5023 1137 5477 1185
rect 5494 1137 5497 1563
rect 5003 1131 5497 1137
rect 5553 1563 6047 1569
rect 5553 1137 5556 1563
rect 5573 1515 6027 1563
rect 5573 1185 5635 1515
rect 5965 1185 6027 1515
rect 5573 1137 6027 1185
rect 6044 1137 6047 1563
rect 5553 1131 6047 1137
rect 6103 1563 6597 1569
rect 6103 1137 6106 1563
rect 6123 1515 6577 1563
rect 6123 1185 6185 1515
rect 6515 1185 6577 1515
rect 6123 1137 6577 1185
rect 6594 1137 6597 1563
rect 6103 1131 6597 1137
rect 6653 1563 7147 1569
rect 6653 1137 6656 1563
rect 6673 1515 7127 1563
rect 6673 1185 6735 1515
rect 7065 1185 7127 1515
rect 6673 1137 7127 1185
rect 7144 1137 7147 1563
rect 6653 1131 7147 1137
rect 7203 1563 7697 1569
rect 7203 1137 7206 1563
rect 7223 1515 7677 1563
rect 7223 1185 7285 1515
rect 7615 1185 7677 1515
rect 7223 1137 7677 1185
rect 7694 1137 7697 1563
rect 7203 1131 7697 1137
rect 7753 1563 8247 1569
rect 7753 1137 7756 1563
rect 7773 1515 8227 1563
rect 7773 1185 7835 1515
rect 8165 1185 8227 1515
rect 7773 1137 8227 1185
rect 8244 1137 8247 1563
rect 7753 1131 8247 1137
rect 8303 1563 8797 1569
rect 8303 1137 8306 1563
rect 8323 1515 8777 1563
rect 8323 1185 8385 1515
rect 8715 1185 8777 1515
rect 8323 1137 8777 1185
rect 8794 1137 8797 1563
rect 8303 1131 8797 1137
rect 8853 1563 9347 1569
rect 8853 1137 8856 1563
rect 8873 1515 9327 1563
rect 8873 1185 8935 1515
rect 9265 1185 9327 1515
rect 8873 1137 9327 1185
rect 9344 1137 9347 1563
rect 8853 1131 9347 1137
rect 9403 1563 9897 1569
rect 9403 1137 9406 1563
rect 9423 1515 9877 1563
rect 9423 1185 9485 1515
rect 9815 1185 9877 1515
rect 9423 1137 9877 1185
rect 9894 1137 9897 1563
rect 9403 1131 9897 1137
rect 9953 1563 10447 1569
rect 9953 1137 9956 1563
rect 9973 1515 10427 1563
rect 9973 1185 10035 1515
rect 10365 1185 10427 1515
rect 9973 1137 10427 1185
rect 10444 1137 10447 1563
rect 9953 1131 10447 1137
rect 10503 1563 10997 1569
rect 10503 1137 10506 1563
rect 10523 1515 10977 1563
rect 10523 1185 10585 1515
rect 10915 1185 10977 1515
rect 10523 1137 10977 1185
rect 10994 1137 10997 1563
rect 10503 1131 10997 1137
rect 11053 1563 11547 1569
rect 11053 1137 11056 1563
rect 11073 1515 11527 1563
rect 11073 1185 11135 1515
rect 11465 1185 11527 1515
rect 11073 1137 11527 1185
rect 11544 1137 11547 1563
rect 11053 1131 11547 1137
rect 11603 1563 12097 1569
rect 11603 1137 11606 1563
rect 11623 1515 12077 1563
rect 11623 1185 11685 1515
rect 12015 1185 12077 1515
rect 11623 1137 12077 1185
rect 12094 1137 12097 1563
rect 11603 1131 12097 1137
rect 12153 1563 12647 1569
rect 12153 1137 12156 1563
rect 12173 1515 12627 1563
rect 12173 1185 12235 1515
rect 12565 1185 12627 1515
rect 12173 1137 12627 1185
rect 12644 1137 12647 1563
rect 12153 1131 12647 1137
rect 12703 1563 13197 1569
rect 12703 1137 12706 1563
rect 12723 1515 13177 1563
rect 12723 1185 12785 1515
rect 13115 1185 13177 1515
rect 12723 1137 13177 1185
rect 13194 1137 13197 1563
rect 12703 1131 13197 1137
rect 13253 1563 13724 1569
rect 13253 1137 13256 1563
rect 13273 1515 13724 1563
rect 13273 1185 13335 1515
rect 13665 1185 13724 1515
rect 13273 1137 13724 1185
rect 13253 1131 13724 1137
rect -474 1126 -26 1131
rect 76 1126 524 1131
rect 626 1126 1074 1131
rect 1176 1126 1624 1131
rect 1726 1126 2174 1131
rect 2276 1126 2724 1131
rect 2826 1126 3274 1131
rect 3376 1126 3824 1131
rect 3926 1126 4374 1131
rect 4476 1126 4924 1131
rect 5026 1126 5474 1131
rect 5576 1126 6024 1131
rect 6126 1126 6574 1131
rect 6676 1126 7124 1131
rect 7226 1126 7674 1131
rect 7776 1126 8224 1131
rect 8326 1126 8774 1131
rect 8876 1126 9324 1131
rect 9426 1126 9874 1131
rect 9976 1126 10424 1131
rect 10526 1126 10974 1131
rect 11076 1126 11524 1131
rect 11626 1126 12074 1131
rect 12176 1126 12624 1131
rect 12726 1126 13174 1131
rect 13276 1126 13724 1131
rect -1025 1100 -725 1119
rect -469 1123 -31 1126
rect -469 1106 -463 1123
rect -37 1106 -31 1123
rect -469 1103 -31 1106
rect 81 1123 519 1126
rect 81 1106 87 1123
rect 513 1106 519 1123
rect 81 1103 519 1106
rect 631 1123 1069 1126
rect 631 1106 637 1123
rect 1063 1106 1069 1123
rect 631 1103 1069 1106
rect 1181 1123 1619 1126
rect 1181 1106 1187 1123
rect 1613 1106 1619 1123
rect 1181 1103 1619 1106
rect 1731 1123 2169 1126
rect 1731 1106 1737 1123
rect 2163 1106 2169 1123
rect 1731 1103 2169 1106
rect 2281 1123 2719 1126
rect 2281 1106 2287 1123
rect 2713 1106 2719 1123
rect 2281 1103 2719 1106
rect 2831 1123 3269 1126
rect 2831 1106 2837 1123
rect 3263 1106 3269 1123
rect 2831 1103 3269 1106
rect 3381 1123 3819 1126
rect 3381 1106 3387 1123
rect 3813 1106 3819 1123
rect 3381 1103 3819 1106
rect 3931 1123 4369 1126
rect 3931 1106 3937 1123
rect 4363 1106 4369 1123
rect 3931 1103 4369 1106
rect 4481 1123 4919 1126
rect 4481 1106 4487 1123
rect 4913 1106 4919 1123
rect 4481 1103 4919 1106
rect 5031 1123 5469 1126
rect 5031 1106 5037 1123
rect 5463 1106 5469 1123
rect 5031 1103 5469 1106
rect 5581 1123 6019 1126
rect 5581 1106 5587 1123
rect 6013 1106 6019 1123
rect 5581 1103 6019 1106
rect 6131 1123 6569 1126
rect 6131 1106 6137 1123
rect 6563 1106 6569 1123
rect 6131 1103 6569 1106
rect 6681 1123 7119 1126
rect 6681 1106 6687 1123
rect 7113 1106 7119 1123
rect 6681 1103 7119 1106
rect 7231 1123 7669 1126
rect 7231 1106 7237 1123
rect 7663 1106 7669 1123
rect 7231 1103 7669 1106
rect 7781 1123 8219 1126
rect 7781 1106 7787 1123
rect 8213 1106 8219 1123
rect 7781 1103 8219 1106
rect 8331 1123 8769 1126
rect 8331 1106 8337 1123
rect 8763 1106 8769 1123
rect 8331 1103 8769 1106
rect 8881 1123 9319 1126
rect 8881 1106 8887 1123
rect 9313 1106 9319 1123
rect 8881 1103 9319 1106
rect 9431 1123 9869 1126
rect 9431 1106 9437 1123
rect 9863 1106 9869 1123
rect 9431 1103 9869 1106
rect 9981 1123 10419 1126
rect 9981 1106 9987 1123
rect 10413 1106 10419 1123
rect 9981 1103 10419 1106
rect 10531 1123 10969 1126
rect 10531 1106 10537 1123
rect 10963 1106 10969 1123
rect 10531 1103 10969 1106
rect 11081 1123 11519 1126
rect 11081 1106 11087 1123
rect 11513 1106 11519 1123
rect 11081 1103 11519 1106
rect 11631 1123 12069 1126
rect 11631 1106 11637 1123
rect 12063 1106 12069 1123
rect 11631 1103 12069 1106
rect 12181 1123 12619 1126
rect 12181 1106 12187 1123
rect 12613 1106 12619 1123
rect 12181 1103 12619 1106
rect 12731 1123 13169 1126
rect 12731 1106 12737 1123
rect 13163 1106 13169 1123
rect 12731 1103 13169 1106
rect 13281 1123 13719 1126
rect 13281 1106 13287 1123
rect 13713 1106 13719 1123
rect 13281 1103 13719 1106
rect 13975 1119 13987 1650
rect 14263 1119 14275 1650
rect 13975 1100 14275 1119
rect -1025 569 -1013 1100
rect -737 569 -725 1100
rect -550 1092 -500 1100
rect -550 1058 -542 1092
rect -508 1058 -500 1092
rect -550 1050 -500 1058
rect 0 1092 50 1100
rect 0 1058 8 1092
rect 42 1058 50 1092
rect 0 1050 50 1058
rect 550 1092 600 1100
rect 550 1058 558 1092
rect 592 1058 600 1092
rect 550 1050 600 1058
rect 1100 1092 1150 1100
rect 1100 1058 1108 1092
rect 1142 1058 1150 1092
rect 1100 1050 1150 1058
rect 1650 1092 1700 1100
rect 1650 1058 1658 1092
rect 1692 1058 1700 1092
rect 1650 1050 1700 1058
rect 2200 1092 2250 1100
rect 2200 1058 2208 1092
rect 2242 1058 2250 1092
rect 2200 1050 2250 1058
rect 2750 1092 2800 1100
rect 2750 1058 2758 1092
rect 2792 1058 2800 1092
rect 2750 1050 2800 1058
rect 3300 1092 3350 1100
rect 3300 1058 3308 1092
rect 3342 1058 3350 1092
rect 3300 1050 3350 1058
rect 3850 1092 3900 1100
rect 3850 1058 3858 1092
rect 3892 1058 3900 1092
rect 3850 1050 3900 1058
rect 4400 1092 4450 1100
rect 4400 1058 4408 1092
rect 4442 1058 4450 1092
rect 4400 1050 4450 1058
rect 4950 1092 5000 1100
rect 4950 1058 4958 1092
rect 4992 1058 5000 1092
rect 4950 1050 5000 1058
rect 5500 1092 5550 1100
rect 5500 1058 5508 1092
rect 5542 1058 5550 1092
rect 5500 1050 5550 1058
rect 6050 1092 6100 1100
rect 6050 1058 6058 1092
rect 6092 1058 6100 1092
rect 6050 1050 6100 1058
rect 6600 1092 6650 1100
rect 6600 1058 6608 1092
rect 6642 1058 6650 1092
rect 6600 1050 6650 1058
rect 7150 1092 7200 1100
rect 7150 1058 7158 1092
rect 7192 1058 7200 1092
rect 7150 1050 7200 1058
rect 7700 1092 7750 1100
rect 7700 1058 7708 1092
rect 7742 1058 7750 1092
rect 7700 1050 7750 1058
rect 8250 1092 8300 1100
rect 8250 1058 8258 1092
rect 8292 1058 8300 1092
rect 8250 1050 8300 1058
rect 8800 1092 8850 1100
rect 8800 1058 8808 1092
rect 8842 1058 8850 1092
rect 8800 1050 8850 1058
rect 9350 1092 9400 1100
rect 9350 1058 9358 1092
rect 9392 1058 9400 1092
rect 9350 1050 9400 1058
rect 9900 1092 9950 1100
rect 9900 1058 9908 1092
rect 9942 1058 9950 1092
rect 9900 1050 9950 1058
rect 10450 1092 10500 1100
rect 10450 1058 10458 1092
rect 10492 1058 10500 1092
rect 10450 1050 10500 1058
rect 11000 1092 11050 1100
rect 11000 1058 11008 1092
rect 11042 1058 11050 1092
rect 11000 1050 11050 1058
rect 11550 1092 11600 1100
rect 11550 1058 11558 1092
rect 11592 1058 11600 1092
rect 11550 1050 11600 1058
rect 12100 1092 12150 1100
rect 12100 1058 12108 1092
rect 12142 1058 12150 1092
rect 12100 1050 12150 1058
rect 12650 1092 12700 1100
rect 12650 1058 12658 1092
rect 12692 1058 12700 1092
rect 12650 1050 12700 1058
rect 13200 1092 13250 1100
rect 13200 1058 13208 1092
rect 13242 1058 13250 1092
rect 13200 1050 13250 1058
rect 13750 1092 13800 1100
rect 13750 1058 13758 1092
rect 13792 1058 13800 1092
rect 13750 1050 13800 1058
rect -469 1044 -31 1047
rect -469 1027 -463 1044
rect -37 1027 -31 1044
rect -469 1024 -31 1027
rect 81 1044 519 1047
rect 81 1027 87 1044
rect 513 1027 519 1044
rect 81 1024 519 1027
rect 631 1044 1069 1047
rect 631 1027 637 1044
rect 1063 1027 1069 1044
rect 631 1024 1069 1027
rect 1181 1044 1619 1047
rect 1181 1027 1187 1044
rect 1613 1027 1619 1044
rect 1181 1024 1619 1027
rect 1731 1044 2169 1047
rect 1731 1027 1737 1044
rect 2163 1027 2169 1044
rect 1731 1024 2169 1027
rect 2281 1044 2719 1047
rect 2281 1027 2287 1044
rect 2713 1027 2719 1044
rect 2281 1024 2719 1027
rect 2831 1044 3269 1047
rect 2831 1027 2837 1044
rect 3263 1027 3269 1044
rect 2831 1024 3269 1027
rect 3381 1044 3819 1047
rect 3381 1027 3387 1044
rect 3813 1027 3819 1044
rect 3381 1024 3819 1027
rect 3931 1044 4369 1047
rect 3931 1027 3937 1044
rect 4363 1027 4369 1044
rect 3931 1024 4369 1027
rect 4481 1044 4919 1047
rect 4481 1027 4487 1044
rect 4913 1027 4919 1044
rect 4481 1024 4919 1027
rect 5031 1044 5469 1047
rect 5031 1027 5037 1044
rect 5463 1027 5469 1044
rect 5031 1024 5469 1027
rect 5581 1044 6019 1047
rect 5581 1027 5587 1044
rect 6013 1027 6019 1044
rect 5581 1024 6019 1027
rect 6131 1044 6569 1047
rect 6131 1027 6137 1044
rect 6563 1027 6569 1044
rect 6131 1024 6569 1027
rect 6681 1044 7119 1047
rect 6681 1027 6687 1044
rect 7113 1027 7119 1044
rect 6681 1024 7119 1027
rect 7231 1044 7669 1047
rect 7231 1027 7237 1044
rect 7663 1027 7669 1044
rect 7231 1024 7669 1027
rect 7781 1044 8219 1047
rect 7781 1027 7787 1044
rect 8213 1027 8219 1044
rect 7781 1024 8219 1027
rect 8331 1044 8769 1047
rect 8331 1027 8337 1044
rect 8763 1027 8769 1044
rect 8331 1024 8769 1027
rect 8881 1044 9319 1047
rect 8881 1027 8887 1044
rect 9313 1027 9319 1044
rect 8881 1024 9319 1027
rect 9431 1044 9869 1047
rect 9431 1027 9437 1044
rect 9863 1027 9869 1044
rect 9431 1024 9869 1027
rect 9981 1044 10419 1047
rect 9981 1027 9987 1044
rect 10413 1027 10419 1044
rect 9981 1024 10419 1027
rect 10531 1044 10969 1047
rect 10531 1027 10537 1044
rect 10963 1027 10969 1044
rect 10531 1024 10969 1027
rect 11081 1044 11519 1047
rect 11081 1027 11087 1044
rect 11513 1027 11519 1044
rect 11081 1024 11519 1027
rect 11631 1044 12069 1047
rect 11631 1027 11637 1044
rect 12063 1027 12069 1044
rect 11631 1024 12069 1027
rect 12181 1044 12619 1047
rect 12181 1027 12187 1044
rect 12613 1027 12619 1044
rect 12181 1024 12619 1027
rect 12731 1044 13169 1047
rect 12731 1027 12737 1044
rect 13163 1027 13169 1044
rect 12731 1024 13169 1027
rect 13281 1044 13719 1047
rect 13281 1027 13287 1044
rect 13713 1027 13719 1044
rect 13281 1024 13719 1027
rect -474 1019 -26 1024
rect 76 1019 524 1024
rect 626 1019 1074 1024
rect 1176 1019 1624 1024
rect 1726 1019 2174 1024
rect 2276 1019 2724 1024
rect 2826 1019 3274 1024
rect 3376 1019 3824 1024
rect 3926 1019 4374 1024
rect 4476 1019 4924 1024
rect 5026 1019 5474 1024
rect 5576 1019 6024 1024
rect 6126 1019 6574 1024
rect 6676 1019 7124 1024
rect 7226 1019 7674 1024
rect 7776 1019 8224 1024
rect 8326 1019 8774 1024
rect 8876 1019 9324 1024
rect 9426 1019 9874 1024
rect 9976 1019 10424 1024
rect 10526 1019 10974 1024
rect 11076 1019 11524 1024
rect 11626 1019 12074 1024
rect 12176 1019 12624 1024
rect 12726 1019 13174 1024
rect 13276 1019 13724 1024
rect -474 1013 -3 1019
rect -474 965 -23 1013
rect -474 635 -415 965
rect -85 635 -23 965
rect -474 587 -23 635
rect -6 587 -3 1013
rect -474 581 -3 587
rect 53 1013 547 1019
rect 53 587 56 1013
rect 73 965 527 1013
rect 73 635 135 965
rect 465 635 527 965
rect 73 587 527 635
rect 544 587 547 1013
rect 53 581 547 587
rect 603 1013 1097 1019
rect 603 587 606 1013
rect 623 965 1077 1013
rect 623 635 685 965
rect 1015 635 1077 965
rect 623 587 1077 635
rect 1094 587 1097 1013
rect 603 581 1097 587
rect 1153 1013 1647 1019
rect 1153 587 1156 1013
rect 1173 965 1627 1013
rect 1173 635 1235 965
rect 1565 635 1627 965
rect 1173 587 1627 635
rect 1644 587 1647 1013
rect 1153 581 1647 587
rect 1703 1013 2197 1019
rect 1703 587 1706 1013
rect 1723 965 2177 1013
rect 1723 635 1785 965
rect 2115 635 2177 965
rect 1723 587 2177 635
rect 2194 587 2197 1013
rect 1703 581 2197 587
rect 2253 1013 2747 1019
rect 2253 587 2256 1013
rect 2273 965 2727 1013
rect 2273 635 2335 965
rect 2665 635 2727 965
rect 2273 587 2727 635
rect 2744 587 2747 1013
rect 2253 581 2747 587
rect 2803 1013 3297 1019
rect 2803 587 2806 1013
rect 2823 965 3277 1013
rect 2823 635 2885 965
rect 3215 635 3277 965
rect 2823 587 3277 635
rect 3294 587 3297 1013
rect 2803 581 3297 587
rect 3353 1013 3847 1019
rect 3353 587 3356 1013
rect 3373 965 3827 1013
rect 3373 635 3435 965
rect 3765 635 3827 965
rect 3373 587 3827 635
rect 3844 587 3847 1013
rect 3353 581 3847 587
rect 3903 1013 4397 1019
rect 3903 587 3906 1013
rect 3923 965 4377 1013
rect 3923 635 3985 965
rect 4315 635 4377 965
rect 3923 587 4377 635
rect 4394 587 4397 1013
rect 3903 581 4397 587
rect 4453 1013 4947 1019
rect 4453 587 4456 1013
rect 4473 965 4927 1013
rect 4473 635 4535 965
rect 4865 635 4927 965
rect 4473 587 4927 635
rect 4944 587 4947 1013
rect 4453 581 4947 587
rect 5003 1013 5497 1019
rect 5003 587 5006 1013
rect 5023 965 5477 1013
rect 5023 635 5085 965
rect 5415 635 5477 965
rect 5023 587 5477 635
rect 5494 587 5497 1013
rect 5003 581 5497 587
rect 5553 1013 6047 1019
rect 5553 587 5556 1013
rect 5573 965 6027 1013
rect 5573 635 5635 965
rect 5965 635 6027 965
rect 5573 587 6027 635
rect 6044 587 6047 1013
rect 5553 581 6047 587
rect 6103 1013 6597 1019
rect 6103 587 6106 1013
rect 6123 965 6577 1013
rect 6123 635 6185 965
rect 6515 635 6577 965
rect 6123 587 6577 635
rect 6594 587 6597 1013
rect 6103 581 6597 587
rect 6653 1013 7147 1019
rect 6653 587 6656 1013
rect 6673 965 7127 1013
rect 6673 635 6735 965
rect 7065 635 7127 965
rect 6673 587 7127 635
rect 7144 587 7147 1013
rect 6653 581 7147 587
rect 7203 1013 7697 1019
rect 7203 587 7206 1013
rect 7223 965 7677 1013
rect 7223 635 7285 965
rect 7615 635 7677 965
rect 7223 587 7677 635
rect 7694 587 7697 1013
rect 7203 581 7697 587
rect 7753 1013 8247 1019
rect 7753 587 7756 1013
rect 7773 965 8227 1013
rect 7773 635 7835 965
rect 8165 635 8227 965
rect 7773 587 8227 635
rect 8244 587 8247 1013
rect 7753 581 8247 587
rect 8303 1013 8797 1019
rect 8303 587 8306 1013
rect 8323 965 8777 1013
rect 8323 635 8385 965
rect 8715 635 8777 965
rect 8323 587 8777 635
rect 8794 587 8797 1013
rect 8303 581 8797 587
rect 8853 1013 9347 1019
rect 8853 587 8856 1013
rect 8873 965 9327 1013
rect 8873 635 8935 965
rect 9265 635 9327 965
rect 8873 587 9327 635
rect 9344 587 9347 1013
rect 8853 581 9347 587
rect 9403 1013 9897 1019
rect 9403 587 9406 1013
rect 9423 965 9877 1013
rect 9423 635 9485 965
rect 9815 635 9877 965
rect 9423 587 9877 635
rect 9894 587 9897 1013
rect 9403 581 9897 587
rect 9953 1013 10447 1019
rect 9953 587 9956 1013
rect 9973 965 10427 1013
rect 9973 635 10035 965
rect 10365 635 10427 965
rect 9973 587 10427 635
rect 10444 587 10447 1013
rect 9953 581 10447 587
rect 10503 1013 10997 1019
rect 10503 587 10506 1013
rect 10523 965 10977 1013
rect 10523 635 10585 965
rect 10915 635 10977 965
rect 10523 587 10977 635
rect 10994 587 10997 1013
rect 10503 581 10997 587
rect 11053 1013 11547 1019
rect 11053 587 11056 1013
rect 11073 965 11527 1013
rect 11073 635 11135 965
rect 11465 635 11527 965
rect 11073 587 11527 635
rect 11544 587 11547 1013
rect 11053 581 11547 587
rect 11603 1013 12097 1019
rect 11603 587 11606 1013
rect 11623 965 12077 1013
rect 11623 635 11685 965
rect 12015 635 12077 965
rect 11623 587 12077 635
rect 12094 587 12097 1013
rect 11603 581 12097 587
rect 12153 1013 12647 1019
rect 12153 587 12156 1013
rect 12173 965 12627 1013
rect 12173 635 12235 965
rect 12565 635 12627 965
rect 12173 587 12627 635
rect 12644 587 12647 1013
rect 12153 581 12647 587
rect 12703 1013 13197 1019
rect 12703 587 12706 1013
rect 12723 965 13177 1013
rect 12723 635 12785 965
rect 13115 635 13177 965
rect 12723 587 13177 635
rect 13194 587 13197 1013
rect 12703 581 13197 587
rect 13253 1013 13724 1019
rect 13253 587 13256 1013
rect 13273 965 13724 1013
rect 13273 635 13335 965
rect 13665 635 13724 965
rect 13273 587 13724 635
rect 13253 581 13724 587
rect -474 576 -26 581
rect 76 576 524 581
rect 626 576 1074 581
rect 1176 576 1624 581
rect 1726 576 2174 581
rect 2276 576 2724 581
rect 2826 576 3274 581
rect 3376 576 3824 581
rect 3926 576 4374 581
rect 4476 576 4924 581
rect 5026 576 5474 581
rect 5576 576 6024 581
rect 6126 576 6574 581
rect 6676 576 7124 581
rect 7226 576 7674 581
rect 7776 576 8224 581
rect 8326 576 8774 581
rect 8876 576 9324 581
rect 9426 576 9874 581
rect 9976 576 10424 581
rect 10526 576 10974 581
rect 11076 576 11524 581
rect 11626 576 12074 581
rect 12176 576 12624 581
rect 12726 576 13174 581
rect 13276 576 13724 581
rect -1025 550 -725 569
rect -469 573 -31 576
rect -469 556 -463 573
rect -37 556 -31 573
rect -469 553 -31 556
rect 81 573 519 576
rect 81 556 87 573
rect 513 556 519 573
rect 81 553 519 556
rect 631 573 1069 576
rect 631 556 637 573
rect 1063 556 1069 573
rect 631 553 1069 556
rect 1181 573 1619 576
rect 1181 556 1187 573
rect 1613 556 1619 573
rect 1181 553 1619 556
rect 1731 573 2169 576
rect 1731 556 1737 573
rect 2163 556 2169 573
rect 1731 553 2169 556
rect 2281 573 2719 576
rect 2281 556 2287 573
rect 2713 556 2719 573
rect 2281 553 2719 556
rect 2831 573 3269 576
rect 2831 556 2837 573
rect 3263 556 3269 573
rect 2831 553 3269 556
rect 3381 573 3819 576
rect 3381 556 3387 573
rect 3813 556 3819 573
rect 3381 553 3819 556
rect 3931 573 4369 576
rect 3931 556 3937 573
rect 4363 556 4369 573
rect 3931 553 4369 556
rect 4481 573 4919 576
rect 4481 556 4487 573
rect 4913 556 4919 573
rect 4481 553 4919 556
rect 5031 573 5469 576
rect 5031 556 5037 573
rect 5463 556 5469 573
rect 5031 553 5469 556
rect 5581 573 6019 576
rect 5581 556 5587 573
rect 6013 556 6019 573
rect 5581 553 6019 556
rect 6131 573 6569 576
rect 6131 556 6137 573
rect 6563 556 6569 573
rect 6131 553 6569 556
rect 6681 573 7119 576
rect 6681 556 6687 573
rect 7113 556 7119 573
rect 6681 553 7119 556
rect 7231 573 7669 576
rect 7231 556 7237 573
rect 7663 556 7669 573
rect 7231 553 7669 556
rect 7781 573 8219 576
rect 7781 556 7787 573
rect 8213 556 8219 573
rect 7781 553 8219 556
rect 8331 573 8769 576
rect 8331 556 8337 573
rect 8763 556 8769 573
rect 8331 553 8769 556
rect 8881 573 9319 576
rect 8881 556 8887 573
rect 9313 556 9319 573
rect 8881 553 9319 556
rect 9431 573 9869 576
rect 9431 556 9437 573
rect 9863 556 9869 573
rect 9431 553 9869 556
rect 9981 573 10419 576
rect 9981 556 9987 573
rect 10413 556 10419 573
rect 9981 553 10419 556
rect 10531 573 10969 576
rect 10531 556 10537 573
rect 10963 556 10969 573
rect 10531 553 10969 556
rect 11081 573 11519 576
rect 11081 556 11087 573
rect 11513 556 11519 573
rect 11081 553 11519 556
rect 11631 573 12069 576
rect 11631 556 11637 573
rect 12063 556 12069 573
rect 11631 553 12069 556
rect 12181 573 12619 576
rect 12181 556 12187 573
rect 12613 556 12619 573
rect 12181 553 12619 556
rect 12731 573 13169 576
rect 12731 556 12737 573
rect 13163 556 13169 573
rect 12731 553 13169 556
rect 13281 573 13719 576
rect 13281 556 13287 573
rect 13713 556 13719 573
rect 13281 553 13719 556
rect 13975 569 13987 1100
rect 14263 569 14275 1100
rect 13975 550 14275 569
rect -1025 19 -1013 550
rect -737 19 -725 550
rect -550 542 -500 550
rect -550 508 -542 542
rect -508 508 -500 542
rect -550 500 -500 508
rect 0 542 50 550
rect 0 508 8 542
rect 42 508 50 542
rect 0 500 50 508
rect 550 542 600 550
rect 550 508 558 542
rect 592 508 600 542
rect 550 500 600 508
rect 1100 542 1150 550
rect 1100 508 1108 542
rect 1142 508 1150 542
rect 1100 500 1150 508
rect 1650 542 1700 550
rect 1650 508 1658 542
rect 1692 508 1700 542
rect 1650 500 1700 508
rect 2200 542 2250 550
rect 2200 508 2208 542
rect 2242 508 2250 542
rect 2200 500 2250 508
rect 2750 542 2800 550
rect 2750 508 2758 542
rect 2792 508 2800 542
rect 2750 500 2800 508
rect 3300 542 3350 550
rect 3300 508 3308 542
rect 3342 508 3350 542
rect 3300 500 3350 508
rect 3850 542 3900 550
rect 3850 508 3858 542
rect 3892 508 3900 542
rect 3850 500 3900 508
rect 4400 542 4450 550
rect 4400 508 4408 542
rect 4442 508 4450 542
rect 4400 500 4450 508
rect 4950 542 5000 550
rect 4950 508 4958 542
rect 4992 508 5000 542
rect 4950 500 5000 508
rect 5500 542 5550 550
rect 5500 508 5508 542
rect 5542 508 5550 542
rect 5500 500 5550 508
rect 6050 542 6100 550
rect 6050 508 6058 542
rect 6092 508 6100 542
rect 6050 500 6100 508
rect 6600 542 6650 550
rect 6600 508 6608 542
rect 6642 508 6650 542
rect 6600 500 6650 508
rect 7150 542 7200 550
rect 7150 508 7158 542
rect 7192 508 7200 542
rect 7150 500 7200 508
rect 7700 542 7750 550
rect 7700 508 7708 542
rect 7742 508 7750 542
rect 7700 500 7750 508
rect 8250 542 8300 550
rect 8250 508 8258 542
rect 8292 508 8300 542
rect 8250 500 8300 508
rect 8800 542 8850 550
rect 8800 508 8808 542
rect 8842 508 8850 542
rect 8800 500 8850 508
rect 9350 542 9400 550
rect 9350 508 9358 542
rect 9392 508 9400 542
rect 9350 500 9400 508
rect 9900 542 9950 550
rect 9900 508 9908 542
rect 9942 508 9950 542
rect 9900 500 9950 508
rect 10450 542 10500 550
rect 10450 508 10458 542
rect 10492 508 10500 542
rect 10450 500 10500 508
rect 11000 542 11050 550
rect 11000 508 11008 542
rect 11042 508 11050 542
rect 11000 500 11050 508
rect 11550 542 11600 550
rect 11550 508 11558 542
rect 11592 508 11600 542
rect 11550 500 11600 508
rect 12100 542 12150 550
rect 12100 508 12108 542
rect 12142 508 12150 542
rect 12100 500 12150 508
rect 12650 542 12700 550
rect 12650 508 12658 542
rect 12692 508 12700 542
rect 12650 500 12700 508
rect 13200 542 13250 550
rect 13200 508 13208 542
rect 13242 508 13250 542
rect 13200 500 13250 508
rect 13750 542 13800 550
rect 13750 508 13758 542
rect 13792 508 13800 542
rect 13750 500 13800 508
rect -469 494 -31 497
rect -469 477 -463 494
rect -37 477 -31 494
rect -469 474 -31 477
rect 81 494 519 497
rect 81 477 87 494
rect 513 477 519 494
rect 81 474 519 477
rect 631 494 1069 497
rect 631 477 637 494
rect 1063 477 1069 494
rect 631 474 1069 477
rect 1181 494 1619 497
rect 1181 477 1187 494
rect 1613 477 1619 494
rect 1181 474 1619 477
rect 1731 494 2169 497
rect 1731 477 1737 494
rect 2163 477 2169 494
rect 1731 474 2169 477
rect 2281 494 2719 497
rect 2281 477 2287 494
rect 2713 477 2719 494
rect 2281 474 2719 477
rect 2831 494 3269 497
rect 2831 477 2837 494
rect 3263 477 3269 494
rect 2831 474 3269 477
rect 3381 494 3819 497
rect 3381 477 3387 494
rect 3813 477 3819 494
rect 3381 474 3819 477
rect 3931 494 4369 497
rect 3931 477 3937 494
rect 4363 477 4369 494
rect 3931 474 4369 477
rect 4481 494 4919 497
rect 4481 477 4487 494
rect 4913 477 4919 494
rect 4481 474 4919 477
rect 5031 494 5469 497
rect 5031 477 5037 494
rect 5463 477 5469 494
rect 5031 474 5469 477
rect 5581 494 6019 497
rect 5581 477 5587 494
rect 6013 477 6019 494
rect 5581 474 6019 477
rect 6131 494 6569 497
rect 6131 477 6137 494
rect 6563 477 6569 494
rect 6131 474 6569 477
rect 6681 494 7119 497
rect 6681 477 6687 494
rect 7113 477 7119 494
rect 6681 474 7119 477
rect 7231 494 7669 497
rect 7231 477 7237 494
rect 7663 477 7669 494
rect 7231 474 7669 477
rect 7781 494 8219 497
rect 7781 477 7787 494
rect 8213 477 8219 494
rect 7781 474 8219 477
rect 8331 494 8769 497
rect 8331 477 8337 494
rect 8763 477 8769 494
rect 8331 474 8769 477
rect 8881 494 9319 497
rect 8881 477 8887 494
rect 9313 477 9319 494
rect 8881 474 9319 477
rect 9431 494 9869 497
rect 9431 477 9437 494
rect 9863 477 9869 494
rect 9431 474 9869 477
rect 9981 494 10419 497
rect 9981 477 9987 494
rect 10413 477 10419 494
rect 9981 474 10419 477
rect 10531 494 10969 497
rect 10531 477 10537 494
rect 10963 477 10969 494
rect 10531 474 10969 477
rect 11081 494 11519 497
rect 11081 477 11087 494
rect 11513 477 11519 494
rect 11081 474 11519 477
rect 11631 494 12069 497
rect 11631 477 11637 494
rect 12063 477 12069 494
rect 11631 474 12069 477
rect 12181 494 12619 497
rect 12181 477 12187 494
rect 12613 477 12619 494
rect 12181 474 12619 477
rect 12731 494 13169 497
rect 12731 477 12737 494
rect 13163 477 13169 494
rect 12731 474 13169 477
rect 13281 494 13719 497
rect 13281 477 13287 494
rect 13713 477 13719 494
rect 13281 474 13719 477
rect -474 469 -26 474
rect 76 469 524 474
rect 626 469 1074 474
rect 1176 469 1624 474
rect 1726 469 2174 474
rect 2276 469 2724 474
rect 2826 469 3274 474
rect 3376 469 3824 474
rect 3926 469 4374 474
rect 4476 469 4924 474
rect 5026 469 5474 474
rect 5576 469 6024 474
rect 6126 469 6574 474
rect 6676 469 7124 474
rect 7226 469 7674 474
rect 7776 469 8224 474
rect 8326 469 8774 474
rect 8876 469 9324 474
rect 9426 469 9874 474
rect 9976 469 10424 474
rect 10526 469 10974 474
rect 11076 469 11524 474
rect 11626 469 12074 474
rect 12176 469 12624 474
rect 12726 469 13174 474
rect 13276 469 13724 474
rect -474 463 -3 469
rect -474 415 -23 463
rect -474 85 -415 415
rect -85 85 -23 415
rect -474 37 -23 85
rect -6 37 -3 463
rect -474 31 -3 37
rect 53 463 547 469
rect 53 37 56 463
rect 73 415 527 463
rect 73 85 135 415
rect 465 85 527 415
rect 73 37 527 85
rect 544 37 547 463
rect 53 31 547 37
rect 603 463 1097 469
rect 603 37 606 463
rect 623 415 1077 463
rect 623 85 685 415
rect 1015 85 1077 415
rect 623 37 1077 85
rect 1094 37 1097 463
rect 603 31 1097 37
rect 1153 463 1647 469
rect 1153 37 1156 463
rect 1173 415 1627 463
rect 1173 85 1235 415
rect 1565 85 1627 415
rect 1173 37 1627 85
rect 1644 37 1647 463
rect 1153 31 1647 37
rect 1703 463 2197 469
rect 1703 37 1706 463
rect 1723 415 2177 463
rect 1723 85 1785 415
rect 2115 85 2177 415
rect 1723 37 2177 85
rect 2194 37 2197 463
rect 1703 31 2197 37
rect 2253 463 2747 469
rect 2253 37 2256 463
rect 2273 415 2727 463
rect 2273 85 2335 415
rect 2665 85 2727 415
rect 2273 37 2727 85
rect 2744 37 2747 463
rect 2253 31 2747 37
rect 2803 463 3297 469
rect 2803 37 2806 463
rect 2823 415 3277 463
rect 2823 85 2885 415
rect 3215 85 3277 415
rect 2823 37 3277 85
rect 3294 37 3297 463
rect 2803 31 3297 37
rect 3353 463 3847 469
rect 3353 37 3356 463
rect 3373 415 3827 463
rect 3373 85 3435 415
rect 3765 85 3827 415
rect 3373 37 3827 85
rect 3844 37 3847 463
rect 3353 31 3847 37
rect 3903 463 4397 469
rect 3903 37 3906 463
rect 3923 415 4377 463
rect 3923 85 3985 415
rect 4315 85 4377 415
rect 3923 37 4377 85
rect 4394 37 4397 463
rect 3903 31 4397 37
rect 4453 463 4947 469
rect 4453 37 4456 463
rect 4473 415 4927 463
rect 4473 85 4535 415
rect 4865 85 4927 415
rect 4473 37 4927 85
rect 4944 37 4947 463
rect 4453 31 4947 37
rect 5003 463 5497 469
rect 5003 37 5006 463
rect 5023 415 5477 463
rect 5023 85 5085 415
rect 5415 85 5477 415
rect 5023 37 5477 85
rect 5494 37 5497 463
rect 5003 31 5497 37
rect 5553 463 6047 469
rect 5553 37 5556 463
rect 5573 415 6027 463
rect 5573 85 5635 415
rect 5965 85 6027 415
rect 5573 37 6027 85
rect 6044 37 6047 463
rect 5553 31 6047 37
rect 6103 463 6597 469
rect 6103 37 6106 463
rect 6123 415 6577 463
rect 6123 85 6185 415
rect 6515 85 6577 415
rect 6123 37 6577 85
rect 6594 37 6597 463
rect 6103 31 6597 37
rect 6653 463 7147 469
rect 6653 37 6656 463
rect 6673 415 7127 463
rect 6673 85 6735 415
rect 7065 85 7127 415
rect 6673 37 7127 85
rect 7144 37 7147 463
rect 6653 31 7147 37
rect 7203 463 7697 469
rect 7203 37 7206 463
rect 7223 415 7677 463
rect 7223 85 7285 415
rect 7615 85 7677 415
rect 7223 37 7677 85
rect 7694 37 7697 463
rect 7203 31 7697 37
rect 7753 463 8247 469
rect 7753 37 7756 463
rect 7773 415 8227 463
rect 7773 85 7835 415
rect 8165 85 8227 415
rect 7773 37 8227 85
rect 8244 37 8247 463
rect 7753 31 8247 37
rect 8303 463 8797 469
rect 8303 37 8306 463
rect 8323 415 8777 463
rect 8323 85 8385 415
rect 8715 85 8777 415
rect 8323 37 8777 85
rect 8794 37 8797 463
rect 8303 31 8797 37
rect 8853 463 9347 469
rect 8853 37 8856 463
rect 8873 415 9327 463
rect 8873 85 8935 415
rect 9265 85 9327 415
rect 8873 37 9327 85
rect 9344 37 9347 463
rect 8853 31 9347 37
rect 9403 463 9897 469
rect 9403 37 9406 463
rect 9423 415 9877 463
rect 9423 85 9485 415
rect 9815 85 9877 415
rect 9423 37 9877 85
rect 9894 37 9897 463
rect 9403 31 9897 37
rect 9953 463 10447 469
rect 9953 37 9956 463
rect 9973 415 10427 463
rect 9973 85 10035 415
rect 10365 85 10427 415
rect 9973 37 10427 85
rect 10444 37 10447 463
rect 9953 31 10447 37
rect 10503 463 10997 469
rect 10503 37 10506 463
rect 10523 415 10977 463
rect 10523 85 10585 415
rect 10915 85 10977 415
rect 10523 37 10977 85
rect 10994 37 10997 463
rect 10503 31 10997 37
rect 11053 463 11547 469
rect 11053 37 11056 463
rect 11073 415 11527 463
rect 11073 85 11135 415
rect 11465 85 11527 415
rect 11073 37 11527 85
rect 11544 37 11547 463
rect 11053 31 11547 37
rect 11603 463 12097 469
rect 11603 37 11606 463
rect 11623 415 12077 463
rect 11623 85 11685 415
rect 12015 85 12077 415
rect 11623 37 12077 85
rect 12094 37 12097 463
rect 11603 31 12097 37
rect 12153 463 12647 469
rect 12153 37 12156 463
rect 12173 415 12627 463
rect 12173 85 12235 415
rect 12565 85 12627 415
rect 12173 37 12627 85
rect 12644 37 12647 463
rect 12153 31 12647 37
rect 12703 463 13197 469
rect 12703 37 12706 463
rect 12723 415 13177 463
rect 12723 85 12785 415
rect 13115 85 13177 415
rect 12723 37 13177 85
rect 13194 37 13197 463
rect 12703 31 13197 37
rect 13253 463 13724 469
rect 13253 37 13256 463
rect 13273 415 13724 463
rect 13273 85 13335 415
rect 13665 85 13724 415
rect 13273 37 13724 85
rect 13253 31 13724 37
rect -474 26 -26 31
rect 76 26 524 31
rect 626 26 1074 31
rect 1176 26 1624 31
rect 1726 26 2174 31
rect 2276 26 2724 31
rect 2826 26 3274 31
rect 3376 26 3824 31
rect 3926 26 4374 31
rect 4476 26 4924 31
rect 5026 26 5474 31
rect 5576 26 6024 31
rect 6126 26 6574 31
rect 6676 26 7124 31
rect 7226 26 7674 31
rect 7776 26 8224 31
rect 8326 26 8774 31
rect 8876 26 9324 31
rect 9426 26 9874 31
rect 9976 26 10424 31
rect 10526 26 10974 31
rect 11076 26 11524 31
rect 11626 26 12074 31
rect 12176 26 12624 31
rect 12726 26 13174 31
rect 13276 26 13724 31
rect -1025 0 -725 19
rect -469 23 -31 26
rect -469 6 -463 23
rect -37 6 -31 23
rect -469 3 -31 6
rect 81 23 519 26
rect 81 6 87 23
rect 513 6 519 23
rect 81 3 519 6
rect 631 23 1069 26
rect 631 6 637 23
rect 1063 6 1069 23
rect 631 3 1069 6
rect 1181 23 1619 26
rect 1181 6 1187 23
rect 1613 6 1619 23
rect 1181 3 1619 6
rect 1731 23 2169 26
rect 1731 6 1737 23
rect 2163 6 2169 23
rect 1731 3 2169 6
rect 2281 23 2719 26
rect 2281 6 2287 23
rect 2713 6 2719 23
rect 2281 3 2719 6
rect 2831 23 3269 26
rect 2831 6 2837 23
rect 3263 6 3269 23
rect 2831 3 3269 6
rect 3381 23 3819 26
rect 3381 6 3387 23
rect 3813 6 3819 23
rect 3381 3 3819 6
rect 3931 23 4369 26
rect 3931 6 3937 23
rect 4363 6 4369 23
rect 3931 3 4369 6
rect 4481 23 4919 26
rect 4481 6 4487 23
rect 4913 6 4919 23
rect 4481 3 4919 6
rect 5031 23 5469 26
rect 5031 6 5037 23
rect 5463 6 5469 23
rect 5031 3 5469 6
rect 5581 23 6019 26
rect 5581 6 5587 23
rect 6013 6 6019 23
rect 5581 3 6019 6
rect 6131 23 6569 26
rect 6131 6 6137 23
rect 6563 6 6569 23
rect 6131 3 6569 6
rect 6681 23 7119 26
rect 6681 6 6687 23
rect 7113 6 7119 23
rect 6681 3 7119 6
rect 7231 23 7669 26
rect 7231 6 7237 23
rect 7663 6 7669 23
rect 7231 3 7669 6
rect 7781 23 8219 26
rect 7781 6 7787 23
rect 8213 6 8219 23
rect 7781 3 8219 6
rect 8331 23 8769 26
rect 8331 6 8337 23
rect 8763 6 8769 23
rect 8331 3 8769 6
rect 8881 23 9319 26
rect 8881 6 8887 23
rect 9313 6 9319 23
rect 8881 3 9319 6
rect 9431 23 9869 26
rect 9431 6 9437 23
rect 9863 6 9869 23
rect 9431 3 9869 6
rect 9981 23 10419 26
rect 9981 6 9987 23
rect 10413 6 10419 23
rect 9981 3 10419 6
rect 10531 23 10969 26
rect 10531 6 10537 23
rect 10963 6 10969 23
rect 10531 3 10969 6
rect 11081 23 11519 26
rect 11081 6 11087 23
rect 11513 6 11519 23
rect 11081 3 11519 6
rect 11631 23 12069 26
rect 11631 6 11637 23
rect 12063 6 12069 23
rect 11631 3 12069 6
rect 12181 23 12619 26
rect 12181 6 12187 23
rect 12613 6 12619 23
rect 12181 3 12619 6
rect 12731 23 13169 26
rect 12731 6 12737 23
rect 13163 6 13169 23
rect 12731 3 13169 6
rect 13281 23 13719 26
rect 13281 6 13287 23
rect 13713 6 13719 23
rect 13281 3 13719 6
rect 13975 19 13987 550
rect 14263 19 14275 550
rect 13975 0 14275 19
rect -1025 -1063 -1013 0
rect -737 -775 -725 0
rect -550 -8 -500 0
rect -550 -42 -542 -8
rect -508 -42 -500 -8
rect -550 -50 -500 -42
rect 0 -8 50 0
rect 0 -42 8 -8
rect 42 -42 50 -8
rect 0 -50 50 -42
rect 550 -8 600 0
rect 550 -42 558 -8
rect 592 -42 600 -8
rect 550 -50 600 -42
rect 1100 -8 1150 0
rect 1100 -42 1108 -8
rect 1142 -42 1150 -8
rect 1100 -50 1150 -42
rect 1650 -8 1700 0
rect 1650 -42 1658 -8
rect 1692 -42 1700 -8
rect 1650 -50 1700 -42
rect 2200 -8 2250 0
rect 2200 -42 2208 -8
rect 2242 -42 2250 -8
rect 2200 -50 2250 -42
rect 2750 -8 2800 0
rect 2750 -42 2758 -8
rect 2792 -42 2800 -8
rect 2750 -50 2800 -42
rect 3300 -8 3350 0
rect 3300 -42 3308 -8
rect 3342 -42 3350 -8
rect 3300 -50 3350 -42
rect 3850 -8 3900 0
rect 3850 -42 3858 -8
rect 3892 -42 3900 -8
rect 3850 -50 3900 -42
rect 4400 -8 4450 0
rect 4400 -42 4408 -8
rect 4442 -42 4450 -8
rect 4400 -50 4450 -42
rect 4950 -8 5000 0
rect 4950 -42 4958 -8
rect 4992 -42 5000 -8
rect 4950 -50 5000 -42
rect 5500 -8 5550 0
rect 5500 -42 5508 -8
rect 5542 -42 5550 -8
rect 5500 -50 5550 -42
rect 6050 -8 6100 0
rect 6050 -42 6058 -8
rect 6092 -42 6100 -8
rect 6050 -50 6100 -42
rect 6600 -8 6650 0
rect 6600 -42 6608 -8
rect 6642 -42 6650 -8
rect 6600 -50 6650 -42
rect 7150 -8 7200 0
rect 7150 -42 7158 -8
rect 7192 -42 7200 -8
rect 7150 -50 7200 -42
rect 7700 -8 7750 0
rect 7700 -42 7708 -8
rect 7742 -42 7750 -8
rect 7700 -50 7750 -42
rect 8250 -8 8300 0
rect 8250 -42 8258 -8
rect 8292 -42 8300 -8
rect 8250 -50 8300 -42
rect 8800 -8 8850 0
rect 8800 -42 8808 -8
rect 8842 -42 8850 -8
rect 8800 -50 8850 -42
rect 9350 -8 9400 0
rect 9350 -42 9358 -8
rect 9392 -42 9400 -8
rect 9350 -50 9400 -42
rect 9900 -8 9950 0
rect 9900 -42 9908 -8
rect 9942 -42 9950 -8
rect 9900 -50 9950 -42
rect 10450 -8 10500 0
rect 10450 -42 10458 -8
rect 10492 -42 10500 -8
rect 10450 -50 10500 -42
rect 11000 -8 11050 0
rect 11000 -42 11008 -8
rect 11042 -42 11050 -8
rect 11000 -50 11050 -42
rect 11550 -8 11600 0
rect 11550 -42 11558 -8
rect 11592 -42 11600 -8
rect 11550 -50 11600 -42
rect 12100 -8 12150 0
rect 12100 -42 12108 -8
rect 12142 -42 12150 -8
rect 12100 -50 12150 -42
rect 12650 -8 12700 0
rect 12650 -42 12658 -8
rect 12692 -42 12700 -8
rect 12650 -50 12700 -42
rect 13200 -8 13250 0
rect 13200 -42 13208 -8
rect 13242 -42 13250 -8
rect 13200 -50 13250 -42
rect 13750 -8 13800 0
rect 13750 -42 13758 -8
rect 13792 -42 13800 -8
rect 13750 -50 13800 -42
rect -469 -56 -31 -53
rect -469 -73 -463 -56
rect -37 -73 -31 -56
rect -469 -76 -31 -73
rect 81 -56 519 -53
rect 81 -73 87 -56
rect 513 -73 519 -56
rect 81 -76 519 -73
rect 631 -56 1069 -53
rect 631 -73 637 -56
rect 1063 -73 1069 -56
rect 631 -76 1069 -73
rect 1181 -56 1619 -53
rect 1181 -73 1187 -56
rect 1613 -73 1619 -56
rect 1181 -76 1619 -73
rect 1731 -56 2169 -53
rect 1731 -73 1737 -56
rect 2163 -73 2169 -56
rect 1731 -76 2169 -73
rect 2281 -56 2719 -53
rect 2281 -73 2287 -56
rect 2713 -73 2719 -56
rect 2281 -76 2719 -73
rect 2831 -56 3269 -53
rect 2831 -73 2837 -56
rect 3263 -73 3269 -56
rect 2831 -76 3269 -73
rect 3381 -56 3819 -53
rect 3381 -73 3387 -56
rect 3813 -73 3819 -56
rect 3381 -76 3819 -73
rect 3931 -56 4369 -53
rect 3931 -73 3937 -56
rect 4363 -73 4369 -56
rect 3931 -76 4369 -73
rect 4481 -56 4919 -53
rect 4481 -73 4487 -56
rect 4913 -73 4919 -56
rect 4481 -76 4919 -73
rect 5031 -56 5469 -53
rect 5031 -73 5037 -56
rect 5463 -73 5469 -56
rect 5031 -76 5469 -73
rect 5581 -56 6019 -53
rect 5581 -73 5587 -56
rect 6013 -73 6019 -56
rect 5581 -76 6019 -73
rect 6131 -56 6569 -53
rect 6131 -73 6137 -56
rect 6563 -73 6569 -56
rect 6131 -76 6569 -73
rect 6681 -56 7119 -53
rect 6681 -73 6687 -56
rect 7113 -73 7119 -56
rect 6681 -76 7119 -73
rect 7231 -56 7669 -53
rect 7231 -73 7237 -56
rect 7663 -73 7669 -56
rect 7231 -76 7669 -73
rect 7781 -56 8219 -53
rect 7781 -73 7787 -56
rect 8213 -73 8219 -56
rect 7781 -76 8219 -73
rect 8331 -56 8769 -53
rect 8331 -73 8337 -56
rect 8763 -73 8769 -56
rect 8331 -76 8769 -73
rect 8881 -56 9319 -53
rect 8881 -73 8887 -56
rect 9313 -73 9319 -56
rect 8881 -76 9319 -73
rect 9431 -56 9869 -53
rect 9431 -73 9437 -56
rect 9863 -73 9869 -56
rect 9431 -76 9869 -73
rect 9981 -56 10419 -53
rect 9981 -73 9987 -56
rect 10413 -73 10419 -56
rect 9981 -76 10419 -73
rect 10531 -56 10969 -53
rect 10531 -73 10537 -56
rect 10963 -73 10969 -56
rect 10531 -76 10969 -73
rect 11081 -56 11519 -53
rect 11081 -73 11087 -56
rect 11513 -73 11519 -56
rect 11081 -76 11519 -73
rect 11631 -56 12069 -53
rect 11631 -73 11637 -56
rect 12063 -73 12069 -56
rect 11631 -76 12069 -73
rect 12181 -56 12619 -53
rect 12181 -73 12187 -56
rect 12613 -73 12619 -56
rect 12181 -76 12619 -73
rect 12731 -56 13169 -53
rect 12731 -73 12737 -56
rect 13163 -73 13169 -56
rect 12731 -76 13169 -73
rect 13281 -56 13719 -53
rect 13281 -73 13287 -56
rect 13713 -73 13719 -56
rect 13281 -76 13719 -73
rect -474 -81 -26 -76
rect 76 -81 524 -76
rect 626 -81 1074 -76
rect 1176 -81 1624 -76
rect 1726 -81 2174 -76
rect 2276 -81 2724 -76
rect 2826 -81 3274 -76
rect 3376 -81 3824 -76
rect 3926 -81 4374 -76
rect 4476 -81 4924 -76
rect 5026 -81 5474 -76
rect 5576 -81 6024 -76
rect 6126 -81 6574 -76
rect 6676 -81 7124 -76
rect 7226 -81 7674 -76
rect 7776 -81 8224 -76
rect 8326 -81 8774 -76
rect 8876 -81 9324 -76
rect 9426 -81 9874 -76
rect 9976 -81 10424 -76
rect 10526 -81 10974 -76
rect 11076 -81 11524 -76
rect 11626 -81 12074 -76
rect 12176 -81 12624 -76
rect 12726 -81 13174 -76
rect 13276 -81 13724 -76
rect -474 -87 -3 -81
rect -474 -135 -23 -87
rect -474 -465 -415 -135
rect -85 -465 -23 -135
rect -474 -513 -23 -465
rect -6 -513 -3 -87
rect -474 -519 -3 -513
rect 53 -87 547 -81
rect 53 -513 56 -87
rect 73 -135 527 -87
rect 73 -465 135 -135
rect 465 -465 527 -135
rect 73 -513 527 -465
rect 544 -513 547 -87
rect 53 -519 547 -513
rect 603 -87 1097 -81
rect 603 -513 606 -87
rect 623 -135 1077 -87
rect 623 -465 685 -135
rect 1015 -465 1077 -135
rect 623 -513 1077 -465
rect 1094 -513 1097 -87
rect 603 -519 1097 -513
rect 1153 -87 1647 -81
rect 1153 -513 1156 -87
rect 1173 -135 1627 -87
rect 1173 -465 1235 -135
rect 1565 -465 1627 -135
rect 1173 -513 1627 -465
rect 1644 -513 1647 -87
rect 1153 -519 1647 -513
rect 1703 -87 2197 -81
rect 1703 -513 1706 -87
rect 1723 -135 2177 -87
rect 1723 -465 1785 -135
rect 2115 -465 2177 -135
rect 1723 -513 2177 -465
rect 2194 -513 2197 -87
rect 1703 -519 2197 -513
rect 2253 -87 2747 -81
rect 2253 -513 2256 -87
rect 2273 -135 2727 -87
rect 2273 -465 2335 -135
rect 2665 -465 2727 -135
rect 2273 -513 2727 -465
rect 2744 -513 2747 -87
rect 2253 -519 2747 -513
rect 2803 -87 3297 -81
rect 2803 -513 2806 -87
rect 2823 -135 3277 -87
rect 2823 -465 2885 -135
rect 3215 -465 3277 -135
rect 2823 -513 3277 -465
rect 3294 -513 3297 -87
rect 2803 -519 3297 -513
rect 3353 -87 3847 -81
rect 3353 -513 3356 -87
rect 3373 -135 3827 -87
rect 3373 -465 3435 -135
rect 3765 -465 3827 -135
rect 3373 -513 3827 -465
rect 3844 -513 3847 -87
rect 3353 -519 3847 -513
rect 3903 -87 4397 -81
rect 3903 -513 3906 -87
rect 3923 -135 4377 -87
rect 3923 -465 3985 -135
rect 4315 -465 4377 -135
rect 3923 -513 4377 -465
rect 4394 -513 4397 -87
rect 3903 -519 4397 -513
rect 4453 -87 4947 -81
rect 4453 -513 4456 -87
rect 4473 -135 4927 -87
rect 4473 -465 4535 -135
rect 4865 -465 4927 -135
rect 4473 -513 4927 -465
rect 4944 -513 4947 -87
rect 4453 -519 4947 -513
rect 5003 -87 5497 -81
rect 5003 -513 5006 -87
rect 5023 -135 5477 -87
rect 5023 -465 5085 -135
rect 5415 -465 5477 -135
rect 5023 -513 5477 -465
rect 5494 -513 5497 -87
rect 5003 -519 5497 -513
rect 5553 -87 6047 -81
rect 5553 -513 5556 -87
rect 5573 -135 6027 -87
rect 5573 -465 5635 -135
rect 5965 -465 6027 -135
rect 5573 -513 6027 -465
rect 6044 -513 6047 -87
rect 5553 -519 6047 -513
rect 6103 -87 6597 -81
rect 6103 -513 6106 -87
rect 6123 -135 6577 -87
rect 6123 -465 6185 -135
rect 6515 -465 6577 -135
rect 6123 -513 6577 -465
rect 6594 -513 6597 -87
rect 6103 -519 6597 -513
rect 6653 -87 7147 -81
rect 6653 -513 6656 -87
rect 6673 -135 7127 -87
rect 6673 -465 6735 -135
rect 7065 -465 7127 -135
rect 6673 -513 7127 -465
rect 7144 -513 7147 -87
rect 6653 -519 7147 -513
rect 7203 -87 7697 -81
rect 7203 -513 7206 -87
rect 7223 -135 7677 -87
rect 7223 -465 7285 -135
rect 7615 -465 7677 -135
rect 7223 -513 7677 -465
rect 7694 -513 7697 -87
rect 7203 -519 7697 -513
rect 7753 -87 8247 -81
rect 7753 -513 7756 -87
rect 7773 -135 8227 -87
rect 7773 -465 7835 -135
rect 8165 -465 8227 -135
rect 7773 -513 8227 -465
rect 8244 -513 8247 -87
rect 7753 -519 8247 -513
rect 8303 -87 8797 -81
rect 8303 -513 8306 -87
rect 8323 -135 8777 -87
rect 8323 -465 8385 -135
rect 8715 -465 8777 -135
rect 8323 -513 8777 -465
rect 8794 -513 8797 -87
rect 8303 -519 8797 -513
rect 8853 -87 9347 -81
rect 8853 -513 8856 -87
rect 8873 -135 9327 -87
rect 8873 -465 8935 -135
rect 9265 -465 9327 -135
rect 8873 -513 9327 -465
rect 9344 -513 9347 -87
rect 8853 -519 9347 -513
rect 9403 -87 9897 -81
rect 9403 -513 9406 -87
rect 9423 -135 9877 -87
rect 9423 -465 9485 -135
rect 9815 -465 9877 -135
rect 9423 -513 9877 -465
rect 9894 -513 9897 -87
rect 9403 -519 9897 -513
rect 9953 -87 10447 -81
rect 9953 -513 9956 -87
rect 9973 -135 10427 -87
rect 9973 -465 10035 -135
rect 10365 -465 10427 -135
rect 9973 -513 10427 -465
rect 10444 -513 10447 -87
rect 9953 -519 10447 -513
rect 10503 -87 10997 -81
rect 10503 -513 10506 -87
rect 10523 -135 10977 -87
rect 10523 -465 10585 -135
rect 10915 -465 10977 -135
rect 10523 -513 10977 -465
rect 10994 -513 10997 -87
rect 10503 -519 10997 -513
rect 11053 -87 11547 -81
rect 11053 -513 11056 -87
rect 11073 -135 11527 -87
rect 11073 -465 11135 -135
rect 11465 -465 11527 -135
rect 11073 -513 11527 -465
rect 11544 -513 11547 -87
rect 11053 -519 11547 -513
rect 11603 -87 12097 -81
rect 11603 -513 11606 -87
rect 11623 -135 12077 -87
rect 11623 -465 11685 -135
rect 12015 -465 12077 -135
rect 11623 -513 12077 -465
rect 12094 -513 12097 -87
rect 11603 -519 12097 -513
rect 12153 -87 12647 -81
rect 12153 -513 12156 -87
rect 12173 -135 12627 -87
rect 12173 -465 12235 -135
rect 12565 -465 12627 -135
rect 12173 -513 12627 -465
rect 12644 -513 12647 -87
rect 12153 -519 12647 -513
rect 12703 -87 13197 -81
rect 12703 -513 12706 -87
rect 12723 -135 13177 -87
rect 12723 -465 12785 -135
rect 13115 -465 13177 -135
rect 12723 -513 13177 -465
rect 13194 -513 13197 -87
rect 12703 -519 13197 -513
rect 13253 -87 13724 -81
rect 13253 -513 13256 -87
rect 13273 -135 13724 -87
rect 13273 -465 13335 -135
rect 13665 -465 13724 -135
rect 13273 -513 13724 -465
rect 13253 -519 13724 -513
rect -474 -524 -26 -519
rect 76 -524 524 -519
rect 626 -524 1074 -519
rect 1176 -524 1624 -519
rect 1726 -524 2174 -519
rect 2276 -524 2724 -519
rect 2826 -524 3274 -519
rect 3376 -524 3824 -519
rect 3926 -524 4374 -519
rect 4476 -524 4924 -519
rect 5026 -524 5474 -519
rect 5576 -524 6024 -519
rect 6126 -524 6574 -519
rect 6676 -524 7124 -519
rect 7226 -524 7674 -519
rect 7776 -524 8224 -519
rect 8326 -524 8774 -519
rect 8876 -524 9324 -519
rect 9426 -524 9874 -519
rect 9976 -524 10424 -519
rect 10526 -524 10974 -519
rect 11076 -524 11524 -519
rect 11626 -524 12074 -519
rect 12176 -524 12624 -519
rect 12726 -524 13174 -519
rect 13276 -524 13724 -519
rect -550 -558 -500 -550
rect -550 -592 -542 -558
rect -508 -592 -500 -558
rect -550 -600 -500 -592
rect 0 -558 50 -550
rect 0 -592 8 -558
rect 42 -592 50 -558
rect 0 -600 50 -592
rect 550 -558 600 -550
rect 550 -592 558 -558
rect 592 -592 600 -558
rect 550 -600 600 -592
rect 1100 -558 1150 -550
rect 1100 -592 1108 -558
rect 1142 -592 1150 -558
rect 1100 -600 1150 -592
rect 1650 -558 1700 -550
rect 1650 -592 1658 -558
rect 1692 -592 1700 -558
rect 1650 -600 1700 -592
rect 2200 -558 2250 -550
rect 2200 -592 2208 -558
rect 2242 -592 2250 -558
rect 2200 -600 2250 -592
rect 2750 -558 2800 -550
rect 2750 -592 2758 -558
rect 2792 -592 2800 -558
rect 2750 -600 2800 -592
rect 3300 -558 3350 -550
rect 3300 -592 3308 -558
rect 3342 -592 3350 -558
rect 3300 -600 3350 -592
rect 3850 -558 3900 -550
rect 3850 -592 3858 -558
rect 3892 -592 3900 -558
rect 3850 -600 3900 -592
rect 4400 -558 4450 -550
rect 4400 -592 4408 -558
rect 4442 -592 4450 -558
rect 4400 -600 4450 -592
rect 4950 -558 5000 -550
rect 4950 -592 4958 -558
rect 4992 -592 5000 -558
rect 4950 -600 5000 -592
rect 5500 -558 5550 -550
rect 5500 -592 5508 -558
rect 5542 -592 5550 -558
rect 5500 -600 5550 -592
rect 6050 -558 6100 -550
rect 6050 -592 6058 -558
rect 6092 -592 6100 -558
rect 6050 -600 6100 -592
rect 6600 -558 6650 -550
rect 6600 -592 6608 -558
rect 6642 -592 6650 -558
rect 6600 -600 6650 -592
rect 7150 -558 7200 -550
rect 7150 -592 7158 -558
rect 7192 -592 7200 -558
rect 7150 -600 7200 -592
rect 7700 -558 7750 -550
rect 7700 -592 7708 -558
rect 7742 -592 7750 -558
rect 7700 -600 7750 -592
rect 8250 -558 8300 -550
rect 8250 -592 8258 -558
rect 8292 -592 8300 -558
rect 8250 -600 8300 -592
rect 8800 -558 8850 -550
rect 8800 -592 8808 -558
rect 8842 -592 8850 -558
rect 8800 -600 8850 -592
rect 9350 -558 9400 -550
rect 9350 -592 9358 -558
rect 9392 -592 9400 -558
rect 9350 -600 9400 -592
rect 9900 -558 9950 -550
rect 9900 -592 9908 -558
rect 9942 -592 9950 -558
rect 9900 -600 9950 -592
rect 10450 -558 10500 -550
rect 10450 -592 10458 -558
rect 10492 -592 10500 -558
rect 10450 -600 10500 -592
rect 11000 -558 11050 -550
rect 11000 -592 11008 -558
rect 11042 -592 11050 -558
rect 11000 -600 11050 -592
rect 11550 -558 11600 -550
rect 11550 -592 11558 -558
rect 11592 -592 11600 -558
rect 11550 -600 11600 -592
rect 12100 -558 12150 -550
rect 12100 -592 12108 -558
rect 12142 -592 12150 -558
rect 12100 -600 12150 -592
rect 12650 -558 12700 -550
rect 12650 -592 12658 -558
rect 12692 -592 12700 -558
rect 12650 -600 12700 -592
rect 13200 -558 13250 -550
rect 13200 -592 13208 -558
rect 13242 -592 13250 -558
rect 13200 -600 13250 -592
rect 13750 -558 13800 -550
rect 13750 -592 13758 -558
rect 13792 -592 13800 -558
rect 13750 -600 13800 -592
rect 13975 -775 13987 0
rect -737 -787 13987 -775
rect -19 -1063 0 -787
rect 531 -1063 550 -787
rect 1081 -1063 1100 -787
rect 1631 -1063 1650 -787
rect 2181 -1063 2200 -787
rect 2731 -1063 2750 -787
rect 3281 -1063 3300 -787
rect 3831 -1063 3850 -787
rect 4381 -1063 4400 -787
rect 4931 -1063 4950 -787
rect 5481 -1063 5500 -787
rect 6031 -1063 6050 -787
rect 6581 -1063 6600 -787
rect 7131 -1063 7150 -787
rect 7681 -1063 7700 -787
rect 8231 -1063 8250 -787
rect 8781 -1063 8800 -787
rect 9331 -1063 9350 -787
rect 9881 -1063 9900 -787
rect 10431 -1063 10450 -787
rect 10981 -1063 11000 -787
rect 11531 -1063 11550 -787
rect 12081 -1063 12100 -787
rect 12631 -1063 12650 -787
rect 13181 -1063 13200 -787
rect 14263 -1063 14275 0
rect -1025 -1075 14275 -1063
rect 14775 -1575 14787 14725
rect -1537 -1587 14787 -1575
rect 18763 -5563 18775 18713
rect -5525 -5575 18775 -5563
<< via1 >>
rect -5513 14737 18763 18713
rect -5513 1117 -1537 14725
rect 88 14025 188 14125
rect 1188 14025 1288 14125
rect 2288 14025 2388 14125
rect 3388 14025 3488 14125
rect 4488 14025 4588 14125
rect 5588 14025 5688 14125
rect 6688 14025 6788 14125
rect 7788 14025 7888 14125
rect 8888 14025 8988 14125
rect 9988 14025 10088 14125
rect 11088 14025 11188 14125
rect 12188 14025 12288 14125
rect 13288 14025 13388 14125
rect -542 13708 -508 13742
rect 8 13708 42 13742
rect 558 13708 592 13742
rect 1108 13708 1142 13742
rect 1658 13708 1692 13742
rect 2208 13708 2242 13742
rect 2758 13708 2792 13742
rect 3308 13708 3342 13742
rect 3858 13708 3892 13742
rect 4408 13708 4442 13742
rect 4958 13708 4992 13742
rect 5508 13708 5542 13742
rect 6058 13708 6092 13742
rect 6608 13708 6642 13742
rect 7158 13708 7192 13742
rect 7708 13708 7742 13742
rect 8258 13708 8292 13742
rect 8808 13708 8842 13742
rect 9358 13708 9392 13742
rect 9908 13708 9942 13742
rect 10458 13708 10492 13742
rect 11008 13708 11042 13742
rect 11558 13708 11592 13742
rect 12108 13708 12142 13742
rect 12658 13708 12692 13742
rect 13208 13708 13242 13742
rect 13758 13708 13792 13742
rect -415 13285 -85 13615
rect 135 13285 465 13615
rect 685 13285 1015 13615
rect 1235 13285 1565 13615
rect 1785 13285 2115 13615
rect 2335 13285 2665 13615
rect 2885 13285 3215 13615
rect 3435 13285 3765 13615
rect 3985 13285 4315 13615
rect 4535 13285 4865 13615
rect 5085 13285 5415 13615
rect 5635 13285 5965 13615
rect 6185 13285 6515 13615
rect 6735 13285 7065 13615
rect 7285 13285 7615 13615
rect 7835 13285 8165 13615
rect 8385 13285 8715 13615
rect 8935 13285 9265 13615
rect 9485 13285 9815 13615
rect 10035 13285 10365 13615
rect 10585 13285 10915 13615
rect 11135 13285 11465 13615
rect 11685 13285 12015 13615
rect 12235 13285 12565 13615
rect 12785 13285 13115 13615
rect 13335 13285 13665 13615
rect 14075 13238 14175 13338
rect -925 13012 -825 13112
rect -542 13158 -508 13192
rect 8 13158 42 13192
rect 558 13158 592 13192
rect 1108 13158 1142 13192
rect 1658 13158 1692 13192
rect 2208 13158 2242 13192
rect 2758 13158 2792 13192
rect 3308 13158 3342 13192
rect 3858 13158 3892 13192
rect 4408 13158 4442 13192
rect 4958 13158 4992 13192
rect 5508 13158 5542 13192
rect 6058 13158 6092 13192
rect 6608 13158 6642 13192
rect 7158 13158 7192 13192
rect 7708 13158 7742 13192
rect 8258 13158 8292 13192
rect 8808 13158 8842 13192
rect 9358 13158 9392 13192
rect 9908 13158 9942 13192
rect 10458 13158 10492 13192
rect 11008 13158 11042 13192
rect 11558 13158 11592 13192
rect 12108 13158 12142 13192
rect 12658 13158 12692 13192
rect 13208 13158 13242 13192
rect 13758 13158 13792 13192
rect -415 12735 -85 13065
rect 135 12735 465 13065
rect 685 12735 1015 13065
rect 1235 12735 1565 13065
rect 1785 12735 2115 13065
rect 2335 12735 2665 13065
rect 2885 12735 3215 13065
rect 3435 12735 3765 13065
rect 3985 12735 4315 13065
rect 4535 12735 4865 13065
rect 5085 12735 5415 13065
rect 5635 12735 5965 13065
rect 6185 12735 6515 13065
rect 6735 12735 7065 13065
rect 7285 12735 7615 13065
rect 7835 12735 8165 13065
rect 8385 12735 8715 13065
rect 8935 12735 9265 13065
rect 9485 12735 9815 13065
rect 10035 12735 10365 13065
rect 10585 12735 10915 13065
rect 11135 12735 11465 13065
rect 11685 12735 12015 13065
rect 12235 12735 12565 13065
rect 12785 12735 13115 13065
rect 13335 12735 13665 13065
rect -542 12608 -508 12642
rect 8 12608 42 12642
rect 558 12608 592 12642
rect 1108 12608 1142 12642
rect 1658 12608 1692 12642
rect 2208 12608 2242 12642
rect 2758 12608 2792 12642
rect 3308 12608 3342 12642
rect 3858 12608 3892 12642
rect 4408 12608 4442 12642
rect 4958 12608 4992 12642
rect 5508 12608 5542 12642
rect 6058 12608 6092 12642
rect 6608 12608 6642 12642
rect 7158 12608 7192 12642
rect 7708 12608 7742 12642
rect 8258 12608 8292 12642
rect 8808 12608 8842 12642
rect 9358 12608 9392 12642
rect 9908 12608 9942 12642
rect 10458 12608 10492 12642
rect 11008 12608 11042 12642
rect 11558 12608 11592 12642
rect 12108 12608 12142 12642
rect 12658 12608 12692 12642
rect 13208 12608 13242 12642
rect 13758 12608 13792 12642
rect -415 12185 -85 12515
rect 135 12185 465 12515
rect 685 12185 1015 12515
rect 1235 12185 1565 12515
rect 1785 12185 2115 12515
rect 2335 12185 2665 12515
rect 2885 12185 3215 12515
rect 3435 12185 3765 12515
rect 3985 12185 4315 12515
rect 4535 12185 4865 12515
rect 5085 12185 5415 12515
rect 5635 12185 5965 12515
rect 6185 12185 6515 12515
rect 6735 12185 7065 12515
rect 7285 12185 7615 12515
rect 7835 12185 8165 12515
rect 8385 12185 8715 12515
rect 8935 12185 9265 12515
rect 9485 12185 9815 12515
rect 10035 12185 10365 12515
rect 10585 12185 10915 12515
rect 11135 12185 11465 12515
rect 11685 12185 12015 12515
rect 12235 12185 12565 12515
rect 12785 12185 13115 12515
rect 13335 12185 13665 12515
rect 14075 12138 14175 12238
rect -925 11912 -825 12012
rect -542 12058 -508 12092
rect 8 12058 42 12092
rect 558 12058 592 12092
rect 1108 12058 1142 12092
rect 1658 12058 1692 12092
rect 2208 12058 2242 12092
rect 2758 12058 2792 12092
rect 3308 12058 3342 12092
rect 3858 12058 3892 12092
rect 4408 12058 4442 12092
rect 4958 12058 4992 12092
rect 5508 12058 5542 12092
rect 6058 12058 6092 12092
rect 6608 12058 6642 12092
rect 7158 12058 7192 12092
rect 7708 12058 7742 12092
rect 8258 12058 8292 12092
rect 8808 12058 8842 12092
rect 9358 12058 9392 12092
rect 9908 12058 9942 12092
rect 10458 12058 10492 12092
rect 11008 12058 11042 12092
rect 11558 12058 11592 12092
rect 12108 12058 12142 12092
rect 12658 12058 12692 12092
rect 13208 12058 13242 12092
rect 13758 12058 13792 12092
rect -415 11635 -85 11965
rect 135 11635 465 11965
rect 685 11635 1015 11965
rect 1235 11635 1565 11965
rect 1785 11635 2115 11965
rect 2335 11635 2665 11965
rect 2885 11635 3215 11965
rect 3435 11635 3765 11965
rect 3985 11635 4315 11965
rect 4535 11635 4865 11965
rect 5085 11635 5415 11965
rect 5635 11635 5965 11965
rect 6185 11635 6515 11965
rect 6735 11635 7065 11965
rect 7285 11635 7615 11965
rect 7835 11635 8165 11965
rect 8385 11635 8715 11965
rect 8935 11635 9265 11965
rect 9485 11635 9815 11965
rect 10035 11635 10365 11965
rect 10585 11635 10915 11965
rect 11135 11635 11465 11965
rect 11685 11635 12015 11965
rect 12235 11635 12565 11965
rect 12785 11635 13115 11965
rect 13335 11635 13665 11965
rect -542 11508 -508 11542
rect 8 11508 42 11542
rect 558 11508 592 11542
rect 1108 11508 1142 11542
rect 1658 11508 1692 11542
rect 2208 11508 2242 11542
rect 2758 11508 2792 11542
rect 3308 11508 3342 11542
rect 3858 11508 3892 11542
rect 4408 11508 4442 11542
rect 4958 11508 4992 11542
rect 5508 11508 5542 11542
rect 6058 11508 6092 11542
rect 6608 11508 6642 11542
rect 7158 11508 7192 11542
rect 7708 11508 7742 11542
rect 8258 11508 8292 11542
rect 8808 11508 8842 11542
rect 9358 11508 9392 11542
rect 9908 11508 9942 11542
rect 10458 11508 10492 11542
rect 11008 11508 11042 11542
rect 11558 11508 11592 11542
rect 12108 11508 12142 11542
rect 12658 11508 12692 11542
rect 13208 11508 13242 11542
rect 13758 11508 13792 11542
rect -415 11085 -85 11415
rect 135 11085 465 11415
rect 685 11085 1015 11415
rect 1235 11085 1565 11415
rect 1785 11085 2115 11415
rect 2335 11085 2665 11415
rect 2885 11085 3215 11415
rect 3435 11085 3765 11415
rect 3985 11085 4315 11415
rect 4535 11085 4865 11415
rect 5085 11085 5415 11415
rect 5635 11085 5965 11415
rect 6185 11085 6515 11415
rect 6735 11085 7065 11415
rect 7285 11085 7615 11415
rect 7835 11085 8165 11415
rect 8385 11085 8715 11415
rect 8935 11085 9265 11415
rect 9485 11085 9815 11415
rect 10035 11085 10365 11415
rect 10585 11085 10915 11415
rect 11135 11085 11465 11415
rect 11685 11085 12015 11415
rect 12235 11085 12565 11415
rect 12785 11085 13115 11415
rect 13335 11085 13665 11415
rect 14075 11038 14175 11138
rect -925 10812 -825 10912
rect -542 10958 -508 10992
rect 8 10958 42 10992
rect 558 10958 592 10992
rect 1108 10958 1142 10992
rect 1658 10958 1692 10992
rect 2208 10958 2242 10992
rect 2758 10958 2792 10992
rect 3308 10958 3342 10992
rect 3858 10958 3892 10992
rect 4408 10958 4442 10992
rect 4958 10958 4992 10992
rect 5508 10958 5542 10992
rect 6058 10958 6092 10992
rect 6608 10958 6642 10992
rect 7158 10958 7192 10992
rect 7708 10958 7742 10992
rect 8258 10958 8292 10992
rect 8808 10958 8842 10992
rect 9358 10958 9392 10992
rect 9908 10958 9942 10992
rect 10458 10958 10492 10992
rect 11008 10958 11042 10992
rect 11558 10958 11592 10992
rect 12108 10958 12142 10992
rect 12658 10958 12692 10992
rect 13208 10958 13242 10992
rect 13758 10958 13792 10992
rect -415 10535 -85 10865
rect 135 10535 465 10865
rect 685 10535 1015 10865
rect 1235 10535 1565 10865
rect 1785 10535 2115 10865
rect 2335 10535 2665 10865
rect 2885 10535 3215 10865
rect 3435 10535 3765 10865
rect 3985 10535 4315 10865
rect 4535 10535 4865 10865
rect 5085 10535 5415 10865
rect 5635 10535 5965 10865
rect 6185 10535 6515 10865
rect 6735 10535 7065 10865
rect 7285 10535 7615 10865
rect 7835 10535 8165 10865
rect 8385 10535 8715 10865
rect 8935 10535 9265 10865
rect 9485 10535 9815 10865
rect 10035 10535 10365 10865
rect 10585 10535 10915 10865
rect 11135 10535 11465 10865
rect 11685 10535 12015 10865
rect 12235 10535 12565 10865
rect 12785 10535 13115 10865
rect 13335 10535 13665 10865
rect -542 10408 -508 10442
rect 8 10408 42 10442
rect 558 10408 592 10442
rect 1108 10408 1142 10442
rect 1658 10408 1692 10442
rect 2208 10408 2242 10442
rect 2758 10408 2792 10442
rect 3308 10408 3342 10442
rect 3858 10408 3892 10442
rect 4408 10408 4442 10442
rect 4958 10408 4992 10442
rect 5508 10408 5542 10442
rect 6058 10408 6092 10442
rect 6608 10408 6642 10442
rect 7158 10408 7192 10442
rect 7708 10408 7742 10442
rect 8258 10408 8292 10442
rect 8808 10408 8842 10442
rect 9358 10408 9392 10442
rect 9908 10408 9942 10442
rect 10458 10408 10492 10442
rect 11008 10408 11042 10442
rect 11558 10408 11592 10442
rect 12108 10408 12142 10442
rect 12658 10408 12692 10442
rect 13208 10408 13242 10442
rect 13758 10408 13792 10442
rect -415 9985 -85 10315
rect 135 9985 465 10315
rect 685 9985 1015 10315
rect 1235 9985 1565 10315
rect 1785 9985 2115 10315
rect 2335 9985 2665 10315
rect 2885 9985 3215 10315
rect 3435 9985 3765 10315
rect 3985 9985 4315 10315
rect 4535 9985 4865 10315
rect 5085 9985 5415 10315
rect 5635 9985 5965 10315
rect 6185 9985 6515 10315
rect 6735 9985 7065 10315
rect 7285 9985 7615 10315
rect 7835 9985 8165 10315
rect 8385 9985 8715 10315
rect 8935 9985 9265 10315
rect 9485 9985 9815 10315
rect 10035 9985 10365 10315
rect 10585 9985 10915 10315
rect 11135 9985 11465 10315
rect 11685 9985 12015 10315
rect 12235 9985 12565 10315
rect 12785 9985 13115 10315
rect 13335 9985 13665 10315
rect 14075 9938 14175 10038
rect -925 9712 -825 9812
rect -542 9858 -508 9892
rect 8 9858 42 9892
rect 558 9858 592 9892
rect 1108 9858 1142 9892
rect 1658 9858 1692 9892
rect 2208 9858 2242 9892
rect 2758 9858 2792 9892
rect 3308 9858 3342 9892
rect 3858 9858 3892 9892
rect 4408 9858 4442 9892
rect 4958 9858 4992 9892
rect 5508 9858 5542 9892
rect 6058 9858 6092 9892
rect 6608 9858 6642 9892
rect 7158 9858 7192 9892
rect 7708 9858 7742 9892
rect 8258 9858 8292 9892
rect 8808 9858 8842 9892
rect 9358 9858 9392 9892
rect 9908 9858 9942 9892
rect 10458 9858 10492 9892
rect 11008 9858 11042 9892
rect 11558 9858 11592 9892
rect 12108 9858 12142 9892
rect 12658 9858 12692 9892
rect 13208 9858 13242 9892
rect 13758 9858 13792 9892
rect -415 9435 -85 9765
rect 135 9435 465 9765
rect 685 9435 1015 9765
rect 1235 9435 1565 9765
rect 1785 9435 2115 9765
rect 2335 9435 2665 9765
rect 2885 9435 3215 9765
rect 3435 9435 3765 9765
rect 3985 9435 4315 9765
rect 4535 9435 4865 9765
rect 5085 9435 5415 9765
rect 5635 9435 5965 9765
rect 6185 9435 6515 9765
rect 6735 9435 7065 9765
rect 7285 9435 7615 9765
rect 7835 9435 8165 9765
rect 8385 9435 8715 9765
rect 8935 9435 9265 9765
rect 9485 9435 9815 9765
rect 10035 9435 10365 9765
rect 10585 9435 10915 9765
rect 11135 9435 11465 9765
rect 11685 9435 12015 9765
rect 12235 9435 12565 9765
rect 12785 9435 13115 9765
rect 13335 9435 13665 9765
rect -542 9308 -508 9342
rect 8 9308 42 9342
rect 558 9308 592 9342
rect 1108 9308 1142 9342
rect 1658 9308 1692 9342
rect 2208 9308 2242 9342
rect 2758 9308 2792 9342
rect 3308 9308 3342 9342
rect 3858 9308 3892 9342
rect 4408 9308 4442 9342
rect 4958 9308 4992 9342
rect 5508 9308 5542 9342
rect 6058 9308 6092 9342
rect 6608 9308 6642 9342
rect 7158 9308 7192 9342
rect 7708 9308 7742 9342
rect 8258 9308 8292 9342
rect 8808 9308 8842 9342
rect 9358 9308 9392 9342
rect 9908 9308 9942 9342
rect 10458 9308 10492 9342
rect 11008 9308 11042 9342
rect 11558 9308 11592 9342
rect 12108 9308 12142 9342
rect 12658 9308 12692 9342
rect 13208 9308 13242 9342
rect 13758 9308 13792 9342
rect -415 8885 -85 9215
rect 135 8885 465 9215
rect 685 8885 1015 9215
rect 1235 8885 1565 9215
rect 1785 8885 2115 9215
rect 2335 8885 2665 9215
rect 2885 8885 3215 9215
rect 3435 8885 3765 9215
rect 3985 8885 4315 9215
rect 4535 8885 4865 9215
rect 5085 8885 5415 9215
rect 5635 8885 5965 9215
rect 6185 8885 6515 9215
rect 6735 8885 7065 9215
rect 7285 8885 7615 9215
rect 7835 8885 8165 9215
rect 8385 8885 8715 9215
rect 8935 8885 9265 9215
rect 9485 8885 9815 9215
rect 10035 8885 10365 9215
rect 10585 8885 10915 9215
rect 11135 8885 11465 9215
rect 11685 8885 12015 9215
rect 12235 8885 12565 9215
rect 12785 8885 13115 9215
rect 13335 8885 13665 9215
rect 14075 8838 14175 8938
rect -925 8612 -825 8712
rect -542 8758 -508 8792
rect 8 8758 42 8792
rect 558 8758 592 8792
rect 1108 8758 1142 8792
rect 1658 8758 1692 8792
rect 2208 8758 2242 8792
rect 2758 8758 2792 8792
rect 3308 8758 3342 8792
rect 3858 8758 3892 8792
rect 4408 8758 4442 8792
rect 4958 8758 4992 8792
rect 5508 8758 5542 8792
rect 6058 8758 6092 8792
rect 6608 8758 6642 8792
rect 7158 8758 7192 8792
rect 7708 8758 7742 8792
rect 8258 8758 8292 8792
rect 8808 8758 8842 8792
rect 9358 8758 9392 8792
rect 9908 8758 9942 8792
rect 10458 8758 10492 8792
rect 11008 8758 11042 8792
rect 11558 8758 11592 8792
rect 12108 8758 12142 8792
rect 12658 8758 12692 8792
rect 13208 8758 13242 8792
rect 13758 8758 13792 8792
rect -415 8335 -85 8665
rect 135 8335 465 8665
rect 685 8335 1015 8665
rect 1235 8335 1565 8665
rect 1785 8335 2115 8665
rect 2335 8335 2665 8665
rect 2885 8335 3215 8665
rect 3435 8335 3765 8665
rect 3985 8335 4315 8665
rect 4535 8335 4865 8665
rect 5085 8335 5415 8665
rect 5635 8335 5965 8665
rect 6185 8335 6515 8665
rect 6735 8335 7065 8665
rect 7285 8335 7615 8665
rect 7835 8335 8165 8665
rect 8385 8335 8715 8665
rect 8935 8335 9265 8665
rect 9485 8335 9815 8665
rect 10035 8335 10365 8665
rect 10585 8335 10915 8665
rect 11135 8335 11465 8665
rect 11685 8335 12015 8665
rect 12235 8335 12565 8665
rect 12785 8335 13115 8665
rect 13335 8335 13665 8665
rect -542 8208 -508 8242
rect 8 8208 42 8242
rect 558 8208 592 8242
rect 1108 8208 1142 8242
rect 1658 8208 1692 8242
rect 2208 8208 2242 8242
rect 2758 8208 2792 8242
rect 3308 8208 3342 8242
rect 3858 8208 3892 8242
rect 4408 8208 4442 8242
rect 4958 8208 4992 8242
rect 5508 8208 5542 8242
rect 6058 8208 6092 8242
rect 6608 8208 6642 8242
rect 7158 8208 7192 8242
rect 7708 8208 7742 8242
rect 8258 8208 8292 8242
rect 8808 8208 8842 8242
rect 9358 8208 9392 8242
rect 9908 8208 9942 8242
rect 10458 8208 10492 8242
rect 11008 8208 11042 8242
rect 11558 8208 11592 8242
rect 12108 8208 12142 8242
rect 12658 8208 12692 8242
rect 13208 8208 13242 8242
rect 13758 8208 13792 8242
rect -415 7785 -85 8115
rect 135 7785 465 8115
rect 685 7785 1015 8115
rect 1235 7785 1565 8115
rect 1785 7785 2115 8115
rect 2335 7785 2665 8115
rect 2885 7785 3215 8115
rect 3435 7785 3765 8115
rect 3985 7785 4315 8115
rect 4535 7785 4865 8115
rect 5085 7785 5415 8115
rect 5635 7785 5965 8115
rect 6185 7785 6515 8115
rect 6735 7785 7065 8115
rect 7285 7785 7615 8115
rect 7835 7785 8165 8115
rect 8385 7785 8715 8115
rect 8935 7785 9265 8115
rect 9485 7785 9815 8115
rect 10035 7785 10365 8115
rect 10585 7785 10915 8115
rect 11135 7785 11465 8115
rect 11685 7785 12015 8115
rect 12235 7785 12565 8115
rect 12785 7785 13115 8115
rect 13335 7785 13665 8115
rect 14075 7738 14175 7838
rect -925 7512 -825 7612
rect -542 7658 -508 7692
rect 8 7658 42 7692
rect 558 7658 592 7692
rect 1108 7658 1142 7692
rect 1658 7658 1692 7692
rect 2208 7658 2242 7692
rect 2758 7658 2792 7692
rect 3308 7658 3342 7692
rect 3858 7658 3892 7692
rect 4408 7658 4442 7692
rect 4958 7658 4992 7692
rect 5508 7658 5542 7692
rect 6058 7658 6092 7692
rect 6608 7658 6642 7692
rect 7158 7658 7192 7692
rect 7708 7658 7742 7692
rect 8258 7658 8292 7692
rect 8808 7658 8842 7692
rect 9358 7658 9392 7692
rect 9908 7658 9942 7692
rect 10458 7658 10492 7692
rect 11008 7658 11042 7692
rect 11558 7658 11592 7692
rect 12108 7658 12142 7692
rect 12658 7658 12692 7692
rect 13208 7658 13242 7692
rect 13758 7658 13792 7692
rect -415 7235 -85 7565
rect 135 7235 465 7565
rect 685 7235 1015 7565
rect 1235 7235 1565 7565
rect 1785 7235 2115 7565
rect 2335 7235 2665 7565
rect 2885 7235 3215 7565
rect 3435 7235 3765 7565
rect 3985 7235 4315 7565
rect 4535 7235 4865 7565
rect 5085 7235 5415 7565
rect 5635 7235 5965 7565
rect 6185 7235 6515 7565
rect 6735 7235 7065 7565
rect 7285 7235 7615 7565
rect 7835 7235 8165 7565
rect 8385 7235 8715 7565
rect 8935 7235 9265 7565
rect 9485 7235 9815 7565
rect 10035 7235 10365 7565
rect 10585 7235 10915 7565
rect 11135 7235 11465 7565
rect 11685 7235 12015 7565
rect 12235 7235 12565 7565
rect 12785 7235 13115 7565
rect 13335 7235 13665 7565
rect -542 7108 -508 7142
rect 8 7108 42 7142
rect 558 7108 592 7142
rect 1108 7108 1142 7142
rect 1658 7108 1692 7142
rect 2208 7108 2242 7142
rect 2758 7108 2792 7142
rect 3308 7108 3342 7142
rect 3858 7108 3892 7142
rect 4408 7108 4442 7142
rect 4958 7108 4992 7142
rect 5508 7108 5542 7142
rect 6058 7108 6092 7142
rect 6608 7108 6642 7142
rect 7158 7108 7192 7142
rect 7708 7108 7742 7142
rect 8258 7108 8292 7142
rect 8808 7108 8842 7142
rect 9358 7108 9392 7142
rect 9908 7108 9942 7142
rect 10458 7108 10492 7142
rect 11008 7108 11042 7142
rect 11558 7108 11592 7142
rect 12108 7108 12142 7142
rect 12658 7108 12692 7142
rect 13208 7108 13242 7142
rect 13758 7108 13792 7142
rect -415 6685 -85 7015
rect 135 6685 465 7015
rect 685 6685 1015 7015
rect 1235 6685 1565 7015
rect 1785 6685 2115 7015
rect 2335 6685 2665 7015
rect 2885 6685 3215 7015
rect 3435 6685 3765 7015
rect 3985 6685 4315 7015
rect 4535 6685 4865 7015
rect 5085 6685 5415 7015
rect 5635 6685 5965 7015
rect 6185 6685 6515 7015
rect 6735 6685 7065 7015
rect 7285 6685 7615 7015
rect 7835 6685 8165 7015
rect 8385 6685 8715 7015
rect 8935 6685 9265 7015
rect 9485 6685 9815 7015
rect 10035 6685 10365 7015
rect 10585 6685 10915 7015
rect 11135 6685 11465 7015
rect 11685 6685 12015 7015
rect 12235 6685 12565 7015
rect 12785 6685 13115 7015
rect 13335 6685 13665 7015
rect 14075 6638 14175 6738
rect -925 6412 -825 6512
rect -542 6558 -508 6592
rect 8 6558 42 6592
rect 558 6558 592 6592
rect 1108 6558 1142 6592
rect 1658 6558 1692 6592
rect 2208 6558 2242 6592
rect 2758 6558 2792 6592
rect 3308 6558 3342 6592
rect 3858 6558 3892 6592
rect 4408 6558 4442 6592
rect 4958 6558 4992 6592
rect 5508 6558 5542 6592
rect 6058 6558 6092 6592
rect 6608 6558 6642 6592
rect 7158 6558 7192 6592
rect 7708 6558 7742 6592
rect 8258 6558 8292 6592
rect 8808 6558 8842 6592
rect 9358 6558 9392 6592
rect 9908 6558 9942 6592
rect 10458 6558 10492 6592
rect 11008 6558 11042 6592
rect 11558 6558 11592 6592
rect 12108 6558 12142 6592
rect 12658 6558 12692 6592
rect 13208 6558 13242 6592
rect 13758 6558 13792 6592
rect -415 6135 -85 6465
rect 135 6135 465 6465
rect 685 6135 1015 6465
rect 1235 6135 1565 6465
rect 1785 6135 2115 6465
rect 2335 6135 2665 6465
rect 2885 6135 3215 6465
rect 3435 6135 3765 6465
rect 3985 6135 4315 6465
rect 4535 6135 4865 6465
rect 5085 6135 5415 6465
rect 5635 6135 5965 6465
rect 6185 6135 6515 6465
rect 6735 6135 7065 6465
rect 7285 6135 7615 6465
rect 7835 6135 8165 6465
rect 8385 6135 8715 6465
rect 8935 6135 9265 6465
rect 9485 6135 9815 6465
rect 10035 6135 10365 6465
rect 10585 6135 10915 6465
rect 11135 6135 11465 6465
rect 11685 6135 12015 6465
rect 12235 6135 12565 6465
rect 12785 6135 13115 6465
rect 13335 6135 13665 6465
rect -542 6008 -508 6042
rect 8 6008 42 6042
rect 558 6008 592 6042
rect 1108 6008 1142 6042
rect 1658 6008 1692 6042
rect 2208 6008 2242 6042
rect 2758 6008 2792 6042
rect 3308 6008 3342 6042
rect 3858 6008 3892 6042
rect 4408 6008 4442 6042
rect 4958 6008 4992 6042
rect 5508 6008 5542 6042
rect 6058 6008 6092 6042
rect 6608 6008 6642 6042
rect 7158 6008 7192 6042
rect 7708 6008 7742 6042
rect 8258 6008 8292 6042
rect 8808 6008 8842 6042
rect 9358 6008 9392 6042
rect 9908 6008 9942 6042
rect 10458 6008 10492 6042
rect 11008 6008 11042 6042
rect 11558 6008 11592 6042
rect 12108 6008 12142 6042
rect 12658 6008 12692 6042
rect 13208 6008 13242 6042
rect 13758 6008 13792 6042
rect -415 5585 -85 5915
rect 135 5585 465 5915
rect 685 5585 1015 5915
rect 1235 5585 1565 5915
rect 1785 5585 2115 5915
rect 2335 5585 2665 5915
rect 2885 5585 3215 5915
rect 3435 5585 3765 5915
rect 3985 5585 4315 5915
rect 4535 5585 4865 5915
rect 5085 5585 5415 5915
rect 5635 5585 5965 5915
rect 6185 5585 6515 5915
rect 6735 5585 7065 5915
rect 7285 5585 7615 5915
rect 7835 5585 8165 5915
rect 8385 5585 8715 5915
rect 8935 5585 9265 5915
rect 9485 5585 9815 5915
rect 10035 5585 10365 5915
rect 10585 5585 10915 5915
rect 11135 5585 11465 5915
rect 11685 5585 12015 5915
rect 12235 5585 12565 5915
rect 12785 5585 13115 5915
rect 13335 5585 13665 5915
rect 14075 5538 14175 5638
rect -925 5312 -825 5412
rect -542 5458 -508 5492
rect 8 5458 42 5492
rect 558 5458 592 5492
rect 1108 5458 1142 5492
rect 1658 5458 1692 5492
rect 2208 5458 2242 5492
rect 2758 5458 2792 5492
rect 3308 5458 3342 5492
rect 3858 5458 3892 5492
rect 4408 5458 4442 5492
rect 4958 5458 4992 5492
rect 5508 5458 5542 5492
rect 6058 5458 6092 5492
rect 6608 5458 6642 5492
rect 7158 5458 7192 5492
rect 7708 5458 7742 5492
rect 8258 5458 8292 5492
rect 8808 5458 8842 5492
rect 9358 5458 9392 5492
rect 9908 5458 9942 5492
rect 10458 5458 10492 5492
rect 11008 5458 11042 5492
rect 11558 5458 11592 5492
rect 12108 5458 12142 5492
rect 12658 5458 12692 5492
rect 13208 5458 13242 5492
rect 13758 5458 13792 5492
rect -415 5035 -85 5365
rect 135 5035 465 5365
rect 685 5035 1015 5365
rect 1235 5035 1565 5365
rect 1785 5035 2115 5365
rect 2335 5035 2665 5365
rect 2885 5035 3215 5365
rect 3435 5035 3765 5365
rect 3985 5035 4315 5365
rect 4535 5035 4865 5365
rect 5085 5035 5415 5365
rect 5635 5035 5965 5365
rect 6185 5035 6515 5365
rect 6735 5035 7065 5365
rect 7285 5035 7615 5365
rect 7835 5035 8165 5365
rect 8385 5035 8715 5365
rect 8935 5035 9265 5365
rect 9485 5035 9815 5365
rect 10035 5035 10365 5365
rect 10585 5035 10915 5365
rect 11135 5035 11465 5365
rect 11685 5035 12015 5365
rect 12235 5035 12565 5365
rect 12785 5035 13115 5365
rect 13335 5035 13665 5365
rect -542 4908 -508 4942
rect 8 4908 42 4942
rect 558 4908 592 4942
rect 1108 4908 1142 4942
rect 1658 4908 1692 4942
rect 2208 4908 2242 4942
rect 2758 4908 2792 4942
rect 3308 4908 3342 4942
rect 3858 4908 3892 4942
rect 4408 4908 4442 4942
rect 4958 4908 4992 4942
rect 5508 4908 5542 4942
rect 6058 4908 6092 4942
rect 6608 4908 6642 4942
rect 7158 4908 7192 4942
rect 7708 4908 7742 4942
rect 8258 4908 8292 4942
rect 8808 4908 8842 4942
rect 9358 4908 9392 4942
rect 9908 4908 9942 4942
rect 10458 4908 10492 4942
rect 11008 4908 11042 4942
rect 11558 4908 11592 4942
rect 12108 4908 12142 4942
rect 12658 4908 12692 4942
rect 13208 4908 13242 4942
rect 13758 4908 13792 4942
rect -415 4485 -85 4815
rect 135 4485 465 4815
rect 685 4485 1015 4815
rect 1235 4485 1565 4815
rect 1785 4485 2115 4815
rect 2335 4485 2665 4815
rect 2885 4485 3215 4815
rect 3435 4485 3765 4815
rect 3985 4485 4315 4815
rect 4535 4485 4865 4815
rect 5085 4485 5415 4815
rect 5635 4485 5965 4815
rect 6185 4485 6515 4815
rect 6735 4485 7065 4815
rect 7285 4485 7615 4815
rect 7835 4485 8165 4815
rect 8385 4485 8715 4815
rect 8935 4485 9265 4815
rect 9485 4485 9815 4815
rect 10035 4485 10365 4815
rect 10585 4485 10915 4815
rect 11135 4485 11465 4815
rect 11685 4485 12015 4815
rect 12235 4485 12565 4815
rect 12785 4485 13115 4815
rect 13335 4485 13665 4815
rect 14075 4438 14175 4538
rect -925 4212 -825 4312
rect -542 4358 -508 4392
rect 8 4358 42 4392
rect 558 4358 592 4392
rect 1108 4358 1142 4392
rect 1658 4358 1692 4392
rect 2208 4358 2242 4392
rect 2758 4358 2792 4392
rect 3308 4358 3342 4392
rect 3858 4358 3892 4392
rect 4408 4358 4442 4392
rect 4958 4358 4992 4392
rect 5508 4358 5542 4392
rect 6058 4358 6092 4392
rect 6608 4358 6642 4392
rect 7158 4358 7192 4392
rect 7708 4358 7742 4392
rect 8258 4358 8292 4392
rect 8808 4358 8842 4392
rect 9358 4358 9392 4392
rect 9908 4358 9942 4392
rect 10458 4358 10492 4392
rect 11008 4358 11042 4392
rect 11558 4358 11592 4392
rect 12108 4358 12142 4392
rect 12658 4358 12692 4392
rect 13208 4358 13242 4392
rect 13758 4358 13792 4392
rect -415 3935 -85 4265
rect 135 3935 465 4265
rect 685 3935 1015 4265
rect 1235 3935 1565 4265
rect 1785 3935 2115 4265
rect 2335 3935 2665 4265
rect 2885 3935 3215 4265
rect 3435 3935 3765 4265
rect 3985 3935 4315 4265
rect 4535 3935 4865 4265
rect 5085 3935 5415 4265
rect 5635 3935 5965 4265
rect 6185 3935 6515 4265
rect 6735 3935 7065 4265
rect 7285 3935 7615 4265
rect 7835 3935 8165 4265
rect 8385 3935 8715 4265
rect 8935 3935 9265 4265
rect 9485 3935 9815 4265
rect 10035 3935 10365 4265
rect 10585 3935 10915 4265
rect 11135 3935 11465 4265
rect 11685 3935 12015 4265
rect 12235 3935 12565 4265
rect 12785 3935 13115 4265
rect 13335 3935 13665 4265
rect -542 3808 -508 3842
rect 8 3808 42 3842
rect 558 3808 592 3842
rect 1108 3808 1142 3842
rect 1658 3808 1692 3842
rect 2208 3808 2242 3842
rect 2758 3808 2792 3842
rect 3308 3808 3342 3842
rect 3858 3808 3892 3842
rect 4408 3808 4442 3842
rect 4958 3808 4992 3842
rect 5508 3808 5542 3842
rect 6058 3808 6092 3842
rect 6608 3808 6642 3842
rect 7158 3808 7192 3842
rect 7708 3808 7742 3842
rect 8258 3808 8292 3842
rect 8808 3808 8842 3842
rect 9358 3808 9392 3842
rect 9908 3808 9942 3842
rect 10458 3808 10492 3842
rect 11008 3808 11042 3842
rect 11558 3808 11592 3842
rect 12108 3808 12142 3842
rect 12658 3808 12692 3842
rect 13208 3808 13242 3842
rect 13758 3808 13792 3842
rect -415 3385 -85 3715
rect 135 3385 465 3715
rect 685 3385 1015 3715
rect 1235 3385 1565 3715
rect 1785 3385 2115 3715
rect 2335 3385 2665 3715
rect 2885 3385 3215 3715
rect 3435 3385 3765 3715
rect 3985 3385 4315 3715
rect 4535 3385 4865 3715
rect 5085 3385 5415 3715
rect 5635 3385 5965 3715
rect 6185 3385 6515 3715
rect 6735 3385 7065 3715
rect 7285 3385 7615 3715
rect 7835 3385 8165 3715
rect 8385 3385 8715 3715
rect 8935 3385 9265 3715
rect 9485 3385 9815 3715
rect 10035 3385 10365 3715
rect 10585 3385 10915 3715
rect 11135 3385 11465 3715
rect 11685 3385 12015 3715
rect 12235 3385 12565 3715
rect 12785 3385 13115 3715
rect 13335 3385 13665 3715
rect 14075 3338 14175 3438
rect -925 3112 -825 3212
rect -542 3258 -508 3292
rect 8 3258 42 3292
rect 558 3258 592 3292
rect 1108 3258 1142 3292
rect 1658 3258 1692 3292
rect 2208 3258 2242 3292
rect 2758 3258 2792 3292
rect 3308 3258 3342 3292
rect 3858 3258 3892 3292
rect 4408 3258 4442 3292
rect 4958 3258 4992 3292
rect 5508 3258 5542 3292
rect 6058 3258 6092 3292
rect 6608 3258 6642 3292
rect 7158 3258 7192 3292
rect 7708 3258 7742 3292
rect 8258 3258 8292 3292
rect 8808 3258 8842 3292
rect 9358 3258 9392 3292
rect 9908 3258 9942 3292
rect 10458 3258 10492 3292
rect 11008 3258 11042 3292
rect 11558 3258 11592 3292
rect 12108 3258 12142 3292
rect 12658 3258 12692 3292
rect 13208 3258 13242 3292
rect 13758 3258 13792 3292
rect -415 2835 -85 3165
rect 135 2835 465 3165
rect 685 2835 1015 3165
rect 1235 2835 1565 3165
rect 1785 2835 2115 3165
rect 2335 2835 2665 3165
rect 2885 2835 3215 3165
rect 3435 2835 3765 3165
rect 3985 2835 4315 3165
rect 4535 2835 4865 3165
rect 5085 2835 5415 3165
rect 5635 2835 5965 3165
rect 6185 2835 6515 3165
rect 6735 2835 7065 3165
rect 7285 2835 7615 3165
rect 7835 2835 8165 3165
rect 8385 2835 8715 3165
rect 8935 2835 9265 3165
rect 9485 2835 9815 3165
rect 10035 2835 10365 3165
rect 10585 2835 10915 3165
rect 11135 2835 11465 3165
rect 11685 2835 12015 3165
rect 12235 2835 12565 3165
rect 12785 2835 13115 3165
rect 13335 2835 13665 3165
rect -542 2708 -508 2742
rect 8 2708 42 2742
rect 558 2708 592 2742
rect 1108 2708 1142 2742
rect 1658 2708 1692 2742
rect 2208 2708 2242 2742
rect 2758 2708 2792 2742
rect 3308 2708 3342 2742
rect 3858 2708 3892 2742
rect 4408 2708 4442 2742
rect 4958 2708 4992 2742
rect 5508 2708 5542 2742
rect 6058 2708 6092 2742
rect 6608 2708 6642 2742
rect 7158 2708 7192 2742
rect 7708 2708 7742 2742
rect 8258 2708 8292 2742
rect 8808 2708 8842 2742
rect 9358 2708 9392 2742
rect 9908 2708 9942 2742
rect 10458 2708 10492 2742
rect 11008 2708 11042 2742
rect 11558 2708 11592 2742
rect 12108 2708 12142 2742
rect 12658 2708 12692 2742
rect 13208 2708 13242 2742
rect 13758 2708 13792 2742
rect -415 2285 -85 2615
rect 135 2285 465 2615
rect 685 2285 1015 2615
rect 1235 2285 1565 2615
rect 1785 2285 2115 2615
rect 2335 2285 2665 2615
rect 2885 2285 3215 2615
rect 3435 2285 3765 2615
rect 3985 2285 4315 2615
rect 4535 2285 4865 2615
rect 5085 2285 5415 2615
rect 5635 2285 5965 2615
rect 6185 2285 6515 2615
rect 6735 2285 7065 2615
rect 7285 2285 7615 2615
rect 7835 2285 8165 2615
rect 8385 2285 8715 2615
rect 8935 2285 9265 2615
rect 9485 2285 9815 2615
rect 10035 2285 10365 2615
rect 10585 2285 10915 2615
rect 11135 2285 11465 2615
rect 11685 2285 12015 2615
rect 12235 2285 12565 2615
rect 12785 2285 13115 2615
rect 13335 2285 13665 2615
rect 14075 2238 14175 2338
rect -925 2012 -825 2112
rect -542 2158 -508 2192
rect 8 2158 42 2192
rect 558 2158 592 2192
rect 1108 2158 1142 2192
rect 1658 2158 1692 2192
rect 2208 2158 2242 2192
rect 2758 2158 2792 2192
rect 3308 2158 3342 2192
rect 3858 2158 3892 2192
rect 4408 2158 4442 2192
rect 4958 2158 4992 2192
rect 5508 2158 5542 2192
rect 6058 2158 6092 2192
rect 6608 2158 6642 2192
rect 7158 2158 7192 2192
rect 7708 2158 7742 2192
rect 8258 2158 8292 2192
rect 8808 2158 8842 2192
rect 9358 2158 9392 2192
rect 9908 2158 9942 2192
rect 10458 2158 10492 2192
rect 11008 2158 11042 2192
rect 11558 2158 11592 2192
rect 12108 2158 12142 2192
rect 12658 2158 12692 2192
rect 13208 2158 13242 2192
rect 13758 2158 13792 2192
rect -415 1735 -85 2065
rect 135 1735 465 2065
rect 685 1735 1015 2065
rect 1235 1735 1565 2065
rect 1785 1735 2115 2065
rect 2335 1735 2665 2065
rect 2885 1735 3215 2065
rect 3435 1735 3765 2065
rect 3985 1735 4315 2065
rect 4535 1735 4865 2065
rect 5085 1735 5415 2065
rect 5635 1735 5965 2065
rect 6185 1735 6515 2065
rect 6735 1735 7065 2065
rect 7285 1735 7615 2065
rect 7835 1735 8165 2065
rect 8385 1735 8715 2065
rect 8935 1735 9265 2065
rect 9485 1735 9815 2065
rect 10035 1735 10365 2065
rect 10585 1735 10915 2065
rect 11135 1735 11465 2065
rect 11685 1735 12015 2065
rect 12235 1735 12565 2065
rect 12785 1735 13115 2065
rect 13335 1735 13665 2065
rect -542 1608 -508 1642
rect 8 1608 42 1642
rect 558 1608 592 1642
rect 1108 1608 1142 1642
rect 1658 1608 1692 1642
rect 2208 1608 2242 1642
rect 2758 1608 2792 1642
rect 3308 1608 3342 1642
rect 3858 1608 3892 1642
rect 4408 1608 4442 1642
rect 4958 1608 4992 1642
rect 5508 1608 5542 1642
rect 6058 1608 6092 1642
rect 6608 1608 6642 1642
rect 7158 1608 7192 1642
rect 7708 1608 7742 1642
rect 8258 1608 8292 1642
rect 8808 1608 8842 1642
rect 9358 1608 9392 1642
rect 9908 1608 9942 1642
rect 10458 1608 10492 1642
rect 11008 1608 11042 1642
rect 11558 1608 11592 1642
rect 12108 1608 12142 1642
rect 12658 1608 12692 1642
rect 13208 1608 13242 1642
rect 13758 1608 13792 1642
rect -415 1185 -85 1515
rect 135 1185 465 1515
rect 685 1185 1015 1515
rect 1235 1185 1565 1515
rect 1785 1185 2115 1515
rect 2335 1185 2665 1515
rect 2885 1185 3215 1515
rect 3435 1185 3765 1515
rect 3985 1185 4315 1515
rect 4535 1185 4865 1515
rect 5085 1185 5415 1515
rect 5635 1185 5965 1515
rect 6185 1185 6515 1515
rect 6735 1185 7065 1515
rect 7285 1185 7615 1515
rect 7835 1185 8165 1515
rect 8385 1185 8715 1515
rect 8935 1185 9265 1515
rect 9485 1185 9815 1515
rect 10035 1185 10365 1515
rect 10585 1185 10915 1515
rect 11135 1185 11465 1515
rect 11685 1185 12015 1515
rect 12235 1185 12565 1515
rect 12785 1185 13115 1515
rect 13335 1185 13665 1515
rect 14075 1138 14175 1238
rect -925 912 -825 1012
rect -542 1058 -508 1092
rect 8 1058 42 1092
rect 558 1058 592 1092
rect 1108 1058 1142 1092
rect 1658 1058 1692 1092
rect 2208 1058 2242 1092
rect 2758 1058 2792 1092
rect 3308 1058 3342 1092
rect 3858 1058 3892 1092
rect 4408 1058 4442 1092
rect 4958 1058 4992 1092
rect 5508 1058 5542 1092
rect 6058 1058 6092 1092
rect 6608 1058 6642 1092
rect 7158 1058 7192 1092
rect 7708 1058 7742 1092
rect 8258 1058 8292 1092
rect 8808 1058 8842 1092
rect 9358 1058 9392 1092
rect 9908 1058 9942 1092
rect 10458 1058 10492 1092
rect 11008 1058 11042 1092
rect 11558 1058 11592 1092
rect 12108 1058 12142 1092
rect 12658 1058 12692 1092
rect 13208 1058 13242 1092
rect 13758 1058 13792 1092
rect -415 635 -85 965
rect 135 635 465 965
rect 685 635 1015 965
rect 1235 635 1565 965
rect 1785 635 2115 965
rect 2335 635 2665 965
rect 2885 635 3215 965
rect 3435 635 3765 965
rect 3985 635 4315 965
rect 4535 635 4865 965
rect 5085 635 5415 965
rect 5635 635 5965 965
rect 6185 635 6515 965
rect 6735 635 7065 965
rect 7285 635 7615 965
rect 7835 635 8165 965
rect 8385 635 8715 965
rect 8935 635 9265 965
rect 9485 635 9815 965
rect 10035 635 10365 965
rect 10585 635 10915 965
rect 11135 635 11465 965
rect 11685 635 12015 965
rect 12235 635 12565 965
rect 12785 635 13115 965
rect 13335 635 13665 965
rect -542 508 -508 542
rect 8 508 42 542
rect 558 508 592 542
rect 1108 508 1142 542
rect 1658 508 1692 542
rect 2208 508 2242 542
rect 2758 508 2792 542
rect 3308 508 3342 542
rect 3858 508 3892 542
rect 4408 508 4442 542
rect 4958 508 4992 542
rect 5508 508 5542 542
rect 6058 508 6092 542
rect 6608 508 6642 542
rect 7158 508 7192 542
rect 7708 508 7742 542
rect 8258 508 8292 542
rect 8808 508 8842 542
rect 9358 508 9392 542
rect 9908 508 9942 542
rect 10458 508 10492 542
rect 11008 508 11042 542
rect 11558 508 11592 542
rect 12108 508 12142 542
rect 12658 508 12692 542
rect 13208 508 13242 542
rect 13758 508 13792 542
rect -415 85 -85 415
rect 135 85 465 415
rect 685 85 1015 415
rect 1235 85 1565 415
rect 1785 85 2115 415
rect 2335 85 2665 415
rect 2885 85 3215 415
rect 3435 85 3765 415
rect 3985 85 4315 415
rect 4535 85 4865 415
rect 5085 85 5415 415
rect 5635 85 5965 415
rect 6185 85 6515 415
rect 6735 85 7065 415
rect 7285 85 7615 415
rect 7835 85 8165 415
rect 8385 85 8715 415
rect 8935 85 9265 415
rect 9485 85 9815 415
rect 10035 85 10365 415
rect 10585 85 10915 415
rect 11135 85 11465 415
rect 11685 85 12015 415
rect 12235 85 12565 415
rect 12785 85 13115 415
rect 13335 85 13665 415
rect 14075 38 14175 138
rect -925 -188 -825 -88
rect -542 -42 -508 -8
rect 8 -42 42 -8
rect 558 -42 592 -8
rect 1108 -42 1142 -8
rect 1658 -42 1692 -8
rect 2208 -42 2242 -8
rect 2758 -42 2792 -8
rect 3308 -42 3342 -8
rect 3858 -42 3892 -8
rect 4408 -42 4442 -8
rect 4958 -42 4992 -8
rect 5508 -42 5542 -8
rect 6058 -42 6092 -8
rect 6608 -42 6642 -8
rect 7158 -42 7192 -8
rect 7708 -42 7742 -8
rect 8258 -42 8292 -8
rect 8808 -42 8842 -8
rect 9358 -42 9392 -8
rect 9908 -42 9942 -8
rect 10458 -42 10492 -8
rect 11008 -42 11042 -8
rect 11558 -42 11592 -8
rect 12108 -42 12142 -8
rect 12658 -42 12692 -8
rect 13208 -42 13242 -8
rect 13758 -42 13792 -8
rect -415 -465 -85 -135
rect 135 -465 465 -135
rect 685 -465 1015 -135
rect 1235 -465 1565 -135
rect 1785 -465 2115 -135
rect 2335 -465 2665 -135
rect 2885 -465 3215 -135
rect 3435 -465 3765 -135
rect 3985 -465 4315 -135
rect 4535 -465 4865 -135
rect 5085 -465 5415 -135
rect 5635 -465 5965 -135
rect 6185 -465 6515 -135
rect 6735 -465 7065 -135
rect 7285 -465 7615 -135
rect 7835 -465 8165 -135
rect 8385 -465 8715 -135
rect 8935 -465 9265 -135
rect 9485 -465 9815 -135
rect 10035 -465 10365 -135
rect 10585 -465 10915 -135
rect 11135 -465 11465 -135
rect 11685 -465 12015 -135
rect 12235 -465 12565 -135
rect 12785 -465 13115 -135
rect 13335 -465 13665 -135
rect -542 -592 -508 -558
rect 8 -592 42 -558
rect 558 -592 592 -558
rect 1108 -592 1142 -558
rect 1658 -592 1692 -558
rect 2208 -592 2242 -558
rect 2758 -592 2792 -558
rect 3308 -592 3342 -558
rect 3858 -592 3892 -558
rect 4408 -592 4442 -558
rect 4958 -592 4992 -558
rect 5508 -592 5542 -558
rect 6058 -592 6092 -558
rect 6608 -592 6642 -558
rect 7158 -592 7192 -558
rect 7708 -592 7742 -558
rect 8258 -592 8292 -558
rect 8808 -592 8842 -558
rect 9358 -592 9392 -558
rect 9908 -592 9942 -558
rect 10458 -592 10492 -558
rect 11008 -592 11042 -558
rect 11558 -592 11592 -558
rect 12108 -592 12142 -558
rect 12658 -592 12692 -558
rect 13208 -592 13242 -558
rect 13758 -592 13792 -558
rect -138 -975 -38 -875
rect 962 -975 1062 -875
rect 2062 -975 2162 -875
rect 3162 -975 3262 -875
rect 4262 -975 4362 -875
rect 5362 -975 5462 -875
rect 6462 -975 6562 -875
rect 7562 -975 7662 -875
rect 8662 -975 8762 -875
rect 9762 -975 9862 -875
rect 10862 -975 10962 -875
rect 11962 -975 12062 -875
rect 13062 -975 13162 -875
rect 14787 -1587 18763 14737
rect -495 -5563 18763 -1587
<< metal2 >>
rect -5525 18713 18775 18725
rect -5525 14737 -5513 18713
rect -5525 14725 14787 14737
rect -5525 1117 -5513 14725
rect -1537 1117 -1525 14725
rect 78 14125 198 14135
rect 78 14025 88 14125
rect 188 14025 198 14125
rect 78 14015 198 14025
rect 1178 14125 1298 14135
rect 1178 14025 1188 14125
rect 1288 14025 1298 14125
rect 1178 14015 1298 14025
rect 2278 14125 2398 14135
rect 2278 14025 2288 14125
rect 2388 14025 2398 14125
rect 2278 14015 2398 14025
rect 3378 14125 3498 14135
rect 3378 14025 3388 14125
rect 3488 14025 3498 14125
rect 3378 14015 3498 14025
rect 4478 14125 4598 14135
rect 4478 14025 4488 14125
rect 4588 14025 4598 14125
rect 4478 14015 4598 14025
rect 5578 14125 5698 14135
rect 5578 14025 5588 14125
rect 5688 14025 5698 14125
rect 5578 14015 5698 14025
rect 6678 14125 6798 14135
rect 6678 14025 6688 14125
rect 6788 14025 6798 14125
rect 6678 14015 6798 14025
rect 7778 14125 7898 14135
rect 7778 14025 7788 14125
rect 7888 14025 7898 14125
rect 7778 14015 7898 14025
rect 8878 14125 8998 14135
rect 8878 14025 8888 14125
rect 8988 14025 8998 14125
rect 8878 14015 8998 14025
rect 9978 14125 10098 14135
rect 9978 14025 9988 14125
rect 10088 14025 10098 14125
rect 9978 14015 10098 14025
rect 11078 14125 11198 14135
rect 11078 14025 11088 14125
rect 11188 14025 11198 14125
rect 11078 14015 11198 14025
rect 12178 14125 12298 14135
rect 12178 14025 12188 14125
rect 12288 14025 12298 14125
rect 12178 14015 12298 14025
rect 13278 14125 13398 14135
rect 13278 14025 13288 14125
rect 13388 14025 13398 14125
rect 13278 14015 13398 14025
rect -725 13742 13975 13925
rect -725 13708 -542 13742
rect -508 13708 8 13742
rect 42 13708 558 13742
rect 592 13708 1108 13742
rect 1142 13708 1658 13742
rect 1692 13708 2208 13742
rect 2242 13708 2758 13742
rect 2792 13708 3308 13742
rect 3342 13708 3858 13742
rect 3892 13708 4408 13742
rect 4442 13708 4958 13742
rect 4992 13708 5508 13742
rect 5542 13708 6058 13742
rect 6092 13708 6608 13742
rect 6642 13708 7158 13742
rect 7192 13708 7708 13742
rect 7742 13708 8258 13742
rect 8292 13708 8808 13742
rect 8842 13708 9358 13742
rect 9392 13708 9908 13742
rect 9942 13708 10458 13742
rect 10492 13708 11008 13742
rect 11042 13708 11558 13742
rect 11592 13708 12108 13742
rect 12142 13708 12658 13742
rect 12692 13708 13208 13742
rect 13242 13708 13758 13742
rect 13792 13708 13975 13742
rect -725 13700 13975 13708
rect -725 13200 -500 13700
rect -425 13615 -75 13625
rect -425 13285 -415 13615
rect -85 13285 -75 13615
rect -425 13275 -75 13285
rect 0 13200 50 13700
rect 125 13615 475 13625
rect 125 13285 135 13615
rect 465 13285 475 13615
rect 125 13275 475 13285
rect 550 13200 600 13700
rect 675 13615 1025 13625
rect 675 13285 685 13615
rect 1015 13285 1025 13615
rect 675 13275 1025 13285
rect 1100 13200 1150 13700
rect 1225 13615 1575 13625
rect 1225 13285 1235 13615
rect 1565 13285 1575 13615
rect 1225 13275 1575 13285
rect 1650 13200 1700 13700
rect 1775 13615 2125 13625
rect 1775 13285 1785 13615
rect 2115 13285 2125 13615
rect 1775 13275 2125 13285
rect 2200 13200 2250 13700
rect 2325 13615 2675 13625
rect 2325 13285 2335 13615
rect 2665 13285 2675 13615
rect 2325 13275 2675 13285
rect 2750 13200 2800 13700
rect 2875 13615 3225 13625
rect 2875 13285 2885 13615
rect 3215 13285 3225 13615
rect 2875 13275 3225 13285
rect 3300 13200 3350 13700
rect 3425 13615 3775 13625
rect 3425 13285 3435 13615
rect 3765 13285 3775 13615
rect 3425 13275 3775 13285
rect 3850 13200 3900 13700
rect 3975 13615 4325 13625
rect 3975 13285 3985 13615
rect 4315 13285 4325 13615
rect 3975 13275 4325 13285
rect 4400 13200 4450 13700
rect 4525 13615 4875 13625
rect 4525 13285 4535 13615
rect 4865 13285 4875 13615
rect 4525 13275 4875 13285
rect 4950 13200 5000 13700
rect 5075 13615 5425 13625
rect 5075 13285 5085 13615
rect 5415 13285 5425 13615
rect 5075 13275 5425 13285
rect 5500 13200 5550 13700
rect 5625 13615 5975 13625
rect 5625 13285 5635 13615
rect 5965 13285 5975 13615
rect 5625 13275 5975 13285
rect 6050 13200 6100 13700
rect 6175 13615 6525 13625
rect 6175 13285 6185 13615
rect 6515 13285 6525 13615
rect 6175 13275 6525 13285
rect 6600 13200 6650 13700
rect 6725 13615 7075 13625
rect 6725 13285 6735 13615
rect 7065 13285 7075 13615
rect 6725 13275 7075 13285
rect 7150 13200 7200 13700
rect 7275 13615 7625 13625
rect 7275 13285 7285 13615
rect 7615 13285 7625 13615
rect 7275 13275 7625 13285
rect 7700 13200 7750 13700
rect 7825 13615 8175 13625
rect 7825 13285 7835 13615
rect 8165 13285 8175 13615
rect 7825 13275 8175 13285
rect 8250 13200 8300 13700
rect 8375 13615 8725 13625
rect 8375 13285 8385 13615
rect 8715 13285 8725 13615
rect 8375 13275 8725 13285
rect 8800 13200 8850 13700
rect 8925 13615 9275 13625
rect 8925 13285 8935 13615
rect 9265 13285 9275 13615
rect 8925 13275 9275 13285
rect 9350 13200 9400 13700
rect 9475 13615 9825 13625
rect 9475 13285 9485 13615
rect 9815 13285 9825 13615
rect 9475 13275 9825 13285
rect 9900 13200 9950 13700
rect 10025 13615 10375 13625
rect 10025 13285 10035 13615
rect 10365 13285 10375 13615
rect 10025 13275 10375 13285
rect 10450 13200 10500 13700
rect 10575 13615 10925 13625
rect 10575 13285 10585 13615
rect 10915 13285 10925 13615
rect 10575 13275 10925 13285
rect 11000 13200 11050 13700
rect 11125 13615 11475 13625
rect 11125 13285 11135 13615
rect 11465 13285 11475 13615
rect 11125 13275 11475 13285
rect 11550 13200 11600 13700
rect 11675 13615 12025 13625
rect 11675 13285 11685 13615
rect 12015 13285 12025 13615
rect 11675 13275 12025 13285
rect 12100 13200 12150 13700
rect 12225 13615 12575 13625
rect 12225 13285 12235 13615
rect 12565 13285 12575 13615
rect 12225 13275 12575 13285
rect 12650 13200 12700 13700
rect 12775 13615 13125 13625
rect 12775 13285 12785 13615
rect 13115 13285 13125 13615
rect 12775 13275 13125 13285
rect 13200 13200 13250 13700
rect 13325 13615 13675 13625
rect 13325 13285 13335 13615
rect 13665 13285 13675 13615
rect 13325 13275 13675 13285
rect 13750 13200 13975 13700
rect 14065 13338 14185 13348
rect 14065 13238 14075 13338
rect 14175 13238 14185 13338
rect 14065 13228 14185 13238
rect -725 13192 13975 13200
rect -725 13158 -542 13192
rect -508 13158 8 13192
rect 42 13158 558 13192
rect 592 13158 1108 13192
rect 1142 13158 1658 13192
rect 1692 13158 2208 13192
rect 2242 13158 2758 13192
rect 2792 13158 3308 13192
rect 3342 13158 3858 13192
rect 3892 13158 4408 13192
rect 4442 13158 4958 13192
rect 4992 13158 5508 13192
rect 5542 13158 6058 13192
rect 6092 13158 6608 13192
rect 6642 13158 7158 13192
rect 7192 13158 7708 13192
rect 7742 13158 8258 13192
rect 8292 13158 8808 13192
rect 8842 13158 9358 13192
rect 9392 13158 9908 13192
rect 9942 13158 10458 13192
rect 10492 13158 11008 13192
rect 11042 13158 11558 13192
rect 11592 13158 12108 13192
rect 12142 13158 12658 13192
rect 12692 13158 13208 13192
rect 13242 13158 13758 13192
rect 13792 13158 13975 13192
rect -725 13150 13975 13158
rect -935 13112 -815 13122
rect -935 13012 -925 13112
rect -825 13012 -815 13112
rect -935 13002 -815 13012
rect -725 12650 -500 13150
rect -425 13065 -75 13075
rect -425 12735 -415 13065
rect -85 12735 -75 13065
rect -425 12725 -75 12735
rect 0 12650 50 13150
rect 125 13065 475 13075
rect 125 12735 135 13065
rect 465 12735 475 13065
rect 125 12725 475 12735
rect 550 12650 600 13150
rect 675 13065 1025 13075
rect 675 12735 685 13065
rect 1015 12735 1025 13065
rect 675 12725 1025 12735
rect 1100 12650 1150 13150
rect 1225 13065 1575 13075
rect 1225 12735 1235 13065
rect 1565 12735 1575 13065
rect 1225 12725 1575 12735
rect 1650 12650 1700 13150
rect 1775 13065 2125 13075
rect 1775 12735 1785 13065
rect 2115 12735 2125 13065
rect 1775 12725 2125 12735
rect 2200 12650 2250 13150
rect 2325 13065 2675 13075
rect 2325 12735 2335 13065
rect 2665 12735 2675 13065
rect 2325 12725 2675 12735
rect 2750 12650 2800 13150
rect 2875 13065 3225 13075
rect 2875 12735 2885 13065
rect 3215 12735 3225 13065
rect 2875 12725 3225 12735
rect 3300 12650 3350 13150
rect 3425 13065 3775 13075
rect 3425 12735 3435 13065
rect 3765 12735 3775 13065
rect 3425 12725 3775 12735
rect 3850 12650 3900 13150
rect 3975 13065 4325 13075
rect 3975 12735 3985 13065
rect 4315 12735 4325 13065
rect 3975 12725 4325 12735
rect 4400 12650 4450 13150
rect 4525 13065 4875 13075
rect 4525 12735 4535 13065
rect 4865 12735 4875 13065
rect 4525 12725 4875 12735
rect 4950 12650 5000 13150
rect 5075 13065 5425 13075
rect 5075 12735 5085 13065
rect 5415 12735 5425 13065
rect 5075 12725 5425 12735
rect 5500 12650 5550 13150
rect 5625 13065 5975 13075
rect 5625 12735 5635 13065
rect 5965 12735 5975 13065
rect 5625 12725 5975 12735
rect 6050 12650 6100 13150
rect 6175 13065 6525 13075
rect 6175 12735 6185 13065
rect 6515 12735 6525 13065
rect 6175 12725 6525 12735
rect 6600 12650 6650 13150
rect 6725 13065 7075 13075
rect 6725 12735 6735 13065
rect 7065 12735 7075 13065
rect 6725 12725 7075 12735
rect 7150 12650 7200 13150
rect 7275 13065 7625 13075
rect 7275 12735 7285 13065
rect 7615 12735 7625 13065
rect 7275 12725 7625 12735
rect 7700 12650 7750 13150
rect 7825 13065 8175 13075
rect 7825 12735 7835 13065
rect 8165 12735 8175 13065
rect 7825 12725 8175 12735
rect 8250 12650 8300 13150
rect 8375 13065 8725 13075
rect 8375 12735 8385 13065
rect 8715 12735 8725 13065
rect 8375 12725 8725 12735
rect 8800 12650 8850 13150
rect 8925 13065 9275 13075
rect 8925 12735 8935 13065
rect 9265 12735 9275 13065
rect 8925 12725 9275 12735
rect 9350 12650 9400 13150
rect 9475 13065 9825 13075
rect 9475 12735 9485 13065
rect 9815 12735 9825 13065
rect 9475 12725 9825 12735
rect 9900 12650 9950 13150
rect 10025 13065 10375 13075
rect 10025 12735 10035 13065
rect 10365 12735 10375 13065
rect 10025 12725 10375 12735
rect 10450 12650 10500 13150
rect 10575 13065 10925 13075
rect 10575 12735 10585 13065
rect 10915 12735 10925 13065
rect 10575 12725 10925 12735
rect 11000 12650 11050 13150
rect 11125 13065 11475 13075
rect 11125 12735 11135 13065
rect 11465 12735 11475 13065
rect 11125 12725 11475 12735
rect 11550 12650 11600 13150
rect 11675 13065 12025 13075
rect 11675 12735 11685 13065
rect 12015 12735 12025 13065
rect 11675 12725 12025 12735
rect 12100 12650 12150 13150
rect 12225 13065 12575 13075
rect 12225 12735 12235 13065
rect 12565 12735 12575 13065
rect 12225 12725 12575 12735
rect 12650 12650 12700 13150
rect 12775 13065 13125 13075
rect 12775 12735 12785 13065
rect 13115 12735 13125 13065
rect 12775 12725 13125 12735
rect 13200 12650 13250 13150
rect 13325 13065 13675 13075
rect 13325 12735 13335 13065
rect 13665 12735 13675 13065
rect 13325 12725 13675 12735
rect 13750 12650 13975 13150
rect -725 12642 13975 12650
rect -725 12608 -542 12642
rect -508 12608 8 12642
rect 42 12608 558 12642
rect 592 12608 1108 12642
rect 1142 12608 1658 12642
rect 1692 12608 2208 12642
rect 2242 12608 2758 12642
rect 2792 12608 3308 12642
rect 3342 12608 3858 12642
rect 3892 12608 4408 12642
rect 4442 12608 4958 12642
rect 4992 12608 5508 12642
rect 5542 12608 6058 12642
rect 6092 12608 6608 12642
rect 6642 12608 7158 12642
rect 7192 12608 7708 12642
rect 7742 12608 8258 12642
rect 8292 12608 8808 12642
rect 8842 12608 9358 12642
rect 9392 12608 9908 12642
rect 9942 12608 10458 12642
rect 10492 12608 11008 12642
rect 11042 12608 11558 12642
rect 11592 12608 12108 12642
rect 12142 12608 12658 12642
rect 12692 12608 13208 12642
rect 13242 12608 13758 12642
rect 13792 12608 13975 12642
rect -725 12600 13975 12608
rect -725 12100 -500 12600
rect -425 12515 -75 12525
rect -425 12185 -415 12515
rect -85 12185 -75 12515
rect -425 12175 -75 12185
rect 0 12100 50 12600
rect 125 12515 475 12525
rect 125 12185 135 12515
rect 465 12185 475 12515
rect 125 12175 475 12185
rect 550 12100 600 12600
rect 675 12515 1025 12525
rect 675 12185 685 12515
rect 1015 12185 1025 12515
rect 675 12175 1025 12185
rect 1100 12100 1150 12600
rect 1225 12515 1575 12525
rect 1225 12185 1235 12515
rect 1565 12185 1575 12515
rect 1225 12175 1575 12185
rect 1650 12100 1700 12600
rect 1775 12515 2125 12525
rect 1775 12185 1785 12515
rect 2115 12185 2125 12515
rect 1775 12175 2125 12185
rect 2200 12100 2250 12600
rect 2325 12515 2675 12525
rect 2325 12185 2335 12515
rect 2665 12185 2675 12515
rect 2325 12175 2675 12185
rect 2750 12100 2800 12600
rect 2875 12515 3225 12525
rect 2875 12185 2885 12515
rect 3215 12185 3225 12515
rect 2875 12175 3225 12185
rect 3300 12100 3350 12600
rect 3425 12515 3775 12525
rect 3425 12185 3435 12515
rect 3765 12185 3775 12515
rect 3425 12175 3775 12185
rect 3850 12100 3900 12600
rect 3975 12515 4325 12525
rect 3975 12185 3985 12515
rect 4315 12185 4325 12515
rect 3975 12175 4325 12185
rect 4400 12100 4450 12600
rect 4525 12515 4875 12525
rect 4525 12185 4535 12515
rect 4865 12185 4875 12515
rect 4525 12175 4875 12185
rect 4950 12100 5000 12600
rect 5075 12515 5425 12525
rect 5075 12185 5085 12515
rect 5415 12185 5425 12515
rect 5075 12175 5425 12185
rect 5500 12100 5550 12600
rect 5625 12515 5975 12525
rect 5625 12185 5635 12515
rect 5965 12185 5975 12515
rect 5625 12175 5975 12185
rect 6050 12100 6100 12600
rect 6175 12515 6525 12525
rect 6175 12185 6185 12515
rect 6515 12185 6525 12515
rect 6175 12175 6525 12185
rect 6600 12100 6650 12600
rect 6725 12515 7075 12525
rect 6725 12185 6735 12515
rect 7065 12185 7075 12515
rect 6725 12175 7075 12185
rect 7150 12100 7200 12600
rect 7275 12515 7625 12525
rect 7275 12185 7285 12515
rect 7615 12185 7625 12515
rect 7275 12175 7625 12185
rect 7700 12100 7750 12600
rect 7825 12515 8175 12525
rect 7825 12185 7835 12515
rect 8165 12185 8175 12515
rect 7825 12175 8175 12185
rect 8250 12100 8300 12600
rect 8375 12515 8725 12525
rect 8375 12185 8385 12515
rect 8715 12185 8725 12515
rect 8375 12175 8725 12185
rect 8800 12100 8850 12600
rect 8925 12515 9275 12525
rect 8925 12185 8935 12515
rect 9265 12185 9275 12515
rect 8925 12175 9275 12185
rect 9350 12100 9400 12600
rect 9475 12515 9825 12525
rect 9475 12185 9485 12515
rect 9815 12185 9825 12515
rect 9475 12175 9825 12185
rect 9900 12100 9950 12600
rect 10025 12515 10375 12525
rect 10025 12185 10035 12515
rect 10365 12185 10375 12515
rect 10025 12175 10375 12185
rect 10450 12100 10500 12600
rect 10575 12515 10925 12525
rect 10575 12185 10585 12515
rect 10915 12185 10925 12515
rect 10575 12175 10925 12185
rect 11000 12100 11050 12600
rect 11125 12515 11475 12525
rect 11125 12185 11135 12515
rect 11465 12185 11475 12515
rect 11125 12175 11475 12185
rect 11550 12100 11600 12600
rect 11675 12515 12025 12525
rect 11675 12185 11685 12515
rect 12015 12185 12025 12515
rect 11675 12175 12025 12185
rect 12100 12100 12150 12600
rect 12225 12515 12575 12525
rect 12225 12185 12235 12515
rect 12565 12185 12575 12515
rect 12225 12175 12575 12185
rect 12650 12100 12700 12600
rect 12775 12515 13125 12525
rect 12775 12185 12785 12515
rect 13115 12185 13125 12515
rect 12775 12175 13125 12185
rect 13200 12100 13250 12600
rect 13325 12515 13675 12525
rect 13325 12185 13335 12515
rect 13665 12185 13675 12515
rect 13325 12175 13675 12185
rect 13750 12100 13975 12600
rect 14065 12238 14185 12248
rect 14065 12138 14075 12238
rect 14175 12138 14185 12238
rect 14065 12128 14185 12138
rect -725 12092 13975 12100
rect -725 12058 -542 12092
rect -508 12058 8 12092
rect 42 12058 558 12092
rect 592 12058 1108 12092
rect 1142 12058 1658 12092
rect 1692 12058 2208 12092
rect 2242 12058 2758 12092
rect 2792 12058 3308 12092
rect 3342 12058 3858 12092
rect 3892 12058 4408 12092
rect 4442 12058 4958 12092
rect 4992 12058 5508 12092
rect 5542 12058 6058 12092
rect 6092 12058 6608 12092
rect 6642 12058 7158 12092
rect 7192 12058 7708 12092
rect 7742 12058 8258 12092
rect 8292 12058 8808 12092
rect 8842 12058 9358 12092
rect 9392 12058 9908 12092
rect 9942 12058 10458 12092
rect 10492 12058 11008 12092
rect 11042 12058 11558 12092
rect 11592 12058 12108 12092
rect 12142 12058 12658 12092
rect 12692 12058 13208 12092
rect 13242 12058 13758 12092
rect 13792 12058 13975 12092
rect -725 12050 13975 12058
rect -935 12012 -815 12022
rect -935 11912 -925 12012
rect -825 11912 -815 12012
rect -935 11902 -815 11912
rect -725 11550 -500 12050
rect -425 11965 -75 11975
rect -425 11635 -415 11965
rect -85 11635 -75 11965
rect -425 11625 -75 11635
rect 0 11550 50 12050
rect 125 11965 475 11975
rect 125 11635 135 11965
rect 465 11635 475 11965
rect 125 11625 475 11635
rect 550 11550 600 12050
rect 675 11965 1025 11975
rect 675 11635 685 11965
rect 1015 11635 1025 11965
rect 675 11625 1025 11635
rect 1100 11550 1150 12050
rect 1225 11965 1575 11975
rect 1225 11635 1235 11965
rect 1565 11635 1575 11965
rect 1225 11625 1575 11635
rect 1650 11550 1700 12050
rect 1775 11965 2125 11975
rect 1775 11635 1785 11965
rect 2115 11635 2125 11965
rect 1775 11625 2125 11635
rect 2200 11550 2250 12050
rect 2325 11965 2675 11975
rect 2325 11635 2335 11965
rect 2665 11635 2675 11965
rect 2325 11625 2675 11635
rect 2750 11550 2800 12050
rect 2875 11965 3225 11975
rect 2875 11635 2885 11965
rect 3215 11635 3225 11965
rect 2875 11625 3225 11635
rect 3300 11550 3350 12050
rect 3425 11965 3775 11975
rect 3425 11635 3435 11965
rect 3765 11635 3775 11965
rect 3425 11625 3775 11635
rect 3850 11550 3900 12050
rect 3975 11965 4325 11975
rect 3975 11635 3985 11965
rect 4315 11635 4325 11965
rect 3975 11625 4325 11635
rect 4400 11550 4450 12050
rect 4525 11965 4875 11975
rect 4525 11635 4535 11965
rect 4865 11635 4875 11965
rect 4525 11625 4875 11635
rect 4950 11550 5000 12050
rect 5075 11965 5425 11975
rect 5075 11635 5085 11965
rect 5415 11635 5425 11965
rect 5075 11625 5425 11635
rect 5500 11550 5550 12050
rect 5625 11965 5975 11975
rect 5625 11635 5635 11965
rect 5965 11635 5975 11965
rect 5625 11625 5975 11635
rect 6050 11550 6100 12050
rect 6175 11965 6525 11975
rect 6175 11635 6185 11965
rect 6515 11635 6525 11965
rect 6175 11625 6525 11635
rect 6600 11550 6650 12050
rect 6725 11965 7075 11975
rect 6725 11635 6735 11965
rect 7065 11635 7075 11965
rect 6725 11625 7075 11635
rect 7150 11550 7200 12050
rect 7275 11965 7625 11975
rect 7275 11635 7285 11965
rect 7615 11635 7625 11965
rect 7275 11625 7625 11635
rect 7700 11550 7750 12050
rect 7825 11965 8175 11975
rect 7825 11635 7835 11965
rect 8165 11635 8175 11965
rect 7825 11625 8175 11635
rect 8250 11550 8300 12050
rect 8375 11965 8725 11975
rect 8375 11635 8385 11965
rect 8715 11635 8725 11965
rect 8375 11625 8725 11635
rect 8800 11550 8850 12050
rect 8925 11965 9275 11975
rect 8925 11635 8935 11965
rect 9265 11635 9275 11965
rect 8925 11625 9275 11635
rect 9350 11550 9400 12050
rect 9475 11965 9825 11975
rect 9475 11635 9485 11965
rect 9815 11635 9825 11965
rect 9475 11625 9825 11635
rect 9900 11550 9950 12050
rect 10025 11965 10375 11975
rect 10025 11635 10035 11965
rect 10365 11635 10375 11965
rect 10025 11625 10375 11635
rect 10450 11550 10500 12050
rect 10575 11965 10925 11975
rect 10575 11635 10585 11965
rect 10915 11635 10925 11965
rect 10575 11625 10925 11635
rect 11000 11550 11050 12050
rect 11125 11965 11475 11975
rect 11125 11635 11135 11965
rect 11465 11635 11475 11965
rect 11125 11625 11475 11635
rect 11550 11550 11600 12050
rect 11675 11965 12025 11975
rect 11675 11635 11685 11965
rect 12015 11635 12025 11965
rect 11675 11625 12025 11635
rect 12100 11550 12150 12050
rect 12225 11965 12575 11975
rect 12225 11635 12235 11965
rect 12565 11635 12575 11965
rect 12225 11625 12575 11635
rect 12650 11550 12700 12050
rect 12775 11965 13125 11975
rect 12775 11635 12785 11965
rect 13115 11635 13125 11965
rect 12775 11625 13125 11635
rect 13200 11550 13250 12050
rect 13325 11965 13675 11975
rect 13325 11635 13335 11965
rect 13665 11635 13675 11965
rect 13325 11625 13675 11635
rect 13750 11550 13975 12050
rect -725 11542 13975 11550
rect -725 11508 -542 11542
rect -508 11508 8 11542
rect 42 11508 558 11542
rect 592 11508 1108 11542
rect 1142 11508 1658 11542
rect 1692 11508 2208 11542
rect 2242 11508 2758 11542
rect 2792 11508 3308 11542
rect 3342 11508 3858 11542
rect 3892 11508 4408 11542
rect 4442 11508 4958 11542
rect 4992 11508 5508 11542
rect 5542 11508 6058 11542
rect 6092 11508 6608 11542
rect 6642 11508 7158 11542
rect 7192 11508 7708 11542
rect 7742 11508 8258 11542
rect 8292 11508 8808 11542
rect 8842 11508 9358 11542
rect 9392 11508 9908 11542
rect 9942 11508 10458 11542
rect 10492 11508 11008 11542
rect 11042 11508 11558 11542
rect 11592 11508 12108 11542
rect 12142 11508 12658 11542
rect 12692 11508 13208 11542
rect 13242 11508 13758 11542
rect 13792 11508 13975 11542
rect -725 11500 13975 11508
rect -725 11000 -500 11500
rect -425 11415 -75 11425
rect -425 11085 -415 11415
rect -85 11085 -75 11415
rect -425 11075 -75 11085
rect 0 11000 50 11500
rect 125 11415 475 11425
rect 125 11085 135 11415
rect 465 11085 475 11415
rect 125 11075 475 11085
rect 550 11000 600 11500
rect 675 11415 1025 11425
rect 675 11085 685 11415
rect 1015 11085 1025 11415
rect 675 11075 1025 11085
rect 1100 11000 1150 11500
rect 1225 11415 1575 11425
rect 1225 11085 1235 11415
rect 1565 11085 1575 11415
rect 1225 11075 1575 11085
rect 1650 11000 1700 11500
rect 1775 11415 2125 11425
rect 1775 11085 1785 11415
rect 2115 11085 2125 11415
rect 1775 11075 2125 11085
rect 2200 11000 2250 11500
rect 2325 11415 2675 11425
rect 2325 11085 2335 11415
rect 2665 11085 2675 11415
rect 2325 11075 2675 11085
rect 2750 11000 2800 11500
rect 2875 11415 3225 11425
rect 2875 11085 2885 11415
rect 3215 11085 3225 11415
rect 2875 11075 3225 11085
rect 3300 11000 3350 11500
rect 3425 11415 3775 11425
rect 3425 11085 3435 11415
rect 3765 11085 3775 11415
rect 3425 11075 3775 11085
rect 3850 11000 3900 11500
rect 3975 11415 4325 11425
rect 3975 11085 3985 11415
rect 4315 11085 4325 11415
rect 3975 11075 4325 11085
rect 4400 11000 4450 11500
rect 4525 11415 4875 11425
rect 4525 11085 4535 11415
rect 4865 11085 4875 11415
rect 4525 11075 4875 11085
rect 4950 11000 5000 11500
rect 5075 11415 5425 11425
rect 5075 11085 5085 11415
rect 5415 11085 5425 11415
rect 5075 11075 5425 11085
rect 5500 11000 5550 11500
rect 5625 11415 5975 11425
rect 5625 11085 5635 11415
rect 5965 11085 5975 11415
rect 5625 11075 5975 11085
rect 6050 11000 6100 11500
rect 6175 11415 6525 11425
rect 6175 11085 6185 11415
rect 6515 11085 6525 11415
rect 6175 11075 6525 11085
rect 6600 11000 6650 11500
rect 6725 11415 7075 11425
rect 6725 11085 6735 11415
rect 7065 11085 7075 11415
rect 6725 11075 7075 11085
rect 7150 11000 7200 11500
rect 7275 11415 7625 11425
rect 7275 11085 7285 11415
rect 7615 11085 7625 11415
rect 7275 11075 7625 11085
rect 7700 11000 7750 11500
rect 7825 11415 8175 11425
rect 7825 11085 7835 11415
rect 8165 11085 8175 11415
rect 7825 11075 8175 11085
rect 8250 11000 8300 11500
rect 8375 11415 8725 11425
rect 8375 11085 8385 11415
rect 8715 11085 8725 11415
rect 8375 11075 8725 11085
rect 8800 11000 8850 11500
rect 8925 11415 9275 11425
rect 8925 11085 8935 11415
rect 9265 11085 9275 11415
rect 8925 11075 9275 11085
rect 9350 11000 9400 11500
rect 9475 11415 9825 11425
rect 9475 11085 9485 11415
rect 9815 11085 9825 11415
rect 9475 11075 9825 11085
rect 9900 11000 9950 11500
rect 10025 11415 10375 11425
rect 10025 11085 10035 11415
rect 10365 11085 10375 11415
rect 10025 11075 10375 11085
rect 10450 11000 10500 11500
rect 10575 11415 10925 11425
rect 10575 11085 10585 11415
rect 10915 11085 10925 11415
rect 10575 11075 10925 11085
rect 11000 11000 11050 11500
rect 11125 11415 11475 11425
rect 11125 11085 11135 11415
rect 11465 11085 11475 11415
rect 11125 11075 11475 11085
rect 11550 11000 11600 11500
rect 11675 11415 12025 11425
rect 11675 11085 11685 11415
rect 12015 11085 12025 11415
rect 11675 11075 12025 11085
rect 12100 11000 12150 11500
rect 12225 11415 12575 11425
rect 12225 11085 12235 11415
rect 12565 11085 12575 11415
rect 12225 11075 12575 11085
rect 12650 11000 12700 11500
rect 12775 11415 13125 11425
rect 12775 11085 12785 11415
rect 13115 11085 13125 11415
rect 12775 11075 13125 11085
rect 13200 11000 13250 11500
rect 13325 11415 13675 11425
rect 13325 11085 13335 11415
rect 13665 11085 13675 11415
rect 13325 11075 13675 11085
rect 13750 11000 13975 11500
rect 14065 11138 14185 11148
rect 14065 11038 14075 11138
rect 14175 11038 14185 11138
rect 14065 11028 14185 11038
rect -725 10992 13975 11000
rect -725 10958 -542 10992
rect -508 10958 8 10992
rect 42 10958 558 10992
rect 592 10958 1108 10992
rect 1142 10958 1658 10992
rect 1692 10958 2208 10992
rect 2242 10958 2758 10992
rect 2792 10958 3308 10992
rect 3342 10958 3858 10992
rect 3892 10958 4408 10992
rect 4442 10958 4958 10992
rect 4992 10958 5508 10992
rect 5542 10958 6058 10992
rect 6092 10958 6608 10992
rect 6642 10958 7158 10992
rect 7192 10958 7708 10992
rect 7742 10958 8258 10992
rect 8292 10958 8808 10992
rect 8842 10958 9358 10992
rect 9392 10958 9908 10992
rect 9942 10958 10458 10992
rect 10492 10958 11008 10992
rect 11042 10958 11558 10992
rect 11592 10958 12108 10992
rect 12142 10958 12658 10992
rect 12692 10958 13208 10992
rect 13242 10958 13758 10992
rect 13792 10958 13975 10992
rect -725 10950 13975 10958
rect -935 10912 -815 10922
rect -935 10812 -925 10912
rect -825 10812 -815 10912
rect -935 10802 -815 10812
rect -725 10450 -500 10950
rect -425 10865 -75 10875
rect -425 10535 -415 10865
rect -85 10535 -75 10865
rect -425 10525 -75 10535
rect 0 10450 50 10950
rect 125 10865 475 10875
rect 125 10535 135 10865
rect 465 10535 475 10865
rect 125 10525 475 10535
rect 550 10450 600 10950
rect 675 10865 1025 10875
rect 675 10535 685 10865
rect 1015 10535 1025 10865
rect 675 10525 1025 10535
rect 1100 10450 1150 10950
rect 1225 10865 1575 10875
rect 1225 10535 1235 10865
rect 1565 10535 1575 10865
rect 1225 10525 1575 10535
rect 1650 10450 1700 10950
rect 1775 10865 2125 10875
rect 1775 10535 1785 10865
rect 2115 10535 2125 10865
rect 1775 10525 2125 10535
rect 2200 10450 2250 10950
rect 2325 10865 2675 10875
rect 2325 10535 2335 10865
rect 2665 10535 2675 10865
rect 2325 10525 2675 10535
rect 2750 10450 2800 10950
rect 2875 10865 3225 10875
rect 2875 10535 2885 10865
rect 3215 10535 3225 10865
rect 2875 10525 3225 10535
rect 3300 10450 3350 10950
rect 3425 10865 3775 10875
rect 3425 10535 3435 10865
rect 3765 10535 3775 10865
rect 3425 10525 3775 10535
rect 3850 10450 3900 10950
rect 3975 10865 4325 10875
rect 3975 10535 3985 10865
rect 4315 10535 4325 10865
rect 3975 10525 4325 10535
rect 4400 10450 4450 10950
rect 4525 10865 4875 10875
rect 4525 10535 4535 10865
rect 4865 10535 4875 10865
rect 4525 10525 4875 10535
rect 4950 10450 5000 10950
rect 5075 10865 5425 10875
rect 5075 10535 5085 10865
rect 5415 10535 5425 10865
rect 5075 10525 5425 10535
rect 5500 10450 5550 10950
rect 5625 10865 5975 10875
rect 5625 10535 5635 10865
rect 5965 10535 5975 10865
rect 5625 10525 5975 10535
rect 6050 10450 6100 10950
rect 6175 10865 6525 10875
rect 6175 10535 6185 10865
rect 6515 10535 6525 10865
rect 6175 10525 6525 10535
rect 6600 10450 6650 10950
rect 6725 10865 7075 10875
rect 6725 10535 6735 10865
rect 7065 10535 7075 10865
rect 6725 10525 7075 10535
rect 7150 10450 7200 10950
rect 7275 10865 7625 10875
rect 7275 10535 7285 10865
rect 7615 10535 7625 10865
rect 7275 10525 7625 10535
rect 7700 10450 7750 10950
rect 7825 10865 8175 10875
rect 7825 10535 7835 10865
rect 8165 10535 8175 10865
rect 7825 10525 8175 10535
rect 8250 10450 8300 10950
rect 8375 10865 8725 10875
rect 8375 10535 8385 10865
rect 8715 10535 8725 10865
rect 8375 10525 8725 10535
rect 8800 10450 8850 10950
rect 8925 10865 9275 10875
rect 8925 10535 8935 10865
rect 9265 10535 9275 10865
rect 8925 10525 9275 10535
rect 9350 10450 9400 10950
rect 9475 10865 9825 10875
rect 9475 10535 9485 10865
rect 9815 10535 9825 10865
rect 9475 10525 9825 10535
rect 9900 10450 9950 10950
rect 10025 10865 10375 10875
rect 10025 10535 10035 10865
rect 10365 10535 10375 10865
rect 10025 10525 10375 10535
rect 10450 10450 10500 10950
rect 10575 10865 10925 10875
rect 10575 10535 10585 10865
rect 10915 10535 10925 10865
rect 10575 10525 10925 10535
rect 11000 10450 11050 10950
rect 11125 10865 11475 10875
rect 11125 10535 11135 10865
rect 11465 10535 11475 10865
rect 11125 10525 11475 10535
rect 11550 10450 11600 10950
rect 11675 10865 12025 10875
rect 11675 10535 11685 10865
rect 12015 10535 12025 10865
rect 11675 10525 12025 10535
rect 12100 10450 12150 10950
rect 12225 10865 12575 10875
rect 12225 10535 12235 10865
rect 12565 10535 12575 10865
rect 12225 10525 12575 10535
rect 12650 10450 12700 10950
rect 12775 10865 13125 10875
rect 12775 10535 12785 10865
rect 13115 10535 13125 10865
rect 12775 10525 13125 10535
rect 13200 10450 13250 10950
rect 13325 10865 13675 10875
rect 13325 10535 13335 10865
rect 13665 10535 13675 10865
rect 13325 10525 13675 10535
rect 13750 10450 13975 10950
rect -725 10442 13975 10450
rect -725 10408 -542 10442
rect -508 10408 8 10442
rect 42 10408 558 10442
rect 592 10408 1108 10442
rect 1142 10408 1658 10442
rect 1692 10408 2208 10442
rect 2242 10408 2758 10442
rect 2792 10408 3308 10442
rect 3342 10408 3858 10442
rect 3892 10408 4408 10442
rect 4442 10408 4958 10442
rect 4992 10408 5508 10442
rect 5542 10408 6058 10442
rect 6092 10408 6608 10442
rect 6642 10408 7158 10442
rect 7192 10408 7708 10442
rect 7742 10408 8258 10442
rect 8292 10408 8808 10442
rect 8842 10408 9358 10442
rect 9392 10408 9908 10442
rect 9942 10408 10458 10442
rect 10492 10408 11008 10442
rect 11042 10408 11558 10442
rect 11592 10408 12108 10442
rect 12142 10408 12658 10442
rect 12692 10408 13208 10442
rect 13242 10408 13758 10442
rect 13792 10408 13975 10442
rect -725 10400 13975 10408
rect -725 9900 -500 10400
rect -425 10315 -75 10325
rect -425 9985 -415 10315
rect -85 9985 -75 10315
rect -425 9975 -75 9985
rect 0 9900 50 10400
rect 125 10315 475 10325
rect 125 9985 135 10315
rect 465 9985 475 10315
rect 125 9975 475 9985
rect 550 9900 600 10400
rect 675 10315 1025 10325
rect 675 9985 685 10315
rect 1015 9985 1025 10315
rect 675 9975 1025 9985
rect 1100 9900 1150 10400
rect 1225 10315 1575 10325
rect 1225 9985 1235 10315
rect 1565 9985 1575 10315
rect 1225 9975 1575 9985
rect 1650 9900 1700 10400
rect 1775 10315 2125 10325
rect 1775 9985 1785 10315
rect 2115 9985 2125 10315
rect 1775 9975 2125 9985
rect 2200 9900 2250 10400
rect 2325 10315 2675 10325
rect 2325 9985 2335 10315
rect 2665 9985 2675 10315
rect 2325 9975 2675 9985
rect 2750 9900 2800 10400
rect 2875 10315 3225 10325
rect 2875 9985 2885 10315
rect 3215 9985 3225 10315
rect 2875 9975 3225 9985
rect 3300 9900 3350 10400
rect 3425 10315 3775 10325
rect 3425 9985 3435 10315
rect 3765 9985 3775 10315
rect 3425 9975 3775 9985
rect 3850 9900 3900 10400
rect 3975 10315 4325 10325
rect 3975 9985 3985 10315
rect 4315 9985 4325 10315
rect 3975 9975 4325 9985
rect 4400 9900 4450 10400
rect 4525 10315 4875 10325
rect 4525 9985 4535 10315
rect 4865 9985 4875 10315
rect 4525 9975 4875 9985
rect 4950 9900 5000 10400
rect 5075 10315 5425 10325
rect 5075 9985 5085 10315
rect 5415 9985 5425 10315
rect 5075 9975 5425 9985
rect 5500 9900 5550 10400
rect 5625 10315 5975 10325
rect 5625 9985 5635 10315
rect 5965 9985 5975 10315
rect 5625 9975 5975 9985
rect 6050 9900 6100 10400
rect 6175 10315 6525 10325
rect 6175 9985 6185 10315
rect 6515 9985 6525 10315
rect 6175 9975 6525 9985
rect 6600 9900 6650 10400
rect 6725 10315 7075 10325
rect 6725 9985 6735 10315
rect 7065 9985 7075 10315
rect 6725 9975 7075 9985
rect 7150 9900 7200 10400
rect 7275 10315 7625 10325
rect 7275 9985 7285 10315
rect 7615 9985 7625 10315
rect 7275 9975 7625 9985
rect 7700 9900 7750 10400
rect 7825 10315 8175 10325
rect 7825 9985 7835 10315
rect 8165 9985 8175 10315
rect 7825 9975 8175 9985
rect 8250 9900 8300 10400
rect 8375 10315 8725 10325
rect 8375 9985 8385 10315
rect 8715 9985 8725 10315
rect 8375 9975 8725 9985
rect 8800 9900 8850 10400
rect 8925 10315 9275 10325
rect 8925 9985 8935 10315
rect 9265 9985 9275 10315
rect 8925 9975 9275 9985
rect 9350 9900 9400 10400
rect 9475 10315 9825 10325
rect 9475 9985 9485 10315
rect 9815 9985 9825 10315
rect 9475 9975 9825 9985
rect 9900 9900 9950 10400
rect 10025 10315 10375 10325
rect 10025 9985 10035 10315
rect 10365 9985 10375 10315
rect 10025 9975 10375 9985
rect 10450 9900 10500 10400
rect 10575 10315 10925 10325
rect 10575 9985 10585 10315
rect 10915 9985 10925 10315
rect 10575 9975 10925 9985
rect 11000 9900 11050 10400
rect 11125 10315 11475 10325
rect 11125 9985 11135 10315
rect 11465 9985 11475 10315
rect 11125 9975 11475 9985
rect 11550 9900 11600 10400
rect 11675 10315 12025 10325
rect 11675 9985 11685 10315
rect 12015 9985 12025 10315
rect 11675 9975 12025 9985
rect 12100 9900 12150 10400
rect 12225 10315 12575 10325
rect 12225 9985 12235 10315
rect 12565 9985 12575 10315
rect 12225 9975 12575 9985
rect 12650 9900 12700 10400
rect 12775 10315 13125 10325
rect 12775 9985 12785 10315
rect 13115 9985 13125 10315
rect 12775 9975 13125 9985
rect 13200 9900 13250 10400
rect 13325 10315 13675 10325
rect 13325 9985 13335 10315
rect 13665 9985 13675 10315
rect 13325 9975 13675 9985
rect 13750 9900 13975 10400
rect 14065 10038 14185 10048
rect 14065 9938 14075 10038
rect 14175 9938 14185 10038
rect 14065 9928 14185 9938
rect -725 9892 13975 9900
rect -725 9858 -542 9892
rect -508 9858 8 9892
rect 42 9858 558 9892
rect 592 9858 1108 9892
rect 1142 9858 1658 9892
rect 1692 9858 2208 9892
rect 2242 9858 2758 9892
rect 2792 9858 3308 9892
rect 3342 9858 3858 9892
rect 3892 9858 4408 9892
rect 4442 9858 4958 9892
rect 4992 9858 5508 9892
rect 5542 9858 6058 9892
rect 6092 9858 6608 9892
rect 6642 9858 7158 9892
rect 7192 9858 7708 9892
rect 7742 9858 8258 9892
rect 8292 9858 8808 9892
rect 8842 9858 9358 9892
rect 9392 9858 9908 9892
rect 9942 9858 10458 9892
rect 10492 9858 11008 9892
rect 11042 9858 11558 9892
rect 11592 9858 12108 9892
rect 12142 9858 12658 9892
rect 12692 9858 13208 9892
rect 13242 9858 13758 9892
rect 13792 9858 13975 9892
rect -725 9850 13975 9858
rect -935 9812 -815 9822
rect -935 9712 -925 9812
rect -825 9712 -815 9812
rect -935 9702 -815 9712
rect -725 9350 -500 9850
rect -425 9765 -75 9775
rect -425 9435 -415 9765
rect -85 9435 -75 9765
rect -425 9425 -75 9435
rect 0 9350 50 9850
rect 125 9765 475 9775
rect 125 9435 135 9765
rect 465 9435 475 9765
rect 125 9425 475 9435
rect 550 9350 600 9850
rect 675 9765 1025 9775
rect 675 9435 685 9765
rect 1015 9435 1025 9765
rect 675 9425 1025 9435
rect 1100 9350 1150 9850
rect 1225 9765 1575 9775
rect 1225 9435 1235 9765
rect 1565 9435 1575 9765
rect 1225 9425 1575 9435
rect 1650 9350 1700 9850
rect 1775 9765 2125 9775
rect 1775 9435 1785 9765
rect 2115 9435 2125 9765
rect 1775 9425 2125 9435
rect 2200 9350 2250 9850
rect 2325 9765 2675 9775
rect 2325 9435 2335 9765
rect 2665 9435 2675 9765
rect 2325 9425 2675 9435
rect 2750 9350 2800 9850
rect 2875 9765 3225 9775
rect 2875 9435 2885 9765
rect 3215 9435 3225 9765
rect 2875 9425 3225 9435
rect 3300 9350 3350 9850
rect 3425 9765 3775 9775
rect 3425 9435 3435 9765
rect 3765 9435 3775 9765
rect 3425 9425 3775 9435
rect 3850 9350 3900 9850
rect 3975 9765 4325 9775
rect 3975 9435 3985 9765
rect 4315 9435 4325 9765
rect 3975 9425 4325 9435
rect 4400 9350 4450 9850
rect 4525 9765 4875 9775
rect 4525 9435 4535 9765
rect 4865 9435 4875 9765
rect 4525 9425 4875 9435
rect 4950 9350 5000 9850
rect 5075 9765 5425 9775
rect 5075 9435 5085 9765
rect 5415 9435 5425 9765
rect 5075 9425 5425 9435
rect 5500 9350 5550 9850
rect 5625 9765 5975 9775
rect 5625 9435 5635 9765
rect 5965 9435 5975 9765
rect 5625 9425 5975 9435
rect 6050 9350 6100 9850
rect 6175 9765 6525 9775
rect 6175 9435 6185 9765
rect 6515 9435 6525 9765
rect 6175 9425 6525 9435
rect 6600 9350 6650 9850
rect 6725 9765 7075 9775
rect 6725 9435 6735 9765
rect 7065 9435 7075 9765
rect 6725 9425 7075 9435
rect 7150 9350 7200 9850
rect 7275 9765 7625 9775
rect 7275 9435 7285 9765
rect 7615 9435 7625 9765
rect 7275 9425 7625 9435
rect 7700 9350 7750 9850
rect 7825 9765 8175 9775
rect 7825 9435 7835 9765
rect 8165 9435 8175 9765
rect 7825 9425 8175 9435
rect 8250 9350 8300 9850
rect 8375 9765 8725 9775
rect 8375 9435 8385 9765
rect 8715 9435 8725 9765
rect 8375 9425 8725 9435
rect 8800 9350 8850 9850
rect 8925 9765 9275 9775
rect 8925 9435 8935 9765
rect 9265 9435 9275 9765
rect 8925 9425 9275 9435
rect 9350 9350 9400 9850
rect 9475 9765 9825 9775
rect 9475 9435 9485 9765
rect 9815 9435 9825 9765
rect 9475 9425 9825 9435
rect 9900 9350 9950 9850
rect 10025 9765 10375 9775
rect 10025 9435 10035 9765
rect 10365 9435 10375 9765
rect 10025 9425 10375 9435
rect 10450 9350 10500 9850
rect 10575 9765 10925 9775
rect 10575 9435 10585 9765
rect 10915 9435 10925 9765
rect 10575 9425 10925 9435
rect 11000 9350 11050 9850
rect 11125 9765 11475 9775
rect 11125 9435 11135 9765
rect 11465 9435 11475 9765
rect 11125 9425 11475 9435
rect 11550 9350 11600 9850
rect 11675 9765 12025 9775
rect 11675 9435 11685 9765
rect 12015 9435 12025 9765
rect 11675 9425 12025 9435
rect 12100 9350 12150 9850
rect 12225 9765 12575 9775
rect 12225 9435 12235 9765
rect 12565 9435 12575 9765
rect 12225 9425 12575 9435
rect 12650 9350 12700 9850
rect 12775 9765 13125 9775
rect 12775 9435 12785 9765
rect 13115 9435 13125 9765
rect 12775 9425 13125 9435
rect 13200 9350 13250 9850
rect 13325 9765 13675 9775
rect 13325 9435 13335 9765
rect 13665 9435 13675 9765
rect 13325 9425 13675 9435
rect 13750 9350 13975 9850
rect -725 9342 13975 9350
rect -725 9308 -542 9342
rect -508 9308 8 9342
rect 42 9308 558 9342
rect 592 9308 1108 9342
rect 1142 9308 1658 9342
rect 1692 9308 2208 9342
rect 2242 9308 2758 9342
rect 2792 9308 3308 9342
rect 3342 9308 3858 9342
rect 3892 9308 4408 9342
rect 4442 9308 4958 9342
rect 4992 9308 5508 9342
rect 5542 9308 6058 9342
rect 6092 9308 6608 9342
rect 6642 9308 7158 9342
rect 7192 9308 7708 9342
rect 7742 9308 8258 9342
rect 8292 9308 8808 9342
rect 8842 9308 9358 9342
rect 9392 9308 9908 9342
rect 9942 9308 10458 9342
rect 10492 9308 11008 9342
rect 11042 9308 11558 9342
rect 11592 9308 12108 9342
rect 12142 9308 12658 9342
rect 12692 9308 13208 9342
rect 13242 9308 13758 9342
rect 13792 9308 13975 9342
rect -725 9300 13975 9308
rect -725 8800 -500 9300
rect -425 9215 -75 9225
rect -425 8885 -415 9215
rect -85 8885 -75 9215
rect -425 8875 -75 8885
rect 0 8800 50 9300
rect 125 9215 475 9225
rect 125 8885 135 9215
rect 465 8885 475 9215
rect 125 8875 475 8885
rect 550 8800 600 9300
rect 675 9215 1025 9225
rect 675 8885 685 9215
rect 1015 8885 1025 9215
rect 675 8875 1025 8885
rect 1100 8800 1150 9300
rect 1225 9215 1575 9225
rect 1225 8885 1235 9215
rect 1565 8885 1575 9215
rect 1225 8875 1575 8885
rect 1650 8800 1700 9300
rect 1775 9215 2125 9225
rect 1775 8885 1785 9215
rect 2115 8885 2125 9215
rect 1775 8875 2125 8885
rect 2200 8800 2250 9300
rect 2325 9215 2675 9225
rect 2325 8885 2335 9215
rect 2665 8885 2675 9215
rect 2325 8875 2675 8885
rect 2750 8800 2800 9300
rect 2875 9215 3225 9225
rect 2875 8885 2885 9215
rect 3215 8885 3225 9215
rect 2875 8875 3225 8885
rect 3300 8800 3350 9300
rect 3425 9215 3775 9225
rect 3425 8885 3435 9215
rect 3765 8885 3775 9215
rect 3425 8875 3775 8885
rect 3850 8800 3900 9300
rect 3975 9215 4325 9225
rect 3975 8885 3985 9215
rect 4315 8885 4325 9215
rect 3975 8875 4325 8885
rect 4400 8800 4450 9300
rect 4525 9215 4875 9225
rect 4525 8885 4535 9215
rect 4865 8885 4875 9215
rect 4525 8875 4875 8885
rect 4950 8800 5000 9300
rect 5075 9215 5425 9225
rect 5075 8885 5085 9215
rect 5415 8885 5425 9215
rect 5075 8875 5425 8885
rect 5500 8800 5550 9300
rect 5625 9215 5975 9225
rect 5625 8885 5635 9215
rect 5965 8885 5975 9215
rect 5625 8875 5975 8885
rect 6050 8800 6100 9300
rect 6175 9215 6525 9225
rect 6175 8885 6185 9215
rect 6515 8885 6525 9215
rect 6175 8875 6525 8885
rect 6600 8800 6650 9300
rect 6725 9215 7075 9225
rect 6725 8885 6735 9215
rect 7065 8885 7075 9215
rect 6725 8875 7075 8885
rect 7150 8800 7200 9300
rect 7275 9215 7625 9225
rect 7275 8885 7285 9215
rect 7615 8885 7625 9215
rect 7275 8875 7625 8885
rect 7700 8800 7750 9300
rect 7825 9215 8175 9225
rect 7825 8885 7835 9215
rect 8165 8885 8175 9215
rect 7825 8875 8175 8885
rect 8250 8800 8300 9300
rect 8375 9215 8725 9225
rect 8375 8885 8385 9215
rect 8715 8885 8725 9215
rect 8375 8875 8725 8885
rect 8800 8800 8850 9300
rect 8925 9215 9275 9225
rect 8925 8885 8935 9215
rect 9265 8885 9275 9215
rect 8925 8875 9275 8885
rect 9350 8800 9400 9300
rect 9475 9215 9825 9225
rect 9475 8885 9485 9215
rect 9815 8885 9825 9215
rect 9475 8875 9825 8885
rect 9900 8800 9950 9300
rect 10025 9215 10375 9225
rect 10025 8885 10035 9215
rect 10365 8885 10375 9215
rect 10025 8875 10375 8885
rect 10450 8800 10500 9300
rect 10575 9215 10925 9225
rect 10575 8885 10585 9215
rect 10915 8885 10925 9215
rect 10575 8875 10925 8885
rect 11000 8800 11050 9300
rect 11125 9215 11475 9225
rect 11125 8885 11135 9215
rect 11465 8885 11475 9215
rect 11125 8875 11475 8885
rect 11550 8800 11600 9300
rect 11675 9215 12025 9225
rect 11675 8885 11685 9215
rect 12015 8885 12025 9215
rect 11675 8875 12025 8885
rect 12100 8800 12150 9300
rect 12225 9215 12575 9225
rect 12225 8885 12235 9215
rect 12565 8885 12575 9215
rect 12225 8875 12575 8885
rect 12650 8800 12700 9300
rect 12775 9215 13125 9225
rect 12775 8885 12785 9215
rect 13115 8885 13125 9215
rect 12775 8875 13125 8885
rect 13200 8800 13250 9300
rect 13325 9215 13675 9225
rect 13325 8885 13335 9215
rect 13665 8885 13675 9215
rect 13325 8875 13675 8885
rect 13750 8800 13975 9300
rect 14065 8938 14185 8948
rect 14065 8838 14075 8938
rect 14175 8838 14185 8938
rect 14065 8828 14185 8838
rect -725 8792 13975 8800
rect -725 8758 -542 8792
rect -508 8758 8 8792
rect 42 8758 558 8792
rect 592 8758 1108 8792
rect 1142 8758 1658 8792
rect 1692 8758 2208 8792
rect 2242 8758 2758 8792
rect 2792 8758 3308 8792
rect 3342 8758 3858 8792
rect 3892 8758 4408 8792
rect 4442 8758 4958 8792
rect 4992 8758 5508 8792
rect 5542 8758 6058 8792
rect 6092 8758 6608 8792
rect 6642 8758 7158 8792
rect 7192 8758 7708 8792
rect 7742 8758 8258 8792
rect 8292 8758 8808 8792
rect 8842 8758 9358 8792
rect 9392 8758 9908 8792
rect 9942 8758 10458 8792
rect 10492 8758 11008 8792
rect 11042 8758 11558 8792
rect 11592 8758 12108 8792
rect 12142 8758 12658 8792
rect 12692 8758 13208 8792
rect 13242 8758 13758 8792
rect 13792 8758 13975 8792
rect -725 8750 13975 8758
rect -935 8712 -815 8722
rect -935 8612 -925 8712
rect -825 8612 -815 8712
rect -935 8602 -815 8612
rect -725 8250 -500 8750
rect -425 8665 -75 8675
rect -425 8335 -415 8665
rect -85 8335 -75 8665
rect -425 8325 -75 8335
rect 0 8250 50 8750
rect 125 8665 475 8675
rect 125 8335 135 8665
rect 465 8335 475 8665
rect 125 8325 475 8335
rect 550 8250 600 8750
rect 675 8665 1025 8675
rect 675 8335 685 8665
rect 1015 8335 1025 8665
rect 675 8325 1025 8335
rect 1100 8250 1150 8750
rect 1225 8665 1575 8675
rect 1225 8335 1235 8665
rect 1565 8335 1575 8665
rect 1225 8325 1575 8335
rect 1650 8250 1700 8750
rect 1775 8665 2125 8675
rect 1775 8335 1785 8665
rect 2115 8335 2125 8665
rect 1775 8325 2125 8335
rect 2200 8250 2250 8750
rect 2325 8665 2675 8675
rect 2325 8335 2335 8665
rect 2665 8335 2675 8665
rect 2325 8325 2675 8335
rect 2750 8250 2800 8750
rect 2875 8665 3225 8675
rect 2875 8335 2885 8665
rect 3215 8335 3225 8665
rect 2875 8325 3225 8335
rect 3300 8250 3350 8750
rect 3425 8665 3775 8675
rect 3425 8335 3435 8665
rect 3765 8335 3775 8665
rect 3425 8325 3775 8335
rect 3850 8250 3900 8750
rect 3975 8665 4325 8675
rect 3975 8335 3985 8665
rect 4315 8335 4325 8665
rect 3975 8325 4325 8335
rect 4400 8250 4450 8750
rect 4525 8665 4875 8675
rect 4525 8335 4535 8665
rect 4865 8335 4875 8665
rect 4525 8325 4875 8335
rect 4950 8250 5000 8750
rect 5075 8665 5425 8675
rect 5075 8335 5085 8665
rect 5415 8335 5425 8665
rect 5075 8325 5425 8335
rect 5500 8250 5550 8750
rect 5625 8665 5975 8675
rect 5625 8335 5635 8665
rect 5965 8335 5975 8665
rect 5625 8325 5975 8335
rect 6050 8250 6100 8750
rect 6175 8665 6525 8675
rect 6175 8335 6185 8665
rect 6515 8335 6525 8665
rect 6175 8325 6525 8335
rect 6600 8250 6650 8750
rect 6725 8665 7075 8675
rect 6725 8335 6735 8665
rect 7065 8335 7075 8665
rect 6725 8325 7075 8335
rect 7150 8250 7200 8750
rect 7275 8665 7625 8675
rect 7275 8335 7285 8665
rect 7615 8335 7625 8665
rect 7275 8325 7625 8335
rect 7700 8250 7750 8750
rect 7825 8665 8175 8675
rect 7825 8335 7835 8665
rect 8165 8335 8175 8665
rect 7825 8325 8175 8335
rect 8250 8250 8300 8750
rect 8375 8665 8725 8675
rect 8375 8335 8385 8665
rect 8715 8335 8725 8665
rect 8375 8325 8725 8335
rect 8800 8250 8850 8750
rect 8925 8665 9275 8675
rect 8925 8335 8935 8665
rect 9265 8335 9275 8665
rect 8925 8325 9275 8335
rect 9350 8250 9400 8750
rect 9475 8665 9825 8675
rect 9475 8335 9485 8665
rect 9815 8335 9825 8665
rect 9475 8325 9825 8335
rect 9900 8250 9950 8750
rect 10025 8665 10375 8675
rect 10025 8335 10035 8665
rect 10365 8335 10375 8665
rect 10025 8325 10375 8335
rect 10450 8250 10500 8750
rect 10575 8665 10925 8675
rect 10575 8335 10585 8665
rect 10915 8335 10925 8665
rect 10575 8325 10925 8335
rect 11000 8250 11050 8750
rect 11125 8665 11475 8675
rect 11125 8335 11135 8665
rect 11465 8335 11475 8665
rect 11125 8325 11475 8335
rect 11550 8250 11600 8750
rect 11675 8665 12025 8675
rect 11675 8335 11685 8665
rect 12015 8335 12025 8665
rect 11675 8325 12025 8335
rect 12100 8250 12150 8750
rect 12225 8665 12575 8675
rect 12225 8335 12235 8665
rect 12565 8335 12575 8665
rect 12225 8325 12575 8335
rect 12650 8250 12700 8750
rect 12775 8665 13125 8675
rect 12775 8335 12785 8665
rect 13115 8335 13125 8665
rect 12775 8325 13125 8335
rect 13200 8250 13250 8750
rect 13325 8665 13675 8675
rect 13325 8335 13335 8665
rect 13665 8335 13675 8665
rect 13325 8325 13675 8335
rect 13750 8250 13975 8750
rect -725 8242 13975 8250
rect -725 8208 -542 8242
rect -508 8208 8 8242
rect 42 8208 558 8242
rect 592 8208 1108 8242
rect 1142 8208 1658 8242
rect 1692 8208 2208 8242
rect 2242 8208 2758 8242
rect 2792 8208 3308 8242
rect 3342 8208 3858 8242
rect 3892 8208 4408 8242
rect 4442 8208 4958 8242
rect 4992 8208 5508 8242
rect 5542 8208 6058 8242
rect 6092 8208 6608 8242
rect 6642 8208 7158 8242
rect 7192 8208 7708 8242
rect 7742 8208 8258 8242
rect 8292 8208 8808 8242
rect 8842 8208 9358 8242
rect 9392 8208 9908 8242
rect 9942 8208 10458 8242
rect 10492 8208 11008 8242
rect 11042 8208 11558 8242
rect 11592 8208 12108 8242
rect 12142 8208 12658 8242
rect 12692 8208 13208 8242
rect 13242 8208 13758 8242
rect 13792 8208 13975 8242
rect -725 8200 13975 8208
rect -725 7700 -500 8200
rect -425 8115 -75 8125
rect -425 7785 -415 8115
rect -85 7785 -75 8115
rect -425 7775 -75 7785
rect 0 7700 50 8200
rect 125 8115 475 8125
rect 125 7785 135 8115
rect 465 7785 475 8115
rect 125 7775 475 7785
rect 550 7700 600 8200
rect 675 8115 1025 8125
rect 675 7785 685 8115
rect 1015 7785 1025 8115
rect 675 7775 1025 7785
rect 1100 7700 1150 8200
rect 1225 8115 1575 8125
rect 1225 7785 1235 8115
rect 1565 7785 1575 8115
rect 1225 7775 1575 7785
rect 1650 7700 1700 8200
rect 1775 8115 2125 8125
rect 1775 7785 1785 8115
rect 2115 7785 2125 8115
rect 1775 7775 2125 7785
rect 2200 7700 2250 8200
rect 2325 8115 2675 8125
rect 2325 7785 2335 8115
rect 2665 7785 2675 8115
rect 2325 7775 2675 7785
rect 2750 7700 2800 8200
rect 2875 8115 3225 8125
rect 2875 7785 2885 8115
rect 3215 7785 3225 8115
rect 2875 7775 3225 7785
rect 3300 7700 3350 8200
rect 3425 8115 3775 8125
rect 3425 7785 3435 8115
rect 3765 7785 3775 8115
rect 3425 7775 3775 7785
rect 3850 7700 3900 8200
rect 3975 8115 4325 8125
rect 3975 7785 3985 8115
rect 4315 7785 4325 8115
rect 3975 7775 4325 7785
rect 4400 7700 4450 8200
rect 4525 8115 4875 8125
rect 4525 7785 4535 8115
rect 4865 7785 4875 8115
rect 4525 7775 4875 7785
rect 4950 7700 5000 8200
rect 5075 8115 5425 8125
rect 5075 7785 5085 8115
rect 5415 7785 5425 8115
rect 5075 7775 5425 7785
rect 5500 7700 5550 8200
rect 5625 8115 5975 8125
rect 5625 7785 5635 8115
rect 5965 7785 5975 8115
rect 5625 7775 5975 7785
rect 6050 7700 6100 8200
rect 6175 8115 6525 8125
rect 6175 7785 6185 8115
rect 6515 7785 6525 8115
rect 6175 7775 6525 7785
rect 6600 7700 6650 8200
rect 6725 8115 7075 8125
rect 6725 7785 6735 8115
rect 7065 7785 7075 8115
rect 6725 7775 7075 7785
rect 7150 7700 7200 8200
rect 7275 8115 7625 8125
rect 7275 7785 7285 8115
rect 7615 7785 7625 8115
rect 7275 7775 7625 7785
rect 7700 7700 7750 8200
rect 7825 8115 8175 8125
rect 7825 7785 7835 8115
rect 8165 7785 8175 8115
rect 7825 7775 8175 7785
rect 8250 7700 8300 8200
rect 8375 8115 8725 8125
rect 8375 7785 8385 8115
rect 8715 7785 8725 8115
rect 8375 7775 8725 7785
rect 8800 7700 8850 8200
rect 8925 8115 9275 8125
rect 8925 7785 8935 8115
rect 9265 7785 9275 8115
rect 8925 7775 9275 7785
rect 9350 7700 9400 8200
rect 9475 8115 9825 8125
rect 9475 7785 9485 8115
rect 9815 7785 9825 8115
rect 9475 7775 9825 7785
rect 9900 7700 9950 8200
rect 10025 8115 10375 8125
rect 10025 7785 10035 8115
rect 10365 7785 10375 8115
rect 10025 7775 10375 7785
rect 10450 7700 10500 8200
rect 10575 8115 10925 8125
rect 10575 7785 10585 8115
rect 10915 7785 10925 8115
rect 10575 7775 10925 7785
rect 11000 7700 11050 8200
rect 11125 8115 11475 8125
rect 11125 7785 11135 8115
rect 11465 7785 11475 8115
rect 11125 7775 11475 7785
rect 11550 7700 11600 8200
rect 11675 8115 12025 8125
rect 11675 7785 11685 8115
rect 12015 7785 12025 8115
rect 11675 7775 12025 7785
rect 12100 7700 12150 8200
rect 12225 8115 12575 8125
rect 12225 7785 12235 8115
rect 12565 7785 12575 8115
rect 12225 7775 12575 7785
rect 12650 7700 12700 8200
rect 12775 8115 13125 8125
rect 12775 7785 12785 8115
rect 13115 7785 13125 8115
rect 12775 7775 13125 7785
rect 13200 7700 13250 8200
rect 13325 8115 13675 8125
rect 13325 7785 13335 8115
rect 13665 7785 13675 8115
rect 13325 7775 13675 7785
rect 13750 7700 13975 8200
rect 14065 7838 14185 7848
rect 14065 7738 14075 7838
rect 14175 7738 14185 7838
rect 14065 7728 14185 7738
rect -725 7692 13975 7700
rect -725 7658 -542 7692
rect -508 7658 8 7692
rect 42 7658 558 7692
rect 592 7658 1108 7692
rect 1142 7658 1658 7692
rect 1692 7658 2208 7692
rect 2242 7658 2758 7692
rect 2792 7658 3308 7692
rect 3342 7658 3858 7692
rect 3892 7658 4408 7692
rect 4442 7658 4958 7692
rect 4992 7658 5508 7692
rect 5542 7658 6058 7692
rect 6092 7658 6608 7692
rect 6642 7658 7158 7692
rect 7192 7658 7708 7692
rect 7742 7658 8258 7692
rect 8292 7658 8808 7692
rect 8842 7658 9358 7692
rect 9392 7658 9908 7692
rect 9942 7658 10458 7692
rect 10492 7658 11008 7692
rect 11042 7658 11558 7692
rect 11592 7658 12108 7692
rect 12142 7658 12658 7692
rect 12692 7658 13208 7692
rect 13242 7658 13758 7692
rect 13792 7658 13975 7692
rect -725 7650 13975 7658
rect -935 7612 -815 7622
rect -935 7512 -925 7612
rect -825 7512 -815 7612
rect -935 7502 -815 7512
rect -725 7150 -500 7650
rect -425 7565 -75 7575
rect -425 7235 -415 7565
rect -85 7235 -75 7565
rect -425 7225 -75 7235
rect 0 7150 50 7650
rect 125 7565 475 7575
rect 125 7235 135 7565
rect 465 7235 475 7565
rect 125 7225 475 7235
rect 550 7150 600 7650
rect 675 7565 1025 7575
rect 675 7235 685 7565
rect 1015 7235 1025 7565
rect 675 7225 1025 7235
rect 1100 7150 1150 7650
rect 1225 7565 1575 7575
rect 1225 7235 1235 7565
rect 1565 7235 1575 7565
rect 1225 7225 1575 7235
rect 1650 7150 1700 7650
rect 1775 7565 2125 7575
rect 1775 7235 1785 7565
rect 2115 7235 2125 7565
rect 1775 7225 2125 7235
rect 2200 7150 2250 7650
rect 2325 7565 2675 7575
rect 2325 7235 2335 7565
rect 2665 7235 2675 7565
rect 2325 7225 2675 7235
rect 2750 7150 2800 7650
rect 2875 7565 3225 7575
rect 2875 7235 2885 7565
rect 3215 7235 3225 7565
rect 2875 7225 3225 7235
rect 3300 7150 3350 7650
rect 3425 7565 3775 7575
rect 3425 7235 3435 7565
rect 3765 7235 3775 7565
rect 3425 7225 3775 7235
rect 3850 7150 3900 7650
rect 3975 7565 4325 7575
rect 3975 7235 3985 7565
rect 4315 7235 4325 7565
rect 3975 7225 4325 7235
rect 4400 7150 4450 7650
rect 4525 7565 4875 7575
rect 4525 7235 4535 7565
rect 4865 7235 4875 7565
rect 4525 7225 4875 7235
rect 4950 7150 5000 7650
rect 5075 7565 5425 7575
rect 5075 7235 5085 7565
rect 5415 7235 5425 7565
rect 5075 7225 5425 7235
rect 5500 7150 5550 7650
rect 5625 7565 5975 7575
rect 5625 7235 5635 7565
rect 5965 7235 5975 7565
rect 5625 7225 5975 7235
rect 6050 7150 6100 7650
rect 6175 7565 6525 7575
rect 6175 7235 6185 7565
rect 6515 7235 6525 7565
rect 6175 7225 6525 7235
rect 6600 7150 6650 7650
rect 6725 7565 7075 7575
rect 6725 7235 6735 7565
rect 7065 7235 7075 7565
rect 6725 7225 7075 7235
rect 7150 7150 7200 7650
rect 7275 7565 7625 7575
rect 7275 7235 7285 7565
rect 7615 7235 7625 7565
rect 7275 7225 7625 7235
rect 7700 7150 7750 7650
rect 7825 7565 8175 7575
rect 7825 7235 7835 7565
rect 8165 7235 8175 7565
rect 7825 7225 8175 7235
rect 8250 7150 8300 7650
rect 8375 7565 8725 7575
rect 8375 7235 8385 7565
rect 8715 7235 8725 7565
rect 8375 7225 8725 7235
rect 8800 7150 8850 7650
rect 8925 7565 9275 7575
rect 8925 7235 8935 7565
rect 9265 7235 9275 7565
rect 8925 7225 9275 7235
rect 9350 7150 9400 7650
rect 9475 7565 9825 7575
rect 9475 7235 9485 7565
rect 9815 7235 9825 7565
rect 9475 7225 9825 7235
rect 9900 7150 9950 7650
rect 10025 7565 10375 7575
rect 10025 7235 10035 7565
rect 10365 7235 10375 7565
rect 10025 7225 10375 7235
rect 10450 7150 10500 7650
rect 10575 7565 10925 7575
rect 10575 7235 10585 7565
rect 10915 7235 10925 7565
rect 10575 7225 10925 7235
rect 11000 7150 11050 7650
rect 11125 7565 11475 7575
rect 11125 7235 11135 7565
rect 11465 7235 11475 7565
rect 11125 7225 11475 7235
rect 11550 7150 11600 7650
rect 11675 7565 12025 7575
rect 11675 7235 11685 7565
rect 12015 7235 12025 7565
rect 11675 7225 12025 7235
rect 12100 7150 12150 7650
rect 12225 7565 12575 7575
rect 12225 7235 12235 7565
rect 12565 7235 12575 7565
rect 12225 7225 12575 7235
rect 12650 7150 12700 7650
rect 12775 7565 13125 7575
rect 12775 7235 12785 7565
rect 13115 7235 13125 7565
rect 12775 7225 13125 7235
rect 13200 7150 13250 7650
rect 13325 7565 13675 7575
rect 13325 7235 13335 7565
rect 13665 7235 13675 7565
rect 13325 7225 13675 7235
rect 13750 7150 13975 7650
rect -725 7142 13975 7150
rect -725 7108 -542 7142
rect -508 7108 8 7142
rect 42 7108 558 7142
rect 592 7108 1108 7142
rect 1142 7108 1658 7142
rect 1692 7108 2208 7142
rect 2242 7108 2758 7142
rect 2792 7108 3308 7142
rect 3342 7108 3858 7142
rect 3892 7108 4408 7142
rect 4442 7108 4958 7142
rect 4992 7108 5508 7142
rect 5542 7108 6058 7142
rect 6092 7108 6608 7142
rect 6642 7108 7158 7142
rect 7192 7108 7708 7142
rect 7742 7108 8258 7142
rect 8292 7108 8808 7142
rect 8842 7108 9358 7142
rect 9392 7108 9908 7142
rect 9942 7108 10458 7142
rect 10492 7108 11008 7142
rect 11042 7108 11558 7142
rect 11592 7108 12108 7142
rect 12142 7108 12658 7142
rect 12692 7108 13208 7142
rect 13242 7108 13758 7142
rect 13792 7108 13975 7142
rect -725 7100 13975 7108
rect -725 6600 -500 7100
rect -425 7015 -75 7025
rect -425 6685 -415 7015
rect -85 6685 -75 7015
rect -425 6675 -75 6685
rect 0 6600 50 7100
rect 125 7015 475 7025
rect 125 6685 135 7015
rect 465 6685 475 7015
rect 125 6675 475 6685
rect 550 6600 600 7100
rect 675 7015 1025 7025
rect 675 6685 685 7015
rect 1015 6685 1025 7015
rect 675 6675 1025 6685
rect 1100 6600 1150 7100
rect 1225 7015 1575 7025
rect 1225 6685 1235 7015
rect 1565 6685 1575 7015
rect 1225 6675 1575 6685
rect 1650 6600 1700 7100
rect 1775 7015 2125 7025
rect 1775 6685 1785 7015
rect 2115 6685 2125 7015
rect 1775 6675 2125 6685
rect 2200 6600 2250 7100
rect 2325 7015 2675 7025
rect 2325 6685 2335 7015
rect 2665 6685 2675 7015
rect 2325 6675 2675 6685
rect 2750 6600 2800 7100
rect 2875 7015 3225 7025
rect 2875 6685 2885 7015
rect 3215 6685 3225 7015
rect 2875 6675 3225 6685
rect 3300 6600 3350 7100
rect 3425 7015 3775 7025
rect 3425 6685 3435 7015
rect 3765 6685 3775 7015
rect 3425 6675 3775 6685
rect 3850 6600 3900 7100
rect 3975 7015 4325 7025
rect 3975 6685 3985 7015
rect 4315 6685 4325 7015
rect 3975 6675 4325 6685
rect 4400 6600 4450 7100
rect 4525 7015 4875 7025
rect 4525 6685 4535 7015
rect 4865 6685 4875 7015
rect 4525 6675 4875 6685
rect 4950 6600 5000 7100
rect 5075 7015 5425 7025
rect 5075 6685 5085 7015
rect 5415 6685 5425 7015
rect 5075 6675 5425 6685
rect 5500 6600 5550 7100
rect 5625 7015 5975 7025
rect 5625 6685 5635 7015
rect 5965 6685 5975 7015
rect 5625 6675 5975 6685
rect 6050 6600 6100 7100
rect 6175 7015 6525 7025
rect 6175 6685 6185 7015
rect 6515 6685 6525 7015
rect 6175 6675 6525 6685
rect 6600 6600 6650 7100
rect 6725 7015 7075 7025
rect 6725 6685 6735 7015
rect 7065 6685 7075 7015
rect 6725 6675 7075 6685
rect 7150 6600 7200 7100
rect 7275 7015 7625 7025
rect 7275 6685 7285 7015
rect 7615 6685 7625 7015
rect 7275 6675 7625 6685
rect 7700 6600 7750 7100
rect 7825 7015 8175 7025
rect 7825 6685 7835 7015
rect 8165 6685 8175 7015
rect 7825 6675 8175 6685
rect 8250 6600 8300 7100
rect 8375 7015 8725 7025
rect 8375 6685 8385 7015
rect 8715 6685 8725 7015
rect 8375 6675 8725 6685
rect 8800 6600 8850 7100
rect 8925 7015 9275 7025
rect 8925 6685 8935 7015
rect 9265 6685 9275 7015
rect 8925 6675 9275 6685
rect 9350 6600 9400 7100
rect 9475 7015 9825 7025
rect 9475 6685 9485 7015
rect 9815 6685 9825 7015
rect 9475 6675 9825 6685
rect 9900 6600 9950 7100
rect 10025 7015 10375 7025
rect 10025 6685 10035 7015
rect 10365 6685 10375 7015
rect 10025 6675 10375 6685
rect 10450 6600 10500 7100
rect 10575 7015 10925 7025
rect 10575 6685 10585 7015
rect 10915 6685 10925 7015
rect 10575 6675 10925 6685
rect 11000 6600 11050 7100
rect 11125 7015 11475 7025
rect 11125 6685 11135 7015
rect 11465 6685 11475 7015
rect 11125 6675 11475 6685
rect 11550 6600 11600 7100
rect 11675 7015 12025 7025
rect 11675 6685 11685 7015
rect 12015 6685 12025 7015
rect 11675 6675 12025 6685
rect 12100 6600 12150 7100
rect 12225 7015 12575 7025
rect 12225 6685 12235 7015
rect 12565 6685 12575 7015
rect 12225 6675 12575 6685
rect 12650 6600 12700 7100
rect 12775 7015 13125 7025
rect 12775 6685 12785 7015
rect 13115 6685 13125 7015
rect 12775 6675 13125 6685
rect 13200 6600 13250 7100
rect 13325 7015 13675 7025
rect 13325 6685 13335 7015
rect 13665 6685 13675 7015
rect 13325 6675 13675 6685
rect 13750 6600 13975 7100
rect 14065 6738 14185 6748
rect 14065 6638 14075 6738
rect 14175 6638 14185 6738
rect 14065 6628 14185 6638
rect -725 6592 13975 6600
rect -725 6558 -542 6592
rect -508 6558 8 6592
rect 42 6558 558 6592
rect 592 6558 1108 6592
rect 1142 6558 1658 6592
rect 1692 6558 2208 6592
rect 2242 6558 2758 6592
rect 2792 6558 3308 6592
rect 3342 6558 3858 6592
rect 3892 6558 4408 6592
rect 4442 6558 4958 6592
rect 4992 6558 5508 6592
rect 5542 6558 6058 6592
rect 6092 6558 6608 6592
rect 6642 6558 7158 6592
rect 7192 6558 7708 6592
rect 7742 6558 8258 6592
rect 8292 6558 8808 6592
rect 8842 6558 9358 6592
rect 9392 6558 9908 6592
rect 9942 6558 10458 6592
rect 10492 6558 11008 6592
rect 11042 6558 11558 6592
rect 11592 6558 12108 6592
rect 12142 6558 12658 6592
rect 12692 6558 13208 6592
rect 13242 6558 13758 6592
rect 13792 6558 13975 6592
rect -725 6550 13975 6558
rect -935 6512 -815 6522
rect -935 6412 -925 6512
rect -825 6412 -815 6512
rect -935 6402 -815 6412
rect -725 6050 -500 6550
rect -425 6465 -75 6475
rect -425 6135 -415 6465
rect -85 6135 -75 6465
rect -425 6125 -75 6135
rect 0 6050 50 6550
rect 125 6465 475 6475
rect 125 6135 135 6465
rect 465 6135 475 6465
rect 125 6125 475 6135
rect 550 6050 600 6550
rect 675 6465 1025 6475
rect 675 6135 685 6465
rect 1015 6135 1025 6465
rect 675 6125 1025 6135
rect 1100 6050 1150 6550
rect 1225 6465 1575 6475
rect 1225 6135 1235 6465
rect 1565 6135 1575 6465
rect 1225 6125 1575 6135
rect 1650 6050 1700 6550
rect 1775 6465 2125 6475
rect 1775 6135 1785 6465
rect 2115 6135 2125 6465
rect 1775 6125 2125 6135
rect 2200 6050 2250 6550
rect 2325 6465 2675 6475
rect 2325 6135 2335 6465
rect 2665 6135 2675 6465
rect 2325 6125 2675 6135
rect 2750 6050 2800 6550
rect 2875 6465 3225 6475
rect 2875 6135 2885 6465
rect 3215 6135 3225 6465
rect 2875 6125 3225 6135
rect 3300 6050 3350 6550
rect 3425 6465 3775 6475
rect 3425 6135 3435 6465
rect 3765 6135 3775 6465
rect 3425 6125 3775 6135
rect 3850 6050 3900 6550
rect 3975 6465 4325 6475
rect 3975 6135 3985 6465
rect 4315 6135 4325 6465
rect 3975 6125 4325 6135
rect 4400 6050 4450 6550
rect 4525 6465 4875 6475
rect 4525 6135 4535 6465
rect 4865 6135 4875 6465
rect 4525 6125 4875 6135
rect 4950 6050 5000 6550
rect 5075 6465 5425 6475
rect 5075 6135 5085 6465
rect 5415 6135 5425 6465
rect 5075 6125 5425 6135
rect 5500 6050 5550 6550
rect 5625 6465 5975 6475
rect 5625 6135 5635 6465
rect 5965 6135 5975 6465
rect 5625 6125 5975 6135
rect 6050 6050 6100 6550
rect 6175 6465 6525 6475
rect 6175 6135 6185 6465
rect 6515 6135 6525 6465
rect 6175 6125 6525 6135
rect 6600 6050 6650 6550
rect 6725 6465 7075 6475
rect 6725 6135 6735 6465
rect 7065 6135 7075 6465
rect 6725 6125 7075 6135
rect 7150 6050 7200 6550
rect 7275 6465 7625 6475
rect 7275 6135 7285 6465
rect 7615 6135 7625 6465
rect 7275 6125 7625 6135
rect 7700 6050 7750 6550
rect 7825 6465 8175 6475
rect 7825 6135 7835 6465
rect 8165 6135 8175 6465
rect 7825 6125 8175 6135
rect 8250 6050 8300 6550
rect 8375 6465 8725 6475
rect 8375 6135 8385 6465
rect 8715 6135 8725 6465
rect 8375 6125 8725 6135
rect 8800 6050 8850 6550
rect 8925 6465 9275 6475
rect 8925 6135 8935 6465
rect 9265 6135 9275 6465
rect 8925 6125 9275 6135
rect 9350 6050 9400 6550
rect 9475 6465 9825 6475
rect 9475 6135 9485 6465
rect 9815 6135 9825 6465
rect 9475 6125 9825 6135
rect 9900 6050 9950 6550
rect 10025 6465 10375 6475
rect 10025 6135 10035 6465
rect 10365 6135 10375 6465
rect 10025 6125 10375 6135
rect 10450 6050 10500 6550
rect 10575 6465 10925 6475
rect 10575 6135 10585 6465
rect 10915 6135 10925 6465
rect 10575 6125 10925 6135
rect 11000 6050 11050 6550
rect 11125 6465 11475 6475
rect 11125 6135 11135 6465
rect 11465 6135 11475 6465
rect 11125 6125 11475 6135
rect 11550 6050 11600 6550
rect 11675 6465 12025 6475
rect 11675 6135 11685 6465
rect 12015 6135 12025 6465
rect 11675 6125 12025 6135
rect 12100 6050 12150 6550
rect 12225 6465 12575 6475
rect 12225 6135 12235 6465
rect 12565 6135 12575 6465
rect 12225 6125 12575 6135
rect 12650 6050 12700 6550
rect 12775 6465 13125 6475
rect 12775 6135 12785 6465
rect 13115 6135 13125 6465
rect 12775 6125 13125 6135
rect 13200 6050 13250 6550
rect 13325 6465 13675 6475
rect 13325 6135 13335 6465
rect 13665 6135 13675 6465
rect 13325 6125 13675 6135
rect 13750 6050 13975 6550
rect -725 6042 13975 6050
rect -725 6008 -542 6042
rect -508 6008 8 6042
rect 42 6008 558 6042
rect 592 6008 1108 6042
rect 1142 6008 1658 6042
rect 1692 6008 2208 6042
rect 2242 6008 2758 6042
rect 2792 6008 3308 6042
rect 3342 6008 3858 6042
rect 3892 6008 4408 6042
rect 4442 6008 4958 6042
rect 4992 6008 5508 6042
rect 5542 6008 6058 6042
rect 6092 6008 6608 6042
rect 6642 6008 7158 6042
rect 7192 6008 7708 6042
rect 7742 6008 8258 6042
rect 8292 6008 8808 6042
rect 8842 6008 9358 6042
rect 9392 6008 9908 6042
rect 9942 6008 10458 6042
rect 10492 6008 11008 6042
rect 11042 6008 11558 6042
rect 11592 6008 12108 6042
rect 12142 6008 12658 6042
rect 12692 6008 13208 6042
rect 13242 6008 13758 6042
rect 13792 6008 13975 6042
rect -725 6000 13975 6008
rect -725 5500 -500 6000
rect -425 5915 -75 5925
rect -425 5585 -415 5915
rect -85 5585 -75 5915
rect -425 5575 -75 5585
rect 0 5500 50 6000
rect 125 5915 475 5925
rect 125 5585 135 5915
rect 465 5585 475 5915
rect 125 5575 475 5585
rect 550 5500 600 6000
rect 675 5915 1025 5925
rect 675 5585 685 5915
rect 1015 5585 1025 5915
rect 675 5575 1025 5585
rect 1100 5500 1150 6000
rect 1225 5915 1575 5925
rect 1225 5585 1235 5915
rect 1565 5585 1575 5915
rect 1225 5575 1575 5585
rect 1650 5500 1700 6000
rect 1775 5915 2125 5925
rect 1775 5585 1785 5915
rect 2115 5585 2125 5915
rect 1775 5575 2125 5585
rect 2200 5500 2250 6000
rect 2325 5915 2675 5925
rect 2325 5585 2335 5915
rect 2665 5585 2675 5915
rect 2325 5575 2675 5585
rect 2750 5500 2800 6000
rect 2875 5915 3225 5925
rect 2875 5585 2885 5915
rect 3215 5585 3225 5915
rect 2875 5575 3225 5585
rect 3300 5500 3350 6000
rect 3425 5915 3775 5925
rect 3425 5585 3435 5915
rect 3765 5585 3775 5915
rect 3425 5575 3775 5585
rect 3850 5500 3900 6000
rect 3975 5915 4325 5925
rect 3975 5585 3985 5915
rect 4315 5585 4325 5915
rect 3975 5575 4325 5585
rect 4400 5500 4450 6000
rect 4525 5915 4875 5925
rect 4525 5585 4535 5915
rect 4865 5585 4875 5915
rect 4525 5575 4875 5585
rect 4950 5500 5000 6000
rect 5075 5915 5425 5925
rect 5075 5585 5085 5915
rect 5415 5585 5425 5915
rect 5075 5575 5425 5585
rect 5500 5500 5550 6000
rect 5625 5915 5975 5925
rect 5625 5585 5635 5915
rect 5965 5585 5975 5915
rect 5625 5575 5975 5585
rect 6050 5500 6100 6000
rect 6175 5915 6525 5925
rect 6175 5585 6185 5915
rect 6515 5585 6525 5915
rect 6175 5575 6525 5585
rect 6600 5500 6650 6000
rect 6725 5915 7075 5925
rect 6725 5585 6735 5915
rect 7065 5585 7075 5915
rect 6725 5575 7075 5585
rect 7150 5500 7200 6000
rect 7275 5915 7625 5925
rect 7275 5585 7285 5915
rect 7615 5585 7625 5915
rect 7275 5575 7625 5585
rect 7700 5500 7750 6000
rect 7825 5915 8175 5925
rect 7825 5585 7835 5915
rect 8165 5585 8175 5915
rect 7825 5575 8175 5585
rect 8250 5500 8300 6000
rect 8375 5915 8725 5925
rect 8375 5585 8385 5915
rect 8715 5585 8725 5915
rect 8375 5575 8725 5585
rect 8800 5500 8850 6000
rect 8925 5915 9275 5925
rect 8925 5585 8935 5915
rect 9265 5585 9275 5915
rect 8925 5575 9275 5585
rect 9350 5500 9400 6000
rect 9475 5915 9825 5925
rect 9475 5585 9485 5915
rect 9815 5585 9825 5915
rect 9475 5575 9825 5585
rect 9900 5500 9950 6000
rect 10025 5915 10375 5925
rect 10025 5585 10035 5915
rect 10365 5585 10375 5915
rect 10025 5575 10375 5585
rect 10450 5500 10500 6000
rect 10575 5915 10925 5925
rect 10575 5585 10585 5915
rect 10915 5585 10925 5915
rect 10575 5575 10925 5585
rect 11000 5500 11050 6000
rect 11125 5915 11475 5925
rect 11125 5585 11135 5915
rect 11465 5585 11475 5915
rect 11125 5575 11475 5585
rect 11550 5500 11600 6000
rect 11675 5915 12025 5925
rect 11675 5585 11685 5915
rect 12015 5585 12025 5915
rect 11675 5575 12025 5585
rect 12100 5500 12150 6000
rect 12225 5915 12575 5925
rect 12225 5585 12235 5915
rect 12565 5585 12575 5915
rect 12225 5575 12575 5585
rect 12650 5500 12700 6000
rect 12775 5915 13125 5925
rect 12775 5585 12785 5915
rect 13115 5585 13125 5915
rect 12775 5575 13125 5585
rect 13200 5500 13250 6000
rect 13325 5915 13675 5925
rect 13325 5585 13335 5915
rect 13665 5585 13675 5915
rect 13325 5575 13675 5585
rect 13750 5500 13975 6000
rect 14065 5638 14185 5648
rect 14065 5538 14075 5638
rect 14175 5538 14185 5638
rect 14065 5528 14185 5538
rect -725 5492 13975 5500
rect -725 5458 -542 5492
rect -508 5458 8 5492
rect 42 5458 558 5492
rect 592 5458 1108 5492
rect 1142 5458 1658 5492
rect 1692 5458 2208 5492
rect 2242 5458 2758 5492
rect 2792 5458 3308 5492
rect 3342 5458 3858 5492
rect 3892 5458 4408 5492
rect 4442 5458 4958 5492
rect 4992 5458 5508 5492
rect 5542 5458 6058 5492
rect 6092 5458 6608 5492
rect 6642 5458 7158 5492
rect 7192 5458 7708 5492
rect 7742 5458 8258 5492
rect 8292 5458 8808 5492
rect 8842 5458 9358 5492
rect 9392 5458 9908 5492
rect 9942 5458 10458 5492
rect 10492 5458 11008 5492
rect 11042 5458 11558 5492
rect 11592 5458 12108 5492
rect 12142 5458 12658 5492
rect 12692 5458 13208 5492
rect 13242 5458 13758 5492
rect 13792 5458 13975 5492
rect -725 5450 13975 5458
rect -935 5412 -815 5422
rect -935 5312 -925 5412
rect -825 5312 -815 5412
rect -935 5302 -815 5312
rect -725 4950 -500 5450
rect -425 5365 -75 5375
rect -425 5035 -415 5365
rect -85 5035 -75 5365
rect -425 5025 -75 5035
rect 0 4950 50 5450
rect 125 5365 475 5375
rect 125 5035 135 5365
rect 465 5035 475 5365
rect 125 5025 475 5035
rect 550 4950 600 5450
rect 675 5365 1025 5375
rect 675 5035 685 5365
rect 1015 5035 1025 5365
rect 675 5025 1025 5035
rect 1100 4950 1150 5450
rect 1225 5365 1575 5375
rect 1225 5035 1235 5365
rect 1565 5035 1575 5365
rect 1225 5025 1575 5035
rect 1650 4950 1700 5450
rect 1775 5365 2125 5375
rect 1775 5035 1785 5365
rect 2115 5035 2125 5365
rect 1775 5025 2125 5035
rect 2200 4950 2250 5450
rect 2325 5365 2675 5375
rect 2325 5035 2335 5365
rect 2665 5035 2675 5365
rect 2325 5025 2675 5035
rect 2750 4950 2800 5450
rect 2875 5365 3225 5375
rect 2875 5035 2885 5365
rect 3215 5035 3225 5365
rect 2875 5025 3225 5035
rect 3300 4950 3350 5450
rect 3425 5365 3775 5375
rect 3425 5035 3435 5365
rect 3765 5035 3775 5365
rect 3425 5025 3775 5035
rect 3850 4950 3900 5450
rect 3975 5365 4325 5375
rect 3975 5035 3985 5365
rect 4315 5035 4325 5365
rect 3975 5025 4325 5035
rect 4400 4950 4450 5450
rect 4525 5365 4875 5375
rect 4525 5035 4535 5365
rect 4865 5035 4875 5365
rect 4525 5025 4875 5035
rect 4950 4950 5000 5450
rect 5075 5365 5425 5375
rect 5075 5035 5085 5365
rect 5415 5035 5425 5365
rect 5075 5025 5425 5035
rect 5500 4950 5550 5450
rect 5625 5365 5975 5375
rect 5625 5035 5635 5365
rect 5965 5035 5975 5365
rect 5625 5025 5975 5035
rect 6050 4950 6100 5450
rect 6175 5365 6525 5375
rect 6175 5035 6185 5365
rect 6515 5035 6525 5365
rect 6175 5025 6525 5035
rect 6600 4950 6650 5450
rect 6725 5365 7075 5375
rect 6725 5035 6735 5365
rect 7065 5035 7075 5365
rect 6725 5025 7075 5035
rect 7150 4950 7200 5450
rect 7275 5365 7625 5375
rect 7275 5035 7285 5365
rect 7615 5035 7625 5365
rect 7275 5025 7625 5035
rect 7700 4950 7750 5450
rect 7825 5365 8175 5375
rect 7825 5035 7835 5365
rect 8165 5035 8175 5365
rect 7825 5025 8175 5035
rect 8250 4950 8300 5450
rect 8375 5365 8725 5375
rect 8375 5035 8385 5365
rect 8715 5035 8725 5365
rect 8375 5025 8725 5035
rect 8800 4950 8850 5450
rect 8925 5365 9275 5375
rect 8925 5035 8935 5365
rect 9265 5035 9275 5365
rect 8925 5025 9275 5035
rect 9350 4950 9400 5450
rect 9475 5365 9825 5375
rect 9475 5035 9485 5365
rect 9815 5035 9825 5365
rect 9475 5025 9825 5035
rect 9900 4950 9950 5450
rect 10025 5365 10375 5375
rect 10025 5035 10035 5365
rect 10365 5035 10375 5365
rect 10025 5025 10375 5035
rect 10450 4950 10500 5450
rect 10575 5365 10925 5375
rect 10575 5035 10585 5365
rect 10915 5035 10925 5365
rect 10575 5025 10925 5035
rect 11000 4950 11050 5450
rect 11125 5365 11475 5375
rect 11125 5035 11135 5365
rect 11465 5035 11475 5365
rect 11125 5025 11475 5035
rect 11550 4950 11600 5450
rect 11675 5365 12025 5375
rect 11675 5035 11685 5365
rect 12015 5035 12025 5365
rect 11675 5025 12025 5035
rect 12100 4950 12150 5450
rect 12225 5365 12575 5375
rect 12225 5035 12235 5365
rect 12565 5035 12575 5365
rect 12225 5025 12575 5035
rect 12650 4950 12700 5450
rect 12775 5365 13125 5375
rect 12775 5035 12785 5365
rect 13115 5035 13125 5365
rect 12775 5025 13125 5035
rect 13200 4950 13250 5450
rect 13325 5365 13675 5375
rect 13325 5035 13335 5365
rect 13665 5035 13675 5365
rect 13325 5025 13675 5035
rect 13750 4950 13975 5450
rect -725 4942 13975 4950
rect -725 4908 -542 4942
rect -508 4908 8 4942
rect 42 4908 558 4942
rect 592 4908 1108 4942
rect 1142 4908 1658 4942
rect 1692 4908 2208 4942
rect 2242 4908 2758 4942
rect 2792 4908 3308 4942
rect 3342 4908 3858 4942
rect 3892 4908 4408 4942
rect 4442 4908 4958 4942
rect 4992 4908 5508 4942
rect 5542 4908 6058 4942
rect 6092 4908 6608 4942
rect 6642 4908 7158 4942
rect 7192 4908 7708 4942
rect 7742 4908 8258 4942
rect 8292 4908 8808 4942
rect 8842 4908 9358 4942
rect 9392 4908 9908 4942
rect 9942 4908 10458 4942
rect 10492 4908 11008 4942
rect 11042 4908 11558 4942
rect 11592 4908 12108 4942
rect 12142 4908 12658 4942
rect 12692 4908 13208 4942
rect 13242 4908 13758 4942
rect 13792 4908 13975 4942
rect -725 4900 13975 4908
rect -725 4400 -500 4900
rect -425 4815 -75 4825
rect -425 4485 -415 4815
rect -85 4485 -75 4815
rect -425 4475 -75 4485
rect 0 4400 50 4900
rect 125 4815 475 4825
rect 125 4485 135 4815
rect 465 4485 475 4815
rect 125 4475 475 4485
rect 550 4400 600 4900
rect 675 4815 1025 4825
rect 675 4485 685 4815
rect 1015 4485 1025 4815
rect 675 4475 1025 4485
rect 1100 4400 1150 4900
rect 1225 4815 1575 4825
rect 1225 4485 1235 4815
rect 1565 4485 1575 4815
rect 1225 4475 1575 4485
rect 1650 4400 1700 4900
rect 1775 4815 2125 4825
rect 1775 4485 1785 4815
rect 2115 4485 2125 4815
rect 1775 4475 2125 4485
rect 2200 4400 2250 4900
rect 2325 4815 2675 4825
rect 2325 4485 2335 4815
rect 2665 4485 2675 4815
rect 2325 4475 2675 4485
rect 2750 4400 2800 4900
rect 2875 4815 3225 4825
rect 2875 4485 2885 4815
rect 3215 4485 3225 4815
rect 2875 4475 3225 4485
rect 3300 4400 3350 4900
rect 3425 4815 3775 4825
rect 3425 4485 3435 4815
rect 3765 4485 3775 4815
rect 3425 4475 3775 4485
rect 3850 4400 3900 4900
rect 3975 4815 4325 4825
rect 3975 4485 3985 4815
rect 4315 4485 4325 4815
rect 3975 4475 4325 4485
rect 4400 4400 4450 4900
rect 4525 4815 4875 4825
rect 4525 4485 4535 4815
rect 4865 4485 4875 4815
rect 4525 4475 4875 4485
rect 4950 4400 5000 4900
rect 5075 4815 5425 4825
rect 5075 4485 5085 4815
rect 5415 4485 5425 4815
rect 5075 4475 5425 4485
rect 5500 4400 5550 4900
rect 5625 4815 5975 4825
rect 5625 4485 5635 4815
rect 5965 4485 5975 4815
rect 5625 4475 5975 4485
rect 6050 4400 6100 4900
rect 6175 4815 6525 4825
rect 6175 4485 6185 4815
rect 6515 4485 6525 4815
rect 6175 4475 6525 4485
rect 6600 4400 6650 4900
rect 6725 4815 7075 4825
rect 6725 4485 6735 4815
rect 7065 4485 7075 4815
rect 6725 4475 7075 4485
rect 7150 4400 7200 4900
rect 7275 4815 7625 4825
rect 7275 4485 7285 4815
rect 7615 4485 7625 4815
rect 7275 4475 7625 4485
rect 7700 4400 7750 4900
rect 7825 4815 8175 4825
rect 7825 4485 7835 4815
rect 8165 4485 8175 4815
rect 7825 4475 8175 4485
rect 8250 4400 8300 4900
rect 8375 4815 8725 4825
rect 8375 4485 8385 4815
rect 8715 4485 8725 4815
rect 8375 4475 8725 4485
rect 8800 4400 8850 4900
rect 8925 4815 9275 4825
rect 8925 4485 8935 4815
rect 9265 4485 9275 4815
rect 8925 4475 9275 4485
rect 9350 4400 9400 4900
rect 9475 4815 9825 4825
rect 9475 4485 9485 4815
rect 9815 4485 9825 4815
rect 9475 4475 9825 4485
rect 9900 4400 9950 4900
rect 10025 4815 10375 4825
rect 10025 4485 10035 4815
rect 10365 4485 10375 4815
rect 10025 4475 10375 4485
rect 10450 4400 10500 4900
rect 10575 4815 10925 4825
rect 10575 4485 10585 4815
rect 10915 4485 10925 4815
rect 10575 4475 10925 4485
rect 11000 4400 11050 4900
rect 11125 4815 11475 4825
rect 11125 4485 11135 4815
rect 11465 4485 11475 4815
rect 11125 4475 11475 4485
rect 11550 4400 11600 4900
rect 11675 4815 12025 4825
rect 11675 4485 11685 4815
rect 12015 4485 12025 4815
rect 11675 4475 12025 4485
rect 12100 4400 12150 4900
rect 12225 4815 12575 4825
rect 12225 4485 12235 4815
rect 12565 4485 12575 4815
rect 12225 4475 12575 4485
rect 12650 4400 12700 4900
rect 12775 4815 13125 4825
rect 12775 4485 12785 4815
rect 13115 4485 13125 4815
rect 12775 4475 13125 4485
rect 13200 4400 13250 4900
rect 13325 4815 13675 4825
rect 13325 4485 13335 4815
rect 13665 4485 13675 4815
rect 13325 4475 13675 4485
rect 13750 4400 13975 4900
rect 14065 4538 14185 4548
rect 14065 4438 14075 4538
rect 14175 4438 14185 4538
rect 14065 4428 14185 4438
rect -725 4392 13975 4400
rect -725 4358 -542 4392
rect -508 4358 8 4392
rect 42 4358 558 4392
rect 592 4358 1108 4392
rect 1142 4358 1658 4392
rect 1692 4358 2208 4392
rect 2242 4358 2758 4392
rect 2792 4358 3308 4392
rect 3342 4358 3858 4392
rect 3892 4358 4408 4392
rect 4442 4358 4958 4392
rect 4992 4358 5508 4392
rect 5542 4358 6058 4392
rect 6092 4358 6608 4392
rect 6642 4358 7158 4392
rect 7192 4358 7708 4392
rect 7742 4358 8258 4392
rect 8292 4358 8808 4392
rect 8842 4358 9358 4392
rect 9392 4358 9908 4392
rect 9942 4358 10458 4392
rect 10492 4358 11008 4392
rect 11042 4358 11558 4392
rect 11592 4358 12108 4392
rect 12142 4358 12658 4392
rect 12692 4358 13208 4392
rect 13242 4358 13758 4392
rect 13792 4358 13975 4392
rect -725 4350 13975 4358
rect -935 4312 -815 4322
rect -935 4212 -925 4312
rect -825 4212 -815 4312
rect -935 4202 -815 4212
rect -725 3850 -500 4350
rect -425 4265 -75 4275
rect -425 3935 -415 4265
rect -85 3935 -75 4265
rect -425 3925 -75 3935
rect 0 3850 50 4350
rect 125 4265 475 4275
rect 125 3935 135 4265
rect 465 3935 475 4265
rect 125 3925 475 3935
rect 550 3850 600 4350
rect 675 4265 1025 4275
rect 675 3935 685 4265
rect 1015 3935 1025 4265
rect 675 3925 1025 3935
rect 1100 3850 1150 4350
rect 1225 4265 1575 4275
rect 1225 3935 1235 4265
rect 1565 3935 1575 4265
rect 1225 3925 1575 3935
rect 1650 3850 1700 4350
rect 1775 4265 2125 4275
rect 1775 3935 1785 4265
rect 2115 3935 2125 4265
rect 1775 3925 2125 3935
rect 2200 3850 2250 4350
rect 2325 4265 2675 4275
rect 2325 3935 2335 4265
rect 2665 3935 2675 4265
rect 2325 3925 2675 3935
rect 2750 3850 2800 4350
rect 2875 4265 3225 4275
rect 2875 3935 2885 4265
rect 3215 3935 3225 4265
rect 2875 3925 3225 3935
rect 3300 3850 3350 4350
rect 3425 4265 3775 4275
rect 3425 3935 3435 4265
rect 3765 3935 3775 4265
rect 3425 3925 3775 3935
rect 3850 3850 3900 4350
rect 3975 4265 4325 4275
rect 3975 3935 3985 4265
rect 4315 3935 4325 4265
rect 3975 3925 4325 3935
rect 4400 3850 4450 4350
rect 4525 4265 4875 4275
rect 4525 3935 4535 4265
rect 4865 3935 4875 4265
rect 4525 3925 4875 3935
rect 4950 3850 5000 4350
rect 5075 4265 5425 4275
rect 5075 3935 5085 4265
rect 5415 3935 5425 4265
rect 5075 3925 5425 3935
rect 5500 3850 5550 4350
rect 5625 4265 5975 4275
rect 5625 3935 5635 4265
rect 5965 3935 5975 4265
rect 5625 3925 5975 3935
rect 6050 3850 6100 4350
rect 6175 4265 6525 4275
rect 6175 3935 6185 4265
rect 6515 3935 6525 4265
rect 6175 3925 6525 3935
rect 6600 3850 6650 4350
rect 6725 4265 7075 4275
rect 6725 3935 6735 4265
rect 7065 3935 7075 4265
rect 6725 3925 7075 3935
rect 7150 3850 7200 4350
rect 7275 4265 7625 4275
rect 7275 3935 7285 4265
rect 7615 3935 7625 4265
rect 7275 3925 7625 3935
rect 7700 3850 7750 4350
rect 7825 4265 8175 4275
rect 7825 3935 7835 4265
rect 8165 3935 8175 4265
rect 7825 3925 8175 3935
rect 8250 3850 8300 4350
rect 8375 4265 8725 4275
rect 8375 3935 8385 4265
rect 8715 3935 8725 4265
rect 8375 3925 8725 3935
rect 8800 3850 8850 4350
rect 8925 4265 9275 4275
rect 8925 3935 8935 4265
rect 9265 3935 9275 4265
rect 8925 3925 9275 3935
rect 9350 3850 9400 4350
rect 9475 4265 9825 4275
rect 9475 3935 9485 4265
rect 9815 3935 9825 4265
rect 9475 3925 9825 3935
rect 9900 3850 9950 4350
rect 10025 4265 10375 4275
rect 10025 3935 10035 4265
rect 10365 3935 10375 4265
rect 10025 3925 10375 3935
rect 10450 3850 10500 4350
rect 10575 4265 10925 4275
rect 10575 3935 10585 4265
rect 10915 3935 10925 4265
rect 10575 3925 10925 3935
rect 11000 3850 11050 4350
rect 11125 4265 11475 4275
rect 11125 3935 11135 4265
rect 11465 3935 11475 4265
rect 11125 3925 11475 3935
rect 11550 3850 11600 4350
rect 11675 4265 12025 4275
rect 11675 3935 11685 4265
rect 12015 3935 12025 4265
rect 11675 3925 12025 3935
rect 12100 3850 12150 4350
rect 12225 4265 12575 4275
rect 12225 3935 12235 4265
rect 12565 3935 12575 4265
rect 12225 3925 12575 3935
rect 12650 3850 12700 4350
rect 12775 4265 13125 4275
rect 12775 3935 12785 4265
rect 13115 3935 13125 4265
rect 12775 3925 13125 3935
rect 13200 3850 13250 4350
rect 13325 4265 13675 4275
rect 13325 3935 13335 4265
rect 13665 3935 13675 4265
rect 13325 3925 13675 3935
rect 13750 3850 13975 4350
rect -725 3842 13975 3850
rect -725 3808 -542 3842
rect -508 3808 8 3842
rect 42 3808 558 3842
rect 592 3808 1108 3842
rect 1142 3808 1658 3842
rect 1692 3808 2208 3842
rect 2242 3808 2758 3842
rect 2792 3808 3308 3842
rect 3342 3808 3858 3842
rect 3892 3808 4408 3842
rect 4442 3808 4958 3842
rect 4992 3808 5508 3842
rect 5542 3808 6058 3842
rect 6092 3808 6608 3842
rect 6642 3808 7158 3842
rect 7192 3808 7708 3842
rect 7742 3808 8258 3842
rect 8292 3808 8808 3842
rect 8842 3808 9358 3842
rect 9392 3808 9908 3842
rect 9942 3808 10458 3842
rect 10492 3808 11008 3842
rect 11042 3808 11558 3842
rect 11592 3808 12108 3842
rect 12142 3808 12658 3842
rect 12692 3808 13208 3842
rect 13242 3808 13758 3842
rect 13792 3808 13975 3842
rect -725 3800 13975 3808
rect -725 3300 -500 3800
rect -425 3715 -75 3725
rect -425 3385 -415 3715
rect -85 3385 -75 3715
rect -425 3375 -75 3385
rect 0 3300 50 3800
rect 125 3715 475 3725
rect 125 3385 135 3715
rect 465 3385 475 3715
rect 125 3375 475 3385
rect 550 3300 600 3800
rect 675 3715 1025 3725
rect 675 3385 685 3715
rect 1015 3385 1025 3715
rect 675 3375 1025 3385
rect 1100 3300 1150 3800
rect 1225 3715 1575 3725
rect 1225 3385 1235 3715
rect 1565 3385 1575 3715
rect 1225 3375 1575 3385
rect 1650 3300 1700 3800
rect 1775 3715 2125 3725
rect 1775 3385 1785 3715
rect 2115 3385 2125 3715
rect 1775 3375 2125 3385
rect 2200 3300 2250 3800
rect 2325 3715 2675 3725
rect 2325 3385 2335 3715
rect 2665 3385 2675 3715
rect 2325 3375 2675 3385
rect 2750 3300 2800 3800
rect 2875 3715 3225 3725
rect 2875 3385 2885 3715
rect 3215 3385 3225 3715
rect 2875 3375 3225 3385
rect 3300 3300 3350 3800
rect 3425 3715 3775 3725
rect 3425 3385 3435 3715
rect 3765 3385 3775 3715
rect 3425 3375 3775 3385
rect 3850 3300 3900 3800
rect 3975 3715 4325 3725
rect 3975 3385 3985 3715
rect 4315 3385 4325 3715
rect 3975 3375 4325 3385
rect 4400 3300 4450 3800
rect 4525 3715 4875 3725
rect 4525 3385 4535 3715
rect 4865 3385 4875 3715
rect 4525 3375 4875 3385
rect 4950 3300 5000 3800
rect 5075 3715 5425 3725
rect 5075 3385 5085 3715
rect 5415 3385 5425 3715
rect 5075 3375 5425 3385
rect 5500 3300 5550 3800
rect 5625 3715 5975 3725
rect 5625 3385 5635 3715
rect 5965 3385 5975 3715
rect 5625 3375 5975 3385
rect 6050 3300 6100 3800
rect 6175 3715 6525 3725
rect 6175 3385 6185 3715
rect 6515 3385 6525 3715
rect 6175 3375 6525 3385
rect 6600 3300 6650 3800
rect 6725 3715 7075 3725
rect 6725 3385 6735 3715
rect 7065 3385 7075 3715
rect 6725 3375 7075 3385
rect 7150 3300 7200 3800
rect 7275 3715 7625 3725
rect 7275 3385 7285 3715
rect 7615 3385 7625 3715
rect 7275 3375 7625 3385
rect 7700 3300 7750 3800
rect 7825 3715 8175 3725
rect 7825 3385 7835 3715
rect 8165 3385 8175 3715
rect 7825 3375 8175 3385
rect 8250 3300 8300 3800
rect 8375 3715 8725 3725
rect 8375 3385 8385 3715
rect 8715 3385 8725 3715
rect 8375 3375 8725 3385
rect 8800 3300 8850 3800
rect 8925 3715 9275 3725
rect 8925 3385 8935 3715
rect 9265 3385 9275 3715
rect 8925 3375 9275 3385
rect 9350 3300 9400 3800
rect 9475 3715 9825 3725
rect 9475 3385 9485 3715
rect 9815 3385 9825 3715
rect 9475 3375 9825 3385
rect 9900 3300 9950 3800
rect 10025 3715 10375 3725
rect 10025 3385 10035 3715
rect 10365 3385 10375 3715
rect 10025 3375 10375 3385
rect 10450 3300 10500 3800
rect 10575 3715 10925 3725
rect 10575 3385 10585 3715
rect 10915 3385 10925 3715
rect 10575 3375 10925 3385
rect 11000 3300 11050 3800
rect 11125 3715 11475 3725
rect 11125 3385 11135 3715
rect 11465 3385 11475 3715
rect 11125 3375 11475 3385
rect 11550 3300 11600 3800
rect 11675 3715 12025 3725
rect 11675 3385 11685 3715
rect 12015 3385 12025 3715
rect 11675 3375 12025 3385
rect 12100 3300 12150 3800
rect 12225 3715 12575 3725
rect 12225 3385 12235 3715
rect 12565 3385 12575 3715
rect 12225 3375 12575 3385
rect 12650 3300 12700 3800
rect 12775 3715 13125 3725
rect 12775 3385 12785 3715
rect 13115 3385 13125 3715
rect 12775 3375 13125 3385
rect 13200 3300 13250 3800
rect 13325 3715 13675 3725
rect 13325 3385 13335 3715
rect 13665 3385 13675 3715
rect 13325 3375 13675 3385
rect 13750 3300 13975 3800
rect 14065 3438 14185 3448
rect 14065 3338 14075 3438
rect 14175 3338 14185 3438
rect 14065 3328 14185 3338
rect -725 3292 13975 3300
rect -725 3258 -542 3292
rect -508 3258 8 3292
rect 42 3258 558 3292
rect 592 3258 1108 3292
rect 1142 3258 1658 3292
rect 1692 3258 2208 3292
rect 2242 3258 2758 3292
rect 2792 3258 3308 3292
rect 3342 3258 3858 3292
rect 3892 3258 4408 3292
rect 4442 3258 4958 3292
rect 4992 3258 5508 3292
rect 5542 3258 6058 3292
rect 6092 3258 6608 3292
rect 6642 3258 7158 3292
rect 7192 3258 7708 3292
rect 7742 3258 8258 3292
rect 8292 3258 8808 3292
rect 8842 3258 9358 3292
rect 9392 3258 9908 3292
rect 9942 3258 10458 3292
rect 10492 3258 11008 3292
rect 11042 3258 11558 3292
rect 11592 3258 12108 3292
rect 12142 3258 12658 3292
rect 12692 3258 13208 3292
rect 13242 3258 13758 3292
rect 13792 3258 13975 3292
rect -725 3250 13975 3258
rect -935 3212 -815 3222
rect -935 3112 -925 3212
rect -825 3112 -815 3212
rect -935 3102 -815 3112
rect -725 2750 -500 3250
rect -425 3165 -75 3175
rect -425 2835 -415 3165
rect -85 2835 -75 3165
rect -425 2825 -75 2835
rect 0 2750 50 3250
rect 125 3165 475 3175
rect 125 2835 135 3165
rect 465 2835 475 3165
rect 125 2825 475 2835
rect 550 2750 600 3250
rect 675 3165 1025 3175
rect 675 2835 685 3165
rect 1015 2835 1025 3165
rect 675 2825 1025 2835
rect 1100 2750 1150 3250
rect 1225 3165 1575 3175
rect 1225 2835 1235 3165
rect 1565 2835 1575 3165
rect 1225 2825 1575 2835
rect 1650 2750 1700 3250
rect 1775 3165 2125 3175
rect 1775 2835 1785 3165
rect 2115 2835 2125 3165
rect 1775 2825 2125 2835
rect 2200 2750 2250 3250
rect 2325 3165 2675 3175
rect 2325 2835 2335 3165
rect 2665 2835 2675 3165
rect 2325 2825 2675 2835
rect 2750 2750 2800 3250
rect 2875 3165 3225 3175
rect 2875 2835 2885 3165
rect 3215 2835 3225 3165
rect 2875 2825 3225 2835
rect 3300 2750 3350 3250
rect 3425 3165 3775 3175
rect 3425 2835 3435 3165
rect 3765 2835 3775 3165
rect 3425 2825 3775 2835
rect 3850 2750 3900 3250
rect 3975 3165 4325 3175
rect 3975 2835 3985 3165
rect 4315 2835 4325 3165
rect 3975 2825 4325 2835
rect 4400 2750 4450 3250
rect 4525 3165 4875 3175
rect 4525 2835 4535 3165
rect 4865 2835 4875 3165
rect 4525 2825 4875 2835
rect 4950 2750 5000 3250
rect 5075 3165 5425 3175
rect 5075 2835 5085 3165
rect 5415 2835 5425 3165
rect 5075 2825 5425 2835
rect 5500 2750 5550 3250
rect 5625 3165 5975 3175
rect 5625 2835 5635 3165
rect 5965 2835 5975 3165
rect 5625 2825 5975 2835
rect 6050 2750 6100 3250
rect 6175 3165 6525 3175
rect 6175 2835 6185 3165
rect 6515 2835 6525 3165
rect 6175 2825 6525 2835
rect 6600 2750 6650 3250
rect 6725 3165 7075 3175
rect 6725 2835 6735 3165
rect 7065 2835 7075 3165
rect 6725 2825 7075 2835
rect 7150 2750 7200 3250
rect 7275 3165 7625 3175
rect 7275 2835 7285 3165
rect 7615 2835 7625 3165
rect 7275 2825 7625 2835
rect 7700 2750 7750 3250
rect 7825 3165 8175 3175
rect 7825 2835 7835 3165
rect 8165 2835 8175 3165
rect 7825 2825 8175 2835
rect 8250 2750 8300 3250
rect 8375 3165 8725 3175
rect 8375 2835 8385 3165
rect 8715 2835 8725 3165
rect 8375 2825 8725 2835
rect 8800 2750 8850 3250
rect 8925 3165 9275 3175
rect 8925 2835 8935 3165
rect 9265 2835 9275 3165
rect 8925 2825 9275 2835
rect 9350 2750 9400 3250
rect 9475 3165 9825 3175
rect 9475 2835 9485 3165
rect 9815 2835 9825 3165
rect 9475 2825 9825 2835
rect 9900 2750 9950 3250
rect 10025 3165 10375 3175
rect 10025 2835 10035 3165
rect 10365 2835 10375 3165
rect 10025 2825 10375 2835
rect 10450 2750 10500 3250
rect 10575 3165 10925 3175
rect 10575 2835 10585 3165
rect 10915 2835 10925 3165
rect 10575 2825 10925 2835
rect 11000 2750 11050 3250
rect 11125 3165 11475 3175
rect 11125 2835 11135 3165
rect 11465 2835 11475 3165
rect 11125 2825 11475 2835
rect 11550 2750 11600 3250
rect 11675 3165 12025 3175
rect 11675 2835 11685 3165
rect 12015 2835 12025 3165
rect 11675 2825 12025 2835
rect 12100 2750 12150 3250
rect 12225 3165 12575 3175
rect 12225 2835 12235 3165
rect 12565 2835 12575 3165
rect 12225 2825 12575 2835
rect 12650 2750 12700 3250
rect 12775 3165 13125 3175
rect 12775 2835 12785 3165
rect 13115 2835 13125 3165
rect 12775 2825 13125 2835
rect 13200 2750 13250 3250
rect 13325 3165 13675 3175
rect 13325 2835 13335 3165
rect 13665 2835 13675 3165
rect 13325 2825 13675 2835
rect 13750 2750 13975 3250
rect -725 2742 13975 2750
rect -725 2708 -542 2742
rect -508 2708 8 2742
rect 42 2708 558 2742
rect 592 2708 1108 2742
rect 1142 2708 1658 2742
rect 1692 2708 2208 2742
rect 2242 2708 2758 2742
rect 2792 2708 3308 2742
rect 3342 2708 3858 2742
rect 3892 2708 4408 2742
rect 4442 2708 4958 2742
rect 4992 2708 5508 2742
rect 5542 2708 6058 2742
rect 6092 2708 6608 2742
rect 6642 2708 7158 2742
rect 7192 2708 7708 2742
rect 7742 2708 8258 2742
rect 8292 2708 8808 2742
rect 8842 2708 9358 2742
rect 9392 2708 9908 2742
rect 9942 2708 10458 2742
rect 10492 2708 11008 2742
rect 11042 2708 11558 2742
rect 11592 2708 12108 2742
rect 12142 2708 12658 2742
rect 12692 2708 13208 2742
rect 13242 2708 13758 2742
rect 13792 2708 13975 2742
rect -725 2700 13975 2708
rect -725 2200 -500 2700
rect -425 2615 -75 2625
rect -425 2285 -415 2615
rect -85 2285 -75 2615
rect -425 2275 -75 2285
rect 0 2200 50 2700
rect 125 2615 475 2625
rect 125 2285 135 2615
rect 465 2285 475 2615
rect 125 2275 475 2285
rect 550 2200 600 2700
rect 675 2615 1025 2625
rect 675 2285 685 2615
rect 1015 2285 1025 2615
rect 675 2275 1025 2285
rect 1100 2200 1150 2700
rect 1225 2615 1575 2625
rect 1225 2285 1235 2615
rect 1565 2285 1575 2615
rect 1225 2275 1575 2285
rect 1650 2200 1700 2700
rect 1775 2615 2125 2625
rect 1775 2285 1785 2615
rect 2115 2285 2125 2615
rect 1775 2275 2125 2285
rect 2200 2200 2250 2700
rect 2325 2615 2675 2625
rect 2325 2285 2335 2615
rect 2665 2285 2675 2615
rect 2325 2275 2675 2285
rect 2750 2200 2800 2700
rect 2875 2615 3225 2625
rect 2875 2285 2885 2615
rect 3215 2285 3225 2615
rect 2875 2275 3225 2285
rect 3300 2200 3350 2700
rect 3425 2615 3775 2625
rect 3425 2285 3435 2615
rect 3765 2285 3775 2615
rect 3425 2275 3775 2285
rect 3850 2200 3900 2700
rect 3975 2615 4325 2625
rect 3975 2285 3985 2615
rect 4315 2285 4325 2615
rect 3975 2275 4325 2285
rect 4400 2200 4450 2700
rect 4525 2615 4875 2625
rect 4525 2285 4535 2615
rect 4865 2285 4875 2615
rect 4525 2275 4875 2285
rect 4950 2200 5000 2700
rect 5075 2615 5425 2625
rect 5075 2285 5085 2615
rect 5415 2285 5425 2615
rect 5075 2275 5425 2285
rect 5500 2200 5550 2700
rect 5625 2615 5975 2625
rect 5625 2285 5635 2615
rect 5965 2285 5975 2615
rect 5625 2275 5975 2285
rect 6050 2200 6100 2700
rect 6175 2615 6525 2625
rect 6175 2285 6185 2615
rect 6515 2285 6525 2615
rect 6175 2275 6525 2285
rect 6600 2200 6650 2700
rect 6725 2615 7075 2625
rect 6725 2285 6735 2615
rect 7065 2285 7075 2615
rect 6725 2275 7075 2285
rect 7150 2200 7200 2700
rect 7275 2615 7625 2625
rect 7275 2285 7285 2615
rect 7615 2285 7625 2615
rect 7275 2275 7625 2285
rect 7700 2200 7750 2700
rect 7825 2615 8175 2625
rect 7825 2285 7835 2615
rect 8165 2285 8175 2615
rect 7825 2275 8175 2285
rect 8250 2200 8300 2700
rect 8375 2615 8725 2625
rect 8375 2285 8385 2615
rect 8715 2285 8725 2615
rect 8375 2275 8725 2285
rect 8800 2200 8850 2700
rect 8925 2615 9275 2625
rect 8925 2285 8935 2615
rect 9265 2285 9275 2615
rect 8925 2275 9275 2285
rect 9350 2200 9400 2700
rect 9475 2615 9825 2625
rect 9475 2285 9485 2615
rect 9815 2285 9825 2615
rect 9475 2275 9825 2285
rect 9900 2200 9950 2700
rect 10025 2615 10375 2625
rect 10025 2285 10035 2615
rect 10365 2285 10375 2615
rect 10025 2275 10375 2285
rect 10450 2200 10500 2700
rect 10575 2615 10925 2625
rect 10575 2285 10585 2615
rect 10915 2285 10925 2615
rect 10575 2275 10925 2285
rect 11000 2200 11050 2700
rect 11125 2615 11475 2625
rect 11125 2285 11135 2615
rect 11465 2285 11475 2615
rect 11125 2275 11475 2285
rect 11550 2200 11600 2700
rect 11675 2615 12025 2625
rect 11675 2285 11685 2615
rect 12015 2285 12025 2615
rect 11675 2275 12025 2285
rect 12100 2200 12150 2700
rect 12225 2615 12575 2625
rect 12225 2285 12235 2615
rect 12565 2285 12575 2615
rect 12225 2275 12575 2285
rect 12650 2200 12700 2700
rect 12775 2615 13125 2625
rect 12775 2285 12785 2615
rect 13115 2285 13125 2615
rect 12775 2275 13125 2285
rect 13200 2200 13250 2700
rect 13325 2615 13675 2625
rect 13325 2285 13335 2615
rect 13665 2285 13675 2615
rect 13325 2275 13675 2285
rect 13750 2200 13975 2700
rect 14065 2338 14185 2348
rect 14065 2238 14075 2338
rect 14175 2238 14185 2338
rect 14065 2228 14185 2238
rect -725 2192 13975 2200
rect -725 2158 -542 2192
rect -508 2158 8 2192
rect 42 2158 558 2192
rect 592 2158 1108 2192
rect 1142 2158 1658 2192
rect 1692 2158 2208 2192
rect 2242 2158 2758 2192
rect 2792 2158 3308 2192
rect 3342 2158 3858 2192
rect 3892 2158 4408 2192
rect 4442 2158 4958 2192
rect 4992 2158 5508 2192
rect 5542 2158 6058 2192
rect 6092 2158 6608 2192
rect 6642 2158 7158 2192
rect 7192 2158 7708 2192
rect 7742 2158 8258 2192
rect 8292 2158 8808 2192
rect 8842 2158 9358 2192
rect 9392 2158 9908 2192
rect 9942 2158 10458 2192
rect 10492 2158 11008 2192
rect 11042 2158 11558 2192
rect 11592 2158 12108 2192
rect 12142 2158 12658 2192
rect 12692 2158 13208 2192
rect 13242 2158 13758 2192
rect 13792 2158 13975 2192
rect -725 2150 13975 2158
rect -935 2112 -815 2122
rect -935 2012 -925 2112
rect -825 2012 -815 2112
rect -935 2002 -815 2012
rect -725 1650 -500 2150
rect -425 2065 -75 2075
rect -425 1735 -415 2065
rect -85 1735 -75 2065
rect -425 1725 -75 1735
rect 0 1650 50 2150
rect 125 2065 475 2075
rect 125 1735 135 2065
rect 465 1735 475 2065
rect 125 1725 475 1735
rect 550 1650 600 2150
rect 675 2065 1025 2075
rect 675 1735 685 2065
rect 1015 1735 1025 2065
rect 675 1725 1025 1735
rect 1100 1650 1150 2150
rect 1225 2065 1575 2075
rect 1225 1735 1235 2065
rect 1565 1735 1575 2065
rect 1225 1725 1575 1735
rect 1650 1650 1700 2150
rect 1775 2065 2125 2075
rect 1775 1735 1785 2065
rect 2115 1735 2125 2065
rect 1775 1725 2125 1735
rect 2200 1650 2250 2150
rect 2325 2065 2675 2075
rect 2325 1735 2335 2065
rect 2665 1735 2675 2065
rect 2325 1725 2675 1735
rect 2750 1650 2800 2150
rect 2875 2065 3225 2075
rect 2875 1735 2885 2065
rect 3215 1735 3225 2065
rect 2875 1725 3225 1735
rect 3300 1650 3350 2150
rect 3425 2065 3775 2075
rect 3425 1735 3435 2065
rect 3765 1735 3775 2065
rect 3425 1725 3775 1735
rect 3850 1650 3900 2150
rect 3975 2065 4325 2075
rect 3975 1735 3985 2065
rect 4315 1735 4325 2065
rect 3975 1725 4325 1735
rect 4400 1650 4450 2150
rect 4525 2065 4875 2075
rect 4525 1735 4535 2065
rect 4865 1735 4875 2065
rect 4525 1725 4875 1735
rect 4950 1650 5000 2150
rect 5075 2065 5425 2075
rect 5075 1735 5085 2065
rect 5415 1735 5425 2065
rect 5075 1725 5425 1735
rect 5500 1650 5550 2150
rect 5625 2065 5975 2075
rect 5625 1735 5635 2065
rect 5965 1735 5975 2065
rect 5625 1725 5975 1735
rect 6050 1650 6100 2150
rect 6175 2065 6525 2075
rect 6175 1735 6185 2065
rect 6515 1735 6525 2065
rect 6175 1725 6525 1735
rect 6600 1650 6650 2150
rect 6725 2065 7075 2075
rect 6725 1735 6735 2065
rect 7065 1735 7075 2065
rect 6725 1725 7075 1735
rect 7150 1650 7200 2150
rect 7275 2065 7625 2075
rect 7275 1735 7285 2065
rect 7615 1735 7625 2065
rect 7275 1725 7625 1735
rect 7700 1650 7750 2150
rect 7825 2065 8175 2075
rect 7825 1735 7835 2065
rect 8165 1735 8175 2065
rect 7825 1725 8175 1735
rect 8250 1650 8300 2150
rect 8375 2065 8725 2075
rect 8375 1735 8385 2065
rect 8715 1735 8725 2065
rect 8375 1725 8725 1735
rect 8800 1650 8850 2150
rect 8925 2065 9275 2075
rect 8925 1735 8935 2065
rect 9265 1735 9275 2065
rect 8925 1725 9275 1735
rect 9350 1650 9400 2150
rect 9475 2065 9825 2075
rect 9475 1735 9485 2065
rect 9815 1735 9825 2065
rect 9475 1725 9825 1735
rect 9900 1650 9950 2150
rect 10025 2065 10375 2075
rect 10025 1735 10035 2065
rect 10365 1735 10375 2065
rect 10025 1725 10375 1735
rect 10450 1650 10500 2150
rect 10575 2065 10925 2075
rect 10575 1735 10585 2065
rect 10915 1735 10925 2065
rect 10575 1725 10925 1735
rect 11000 1650 11050 2150
rect 11125 2065 11475 2075
rect 11125 1735 11135 2065
rect 11465 1735 11475 2065
rect 11125 1725 11475 1735
rect 11550 1650 11600 2150
rect 11675 2065 12025 2075
rect 11675 1735 11685 2065
rect 12015 1735 12025 2065
rect 11675 1725 12025 1735
rect 12100 1650 12150 2150
rect 12225 2065 12575 2075
rect 12225 1735 12235 2065
rect 12565 1735 12575 2065
rect 12225 1725 12575 1735
rect 12650 1650 12700 2150
rect 12775 2065 13125 2075
rect 12775 1735 12785 2065
rect 13115 1735 13125 2065
rect 12775 1725 13125 1735
rect 13200 1650 13250 2150
rect 13325 2065 13675 2075
rect 13325 1735 13335 2065
rect 13665 1735 13675 2065
rect 13325 1725 13675 1735
rect 13750 1650 13975 2150
rect -725 1642 13975 1650
rect -725 1608 -542 1642
rect -508 1608 8 1642
rect 42 1608 558 1642
rect 592 1608 1108 1642
rect 1142 1608 1658 1642
rect 1692 1608 2208 1642
rect 2242 1608 2758 1642
rect 2792 1608 3308 1642
rect 3342 1608 3858 1642
rect 3892 1608 4408 1642
rect 4442 1608 4958 1642
rect 4992 1608 5508 1642
rect 5542 1608 6058 1642
rect 6092 1608 6608 1642
rect 6642 1608 7158 1642
rect 7192 1608 7708 1642
rect 7742 1608 8258 1642
rect 8292 1608 8808 1642
rect 8842 1608 9358 1642
rect 9392 1608 9908 1642
rect 9942 1608 10458 1642
rect 10492 1608 11008 1642
rect 11042 1608 11558 1642
rect 11592 1608 12108 1642
rect 12142 1608 12658 1642
rect 12692 1608 13208 1642
rect 13242 1608 13758 1642
rect 13792 1608 13975 1642
rect -725 1600 13975 1608
rect -725 1100 -500 1600
rect -425 1515 -75 1525
rect -425 1185 -415 1515
rect -85 1185 -75 1515
rect -425 1175 -75 1185
rect 0 1100 50 1600
rect 125 1515 475 1525
rect 125 1185 135 1515
rect 465 1185 475 1515
rect 125 1175 475 1185
rect 550 1100 600 1600
rect 675 1515 1025 1525
rect 675 1185 685 1515
rect 1015 1185 1025 1515
rect 675 1175 1025 1185
rect 1100 1100 1150 1600
rect 1225 1515 1575 1525
rect 1225 1185 1235 1515
rect 1565 1185 1575 1515
rect 1225 1175 1575 1185
rect 1650 1100 1700 1600
rect 1775 1515 2125 1525
rect 1775 1185 1785 1515
rect 2115 1185 2125 1515
rect 1775 1175 2125 1185
rect 2200 1100 2250 1600
rect 2325 1515 2675 1525
rect 2325 1185 2335 1515
rect 2665 1185 2675 1515
rect 2325 1175 2675 1185
rect 2750 1100 2800 1600
rect 2875 1515 3225 1525
rect 2875 1185 2885 1515
rect 3215 1185 3225 1515
rect 2875 1175 3225 1185
rect 3300 1100 3350 1600
rect 3425 1515 3775 1525
rect 3425 1185 3435 1515
rect 3765 1185 3775 1515
rect 3425 1175 3775 1185
rect 3850 1100 3900 1600
rect 3975 1515 4325 1525
rect 3975 1185 3985 1515
rect 4315 1185 4325 1515
rect 3975 1175 4325 1185
rect 4400 1100 4450 1600
rect 4525 1515 4875 1525
rect 4525 1185 4535 1515
rect 4865 1185 4875 1515
rect 4525 1175 4875 1185
rect 4950 1100 5000 1600
rect 5075 1515 5425 1525
rect 5075 1185 5085 1515
rect 5415 1185 5425 1515
rect 5075 1175 5425 1185
rect 5500 1100 5550 1600
rect 5625 1515 5975 1525
rect 5625 1185 5635 1515
rect 5965 1185 5975 1515
rect 5625 1175 5975 1185
rect 6050 1100 6100 1600
rect 6175 1515 6525 1525
rect 6175 1185 6185 1515
rect 6515 1185 6525 1515
rect 6175 1175 6525 1185
rect 6600 1100 6650 1600
rect 6725 1515 7075 1525
rect 6725 1185 6735 1515
rect 7065 1185 7075 1515
rect 6725 1175 7075 1185
rect 7150 1100 7200 1600
rect 7275 1515 7625 1525
rect 7275 1185 7285 1515
rect 7615 1185 7625 1515
rect 7275 1175 7625 1185
rect 7700 1100 7750 1600
rect 7825 1515 8175 1525
rect 7825 1185 7835 1515
rect 8165 1185 8175 1515
rect 7825 1175 8175 1185
rect 8250 1100 8300 1600
rect 8375 1515 8725 1525
rect 8375 1185 8385 1515
rect 8715 1185 8725 1515
rect 8375 1175 8725 1185
rect 8800 1100 8850 1600
rect 8925 1515 9275 1525
rect 8925 1185 8935 1515
rect 9265 1185 9275 1515
rect 8925 1175 9275 1185
rect 9350 1100 9400 1600
rect 9475 1515 9825 1525
rect 9475 1185 9485 1515
rect 9815 1185 9825 1515
rect 9475 1175 9825 1185
rect 9900 1100 9950 1600
rect 10025 1515 10375 1525
rect 10025 1185 10035 1515
rect 10365 1185 10375 1515
rect 10025 1175 10375 1185
rect 10450 1100 10500 1600
rect 10575 1515 10925 1525
rect 10575 1185 10585 1515
rect 10915 1185 10925 1515
rect 10575 1175 10925 1185
rect 11000 1100 11050 1600
rect 11125 1515 11475 1525
rect 11125 1185 11135 1515
rect 11465 1185 11475 1515
rect 11125 1175 11475 1185
rect 11550 1100 11600 1600
rect 11675 1515 12025 1525
rect 11675 1185 11685 1515
rect 12015 1185 12025 1515
rect 11675 1175 12025 1185
rect 12100 1100 12150 1600
rect 12225 1515 12575 1525
rect 12225 1185 12235 1515
rect 12565 1185 12575 1515
rect 12225 1175 12575 1185
rect 12650 1100 12700 1600
rect 12775 1515 13125 1525
rect 12775 1185 12785 1515
rect 13115 1185 13125 1515
rect 12775 1175 13125 1185
rect 13200 1100 13250 1600
rect 13325 1515 13675 1525
rect 13325 1185 13335 1515
rect 13665 1185 13675 1515
rect 13325 1175 13675 1185
rect 13750 1100 13975 1600
rect 14065 1238 14185 1248
rect 14065 1138 14075 1238
rect 14175 1138 14185 1238
rect 14065 1128 14185 1138
rect -725 1092 13975 1100
rect -725 1058 -542 1092
rect -508 1058 8 1092
rect 42 1058 558 1092
rect 592 1058 1108 1092
rect 1142 1058 1658 1092
rect 1692 1058 2208 1092
rect 2242 1058 2758 1092
rect 2792 1058 3308 1092
rect 3342 1058 3858 1092
rect 3892 1058 4408 1092
rect 4442 1058 4958 1092
rect 4992 1058 5508 1092
rect 5542 1058 6058 1092
rect 6092 1058 6608 1092
rect 6642 1058 7158 1092
rect 7192 1058 7708 1092
rect 7742 1058 8258 1092
rect 8292 1058 8808 1092
rect 8842 1058 9358 1092
rect 9392 1058 9908 1092
rect 9942 1058 10458 1092
rect 10492 1058 11008 1092
rect 11042 1058 11558 1092
rect 11592 1058 12108 1092
rect 12142 1058 12658 1092
rect 12692 1058 13208 1092
rect 13242 1058 13758 1092
rect 13792 1058 13975 1092
rect -725 1050 13975 1058
rect -935 1012 -815 1022
rect -935 912 -925 1012
rect -825 912 -815 1012
rect -935 902 -815 912
rect -725 550 -500 1050
rect -425 965 -75 975
rect -425 635 -415 965
rect -85 635 -75 965
rect -425 625 -75 635
rect 0 550 50 1050
rect 125 965 475 975
rect 125 635 135 965
rect 465 635 475 965
rect 125 625 475 635
rect 550 550 600 1050
rect 675 965 1025 975
rect 675 635 685 965
rect 1015 635 1025 965
rect 675 625 1025 635
rect 1100 550 1150 1050
rect 1225 965 1575 975
rect 1225 635 1235 965
rect 1565 635 1575 965
rect 1225 625 1575 635
rect 1650 550 1700 1050
rect 1775 965 2125 975
rect 1775 635 1785 965
rect 2115 635 2125 965
rect 1775 625 2125 635
rect 2200 550 2250 1050
rect 2325 965 2675 975
rect 2325 635 2335 965
rect 2665 635 2675 965
rect 2325 625 2675 635
rect 2750 550 2800 1050
rect 2875 965 3225 975
rect 2875 635 2885 965
rect 3215 635 3225 965
rect 2875 625 3225 635
rect 3300 550 3350 1050
rect 3425 965 3775 975
rect 3425 635 3435 965
rect 3765 635 3775 965
rect 3425 625 3775 635
rect 3850 550 3900 1050
rect 3975 965 4325 975
rect 3975 635 3985 965
rect 4315 635 4325 965
rect 3975 625 4325 635
rect 4400 550 4450 1050
rect 4525 965 4875 975
rect 4525 635 4535 965
rect 4865 635 4875 965
rect 4525 625 4875 635
rect 4950 550 5000 1050
rect 5075 965 5425 975
rect 5075 635 5085 965
rect 5415 635 5425 965
rect 5075 625 5425 635
rect 5500 550 5550 1050
rect 5625 965 5975 975
rect 5625 635 5635 965
rect 5965 635 5975 965
rect 5625 625 5975 635
rect 6050 550 6100 1050
rect 6175 965 6525 975
rect 6175 635 6185 965
rect 6515 635 6525 965
rect 6175 625 6525 635
rect 6600 550 6650 1050
rect 6725 965 7075 975
rect 6725 635 6735 965
rect 7065 635 7075 965
rect 6725 625 7075 635
rect 7150 550 7200 1050
rect 7275 965 7625 975
rect 7275 635 7285 965
rect 7615 635 7625 965
rect 7275 625 7625 635
rect 7700 550 7750 1050
rect 7825 965 8175 975
rect 7825 635 7835 965
rect 8165 635 8175 965
rect 7825 625 8175 635
rect 8250 550 8300 1050
rect 8375 965 8725 975
rect 8375 635 8385 965
rect 8715 635 8725 965
rect 8375 625 8725 635
rect 8800 550 8850 1050
rect 8925 965 9275 975
rect 8925 635 8935 965
rect 9265 635 9275 965
rect 8925 625 9275 635
rect 9350 550 9400 1050
rect 9475 965 9825 975
rect 9475 635 9485 965
rect 9815 635 9825 965
rect 9475 625 9825 635
rect 9900 550 9950 1050
rect 10025 965 10375 975
rect 10025 635 10035 965
rect 10365 635 10375 965
rect 10025 625 10375 635
rect 10450 550 10500 1050
rect 10575 965 10925 975
rect 10575 635 10585 965
rect 10915 635 10925 965
rect 10575 625 10925 635
rect 11000 550 11050 1050
rect 11125 965 11475 975
rect 11125 635 11135 965
rect 11465 635 11475 965
rect 11125 625 11475 635
rect 11550 550 11600 1050
rect 11675 965 12025 975
rect 11675 635 11685 965
rect 12015 635 12025 965
rect 11675 625 12025 635
rect 12100 550 12150 1050
rect 12225 965 12575 975
rect 12225 635 12235 965
rect 12565 635 12575 965
rect 12225 625 12575 635
rect 12650 550 12700 1050
rect 12775 965 13125 975
rect 12775 635 12785 965
rect 13115 635 13125 965
rect 12775 625 13125 635
rect 13200 550 13250 1050
rect 13325 965 13675 975
rect 13325 635 13335 965
rect 13665 635 13675 965
rect 13325 625 13675 635
rect 13750 550 13975 1050
rect -725 542 13975 550
rect -725 508 -542 542
rect -508 508 8 542
rect 42 508 558 542
rect 592 508 1108 542
rect 1142 508 1658 542
rect 1692 508 2208 542
rect 2242 508 2758 542
rect 2792 508 3308 542
rect 3342 508 3858 542
rect 3892 508 4408 542
rect 4442 508 4958 542
rect 4992 508 5508 542
rect 5542 508 6058 542
rect 6092 508 6608 542
rect 6642 508 7158 542
rect 7192 508 7708 542
rect 7742 508 8258 542
rect 8292 508 8808 542
rect 8842 508 9358 542
rect 9392 508 9908 542
rect 9942 508 10458 542
rect 10492 508 11008 542
rect 11042 508 11558 542
rect 11592 508 12108 542
rect 12142 508 12658 542
rect 12692 508 13208 542
rect 13242 508 13758 542
rect 13792 508 13975 542
rect -725 500 13975 508
rect -725 0 -500 500
rect -425 415 -75 425
rect -425 85 -415 415
rect -85 85 -75 415
rect -425 75 -75 85
rect 0 0 50 500
rect 125 415 475 425
rect 125 85 135 415
rect 465 85 475 415
rect 125 75 475 85
rect 550 0 600 500
rect 675 415 1025 425
rect 675 85 685 415
rect 1015 85 1025 415
rect 675 75 1025 85
rect 1100 0 1150 500
rect 1225 415 1575 425
rect 1225 85 1235 415
rect 1565 85 1575 415
rect 1225 75 1575 85
rect 1650 0 1700 500
rect 1775 415 2125 425
rect 1775 85 1785 415
rect 2115 85 2125 415
rect 1775 75 2125 85
rect 2200 0 2250 500
rect 2325 415 2675 425
rect 2325 85 2335 415
rect 2665 85 2675 415
rect 2325 75 2675 85
rect 2750 0 2800 500
rect 2875 415 3225 425
rect 2875 85 2885 415
rect 3215 85 3225 415
rect 2875 75 3225 85
rect 3300 0 3350 500
rect 3425 415 3775 425
rect 3425 85 3435 415
rect 3765 85 3775 415
rect 3425 75 3775 85
rect 3850 0 3900 500
rect 3975 415 4325 425
rect 3975 85 3985 415
rect 4315 85 4325 415
rect 3975 75 4325 85
rect 4400 0 4450 500
rect 4525 415 4875 425
rect 4525 85 4535 415
rect 4865 85 4875 415
rect 4525 75 4875 85
rect 4950 0 5000 500
rect 5075 415 5425 425
rect 5075 85 5085 415
rect 5415 85 5425 415
rect 5075 75 5425 85
rect 5500 0 5550 500
rect 5625 415 5975 425
rect 5625 85 5635 415
rect 5965 85 5975 415
rect 5625 75 5975 85
rect 6050 0 6100 500
rect 6175 415 6525 425
rect 6175 85 6185 415
rect 6515 85 6525 415
rect 6175 75 6525 85
rect 6600 0 6650 500
rect 6725 415 7075 425
rect 6725 85 6735 415
rect 7065 85 7075 415
rect 6725 75 7075 85
rect 7150 0 7200 500
rect 7275 415 7625 425
rect 7275 85 7285 415
rect 7615 85 7625 415
rect 7275 75 7625 85
rect 7700 0 7750 500
rect 7825 415 8175 425
rect 7825 85 7835 415
rect 8165 85 8175 415
rect 7825 75 8175 85
rect 8250 0 8300 500
rect 8375 415 8725 425
rect 8375 85 8385 415
rect 8715 85 8725 415
rect 8375 75 8725 85
rect 8800 0 8850 500
rect 8925 415 9275 425
rect 8925 85 8935 415
rect 9265 85 9275 415
rect 8925 75 9275 85
rect 9350 0 9400 500
rect 9475 415 9825 425
rect 9475 85 9485 415
rect 9815 85 9825 415
rect 9475 75 9825 85
rect 9900 0 9950 500
rect 10025 415 10375 425
rect 10025 85 10035 415
rect 10365 85 10375 415
rect 10025 75 10375 85
rect 10450 0 10500 500
rect 10575 415 10925 425
rect 10575 85 10585 415
rect 10915 85 10925 415
rect 10575 75 10925 85
rect 11000 0 11050 500
rect 11125 415 11475 425
rect 11125 85 11135 415
rect 11465 85 11475 415
rect 11125 75 11475 85
rect 11550 0 11600 500
rect 11675 415 12025 425
rect 11675 85 11685 415
rect 12015 85 12025 415
rect 11675 75 12025 85
rect 12100 0 12150 500
rect 12225 415 12575 425
rect 12225 85 12235 415
rect 12565 85 12575 415
rect 12225 75 12575 85
rect 12650 0 12700 500
rect 12775 415 13125 425
rect 12775 85 12785 415
rect 13115 85 13125 415
rect 12775 75 13125 85
rect 13200 0 13250 500
rect 13325 415 13675 425
rect 13325 85 13335 415
rect 13665 85 13675 415
rect 13325 75 13675 85
rect 13750 0 13975 500
rect 14065 138 14185 148
rect 14065 38 14075 138
rect 14175 38 14185 138
rect 14065 28 14185 38
rect -725 -8 13975 0
rect -725 -42 -542 -8
rect -508 -42 8 -8
rect 42 -42 558 -8
rect 592 -42 1108 -8
rect 1142 -42 1658 -8
rect 1692 -42 2208 -8
rect 2242 -42 2758 -8
rect 2792 -42 3308 -8
rect 3342 -42 3858 -8
rect 3892 -42 4408 -8
rect 4442 -42 4958 -8
rect 4992 -42 5508 -8
rect 5542 -42 6058 -8
rect 6092 -42 6608 -8
rect 6642 -42 7158 -8
rect 7192 -42 7708 -8
rect 7742 -42 8258 -8
rect 8292 -42 8808 -8
rect 8842 -42 9358 -8
rect 9392 -42 9908 -8
rect 9942 -42 10458 -8
rect 10492 -42 11008 -8
rect 11042 -42 11558 -8
rect 11592 -42 12108 -8
rect 12142 -42 12658 -8
rect 12692 -42 13208 -8
rect 13242 -42 13758 -8
rect 13792 -42 13975 -8
rect -725 -50 13975 -42
rect -935 -88 -815 -78
rect -935 -188 -925 -88
rect -825 -188 -815 -88
rect -935 -198 -815 -188
rect -725 -550 -500 -50
rect -425 -135 -75 -125
rect -425 -465 -415 -135
rect -85 -465 -75 -135
rect -425 -475 -75 -465
rect 0 -550 50 -50
rect 125 -135 475 -125
rect 125 -465 135 -135
rect 465 -465 475 -135
rect 125 -475 475 -465
rect 550 -550 600 -50
rect 675 -135 1025 -125
rect 675 -465 685 -135
rect 1015 -465 1025 -135
rect 675 -475 1025 -465
rect 1100 -550 1150 -50
rect 1225 -135 1575 -125
rect 1225 -465 1235 -135
rect 1565 -465 1575 -135
rect 1225 -475 1575 -465
rect 1650 -550 1700 -50
rect 1775 -135 2125 -125
rect 1775 -465 1785 -135
rect 2115 -465 2125 -135
rect 1775 -475 2125 -465
rect 2200 -550 2250 -50
rect 2325 -135 2675 -125
rect 2325 -465 2335 -135
rect 2665 -465 2675 -135
rect 2325 -475 2675 -465
rect 2750 -550 2800 -50
rect 2875 -135 3225 -125
rect 2875 -465 2885 -135
rect 3215 -465 3225 -135
rect 2875 -475 3225 -465
rect 3300 -550 3350 -50
rect 3425 -135 3775 -125
rect 3425 -465 3435 -135
rect 3765 -465 3775 -135
rect 3425 -475 3775 -465
rect 3850 -550 3900 -50
rect 3975 -135 4325 -125
rect 3975 -465 3985 -135
rect 4315 -465 4325 -135
rect 3975 -475 4325 -465
rect 4400 -550 4450 -50
rect 4525 -135 4875 -125
rect 4525 -465 4535 -135
rect 4865 -465 4875 -135
rect 4525 -475 4875 -465
rect 4950 -550 5000 -50
rect 5075 -135 5425 -125
rect 5075 -465 5085 -135
rect 5415 -465 5425 -135
rect 5075 -475 5425 -465
rect 5500 -550 5550 -50
rect 5625 -135 5975 -125
rect 5625 -465 5635 -135
rect 5965 -465 5975 -135
rect 5625 -475 5975 -465
rect 6050 -550 6100 -50
rect 6175 -135 6525 -125
rect 6175 -465 6185 -135
rect 6515 -465 6525 -135
rect 6175 -475 6525 -465
rect 6600 -550 6650 -50
rect 6725 -135 7075 -125
rect 6725 -465 6735 -135
rect 7065 -465 7075 -135
rect 6725 -475 7075 -465
rect 7150 -550 7200 -50
rect 7275 -135 7625 -125
rect 7275 -465 7285 -135
rect 7615 -465 7625 -135
rect 7275 -475 7625 -465
rect 7700 -550 7750 -50
rect 7825 -135 8175 -125
rect 7825 -465 7835 -135
rect 8165 -465 8175 -135
rect 7825 -475 8175 -465
rect 8250 -550 8300 -50
rect 8375 -135 8725 -125
rect 8375 -465 8385 -135
rect 8715 -465 8725 -135
rect 8375 -475 8725 -465
rect 8800 -550 8850 -50
rect 8925 -135 9275 -125
rect 8925 -465 8935 -135
rect 9265 -465 9275 -135
rect 8925 -475 9275 -465
rect 9350 -550 9400 -50
rect 9475 -135 9825 -125
rect 9475 -465 9485 -135
rect 9815 -465 9825 -135
rect 9475 -475 9825 -465
rect 9900 -550 9950 -50
rect 10025 -135 10375 -125
rect 10025 -465 10035 -135
rect 10365 -465 10375 -135
rect 10025 -475 10375 -465
rect 10450 -550 10500 -50
rect 10575 -135 10925 -125
rect 10575 -465 10585 -135
rect 10915 -465 10925 -135
rect 10575 -475 10925 -465
rect 11000 -550 11050 -50
rect 11125 -135 11475 -125
rect 11125 -465 11135 -135
rect 11465 -465 11475 -135
rect 11125 -475 11475 -465
rect 11550 -550 11600 -50
rect 11675 -135 12025 -125
rect 11675 -465 11685 -135
rect 12015 -465 12025 -135
rect 11675 -475 12025 -465
rect 12100 -550 12150 -50
rect 12225 -135 12575 -125
rect 12225 -465 12235 -135
rect 12565 -465 12575 -135
rect 12225 -475 12575 -465
rect 12650 -550 12700 -50
rect 12775 -135 13125 -125
rect 12775 -465 12785 -135
rect 13115 -465 13125 -135
rect 12775 -475 13125 -465
rect 13200 -550 13250 -50
rect 13325 -135 13675 -125
rect 13325 -465 13335 -135
rect 13665 -465 13675 -135
rect 13325 -475 13675 -465
rect 13750 -550 13975 -50
rect -725 -558 13975 -550
rect -725 -592 -542 -558
rect -508 -592 8 -558
rect 42 -592 558 -558
rect 592 -592 1108 -558
rect 1142 -592 1658 -558
rect 1692 -592 2208 -558
rect 2242 -592 2758 -558
rect 2792 -592 3308 -558
rect 3342 -592 3858 -558
rect 3892 -592 4408 -558
rect 4442 -592 4958 -558
rect 4992 -592 5508 -558
rect 5542 -592 6058 -558
rect 6092 -592 6608 -558
rect 6642 -592 7158 -558
rect 7192 -592 7708 -558
rect 7742 -592 8258 -558
rect 8292 -592 8808 -558
rect 8842 -592 9358 -558
rect 9392 -592 9908 -558
rect 9942 -592 10458 -558
rect 10492 -592 11008 -558
rect 11042 -592 11558 -558
rect 11592 -592 12108 -558
rect 12142 -592 12658 -558
rect 12692 -592 13208 -558
rect 13242 -592 13758 -558
rect 13792 -592 13975 -558
rect -725 -775 13975 -592
rect -148 -875 -28 -865
rect -148 -975 -138 -875
rect -38 -975 -28 -875
rect -148 -985 -28 -975
rect 952 -875 1072 -865
rect 952 -975 962 -875
rect 1062 -975 1072 -875
rect 952 -985 1072 -975
rect 2052 -875 2172 -865
rect 2052 -975 2062 -875
rect 2162 -975 2172 -875
rect 2052 -985 2172 -975
rect 3152 -875 3272 -865
rect 3152 -975 3162 -875
rect 3262 -975 3272 -875
rect 3152 -985 3272 -975
rect 4252 -875 4372 -865
rect 4252 -975 4262 -875
rect 4362 -975 4372 -875
rect 4252 -985 4372 -975
rect 5352 -875 5472 -865
rect 5352 -975 5362 -875
rect 5462 -975 5472 -875
rect 5352 -985 5472 -975
rect 6452 -875 6572 -865
rect 6452 -975 6462 -875
rect 6562 -975 6572 -875
rect 6452 -985 6572 -975
rect 7552 -875 7672 -865
rect 7552 -975 7562 -875
rect 7662 -975 7672 -875
rect 7552 -985 7672 -975
rect 8652 -875 8772 -865
rect 8652 -975 8662 -875
rect 8762 -975 8772 -875
rect 8652 -985 8772 -975
rect 9752 -875 9872 -865
rect 9752 -975 9762 -875
rect 9862 -975 9872 -875
rect 9752 -985 9872 -975
rect 10852 -875 10972 -865
rect 10852 -975 10862 -875
rect 10962 -975 10972 -875
rect 10852 -985 10972 -975
rect 11952 -875 12072 -865
rect 11952 -975 11962 -875
rect 12062 -975 12072 -875
rect 11952 -985 12072 -975
rect 13052 -875 13172 -865
rect 13052 -975 13062 -875
rect 13162 -975 13172 -875
rect 13052 -985 13172 -975
rect 14775 -1575 14787 14725
rect -507 -1587 14787 -1575
rect -507 -5563 -495 -1587
rect 18763 -5563 18775 18713
rect -507 -5575 18775 -5563
<< via2 >>
rect 88 14025 188 14125
rect 1188 14025 1288 14125
rect 2288 14025 2388 14125
rect 3388 14025 3488 14125
rect 4488 14025 4588 14125
rect 5588 14025 5688 14125
rect 6688 14025 6788 14125
rect 7788 14025 7888 14125
rect 8888 14025 8988 14125
rect 9988 14025 10088 14125
rect 11088 14025 11188 14125
rect 12188 14025 12288 14125
rect 13288 14025 13388 14125
rect -310 13390 -190 13510
rect 240 13390 360 13510
rect 790 13390 910 13510
rect 1340 13390 1460 13510
rect 1890 13390 2010 13510
rect 2440 13390 2560 13510
rect 2990 13390 3110 13510
rect 3540 13390 3660 13510
rect 4090 13390 4210 13510
rect 4640 13390 4760 13510
rect 5190 13390 5310 13510
rect 5740 13390 5860 13510
rect 6290 13390 6410 13510
rect 6840 13390 6960 13510
rect 7390 13390 7510 13510
rect 7940 13390 8060 13510
rect 8490 13390 8610 13510
rect 9040 13390 9160 13510
rect 9590 13390 9710 13510
rect 10140 13390 10260 13510
rect 10690 13390 10810 13510
rect 11240 13390 11360 13510
rect 11790 13390 11910 13510
rect 12340 13390 12460 13510
rect 12890 13390 13010 13510
rect 13440 13390 13560 13510
rect 14075 13238 14175 13338
rect -925 13012 -825 13112
rect -310 12840 -190 12960
rect 240 12840 360 12960
rect 790 12840 910 12960
rect 1340 12840 1460 12960
rect 1890 12840 2010 12960
rect 2440 12840 2560 12960
rect 2990 12840 3110 12960
rect 3540 12840 3660 12960
rect 4090 12840 4210 12960
rect 4640 12840 4760 12960
rect 5190 12840 5310 12960
rect 5740 12840 5860 12960
rect 6290 12840 6410 12960
rect 6840 12840 6960 12960
rect 7390 12840 7510 12960
rect 7940 12840 8060 12960
rect 8490 12840 8610 12960
rect 9040 12840 9160 12960
rect 9590 12840 9710 12960
rect 10140 12840 10260 12960
rect 10690 12840 10810 12960
rect 11240 12840 11360 12960
rect 11790 12840 11910 12960
rect 12340 12840 12460 12960
rect 12890 12840 13010 12960
rect 13440 12840 13560 12960
rect -310 12290 -190 12410
rect 240 12290 360 12410
rect 790 12290 910 12410
rect 1340 12290 1460 12410
rect 1890 12290 2010 12410
rect 2440 12290 2560 12410
rect 2990 12290 3110 12410
rect 3540 12290 3660 12410
rect 4090 12290 4210 12410
rect 4640 12290 4760 12410
rect 5190 12290 5310 12410
rect 5740 12290 5860 12410
rect 6290 12290 6410 12410
rect 6840 12290 6960 12410
rect 7390 12290 7510 12410
rect 7940 12290 8060 12410
rect 8490 12290 8610 12410
rect 9040 12290 9160 12410
rect 9590 12290 9710 12410
rect 10140 12290 10260 12410
rect 10690 12290 10810 12410
rect 11240 12290 11360 12410
rect 11790 12290 11910 12410
rect 12340 12290 12460 12410
rect 12890 12290 13010 12410
rect 13440 12290 13560 12410
rect 14075 12138 14175 12238
rect -925 11912 -825 12012
rect -310 11740 -190 11860
rect 240 11740 360 11860
rect 790 11740 910 11860
rect 1340 11740 1460 11860
rect 1890 11740 2010 11860
rect 2440 11740 2560 11860
rect 2990 11740 3110 11860
rect 3540 11740 3660 11860
rect 4090 11740 4210 11860
rect 4640 11740 4760 11860
rect 5190 11740 5310 11860
rect 5740 11740 5860 11860
rect 6290 11740 6410 11860
rect 6840 11740 6960 11860
rect 7390 11740 7510 11860
rect 7940 11740 8060 11860
rect 8490 11740 8610 11860
rect 9040 11740 9160 11860
rect 9590 11740 9710 11860
rect 10140 11740 10260 11860
rect 10690 11740 10810 11860
rect 11240 11740 11360 11860
rect 11790 11740 11910 11860
rect 12340 11740 12460 11860
rect 12890 11740 13010 11860
rect 13440 11740 13560 11860
rect -310 11190 -190 11310
rect 240 11190 360 11310
rect 790 11190 910 11310
rect 1340 11190 1460 11310
rect 1890 11190 2010 11310
rect 2440 11190 2560 11310
rect 2990 11190 3110 11310
rect 3540 11190 3660 11310
rect 4090 11190 4210 11310
rect 4640 11190 4760 11310
rect 5190 11190 5310 11310
rect 5740 11190 5860 11310
rect 6290 11190 6410 11310
rect 6840 11190 6960 11310
rect 7390 11190 7510 11310
rect 7940 11190 8060 11310
rect 8490 11190 8610 11310
rect 9040 11190 9160 11310
rect 9590 11190 9710 11310
rect 10140 11190 10260 11310
rect 10690 11190 10810 11310
rect 11240 11190 11360 11310
rect 11790 11190 11910 11310
rect 12340 11190 12460 11310
rect 12890 11190 13010 11310
rect 13440 11190 13560 11310
rect 14075 11038 14175 11138
rect -925 10812 -825 10912
rect -310 10640 -190 10760
rect 240 10640 360 10760
rect 790 10640 910 10760
rect 1340 10640 1460 10760
rect 1890 10640 2010 10760
rect 2440 10640 2560 10760
rect 2990 10640 3110 10760
rect 3540 10640 3660 10760
rect 4090 10640 4210 10760
rect 4640 10640 4760 10760
rect 5190 10640 5310 10760
rect 5740 10640 5860 10760
rect 6290 10640 6410 10760
rect 6840 10640 6960 10760
rect 7390 10640 7510 10760
rect 7940 10640 8060 10760
rect 8490 10640 8610 10760
rect 9040 10640 9160 10760
rect 9590 10640 9710 10760
rect 10140 10640 10260 10760
rect 10690 10640 10810 10760
rect 11240 10640 11360 10760
rect 11790 10640 11910 10760
rect 12340 10640 12460 10760
rect 12890 10640 13010 10760
rect 13440 10640 13560 10760
rect -310 10090 -190 10210
rect 240 10090 360 10210
rect 790 10090 910 10210
rect 1340 10090 1460 10210
rect 1890 10090 2010 10210
rect 2440 10090 2560 10210
rect 2990 10090 3110 10210
rect 3540 10090 3660 10210
rect 4090 10090 4210 10210
rect 4640 10090 4760 10210
rect 5190 10090 5310 10210
rect 5740 10090 5860 10210
rect 6290 10090 6410 10210
rect 6840 10090 6960 10210
rect 7390 10090 7510 10210
rect 7940 10090 8060 10210
rect 8490 10090 8610 10210
rect 9040 10090 9160 10210
rect 9590 10090 9710 10210
rect 10140 10090 10260 10210
rect 10690 10090 10810 10210
rect 11240 10090 11360 10210
rect 11790 10090 11910 10210
rect 12340 10090 12460 10210
rect 12890 10090 13010 10210
rect 13440 10090 13560 10210
rect 14075 9938 14175 10038
rect -925 9712 -825 9812
rect -310 9540 -190 9660
rect 240 9540 360 9660
rect 790 9540 910 9660
rect 1340 9540 1460 9660
rect 1890 9540 2010 9660
rect 2440 9540 2560 9660
rect 2990 9540 3110 9660
rect 3540 9540 3660 9660
rect 4090 9540 4210 9660
rect 4640 9540 4760 9660
rect 5190 9540 5310 9660
rect 5740 9540 5860 9660
rect 6290 9540 6410 9660
rect 6840 9540 6960 9660
rect 7390 9540 7510 9660
rect 7940 9540 8060 9660
rect 8490 9540 8610 9660
rect 9040 9540 9160 9660
rect 9590 9540 9710 9660
rect 10140 9540 10260 9660
rect 10690 9540 10810 9660
rect 11240 9540 11360 9660
rect 11790 9540 11910 9660
rect 12340 9540 12460 9660
rect 12890 9540 13010 9660
rect 13440 9540 13560 9660
rect -310 8990 -190 9110
rect 240 8990 360 9110
rect 790 8990 910 9110
rect 1340 8990 1460 9110
rect 1890 8990 2010 9110
rect 2440 8990 2560 9110
rect 2990 8990 3110 9110
rect 3540 8990 3660 9110
rect 4090 8990 4210 9110
rect 4640 8990 4760 9110
rect 5190 8990 5310 9110
rect 5740 8990 5860 9110
rect 6290 8990 6410 9110
rect 6840 8990 6960 9110
rect 7390 8990 7510 9110
rect 7940 8990 8060 9110
rect 8490 8990 8610 9110
rect 9040 8990 9160 9110
rect 9590 8990 9710 9110
rect 10140 8990 10260 9110
rect 10690 8990 10810 9110
rect 11240 8990 11360 9110
rect 11790 8990 11910 9110
rect 12340 8990 12460 9110
rect 12890 8990 13010 9110
rect 13440 8990 13560 9110
rect 14075 8838 14175 8938
rect -925 8612 -825 8712
rect -310 8440 -190 8560
rect 240 8440 360 8560
rect 790 8440 910 8560
rect 1340 8440 1460 8560
rect 1890 8440 2010 8560
rect 2440 8440 2560 8560
rect 2990 8440 3110 8560
rect 3540 8440 3660 8560
rect 4090 8440 4210 8560
rect 4640 8440 4760 8560
rect 5190 8440 5310 8560
rect 5740 8440 5860 8560
rect 6290 8440 6410 8560
rect 6840 8440 6960 8560
rect 7390 8440 7510 8560
rect 7940 8440 8060 8560
rect 8490 8440 8610 8560
rect 9040 8440 9160 8560
rect 9590 8440 9710 8560
rect 10140 8440 10260 8560
rect 10690 8440 10810 8560
rect 11240 8440 11360 8560
rect 11790 8440 11910 8560
rect 12340 8440 12460 8560
rect 12890 8440 13010 8560
rect 13440 8440 13560 8560
rect -310 7890 -190 8010
rect 240 7890 360 8010
rect 790 7890 910 8010
rect 1340 7890 1460 8010
rect 1890 7890 2010 8010
rect 2440 7890 2560 8010
rect 2990 7890 3110 8010
rect 3540 7890 3660 8010
rect 4090 7890 4210 8010
rect 4640 7890 4760 8010
rect 5190 7890 5310 8010
rect 5740 7890 5860 8010
rect 6290 7890 6410 8010
rect 6840 7890 6960 8010
rect 7390 7890 7510 8010
rect 7940 7890 8060 8010
rect 8490 7890 8610 8010
rect 9040 7890 9160 8010
rect 9590 7890 9710 8010
rect 10140 7890 10260 8010
rect 10690 7890 10810 8010
rect 11240 7890 11360 8010
rect 11790 7890 11910 8010
rect 12340 7890 12460 8010
rect 12890 7890 13010 8010
rect 13440 7890 13560 8010
rect 14075 7738 14175 7838
rect -925 7512 -825 7612
rect -310 7340 -190 7460
rect 240 7340 360 7460
rect 790 7340 910 7460
rect 1340 7340 1460 7460
rect 1890 7340 2010 7460
rect 2440 7340 2560 7460
rect 2990 7340 3110 7460
rect 3540 7340 3660 7460
rect 4090 7340 4210 7460
rect 4640 7340 4760 7460
rect 5190 7340 5310 7460
rect 5740 7340 5860 7460
rect 6290 7340 6410 7460
rect 6840 7340 6960 7460
rect 7390 7340 7510 7460
rect 7940 7340 8060 7460
rect 8490 7340 8610 7460
rect 9040 7340 9160 7460
rect 9590 7340 9710 7460
rect 10140 7340 10260 7460
rect 10690 7340 10810 7460
rect 11240 7340 11360 7460
rect 11790 7340 11910 7460
rect 12340 7340 12460 7460
rect 12890 7340 13010 7460
rect 13440 7340 13560 7460
rect -310 6790 -190 6910
rect 240 6790 360 6910
rect 790 6790 910 6910
rect 1340 6790 1460 6910
rect 1890 6790 2010 6910
rect 2440 6790 2560 6910
rect 2990 6790 3110 6910
rect 3540 6790 3660 6910
rect 4090 6790 4210 6910
rect 4640 6790 4760 6910
rect 5190 6790 5310 6910
rect 5740 6790 5860 6910
rect 6290 6790 6410 6910
rect 6840 6790 6960 6910
rect 7390 6790 7510 6910
rect 7940 6790 8060 6910
rect 8490 6790 8610 6910
rect 9040 6790 9160 6910
rect 9590 6790 9710 6910
rect 10140 6790 10260 6910
rect 10690 6790 10810 6910
rect 11240 6790 11360 6910
rect 11790 6790 11910 6910
rect 12340 6790 12460 6910
rect 12890 6790 13010 6910
rect 13440 6790 13560 6910
rect 14075 6638 14175 6738
rect -925 6412 -825 6512
rect -310 6240 -190 6360
rect 240 6240 360 6360
rect 790 6240 910 6360
rect 1340 6240 1460 6360
rect 1890 6240 2010 6360
rect 2440 6240 2560 6360
rect 2990 6240 3110 6360
rect 3540 6240 3660 6360
rect 4090 6240 4210 6360
rect 4640 6240 4760 6360
rect 5190 6240 5310 6360
rect 5740 6240 5860 6360
rect 6290 6240 6410 6360
rect 6840 6240 6960 6360
rect 7390 6240 7510 6360
rect 7940 6240 8060 6360
rect 8490 6240 8610 6360
rect 9040 6240 9160 6360
rect 9590 6240 9710 6360
rect 10140 6240 10260 6360
rect 10690 6240 10810 6360
rect 11240 6240 11360 6360
rect 11790 6240 11910 6360
rect 12340 6240 12460 6360
rect 12890 6240 13010 6360
rect 13440 6240 13560 6360
rect -310 5690 -190 5810
rect 240 5690 360 5810
rect 790 5690 910 5810
rect 1340 5690 1460 5810
rect 1890 5690 2010 5810
rect 2440 5690 2560 5810
rect 2990 5690 3110 5810
rect 3540 5690 3660 5810
rect 4090 5690 4210 5810
rect 4640 5690 4760 5810
rect 5190 5690 5310 5810
rect 5740 5690 5860 5810
rect 6290 5690 6410 5810
rect 6840 5690 6960 5810
rect 7390 5690 7510 5810
rect 7940 5690 8060 5810
rect 8490 5690 8610 5810
rect 9040 5690 9160 5810
rect 9590 5690 9710 5810
rect 10140 5690 10260 5810
rect 10690 5690 10810 5810
rect 11240 5690 11360 5810
rect 11790 5690 11910 5810
rect 12340 5690 12460 5810
rect 12890 5690 13010 5810
rect 13440 5690 13560 5810
rect 14075 5538 14175 5638
rect -925 5312 -825 5412
rect -310 5140 -190 5260
rect 240 5140 360 5260
rect 790 5140 910 5260
rect 1340 5140 1460 5260
rect 1890 5140 2010 5260
rect 2440 5140 2560 5260
rect 2990 5140 3110 5260
rect 3540 5140 3660 5260
rect 4090 5140 4210 5260
rect 4640 5140 4760 5260
rect 5190 5140 5310 5260
rect 5740 5140 5860 5260
rect 6290 5140 6410 5260
rect 6840 5140 6960 5260
rect 7390 5140 7510 5260
rect 7940 5140 8060 5260
rect 8490 5140 8610 5260
rect 9040 5140 9160 5260
rect 9590 5140 9710 5260
rect 10140 5140 10260 5260
rect 10690 5140 10810 5260
rect 11240 5140 11360 5260
rect 11790 5140 11910 5260
rect 12340 5140 12460 5260
rect 12890 5140 13010 5260
rect 13440 5140 13560 5260
rect -310 4590 -190 4710
rect 240 4590 360 4710
rect 790 4590 910 4710
rect 1340 4590 1460 4710
rect 1890 4590 2010 4710
rect 2440 4590 2560 4710
rect 2990 4590 3110 4710
rect 3540 4590 3660 4710
rect 4090 4590 4210 4710
rect 4640 4590 4760 4710
rect 5190 4590 5310 4710
rect 5740 4590 5860 4710
rect 6290 4590 6410 4710
rect 6840 4590 6960 4710
rect 7390 4590 7510 4710
rect 7940 4590 8060 4710
rect 8490 4590 8610 4710
rect 9040 4590 9160 4710
rect 9590 4590 9710 4710
rect 10140 4590 10260 4710
rect 10690 4590 10810 4710
rect 11240 4590 11360 4710
rect 11790 4590 11910 4710
rect 12340 4590 12460 4710
rect 12890 4590 13010 4710
rect 13440 4590 13560 4710
rect 14075 4438 14175 4538
rect -925 4212 -825 4312
rect -310 4040 -190 4160
rect 240 4040 360 4160
rect 790 4040 910 4160
rect 1340 4040 1460 4160
rect 1890 4040 2010 4160
rect 2440 4040 2560 4160
rect 2990 4040 3110 4160
rect 3540 4040 3660 4160
rect 4090 4040 4210 4160
rect 4640 4040 4760 4160
rect 5190 4040 5310 4160
rect 5740 4040 5860 4160
rect 6290 4040 6410 4160
rect 6840 4040 6960 4160
rect 7390 4040 7510 4160
rect 7940 4040 8060 4160
rect 8490 4040 8610 4160
rect 9040 4040 9160 4160
rect 9590 4040 9710 4160
rect 10140 4040 10260 4160
rect 10690 4040 10810 4160
rect 11240 4040 11360 4160
rect 11790 4040 11910 4160
rect 12340 4040 12460 4160
rect 12890 4040 13010 4160
rect 13440 4040 13560 4160
rect -310 3490 -190 3610
rect 240 3490 360 3610
rect 790 3490 910 3610
rect 1340 3490 1460 3610
rect 1890 3490 2010 3610
rect 2440 3490 2560 3610
rect 2990 3490 3110 3610
rect 3540 3490 3660 3610
rect 4090 3490 4210 3610
rect 4640 3490 4760 3610
rect 5190 3490 5310 3610
rect 5740 3490 5860 3610
rect 6290 3490 6410 3610
rect 6840 3490 6960 3610
rect 7390 3490 7510 3610
rect 7940 3490 8060 3610
rect 8490 3490 8610 3610
rect 9040 3490 9160 3610
rect 9590 3490 9710 3610
rect 10140 3490 10260 3610
rect 10690 3490 10810 3610
rect 11240 3490 11360 3610
rect 11790 3490 11910 3610
rect 12340 3490 12460 3610
rect 12890 3490 13010 3610
rect 13440 3490 13560 3610
rect 14075 3338 14175 3438
rect -925 3112 -825 3212
rect -310 2940 -190 3060
rect 240 2940 360 3060
rect 790 2940 910 3060
rect 1340 2940 1460 3060
rect 1890 2940 2010 3060
rect 2440 2940 2560 3060
rect 2990 2940 3110 3060
rect 3540 2940 3660 3060
rect 4090 2940 4210 3060
rect 4640 2940 4760 3060
rect 5190 2940 5310 3060
rect 5740 2940 5860 3060
rect 6290 2940 6410 3060
rect 6840 2940 6960 3060
rect 7390 2940 7510 3060
rect 7940 2940 8060 3060
rect 8490 2940 8610 3060
rect 9040 2940 9160 3060
rect 9590 2940 9710 3060
rect 10140 2940 10260 3060
rect 10690 2940 10810 3060
rect 11240 2940 11360 3060
rect 11790 2940 11910 3060
rect 12340 2940 12460 3060
rect 12890 2940 13010 3060
rect 13440 2940 13560 3060
rect -310 2390 -190 2510
rect 240 2390 360 2510
rect 790 2390 910 2510
rect 1340 2390 1460 2510
rect 1890 2390 2010 2510
rect 2440 2390 2560 2510
rect 2990 2390 3110 2510
rect 3540 2390 3660 2510
rect 4090 2390 4210 2510
rect 4640 2390 4760 2510
rect 5190 2390 5310 2510
rect 5740 2390 5860 2510
rect 6290 2390 6410 2510
rect 6840 2390 6960 2510
rect 7390 2390 7510 2510
rect 7940 2390 8060 2510
rect 8490 2390 8610 2510
rect 9040 2390 9160 2510
rect 9590 2390 9710 2510
rect 10140 2390 10260 2510
rect 10690 2390 10810 2510
rect 11240 2390 11360 2510
rect 11790 2390 11910 2510
rect 12340 2390 12460 2510
rect 12890 2390 13010 2510
rect 13440 2390 13560 2510
rect 14075 2238 14175 2338
rect -925 2012 -825 2112
rect -310 1840 -190 1960
rect 240 1840 360 1960
rect 790 1840 910 1960
rect 1340 1840 1460 1960
rect 1890 1840 2010 1960
rect 2440 1840 2560 1960
rect 2990 1840 3110 1960
rect 3540 1840 3660 1960
rect 4090 1840 4210 1960
rect 4640 1840 4760 1960
rect 5190 1840 5310 1960
rect 5740 1840 5860 1960
rect 6290 1840 6410 1960
rect 6840 1840 6960 1960
rect 7390 1840 7510 1960
rect 7940 1840 8060 1960
rect 8490 1840 8610 1960
rect 9040 1840 9160 1960
rect 9590 1840 9710 1960
rect 10140 1840 10260 1960
rect 10690 1840 10810 1960
rect 11240 1840 11360 1960
rect 11790 1840 11910 1960
rect 12340 1840 12460 1960
rect 12890 1840 13010 1960
rect 13440 1840 13560 1960
rect -310 1290 -190 1410
rect 240 1290 360 1410
rect 790 1290 910 1410
rect 1340 1290 1460 1410
rect 1890 1290 2010 1410
rect 2440 1290 2560 1410
rect 2990 1290 3110 1410
rect 3540 1290 3660 1410
rect 4090 1290 4210 1410
rect 4640 1290 4760 1410
rect 5190 1290 5310 1410
rect 5740 1290 5860 1410
rect 6290 1290 6410 1410
rect 6840 1290 6960 1410
rect 7390 1290 7510 1410
rect 7940 1290 8060 1410
rect 8490 1290 8610 1410
rect 9040 1290 9160 1410
rect 9590 1290 9710 1410
rect 10140 1290 10260 1410
rect 10690 1290 10810 1410
rect 11240 1290 11360 1410
rect 11790 1290 11910 1410
rect 12340 1290 12460 1410
rect 12890 1290 13010 1410
rect 13440 1290 13560 1410
rect 14075 1138 14175 1238
rect -925 912 -825 1012
rect -310 740 -190 860
rect 240 740 360 860
rect 790 740 910 860
rect 1340 740 1460 860
rect 1890 740 2010 860
rect 2440 740 2560 860
rect 2990 740 3110 860
rect 3540 740 3660 860
rect 4090 740 4210 860
rect 4640 740 4760 860
rect 5190 740 5310 860
rect 5740 740 5860 860
rect 6290 740 6410 860
rect 6840 740 6960 860
rect 7390 740 7510 860
rect 7940 740 8060 860
rect 8490 740 8610 860
rect 9040 740 9160 860
rect 9590 740 9710 860
rect 10140 740 10260 860
rect 10690 740 10810 860
rect 11240 740 11360 860
rect 11790 740 11910 860
rect 12340 740 12460 860
rect 12890 740 13010 860
rect 13440 740 13560 860
rect -310 190 -190 310
rect 240 190 360 310
rect 790 190 910 310
rect 1340 190 1460 310
rect 1890 190 2010 310
rect 2440 190 2560 310
rect 2990 190 3110 310
rect 3540 190 3660 310
rect 4090 190 4210 310
rect 4640 190 4760 310
rect 5190 190 5310 310
rect 5740 190 5860 310
rect 6290 190 6410 310
rect 6840 190 6960 310
rect 7390 190 7510 310
rect 7940 190 8060 310
rect 8490 190 8610 310
rect 9040 190 9160 310
rect 9590 190 9710 310
rect 10140 190 10260 310
rect 10690 190 10810 310
rect 11240 190 11360 310
rect 11790 190 11910 310
rect 12340 190 12460 310
rect 12890 190 13010 310
rect 13440 190 13560 310
rect 14075 38 14175 138
rect -925 -188 -825 -88
rect -310 -360 -190 -240
rect 240 -360 360 -240
rect 790 -360 910 -240
rect 1340 -360 1460 -240
rect 1890 -360 2010 -240
rect 2440 -360 2560 -240
rect 2990 -360 3110 -240
rect 3540 -360 3660 -240
rect 4090 -360 4210 -240
rect 4640 -360 4760 -240
rect 5190 -360 5310 -240
rect 5740 -360 5860 -240
rect 6290 -360 6410 -240
rect 6840 -360 6960 -240
rect 7390 -360 7510 -240
rect 7940 -360 8060 -240
rect 8490 -360 8610 -240
rect 9040 -360 9160 -240
rect 9590 -360 9710 -240
rect 10140 -360 10260 -240
rect 10690 -360 10810 -240
rect 11240 -360 11360 -240
rect 11790 -360 11910 -240
rect 12340 -360 12460 -240
rect 12890 -360 13010 -240
rect 13440 -360 13560 -240
rect -138 -975 -38 -875
rect 962 -975 1062 -875
rect 2062 -975 2162 -875
rect 3162 -975 3262 -875
rect 4262 -975 4362 -875
rect 5362 -975 5462 -875
rect 6462 -975 6562 -875
rect 7562 -975 7662 -875
rect 8662 -975 8762 -875
rect 9762 -975 9862 -875
rect 10862 -975 10962 -875
rect 11962 -975 12062 -875
rect 13062 -975 13162 -875
<< metal3 >>
rect -2525 14725 13775 15725
rect -2525 13838 -1525 14725
rect -638 13838 -186 14725
rect -2525 13514 -186 13838
rect -88 14125 364 14225
rect -88 14025 88 14125
rect 188 14025 364 14125
rect -88 13612 364 14025
rect 462 13612 914 14725
rect 1012 14125 1464 14225
rect 1012 14025 1188 14125
rect 1288 14025 1464 14125
rect 1012 13612 1464 14025
rect 1562 13612 2014 14725
rect 2112 14125 2564 14225
rect 2112 14025 2288 14125
rect 2388 14025 2564 14125
rect 2112 13612 2564 14025
rect 2662 13612 3114 14725
rect 3212 14125 3664 14225
rect 3212 14025 3388 14125
rect 3488 14025 3664 14125
rect 3212 13612 3664 14025
rect 3762 13612 4214 14725
rect 4312 14125 4764 14225
rect 4312 14025 4488 14125
rect 4588 14025 4764 14125
rect 4312 13612 4764 14025
rect 4862 13612 5314 14725
rect 5412 14125 5864 14225
rect 5412 14025 5588 14125
rect 5688 14025 5864 14125
rect 5412 13612 5864 14025
rect 5962 13612 6414 14725
rect 6512 14125 6964 14225
rect 6512 14025 6688 14125
rect 6788 14025 6964 14125
rect 6512 13612 6964 14025
rect 7062 13612 7514 14725
rect 7612 14125 8064 14225
rect 7612 14025 7788 14125
rect 7888 14025 8064 14125
rect 7612 13612 8064 14025
rect 8162 13612 8614 14725
rect 8712 14125 9164 14225
rect 8712 14025 8888 14125
rect 8988 14025 9164 14125
rect 8712 13612 9164 14025
rect 9262 13612 9714 14725
rect 9812 14125 10264 14225
rect 9812 14025 9988 14125
rect 10088 14025 10264 14125
rect 9812 13612 10264 14025
rect 10362 13612 10814 14725
rect 10912 14125 11364 14225
rect 10912 14025 11088 14125
rect 11188 14025 11364 14125
rect 10912 13612 11364 14025
rect 11462 13612 11914 14725
rect 12012 14125 12464 14225
rect 12012 14025 12188 14125
rect 12288 14025 12464 14125
rect 12012 13612 12464 14025
rect 12562 13612 13014 14725
rect 13112 14125 13564 14225
rect 13112 14025 13288 14125
rect 13388 14025 13564 14125
rect 13112 13612 13564 14025
tri -186 13514 -88 13612 sw
tri -88 13514 10 13612 ne
rect 10 13514 364 13612
tri 364 13514 462 13612 sw
tri 462 13514 560 13612 ne
rect 560 13514 914 13612
tri 914 13514 1012 13612 sw
tri 1012 13514 1110 13612 ne
rect 1110 13514 1464 13612
tri 1464 13514 1562 13612 sw
tri 1562 13514 1660 13612 ne
rect 1660 13514 2014 13612
tri 2014 13514 2112 13612 sw
tri 2112 13514 2210 13612 ne
rect 2210 13514 2564 13612
tri 2564 13514 2662 13612 sw
tri 2662 13514 2760 13612 ne
rect 2760 13514 3114 13612
tri 3114 13514 3212 13612 sw
tri 3212 13514 3310 13612 ne
rect 3310 13514 3664 13612
tri 3664 13514 3762 13612 sw
tri 3762 13514 3860 13612 ne
rect 3860 13514 4214 13612
tri 4214 13514 4312 13612 sw
tri 4312 13514 4410 13612 ne
rect 4410 13514 4764 13612
tri 4764 13514 4862 13612 sw
tri 4862 13514 4960 13612 ne
rect 4960 13514 5314 13612
tri 5314 13514 5412 13612 sw
tri 5412 13514 5510 13612 ne
rect 5510 13514 5864 13612
tri 5864 13514 5962 13612 sw
tri 5962 13514 6060 13612 ne
rect 6060 13514 6414 13612
tri 6414 13514 6512 13612 sw
tri 6512 13514 6610 13612 ne
rect 6610 13514 6964 13612
tri 6964 13514 7062 13612 sw
tri 7062 13514 7160 13612 ne
rect 7160 13514 7514 13612
tri 7514 13514 7612 13612 sw
tri 7612 13514 7710 13612 ne
rect 7710 13514 8064 13612
tri 8064 13514 8162 13612 sw
tri 8162 13514 8260 13612 ne
rect 8260 13514 8614 13612
tri 8614 13514 8712 13612 sw
tri 8712 13514 8810 13612 ne
rect 8810 13514 9164 13612
tri 9164 13514 9262 13612 sw
tri 9262 13514 9360 13612 ne
rect 9360 13514 9714 13612
tri 9714 13514 9812 13612 sw
tri 9812 13514 9910 13612 ne
rect 9910 13514 10264 13612
tri 10264 13514 10362 13612 sw
tri 10362 13514 10460 13612 ne
rect 10460 13514 10814 13612
tri 10814 13514 10912 13612 sw
tri 10912 13514 11010 13612 ne
rect 11010 13514 11364 13612
tri 11364 13514 11462 13612 sw
tri 11462 13514 11560 13612 ne
rect 11560 13514 11914 13612
tri 11914 13514 12012 13612 sw
tri 12012 13514 12110 13612 ne
rect 12110 13514 12464 13612
tri 12464 13514 12562 13612 sw
tri 12562 13514 12660 13612 ne
rect 12660 13514 13014 13612
tri 13014 13514 13112 13612 sw
tri 13112 13514 13210 13612 ne
rect 13210 13514 13564 13612
tri 13564 13514 13662 13612 sw
rect 14775 13514 15775 13725
rect -2525 13510 -88 13514
rect -2525 13390 -310 13510
rect -190 13426 -88 13510
tri -88 13426 0 13514 sw
tri 10 13426 98 13514 ne
rect 98 13510 462 13514
rect 98 13426 240 13510
rect -190 13390 0 13426
rect -2525 13386 0 13390
tri 0 13386 40 13426 sw
tri 98 13386 138 13426 ne
rect 138 13390 240 13426
rect 360 13426 462 13510
tri 462 13426 550 13514 sw
tri 560 13426 648 13514 ne
rect 648 13510 1012 13514
rect 648 13426 790 13510
rect 360 13390 550 13426
rect 138 13386 550 13390
tri 550 13386 590 13426 sw
tri 648 13386 688 13426 ne
rect 688 13390 790 13426
rect 910 13426 1012 13510
tri 1012 13426 1100 13514 sw
tri 1110 13426 1198 13514 ne
rect 1198 13510 1562 13514
rect 1198 13426 1340 13510
rect 910 13390 1100 13426
rect 688 13386 1100 13390
tri 1100 13386 1140 13426 sw
tri 1198 13386 1238 13426 ne
rect 1238 13390 1340 13426
rect 1460 13426 1562 13510
tri 1562 13426 1650 13514 sw
tri 1660 13426 1748 13514 ne
rect 1748 13510 2112 13514
rect 1748 13426 1890 13510
rect 1460 13390 1650 13426
rect 1238 13386 1650 13390
tri 1650 13386 1690 13426 sw
tri 1748 13386 1788 13426 ne
rect 1788 13390 1890 13426
rect 2010 13426 2112 13510
tri 2112 13426 2200 13514 sw
tri 2210 13426 2298 13514 ne
rect 2298 13510 2662 13514
rect 2298 13426 2440 13510
rect 2010 13390 2200 13426
rect 1788 13386 2200 13390
tri 2200 13386 2240 13426 sw
tri 2298 13386 2338 13426 ne
rect 2338 13390 2440 13426
rect 2560 13426 2662 13510
tri 2662 13426 2750 13514 sw
tri 2760 13426 2848 13514 ne
rect 2848 13510 3212 13514
rect 2848 13426 2990 13510
rect 2560 13390 2750 13426
rect 2338 13386 2750 13390
tri 2750 13386 2790 13426 sw
tri 2848 13386 2888 13426 ne
rect 2888 13390 2990 13426
rect 3110 13426 3212 13510
tri 3212 13426 3300 13514 sw
tri 3310 13426 3398 13514 ne
rect 3398 13510 3762 13514
rect 3398 13426 3540 13510
rect 3110 13390 3300 13426
rect 2888 13386 3300 13390
tri 3300 13386 3340 13426 sw
tri 3398 13386 3438 13426 ne
rect 3438 13390 3540 13426
rect 3660 13426 3762 13510
tri 3762 13426 3850 13514 sw
tri 3860 13426 3948 13514 ne
rect 3948 13510 4312 13514
rect 3948 13426 4090 13510
rect 3660 13390 3850 13426
rect 3438 13386 3850 13390
tri 3850 13386 3890 13426 sw
tri 3948 13386 3988 13426 ne
rect 3988 13390 4090 13426
rect 4210 13426 4312 13510
tri 4312 13426 4400 13514 sw
tri 4410 13426 4498 13514 ne
rect 4498 13510 4862 13514
rect 4498 13426 4640 13510
rect 4210 13390 4400 13426
rect 3988 13386 4400 13390
tri 4400 13386 4440 13426 sw
tri 4498 13386 4538 13426 ne
rect 4538 13390 4640 13426
rect 4760 13426 4862 13510
tri 4862 13426 4950 13514 sw
tri 4960 13426 5048 13514 ne
rect 5048 13510 5412 13514
rect 5048 13426 5190 13510
rect 4760 13390 4950 13426
rect 4538 13386 4950 13390
tri 4950 13386 4990 13426 sw
tri 5048 13386 5088 13426 ne
rect 5088 13390 5190 13426
rect 5310 13426 5412 13510
tri 5412 13426 5500 13514 sw
tri 5510 13426 5598 13514 ne
rect 5598 13510 5962 13514
rect 5598 13426 5740 13510
rect 5310 13390 5500 13426
rect 5088 13386 5500 13390
tri 5500 13386 5540 13426 sw
tri 5598 13386 5638 13426 ne
rect 5638 13390 5740 13426
rect 5860 13426 5962 13510
tri 5962 13426 6050 13514 sw
tri 6060 13426 6148 13514 ne
rect 6148 13510 6512 13514
rect 6148 13426 6290 13510
rect 5860 13390 6050 13426
rect 5638 13386 6050 13390
tri 6050 13386 6090 13426 sw
tri 6148 13386 6188 13426 ne
rect 6188 13390 6290 13426
rect 6410 13426 6512 13510
tri 6512 13426 6600 13514 sw
tri 6610 13426 6698 13514 ne
rect 6698 13510 7062 13514
rect 6698 13426 6840 13510
rect 6410 13390 6600 13426
rect 6188 13386 6600 13390
tri 6600 13386 6640 13426 sw
tri 6698 13386 6738 13426 ne
rect 6738 13390 6840 13426
rect 6960 13426 7062 13510
tri 7062 13426 7150 13514 sw
tri 7160 13426 7248 13514 ne
rect 7248 13510 7612 13514
rect 7248 13426 7390 13510
rect 6960 13390 7150 13426
rect 6738 13386 7150 13390
tri 7150 13386 7190 13426 sw
tri 7248 13386 7288 13426 ne
rect 7288 13390 7390 13426
rect 7510 13426 7612 13510
tri 7612 13426 7700 13514 sw
tri 7710 13426 7798 13514 ne
rect 7798 13510 8162 13514
rect 7798 13426 7940 13510
rect 7510 13390 7700 13426
rect 7288 13386 7700 13390
tri 7700 13386 7740 13426 sw
tri 7798 13386 7838 13426 ne
rect 7838 13390 7940 13426
rect 8060 13426 8162 13510
tri 8162 13426 8250 13514 sw
tri 8260 13426 8348 13514 ne
rect 8348 13510 8712 13514
rect 8348 13426 8490 13510
rect 8060 13390 8250 13426
rect 7838 13386 8250 13390
tri 8250 13386 8290 13426 sw
tri 8348 13386 8388 13426 ne
rect 8388 13390 8490 13426
rect 8610 13426 8712 13510
tri 8712 13426 8800 13514 sw
tri 8810 13426 8898 13514 ne
rect 8898 13510 9262 13514
rect 8898 13426 9040 13510
rect 8610 13390 8800 13426
rect 8388 13386 8800 13390
tri 8800 13386 8840 13426 sw
tri 8898 13386 8938 13426 ne
rect 8938 13390 9040 13426
rect 9160 13426 9262 13510
tri 9262 13426 9350 13514 sw
tri 9360 13426 9448 13514 ne
rect 9448 13510 9812 13514
rect 9448 13426 9590 13510
rect 9160 13390 9350 13426
rect 8938 13386 9350 13390
tri 9350 13386 9390 13426 sw
tri 9448 13386 9488 13426 ne
rect 9488 13390 9590 13426
rect 9710 13426 9812 13510
tri 9812 13426 9900 13514 sw
tri 9910 13426 9998 13514 ne
rect 9998 13510 10362 13514
rect 9998 13426 10140 13510
rect 9710 13390 9900 13426
rect 9488 13386 9900 13390
tri 9900 13386 9940 13426 sw
tri 9998 13386 10038 13426 ne
rect 10038 13390 10140 13426
rect 10260 13426 10362 13510
tri 10362 13426 10450 13514 sw
tri 10460 13426 10548 13514 ne
rect 10548 13510 10912 13514
rect 10548 13426 10690 13510
rect 10260 13390 10450 13426
rect 10038 13386 10450 13390
tri 10450 13386 10490 13426 sw
tri 10548 13386 10588 13426 ne
rect 10588 13390 10690 13426
rect 10810 13426 10912 13510
tri 10912 13426 11000 13514 sw
tri 11010 13426 11098 13514 ne
rect 11098 13510 11462 13514
rect 11098 13426 11240 13510
rect 10810 13390 11000 13426
rect 10588 13386 11000 13390
tri 11000 13386 11040 13426 sw
tri 11098 13386 11138 13426 ne
rect 11138 13390 11240 13426
rect 11360 13426 11462 13510
tri 11462 13426 11550 13514 sw
tri 11560 13426 11648 13514 ne
rect 11648 13510 12012 13514
rect 11648 13426 11790 13510
rect 11360 13390 11550 13426
rect 11138 13386 11550 13390
tri 11550 13386 11590 13426 sw
tri 11648 13386 11688 13426 ne
rect 11688 13390 11790 13426
rect 11910 13426 12012 13510
tri 12012 13426 12100 13514 sw
tri 12110 13426 12198 13514 ne
rect 12198 13510 12562 13514
rect 12198 13426 12340 13510
rect 11910 13390 12100 13426
rect 11688 13386 12100 13390
tri 12100 13386 12140 13426 sw
tri 12198 13386 12238 13426 ne
rect 12238 13390 12340 13426
rect 12460 13426 12562 13510
tri 12562 13426 12650 13514 sw
tri 12660 13426 12748 13514 ne
rect 12748 13510 13112 13514
rect 12748 13426 12890 13510
rect 12460 13390 12650 13426
rect 12238 13386 12650 13390
tri 12650 13386 12690 13426 sw
tri 12748 13386 12788 13426 ne
rect 12788 13390 12890 13426
rect 13010 13426 13112 13510
tri 13112 13426 13200 13514 sw
tri 13210 13426 13298 13514 ne
rect 13298 13510 15775 13514
rect 13298 13426 13440 13510
rect 13010 13390 13200 13426
rect 12788 13386 13200 13390
rect -2525 12738 -1525 13386
tri -412 13288 -314 13386 ne
rect -314 13288 40 13386
tri 40 13288 138 13386 sw
tri 138 13288 236 13386 ne
rect 236 13288 590 13386
tri 590 13288 688 13386 sw
tri 688 13288 786 13386 ne
rect 786 13288 1140 13386
tri 1140 13288 1238 13386 sw
tri 1238 13288 1336 13386 ne
rect 1336 13288 1690 13386
tri 1690 13288 1788 13386 sw
tri 1788 13288 1886 13386 ne
rect 1886 13288 2240 13386
tri 2240 13288 2338 13386 sw
tri 2338 13288 2436 13386 ne
rect 2436 13288 2790 13386
tri 2790 13288 2888 13386 sw
tri 2888 13288 2986 13386 ne
rect 2986 13288 3340 13386
tri 3340 13288 3438 13386 sw
tri 3438 13288 3536 13386 ne
rect 3536 13288 3890 13386
tri 3890 13288 3988 13386 sw
tri 3988 13288 4086 13386 ne
rect 4086 13288 4440 13386
tri 4440 13288 4538 13386 sw
tri 4538 13288 4636 13386 ne
rect 4636 13288 4990 13386
tri 4990 13288 5088 13386 sw
tri 5088 13288 5186 13386 ne
rect 5186 13288 5540 13386
tri 5540 13288 5638 13386 sw
tri 5638 13288 5736 13386 ne
rect 5736 13288 6090 13386
tri 6090 13288 6188 13386 sw
tri 6188 13288 6286 13386 ne
rect 6286 13288 6640 13386
tri 6640 13288 6738 13386 sw
tri 6738 13288 6836 13386 ne
rect 6836 13288 7190 13386
tri 7190 13288 7288 13386 sw
tri 7288 13288 7386 13386 ne
rect 7386 13288 7740 13386
tri 7740 13288 7838 13386 sw
tri 7838 13288 7936 13386 ne
rect 7936 13288 8290 13386
tri 8290 13288 8388 13386 sw
tri 8388 13288 8486 13386 ne
rect 8486 13288 8840 13386
tri 8840 13288 8938 13386 sw
tri 8938 13288 9036 13386 ne
rect 9036 13288 9390 13386
tri 9390 13288 9488 13386 sw
tri 9488 13288 9586 13386 ne
rect 9586 13288 9940 13386
tri 9940 13288 10038 13386 sw
tri 10038 13288 10136 13386 ne
rect 10136 13288 10490 13386
tri 10490 13288 10588 13386 sw
tri 10588 13288 10686 13386 ne
rect 10686 13288 11040 13386
tri 11040 13288 11138 13386 sw
tri 11138 13288 11236 13386 ne
rect 11236 13288 11590 13386
tri 11590 13288 11688 13386 sw
tri 11688 13288 11786 13386 ne
rect 11786 13288 12140 13386
tri 12140 13288 12238 13386 sw
tri 12238 13288 12336 13386 ne
rect 12336 13288 12690 13386
tri 12690 13288 12788 13386 sw
tri 12788 13288 12886 13386 ne
rect 12886 13338 13200 13386
tri 13200 13338 13288 13426 sw
tri 13298 13338 13386 13426 ne
rect 13386 13390 13440 13426
rect 13560 13390 15775 13510
rect 13386 13338 15775 13390
rect 12886 13288 13288 13338
rect -1025 13200 -412 13288
tri -412 13200 -324 13288 sw
tri -314 13200 -226 13288 ne
rect -226 13200 138 13288
tri 138 13200 226 13288 sw
tri 236 13200 324 13288 ne
rect 324 13200 688 13288
tri 688 13200 776 13288 sw
tri 786 13200 874 13288 ne
rect 874 13200 1238 13288
tri 1238 13200 1326 13288 sw
tri 1336 13200 1424 13288 ne
rect 1424 13200 1788 13288
tri 1788 13200 1876 13288 sw
tri 1886 13200 1974 13288 ne
rect 1974 13200 2338 13288
tri 2338 13200 2426 13288 sw
tri 2436 13200 2524 13288 ne
rect 2524 13200 2888 13288
tri 2888 13200 2976 13288 sw
tri 2986 13200 3074 13288 ne
rect 3074 13200 3438 13288
tri 3438 13200 3526 13288 sw
tri 3536 13200 3624 13288 ne
rect 3624 13200 3988 13288
tri 3988 13200 4076 13288 sw
tri 4086 13200 4174 13288 ne
rect 4174 13200 4538 13288
tri 4538 13200 4626 13288 sw
tri 4636 13200 4724 13288 ne
rect 4724 13200 5088 13288
tri 5088 13200 5176 13288 sw
tri 5186 13200 5274 13288 ne
rect 5274 13200 5638 13288
tri 5638 13200 5726 13288 sw
tri 5736 13200 5824 13288 ne
rect 5824 13200 6188 13288
tri 6188 13200 6276 13288 sw
tri 6286 13200 6374 13288 ne
rect 6374 13200 6738 13288
tri 6738 13200 6826 13288 sw
tri 6836 13200 6924 13288 ne
rect 6924 13200 7288 13288
tri 7288 13200 7376 13288 sw
tri 7386 13200 7474 13288 ne
rect 7474 13200 7838 13288
tri 7838 13200 7926 13288 sw
tri 7936 13200 8024 13288 ne
rect 8024 13200 8388 13288
tri 8388 13200 8476 13288 sw
tri 8486 13200 8574 13288 ne
rect 8574 13200 8938 13288
tri 8938 13200 9026 13288 sw
tri 9036 13200 9124 13288 ne
rect 9124 13200 9488 13288
tri 9488 13200 9576 13288 sw
tri 9586 13200 9674 13288 ne
rect 9674 13200 10038 13288
tri 10038 13200 10126 13288 sw
tri 10136 13200 10224 13288 ne
rect 10224 13200 10588 13288
tri 10588 13200 10676 13288 sw
tri 10686 13200 10774 13288 ne
rect 10774 13200 11138 13288
tri 11138 13200 11226 13288 sw
tri 11236 13200 11324 13288 ne
rect 11324 13200 11688 13288
tri 11688 13200 11776 13288 sw
tri 11786 13200 11874 13288 ne
rect 11874 13200 12238 13288
tri 12238 13200 12326 13288 sw
tri 12336 13200 12424 13288 ne
rect 12424 13200 12788 13288
tri 12788 13200 12876 13288 sw
tri 12886 13200 12974 13288 ne
rect 12974 13258 13288 13288
tri 13288 13258 13368 13338 sw
tri 13386 13258 13466 13338 ne
rect 13466 13258 14075 13338
rect 12974 13200 13368 13258
rect -1025 13160 -324 13200
tri -324 13160 -284 13200 sw
tri -226 13160 -186 13200 ne
rect -186 13160 226 13200
tri 226 13160 266 13200 sw
tri 324 13160 364 13200 ne
rect 364 13160 776 13200
tri 776 13160 816 13200 sw
tri 874 13160 914 13200 ne
rect 914 13160 1326 13200
tri 1326 13160 1366 13200 sw
tri 1424 13160 1464 13200 ne
rect 1464 13160 1876 13200
tri 1876 13160 1916 13200 sw
tri 1974 13160 2014 13200 ne
rect 2014 13160 2426 13200
tri 2426 13160 2466 13200 sw
tri 2524 13160 2564 13200 ne
rect 2564 13160 2976 13200
tri 2976 13160 3016 13200 sw
tri 3074 13160 3114 13200 ne
rect 3114 13160 3526 13200
tri 3526 13160 3566 13200 sw
tri 3624 13160 3664 13200 ne
rect 3664 13160 4076 13200
tri 4076 13160 4116 13200 sw
tri 4174 13160 4214 13200 ne
rect 4214 13160 4626 13200
tri 4626 13160 4666 13200 sw
tri 4724 13160 4764 13200 ne
rect 4764 13160 5176 13200
tri 5176 13160 5216 13200 sw
tri 5274 13160 5314 13200 ne
rect 5314 13160 5726 13200
tri 5726 13160 5766 13200 sw
tri 5824 13160 5864 13200 ne
rect 5864 13160 6276 13200
tri 6276 13160 6316 13200 sw
tri 6374 13160 6414 13200 ne
rect 6414 13160 6826 13200
tri 6826 13160 6866 13200 sw
tri 6924 13160 6964 13200 ne
rect 6964 13160 7376 13200
tri 7376 13160 7416 13200 sw
tri 7474 13160 7514 13200 ne
rect 7514 13160 7926 13200
tri 7926 13160 7966 13200 sw
tri 8024 13160 8064 13200 ne
rect 8064 13160 8476 13200
tri 8476 13160 8516 13200 sw
tri 8574 13160 8614 13200 ne
rect 8614 13160 9026 13200
tri 9026 13160 9066 13200 sw
tri 9124 13160 9164 13200 ne
rect 9164 13160 9576 13200
tri 9576 13160 9616 13200 sw
tri 9674 13160 9714 13200 ne
rect 9714 13160 10126 13200
tri 10126 13160 10166 13200 sw
tri 10224 13160 10264 13200 ne
rect 10264 13160 10676 13200
tri 10676 13160 10716 13200 sw
tri 10774 13160 10814 13200 ne
rect 10814 13160 11226 13200
tri 11226 13160 11266 13200 sw
tri 11324 13160 11364 13200 ne
rect 11364 13160 11776 13200
tri 11776 13160 11816 13200 sw
tri 11874 13160 11914 13200 ne
rect 11914 13160 12326 13200
tri 12326 13160 12366 13200 sw
tri 12424 13160 12464 13200 ne
rect 12464 13160 12876 13200
tri 12876 13160 12916 13200 sw
tri 12974 13160 13014 13200 ne
rect 13014 13160 13368 13200
tri 13368 13160 13466 13258 sw
tri 13466 13160 13564 13258 ne
rect 13564 13238 14075 13258
rect 14175 13238 15775 13338
rect 13564 13160 15775 13238
rect -1025 13112 -284 13160
rect -1025 13012 -925 13112
rect -825 13062 -284 13112
tri -284 13062 -186 13160 sw
tri -186 13062 -88 13160 ne
rect -88 13062 266 13160
tri 266 13062 364 13160 sw
tri 364 13062 462 13160 ne
rect 462 13062 816 13160
tri 816 13062 914 13160 sw
tri 914 13062 1012 13160 ne
rect 1012 13062 1366 13160
tri 1366 13062 1464 13160 sw
tri 1464 13062 1562 13160 ne
rect 1562 13062 1916 13160
tri 1916 13062 2014 13160 sw
tri 2014 13062 2112 13160 ne
rect 2112 13062 2466 13160
tri 2466 13062 2564 13160 sw
tri 2564 13062 2662 13160 ne
rect 2662 13062 3016 13160
tri 3016 13062 3114 13160 sw
tri 3114 13062 3212 13160 ne
rect 3212 13062 3566 13160
tri 3566 13062 3664 13160 sw
tri 3664 13062 3762 13160 ne
rect 3762 13062 4116 13160
tri 4116 13062 4214 13160 sw
tri 4214 13062 4312 13160 ne
rect 4312 13062 4666 13160
tri 4666 13062 4764 13160 sw
tri 4764 13062 4862 13160 ne
rect 4862 13062 5216 13160
tri 5216 13062 5314 13160 sw
tri 5314 13062 5412 13160 ne
rect 5412 13062 5766 13160
tri 5766 13062 5864 13160 sw
tri 5864 13062 5962 13160 ne
rect 5962 13062 6316 13160
tri 6316 13062 6414 13160 sw
tri 6414 13062 6512 13160 ne
rect 6512 13062 6866 13160
tri 6866 13062 6964 13160 sw
tri 6964 13062 7062 13160 ne
rect 7062 13062 7416 13160
tri 7416 13062 7514 13160 sw
tri 7514 13062 7612 13160 ne
rect 7612 13062 7966 13160
tri 7966 13062 8064 13160 sw
tri 8064 13062 8162 13160 ne
rect 8162 13062 8516 13160
tri 8516 13062 8614 13160 sw
tri 8614 13062 8712 13160 ne
rect 8712 13062 9066 13160
tri 9066 13062 9164 13160 sw
tri 9164 13062 9262 13160 ne
rect 9262 13062 9616 13160
tri 9616 13062 9714 13160 sw
tri 9714 13062 9812 13160 ne
rect 9812 13062 10166 13160
tri 10166 13062 10264 13160 sw
tri 10264 13062 10362 13160 ne
rect 10362 13062 10716 13160
tri 10716 13062 10814 13160 sw
tri 10814 13062 10912 13160 ne
rect 10912 13062 11266 13160
tri 11266 13062 11364 13160 sw
tri 11364 13062 11462 13160 ne
rect 11462 13062 11816 13160
tri 11816 13062 11914 13160 sw
tri 11914 13062 12012 13160 ne
rect 12012 13062 12366 13160
tri 12366 13062 12464 13160 sw
tri 12464 13062 12562 13160 ne
rect 12562 13062 12916 13160
tri 12916 13062 13014 13160 sw
tri 13014 13062 13112 13160 ne
rect 13112 13062 13466 13160
tri 13466 13062 13564 13160 sw
tri 13564 13062 13662 13160 ne
rect 13662 13062 15775 13160
rect -825 13012 -186 13062
rect -1025 12964 -186 13012
tri -186 12964 -88 13062 sw
tri -88 12964 10 13062 ne
rect 10 12964 364 13062
tri 364 12964 462 13062 sw
tri 462 12964 560 13062 ne
rect 560 12964 914 13062
tri 914 12964 1012 13062 sw
tri 1012 12964 1110 13062 ne
rect 1110 12964 1464 13062
tri 1464 12964 1562 13062 sw
tri 1562 12964 1660 13062 ne
rect 1660 12964 2014 13062
tri 2014 12964 2112 13062 sw
tri 2112 12964 2210 13062 ne
rect 2210 12964 2564 13062
tri 2564 12964 2662 13062 sw
tri 2662 12964 2760 13062 ne
rect 2760 12964 3114 13062
tri 3114 12964 3212 13062 sw
tri 3212 12964 3310 13062 ne
rect 3310 12964 3664 13062
tri 3664 12964 3762 13062 sw
tri 3762 12964 3860 13062 ne
rect 3860 12964 4214 13062
tri 4214 12964 4312 13062 sw
tri 4312 12964 4410 13062 ne
rect 4410 12964 4764 13062
tri 4764 12964 4862 13062 sw
tri 4862 12964 4960 13062 ne
rect 4960 12964 5314 13062
tri 5314 12964 5412 13062 sw
tri 5412 12964 5510 13062 ne
rect 5510 12964 5864 13062
tri 5864 12964 5962 13062 sw
tri 5962 12964 6060 13062 ne
rect 6060 12964 6414 13062
tri 6414 12964 6512 13062 sw
tri 6512 12964 6610 13062 ne
rect 6610 12964 6964 13062
tri 6964 12964 7062 13062 sw
tri 7062 12964 7160 13062 ne
rect 7160 12964 7514 13062
tri 7514 12964 7612 13062 sw
tri 7612 12964 7710 13062 ne
rect 7710 12964 8064 13062
tri 8064 12964 8162 13062 sw
tri 8162 12964 8260 13062 ne
rect 8260 12964 8614 13062
tri 8614 12964 8712 13062 sw
tri 8712 12964 8810 13062 ne
rect 8810 12964 9164 13062
tri 9164 12964 9262 13062 sw
tri 9262 12964 9360 13062 ne
rect 9360 12964 9714 13062
tri 9714 12964 9812 13062 sw
tri 9812 12964 9910 13062 ne
rect 9910 12964 10264 13062
tri 10264 12964 10362 13062 sw
tri 10362 12964 10460 13062 ne
rect 10460 12964 10814 13062
tri 10814 12964 10912 13062 sw
tri 10912 12964 11010 13062 ne
rect 11010 12964 11364 13062
tri 11364 12964 11462 13062 sw
tri 11462 12964 11560 13062 ne
rect 11560 12964 11914 13062
tri 11914 12964 12012 13062 sw
tri 12012 12964 12110 13062 ne
rect 12110 12964 12464 13062
tri 12464 12964 12562 13062 sw
tri 12562 12964 12660 13062 ne
rect 12660 12964 13014 13062
tri 13014 12964 13112 13062 sw
tri 13112 12964 13210 13062 ne
rect 13210 12964 13564 13062
tri 13564 12964 13662 13062 sw
rect -1025 12960 -88 12964
rect -1025 12840 -310 12960
rect -190 12876 -88 12960
tri -88 12876 0 12964 sw
tri 10 12876 98 12964 ne
rect 98 12960 462 12964
rect 98 12876 240 12960
rect -190 12840 0 12876
rect -1025 12836 0 12840
tri 0 12836 40 12876 sw
tri 98 12836 138 12876 ne
rect 138 12840 240 12876
rect 360 12876 462 12960
tri 462 12876 550 12964 sw
tri 560 12876 648 12964 ne
rect 648 12960 1012 12964
rect 648 12876 790 12960
rect 360 12840 550 12876
rect 138 12836 550 12840
tri -412 12738 -314 12836 ne
rect -314 12738 40 12836
tri 40 12738 138 12836 sw
tri 138 12738 236 12836 ne
rect 236 12788 550 12836
tri 550 12788 638 12876 sw
tri 648 12788 736 12876 ne
rect 736 12840 790 12876
rect 910 12876 1012 12960
tri 1012 12876 1100 12964 sw
tri 1110 12876 1198 12964 ne
rect 1198 12960 1562 12964
rect 1198 12876 1340 12960
rect 910 12840 1100 12876
rect 736 12836 1100 12840
tri 1100 12836 1140 12876 sw
tri 1198 12836 1238 12876 ne
rect 1238 12840 1340 12876
rect 1460 12876 1562 12960
tri 1562 12876 1650 12964 sw
tri 1660 12876 1748 12964 ne
rect 1748 12960 2112 12964
rect 1748 12876 1890 12960
rect 1460 12840 1650 12876
rect 1238 12836 1650 12840
rect 736 12788 1140 12836
rect 236 12738 638 12788
rect -2525 12650 -412 12738
tri -412 12650 -324 12738 sw
tri -314 12650 -226 12738 ne
rect -226 12650 138 12738
tri 138 12650 226 12738 sw
tri 236 12650 324 12738 ne
rect 324 12708 638 12738
tri 638 12708 718 12788 sw
tri 736 12708 816 12788 ne
rect 816 12738 1140 12788
tri 1140 12738 1238 12836 sw
tri 1238 12738 1336 12836 ne
rect 1336 12788 1650 12836
tri 1650 12788 1738 12876 sw
tri 1748 12788 1836 12876 ne
rect 1836 12840 1890 12876
rect 2010 12876 2112 12960
tri 2112 12876 2200 12964 sw
tri 2210 12876 2298 12964 ne
rect 2298 12960 2662 12964
rect 2298 12876 2440 12960
rect 2010 12840 2200 12876
rect 1836 12836 2200 12840
tri 2200 12836 2240 12876 sw
tri 2298 12836 2338 12876 ne
rect 2338 12840 2440 12876
rect 2560 12876 2662 12960
tri 2662 12876 2750 12964 sw
tri 2760 12876 2848 12964 ne
rect 2848 12960 3212 12964
rect 2848 12876 2990 12960
rect 2560 12840 2750 12876
rect 2338 12836 2750 12840
rect 1836 12788 2240 12836
rect 1336 12738 1738 12788
rect 816 12708 1238 12738
rect 324 12650 718 12708
rect -2525 12610 -324 12650
tri -324 12610 -284 12650 sw
tri -226 12610 -186 12650 ne
rect -186 12610 226 12650
tri 226 12610 266 12650 sw
tri 324 12610 364 12650 ne
rect 364 12610 718 12650
tri 718 12610 816 12708 sw
tri 816 12610 914 12708 ne
rect 914 12650 1238 12708
tri 1238 12650 1326 12738 sw
tri 1336 12650 1424 12738 ne
rect 1424 12708 1738 12738
tri 1738 12708 1818 12788 sw
tri 1836 12708 1916 12788 ne
rect 1916 12738 2240 12788
tri 2240 12738 2338 12836 sw
tri 2338 12738 2436 12836 ne
rect 2436 12788 2750 12836
tri 2750 12788 2838 12876 sw
tri 2848 12788 2936 12876 ne
rect 2936 12840 2990 12876
rect 3110 12876 3212 12960
tri 3212 12876 3300 12964 sw
tri 3310 12876 3398 12964 ne
rect 3398 12960 3762 12964
rect 3398 12876 3540 12960
rect 3110 12840 3300 12876
rect 2936 12836 3300 12840
tri 3300 12836 3340 12876 sw
tri 3398 12836 3438 12876 ne
rect 3438 12840 3540 12876
rect 3660 12876 3762 12960
tri 3762 12876 3850 12964 sw
tri 3860 12876 3948 12964 ne
rect 3948 12960 4312 12964
rect 3948 12876 4090 12960
rect 3660 12840 3850 12876
rect 3438 12836 3850 12840
rect 2936 12788 3340 12836
rect 2436 12738 2838 12788
rect 1916 12708 2338 12738
rect 1424 12650 1818 12708
rect 914 12610 1326 12650
tri 1326 12610 1366 12650 sw
tri 1424 12610 1464 12650 ne
rect 1464 12610 1818 12650
tri 1818 12610 1916 12708 sw
tri 1916 12610 2014 12708 ne
rect 2014 12650 2338 12708
tri 2338 12650 2426 12738 sw
tri 2436 12650 2524 12738 ne
rect 2524 12708 2838 12738
tri 2838 12708 2918 12788 sw
tri 2936 12708 3016 12788 ne
rect 3016 12738 3340 12788
tri 3340 12738 3438 12836 sw
tri 3438 12738 3536 12836 ne
rect 3536 12788 3850 12836
tri 3850 12788 3938 12876 sw
tri 3948 12788 4036 12876 ne
rect 4036 12840 4090 12876
rect 4210 12876 4312 12960
tri 4312 12876 4400 12964 sw
tri 4410 12876 4498 12964 ne
rect 4498 12960 4862 12964
rect 4498 12876 4640 12960
rect 4210 12840 4400 12876
rect 4036 12836 4400 12840
tri 4400 12836 4440 12876 sw
tri 4498 12836 4538 12876 ne
rect 4538 12840 4640 12876
rect 4760 12876 4862 12960
tri 4862 12876 4950 12964 sw
tri 4960 12876 5048 12964 ne
rect 5048 12960 5412 12964
rect 5048 12876 5190 12960
rect 4760 12840 4950 12876
rect 4538 12836 4950 12840
rect 4036 12788 4440 12836
rect 3536 12738 3938 12788
rect 3016 12708 3438 12738
rect 2524 12650 2918 12708
rect 2014 12610 2426 12650
tri 2426 12610 2466 12650 sw
tri 2524 12610 2564 12650 ne
rect 2564 12610 2918 12650
tri 2918 12610 3016 12708 sw
tri 3016 12610 3114 12708 ne
rect 3114 12650 3438 12708
tri 3438 12650 3526 12738 sw
tri 3536 12650 3624 12738 ne
rect 3624 12708 3938 12738
tri 3938 12708 4018 12788 sw
tri 4036 12708 4116 12788 ne
rect 4116 12738 4440 12788
tri 4440 12738 4538 12836 sw
tri 4538 12738 4636 12836 ne
rect 4636 12788 4950 12836
tri 4950 12788 5038 12876 sw
tri 5048 12788 5136 12876 ne
rect 5136 12840 5190 12876
rect 5310 12876 5412 12960
tri 5412 12876 5500 12964 sw
tri 5510 12876 5598 12964 ne
rect 5598 12960 5962 12964
rect 5598 12876 5740 12960
rect 5310 12840 5500 12876
rect 5136 12836 5500 12840
tri 5500 12836 5540 12876 sw
tri 5598 12836 5638 12876 ne
rect 5638 12840 5740 12876
rect 5860 12876 5962 12960
tri 5962 12876 6050 12964 sw
tri 6060 12876 6148 12964 ne
rect 6148 12960 6512 12964
rect 6148 12876 6290 12960
rect 5860 12840 6050 12876
rect 5638 12836 6050 12840
rect 5136 12788 5540 12836
rect 4636 12738 5038 12788
rect 4116 12708 4538 12738
rect 3624 12650 4018 12708
rect 3114 12610 3526 12650
tri 3526 12610 3566 12650 sw
tri 3624 12610 3664 12650 ne
rect 3664 12610 4018 12650
tri 4018 12610 4116 12708 sw
tri 4116 12610 4214 12708 ne
rect 4214 12650 4538 12708
tri 4538 12650 4626 12738 sw
tri 4636 12650 4724 12738 ne
rect 4724 12708 5038 12738
tri 5038 12708 5118 12788 sw
tri 5136 12708 5216 12788 ne
rect 5216 12738 5540 12788
tri 5540 12738 5638 12836 sw
tri 5638 12738 5736 12836 ne
rect 5736 12788 6050 12836
tri 6050 12788 6138 12876 sw
tri 6148 12788 6236 12876 ne
rect 6236 12840 6290 12876
rect 6410 12876 6512 12960
tri 6512 12876 6600 12964 sw
tri 6610 12876 6698 12964 ne
rect 6698 12960 7062 12964
rect 6698 12876 6840 12960
rect 6410 12840 6600 12876
rect 6236 12836 6600 12840
tri 6600 12836 6640 12876 sw
tri 6698 12836 6738 12876 ne
rect 6738 12840 6840 12876
rect 6960 12876 7062 12960
tri 7062 12876 7150 12964 sw
tri 7160 12876 7248 12964 ne
rect 7248 12960 7612 12964
rect 7248 12876 7390 12960
rect 6960 12840 7150 12876
rect 6738 12836 7150 12840
rect 6236 12788 6640 12836
rect 5736 12738 6138 12788
rect 5216 12708 5638 12738
rect 4724 12650 5118 12708
rect 4214 12610 4626 12650
tri 4626 12610 4666 12650 sw
tri 4724 12610 4764 12650 ne
rect 4764 12610 5118 12650
tri 5118 12610 5216 12708 sw
tri 5216 12610 5314 12708 ne
rect 5314 12650 5638 12708
tri 5638 12650 5726 12738 sw
tri 5736 12650 5824 12738 ne
rect 5824 12708 6138 12738
tri 6138 12708 6218 12788 sw
tri 6236 12708 6316 12788 ne
rect 6316 12738 6640 12788
tri 6640 12738 6738 12836 sw
tri 6738 12738 6836 12836 ne
rect 6836 12788 7150 12836
tri 7150 12788 7238 12876 sw
tri 7248 12788 7336 12876 ne
rect 7336 12840 7390 12876
rect 7510 12876 7612 12960
tri 7612 12876 7700 12964 sw
tri 7710 12876 7798 12964 ne
rect 7798 12960 8162 12964
rect 7798 12876 7940 12960
rect 7510 12840 7700 12876
rect 7336 12836 7700 12840
tri 7700 12836 7740 12876 sw
tri 7798 12836 7838 12876 ne
rect 7838 12840 7940 12876
rect 8060 12876 8162 12960
tri 8162 12876 8250 12964 sw
tri 8260 12876 8348 12964 ne
rect 8348 12960 8712 12964
rect 8348 12876 8490 12960
rect 8060 12840 8250 12876
rect 7838 12836 8250 12840
rect 7336 12788 7740 12836
rect 6836 12738 7238 12788
rect 6316 12708 6738 12738
rect 5824 12650 6218 12708
rect 5314 12610 5726 12650
tri 5726 12610 5766 12650 sw
tri 5824 12610 5864 12650 ne
rect 5864 12610 6218 12650
tri 6218 12610 6316 12708 sw
tri 6316 12610 6414 12708 ne
rect 6414 12650 6738 12708
tri 6738 12650 6826 12738 sw
tri 6836 12650 6924 12738 ne
rect 6924 12708 7238 12738
tri 7238 12708 7318 12788 sw
tri 7336 12708 7416 12788 ne
rect 7416 12738 7740 12788
tri 7740 12738 7838 12836 sw
tri 7838 12738 7936 12836 ne
rect 7936 12788 8250 12836
tri 8250 12788 8338 12876 sw
tri 8348 12788 8436 12876 ne
rect 8436 12840 8490 12876
rect 8610 12876 8712 12960
tri 8712 12876 8800 12964 sw
tri 8810 12876 8898 12964 ne
rect 8898 12960 9262 12964
rect 8898 12876 9040 12960
rect 8610 12840 8800 12876
rect 8436 12836 8800 12840
tri 8800 12836 8840 12876 sw
tri 8898 12836 8938 12876 ne
rect 8938 12840 9040 12876
rect 9160 12876 9262 12960
tri 9262 12876 9350 12964 sw
tri 9360 12876 9448 12964 ne
rect 9448 12960 9812 12964
rect 9448 12876 9590 12960
rect 9160 12840 9350 12876
rect 8938 12836 9350 12840
rect 8436 12788 8840 12836
rect 7936 12738 8338 12788
rect 7416 12708 7838 12738
rect 6924 12650 7318 12708
rect 6414 12610 6826 12650
tri 6826 12610 6866 12650 sw
tri 6924 12610 6964 12650 ne
rect 6964 12610 7318 12650
tri 7318 12610 7416 12708 sw
tri 7416 12610 7514 12708 ne
rect 7514 12650 7838 12708
tri 7838 12650 7926 12738 sw
tri 7936 12650 8024 12738 ne
rect 8024 12708 8338 12738
tri 8338 12708 8418 12788 sw
tri 8436 12708 8516 12788 ne
rect 8516 12738 8840 12788
tri 8840 12738 8938 12836 sw
tri 8938 12738 9036 12836 ne
rect 9036 12788 9350 12836
tri 9350 12788 9438 12876 sw
tri 9448 12788 9536 12876 ne
rect 9536 12840 9590 12876
rect 9710 12876 9812 12960
tri 9812 12876 9900 12964 sw
tri 9910 12876 9998 12964 ne
rect 9998 12960 10362 12964
rect 9998 12876 10140 12960
rect 9710 12840 9900 12876
rect 9536 12836 9900 12840
tri 9900 12836 9940 12876 sw
tri 9998 12836 10038 12876 ne
rect 10038 12840 10140 12876
rect 10260 12876 10362 12960
tri 10362 12876 10450 12964 sw
tri 10460 12876 10548 12964 ne
rect 10548 12960 10912 12964
rect 10548 12876 10690 12960
rect 10260 12840 10450 12876
rect 10038 12836 10450 12840
rect 9536 12788 9940 12836
rect 9036 12738 9438 12788
rect 8516 12708 8938 12738
rect 8024 12650 8418 12708
rect 7514 12610 7926 12650
tri 7926 12610 7966 12650 sw
tri 8024 12610 8064 12650 ne
rect 8064 12610 8418 12650
tri 8418 12610 8516 12708 sw
tri 8516 12610 8614 12708 ne
rect 8614 12650 8938 12708
tri 8938 12650 9026 12738 sw
tri 9036 12650 9124 12738 ne
rect 9124 12708 9438 12738
tri 9438 12708 9518 12788 sw
tri 9536 12708 9616 12788 ne
rect 9616 12738 9940 12788
tri 9940 12738 10038 12836 sw
tri 10038 12738 10136 12836 ne
rect 10136 12788 10450 12836
tri 10450 12788 10538 12876 sw
tri 10548 12788 10636 12876 ne
rect 10636 12840 10690 12876
rect 10810 12876 10912 12960
tri 10912 12876 11000 12964 sw
tri 11010 12876 11098 12964 ne
rect 11098 12960 11462 12964
rect 11098 12876 11240 12960
rect 10810 12840 11000 12876
rect 10636 12836 11000 12840
tri 11000 12836 11040 12876 sw
tri 11098 12836 11138 12876 ne
rect 11138 12840 11240 12876
rect 11360 12876 11462 12960
tri 11462 12876 11550 12964 sw
tri 11560 12876 11648 12964 ne
rect 11648 12960 12012 12964
rect 11648 12876 11790 12960
rect 11360 12840 11550 12876
rect 11138 12836 11550 12840
rect 10636 12788 11040 12836
rect 10136 12738 10538 12788
rect 9616 12708 10038 12738
rect 9124 12650 9518 12708
rect 8614 12610 9026 12650
tri 9026 12610 9066 12650 sw
tri 9124 12610 9164 12650 ne
rect 9164 12610 9518 12650
tri 9518 12610 9616 12708 sw
tri 9616 12610 9714 12708 ne
rect 9714 12650 10038 12708
tri 10038 12650 10126 12738 sw
tri 10136 12650 10224 12738 ne
rect 10224 12708 10538 12738
tri 10538 12708 10618 12788 sw
tri 10636 12708 10716 12788 ne
rect 10716 12738 11040 12788
tri 11040 12738 11138 12836 sw
tri 11138 12738 11236 12836 ne
rect 11236 12788 11550 12836
tri 11550 12788 11638 12876 sw
tri 11648 12788 11736 12876 ne
rect 11736 12840 11790 12876
rect 11910 12876 12012 12960
tri 12012 12876 12100 12964 sw
tri 12110 12876 12198 12964 ne
rect 12198 12960 12562 12964
rect 12198 12876 12340 12960
rect 11910 12840 12100 12876
rect 11736 12836 12100 12840
tri 12100 12836 12140 12876 sw
tri 12198 12836 12238 12876 ne
rect 12238 12840 12340 12876
rect 12460 12876 12562 12960
tri 12562 12876 12650 12964 sw
tri 12660 12876 12748 12964 ne
rect 12748 12960 13112 12964
rect 12748 12876 12890 12960
rect 12460 12840 12650 12876
rect 12238 12836 12650 12840
rect 11736 12788 12140 12836
rect 11236 12738 11638 12788
rect 10716 12708 11138 12738
rect 10224 12650 10618 12708
rect 9714 12610 10126 12650
tri 10126 12610 10166 12650 sw
tri 10224 12610 10264 12650 ne
rect 10264 12610 10618 12650
tri 10618 12610 10716 12708 sw
tri 10716 12610 10814 12708 ne
rect 10814 12650 11138 12708
tri 11138 12650 11226 12738 sw
tri 11236 12650 11324 12738 ne
rect 11324 12708 11638 12738
tri 11638 12708 11718 12788 sw
tri 11736 12708 11816 12788 ne
rect 11816 12738 12140 12788
tri 12140 12738 12238 12836 sw
tri 12238 12738 12336 12836 ne
rect 12336 12788 12650 12836
tri 12650 12788 12738 12876 sw
tri 12748 12788 12836 12876 ne
rect 12836 12840 12890 12876
rect 13010 12876 13112 12960
tri 13112 12876 13200 12964 sw
tri 13210 12876 13298 12964 ne
rect 13298 12960 14275 12964
rect 13298 12876 13440 12960
rect 13010 12840 13200 12876
rect 12836 12836 13200 12840
tri 13200 12836 13240 12876 sw
tri 13298 12836 13338 12876 ne
rect 13338 12840 13440 12876
rect 13560 12840 14275 12960
rect 13338 12836 14275 12840
rect 12836 12788 13240 12836
rect 12336 12738 12738 12788
rect 11816 12708 12238 12738
rect 11324 12650 11718 12708
rect 10814 12610 11226 12650
tri 11226 12610 11266 12650 sw
tri 11324 12610 11364 12650 ne
rect 11364 12610 11718 12650
tri 11718 12610 11816 12708 sw
tri 11816 12610 11914 12708 ne
rect 11914 12650 12238 12708
tri 12238 12650 12326 12738 sw
tri 12336 12650 12424 12738 ne
rect 12424 12708 12738 12738
tri 12738 12708 12818 12788 sw
tri 12836 12708 12916 12788 ne
rect 12916 12738 13240 12788
tri 13240 12738 13338 12836 sw
tri 13338 12738 13436 12836 ne
rect 13436 12738 14275 12836
rect 12916 12708 13338 12738
rect 12424 12650 12818 12708
rect 11914 12610 12326 12650
tri 12326 12610 12366 12650 sw
tri 12424 12610 12464 12650 ne
rect 12464 12610 12818 12650
tri 12818 12610 12916 12708 sw
tri 12916 12610 13014 12708 ne
rect 13014 12650 13338 12708
tri 13338 12650 13426 12738 sw
tri 13436 12650 13524 12738 ne
rect 13524 12650 14275 12738
rect 13014 12610 13426 12650
tri 13426 12610 13466 12650 sw
tri 13524 12610 13564 12650 ne
rect 13564 12610 14275 12650
rect -2525 12512 -284 12610
tri -284 12512 -186 12610 sw
tri -186 12512 -88 12610 ne
rect -88 12512 266 12610
tri 266 12512 364 12610 sw
tri 364 12512 462 12610 ne
rect 462 12512 816 12610
tri 816 12512 914 12610 sw
tri 914 12512 1012 12610 ne
rect 1012 12512 1366 12610
tri 1366 12512 1464 12610 sw
tri 1464 12512 1562 12610 ne
rect 1562 12512 1916 12610
tri 1916 12512 2014 12610 sw
tri 2014 12512 2112 12610 ne
rect 2112 12512 2466 12610
tri 2466 12512 2564 12610 sw
tri 2564 12512 2662 12610 ne
rect 2662 12512 3016 12610
tri 3016 12512 3114 12610 sw
tri 3114 12512 3212 12610 ne
rect 3212 12512 3566 12610
tri 3566 12512 3664 12610 sw
tri 3664 12512 3762 12610 ne
rect 3762 12512 4116 12610
tri 4116 12512 4214 12610 sw
tri 4214 12512 4312 12610 ne
rect 4312 12512 4666 12610
tri 4666 12512 4764 12610 sw
tri 4764 12512 4862 12610 ne
rect 4862 12512 5216 12610
tri 5216 12512 5314 12610 sw
tri 5314 12512 5412 12610 ne
rect 5412 12512 5766 12610
tri 5766 12512 5864 12610 sw
tri 5864 12512 5962 12610 ne
rect 5962 12512 6316 12610
tri 6316 12512 6414 12610 sw
tri 6414 12512 6512 12610 ne
rect 6512 12512 6866 12610
tri 6866 12512 6964 12610 sw
tri 6964 12512 7062 12610 ne
rect 7062 12512 7416 12610
tri 7416 12512 7514 12610 sw
tri 7514 12512 7612 12610 ne
rect 7612 12512 7966 12610
tri 7966 12512 8064 12610 sw
tri 8064 12512 8162 12610 ne
rect 8162 12512 8516 12610
tri 8516 12512 8614 12610 sw
tri 8614 12512 8712 12610 ne
rect 8712 12512 9066 12610
tri 9066 12512 9164 12610 sw
tri 9164 12512 9262 12610 ne
rect 9262 12512 9616 12610
tri 9616 12512 9714 12610 sw
tri 9714 12512 9812 12610 ne
rect 9812 12512 10166 12610
tri 10166 12512 10264 12610 sw
tri 10264 12512 10362 12610 ne
rect 10362 12512 10716 12610
tri 10716 12512 10814 12610 sw
tri 10814 12512 10912 12610 ne
rect 10912 12512 11266 12610
tri 11266 12512 11364 12610 sw
tri 11364 12512 11462 12610 ne
rect 11462 12512 11816 12610
tri 11816 12512 11914 12610 sw
tri 11914 12512 12012 12610 ne
rect 12012 12512 12366 12610
tri 12366 12512 12464 12610 sw
tri 12464 12512 12562 12610 ne
rect 12562 12512 12916 12610
tri 12916 12512 13014 12610 sw
tri 13014 12512 13112 12610 ne
rect 13112 12512 13466 12610
tri 13466 12512 13564 12610 sw
tri 13564 12512 13662 12610 ne
rect 13662 12512 14275 12610
rect -2525 12414 -186 12512
tri -186 12414 -88 12512 sw
tri -88 12414 10 12512 ne
rect 10 12414 364 12512
tri 364 12414 462 12512 sw
tri 462 12414 560 12512 ne
rect 560 12414 914 12512
tri 914 12414 1012 12512 sw
tri 1012 12414 1110 12512 ne
rect 1110 12414 1464 12512
tri 1464 12414 1562 12512 sw
tri 1562 12414 1660 12512 ne
rect 1660 12414 2014 12512
tri 2014 12414 2112 12512 sw
tri 2112 12414 2210 12512 ne
rect 2210 12414 2564 12512
tri 2564 12414 2662 12512 sw
tri 2662 12414 2760 12512 ne
rect 2760 12414 3114 12512
tri 3114 12414 3212 12512 sw
tri 3212 12414 3310 12512 ne
rect 3310 12414 3664 12512
tri 3664 12414 3762 12512 sw
tri 3762 12414 3860 12512 ne
rect 3860 12414 4214 12512
tri 4214 12414 4312 12512 sw
tri 4312 12414 4410 12512 ne
rect 4410 12414 4764 12512
tri 4764 12414 4862 12512 sw
tri 4862 12414 4960 12512 ne
rect 4960 12414 5314 12512
tri 5314 12414 5412 12512 sw
tri 5412 12414 5510 12512 ne
rect 5510 12414 5864 12512
tri 5864 12414 5962 12512 sw
tri 5962 12414 6060 12512 ne
rect 6060 12414 6414 12512
tri 6414 12414 6512 12512 sw
tri 6512 12414 6610 12512 ne
rect 6610 12414 6964 12512
tri 6964 12414 7062 12512 sw
tri 7062 12414 7160 12512 ne
rect 7160 12414 7514 12512
tri 7514 12414 7612 12512 sw
tri 7612 12414 7710 12512 ne
rect 7710 12414 8064 12512
tri 8064 12414 8162 12512 sw
tri 8162 12414 8260 12512 ne
rect 8260 12414 8614 12512
tri 8614 12414 8712 12512 sw
tri 8712 12414 8810 12512 ne
rect 8810 12414 9164 12512
tri 9164 12414 9262 12512 sw
tri 9262 12414 9360 12512 ne
rect 9360 12414 9714 12512
tri 9714 12414 9812 12512 sw
tri 9812 12414 9910 12512 ne
rect 9910 12414 10264 12512
tri 10264 12414 10362 12512 sw
tri 10362 12414 10460 12512 ne
rect 10460 12414 10814 12512
tri 10814 12414 10912 12512 sw
tri 10912 12414 11010 12512 ne
rect 11010 12414 11364 12512
tri 11364 12414 11462 12512 sw
tri 11462 12414 11560 12512 ne
rect 11560 12414 11914 12512
tri 11914 12414 12012 12512 sw
tri 12012 12414 12110 12512 ne
rect 12110 12414 12464 12512
tri 12464 12414 12562 12512 sw
tri 12562 12414 12660 12512 ne
rect 12660 12414 13014 12512
tri 13014 12414 13112 12512 sw
tri 13112 12414 13210 12512 ne
rect 13210 12414 13564 12512
tri 13564 12414 13662 12512 sw
rect 14775 12414 15775 13062
rect -2525 12410 -88 12414
rect -2525 12290 -310 12410
rect -190 12326 -88 12410
tri -88 12326 0 12414 sw
tri 10 12326 98 12414 ne
rect 98 12410 462 12414
rect 98 12326 240 12410
rect -190 12290 0 12326
rect -2525 12286 0 12290
rect -2525 11638 -1525 12286
tri -412 12188 -314 12286 ne
rect -314 12238 0 12286
tri 0 12238 88 12326 sw
tri 98 12238 186 12326 ne
rect 186 12290 240 12326
rect 360 12326 462 12410
tri 462 12326 550 12414 sw
tri 560 12326 648 12414 ne
rect 648 12410 1012 12414
rect 648 12326 790 12410
rect 360 12290 550 12326
rect 186 12286 550 12290
tri 550 12286 590 12326 sw
tri 648 12286 688 12326 ne
rect 688 12290 790 12326
rect 910 12326 1012 12410
tri 1012 12326 1100 12414 sw
tri 1110 12326 1198 12414 ne
rect 1198 12410 1562 12414
rect 1198 12326 1340 12410
rect 910 12290 1100 12326
rect 688 12286 1100 12290
rect 186 12238 590 12286
rect -314 12188 88 12238
rect -1025 12100 -412 12188
tri -412 12100 -324 12188 sw
tri -314 12100 -226 12188 ne
rect -226 12158 88 12188
tri 88 12158 168 12238 sw
tri 186 12158 266 12238 ne
rect 266 12188 590 12238
tri 590 12188 688 12286 sw
tri 688 12188 786 12286 ne
rect 786 12238 1100 12286
tri 1100 12238 1188 12326 sw
tri 1198 12238 1286 12326 ne
rect 1286 12290 1340 12326
rect 1460 12326 1562 12410
tri 1562 12326 1650 12414 sw
tri 1660 12326 1748 12414 ne
rect 1748 12410 2112 12414
rect 1748 12326 1890 12410
rect 1460 12290 1650 12326
rect 1286 12286 1650 12290
tri 1650 12286 1690 12326 sw
tri 1748 12286 1788 12326 ne
rect 1788 12290 1890 12326
rect 2010 12326 2112 12410
tri 2112 12326 2200 12414 sw
tri 2210 12326 2298 12414 ne
rect 2298 12410 2662 12414
rect 2298 12326 2440 12410
rect 2010 12290 2200 12326
rect 1788 12286 2200 12290
rect 1286 12238 1690 12286
rect 786 12188 1188 12238
rect 266 12158 688 12188
rect -226 12100 168 12158
rect -1025 12060 -324 12100
tri -324 12060 -284 12100 sw
tri -226 12060 -186 12100 ne
rect -186 12060 168 12100
tri 168 12060 266 12158 sw
tri 266 12060 364 12158 ne
rect 364 12100 688 12158
tri 688 12100 776 12188 sw
tri 786 12100 874 12188 ne
rect 874 12158 1188 12188
tri 1188 12158 1268 12238 sw
tri 1286 12158 1366 12238 ne
rect 1366 12188 1690 12238
tri 1690 12188 1788 12286 sw
tri 1788 12188 1886 12286 ne
rect 1886 12238 2200 12286
tri 2200 12238 2288 12326 sw
tri 2298 12238 2386 12326 ne
rect 2386 12290 2440 12326
rect 2560 12326 2662 12410
tri 2662 12326 2750 12414 sw
tri 2760 12326 2848 12414 ne
rect 2848 12410 3212 12414
rect 2848 12326 2990 12410
rect 2560 12290 2750 12326
rect 2386 12286 2750 12290
tri 2750 12286 2790 12326 sw
tri 2848 12286 2888 12326 ne
rect 2888 12290 2990 12326
rect 3110 12326 3212 12410
tri 3212 12326 3300 12414 sw
tri 3310 12326 3398 12414 ne
rect 3398 12410 3762 12414
rect 3398 12326 3540 12410
rect 3110 12290 3300 12326
rect 2888 12286 3300 12290
rect 2386 12238 2790 12286
rect 1886 12188 2288 12238
rect 1366 12158 1788 12188
rect 874 12100 1268 12158
rect 364 12060 776 12100
tri 776 12060 816 12100 sw
tri 874 12060 914 12100 ne
rect 914 12060 1268 12100
tri 1268 12060 1366 12158 sw
tri 1366 12060 1464 12158 ne
rect 1464 12100 1788 12158
tri 1788 12100 1876 12188 sw
tri 1886 12100 1974 12188 ne
rect 1974 12158 2288 12188
tri 2288 12158 2368 12238 sw
tri 2386 12158 2466 12238 ne
rect 2466 12188 2790 12238
tri 2790 12188 2888 12286 sw
tri 2888 12188 2986 12286 ne
rect 2986 12238 3300 12286
tri 3300 12238 3388 12326 sw
tri 3398 12238 3486 12326 ne
rect 3486 12290 3540 12326
rect 3660 12326 3762 12410
tri 3762 12326 3850 12414 sw
tri 3860 12326 3948 12414 ne
rect 3948 12410 4312 12414
rect 3948 12326 4090 12410
rect 3660 12290 3850 12326
rect 3486 12286 3850 12290
tri 3850 12286 3890 12326 sw
tri 3948 12286 3988 12326 ne
rect 3988 12290 4090 12326
rect 4210 12326 4312 12410
tri 4312 12326 4400 12414 sw
tri 4410 12326 4498 12414 ne
rect 4498 12410 4862 12414
rect 4498 12326 4640 12410
rect 4210 12290 4400 12326
rect 3988 12286 4400 12290
rect 3486 12238 3890 12286
rect 2986 12188 3388 12238
rect 2466 12158 2888 12188
rect 1974 12100 2368 12158
rect 1464 12060 1876 12100
tri 1876 12060 1916 12100 sw
tri 1974 12060 2014 12100 ne
rect 2014 12060 2368 12100
tri 2368 12060 2466 12158 sw
tri 2466 12060 2564 12158 ne
rect 2564 12100 2888 12158
tri 2888 12100 2976 12188 sw
tri 2986 12100 3074 12188 ne
rect 3074 12158 3388 12188
tri 3388 12158 3468 12238 sw
tri 3486 12158 3566 12238 ne
rect 3566 12188 3890 12238
tri 3890 12188 3988 12286 sw
tri 3988 12188 4086 12286 ne
rect 4086 12238 4400 12286
tri 4400 12238 4488 12326 sw
tri 4498 12238 4586 12326 ne
rect 4586 12290 4640 12326
rect 4760 12326 4862 12410
tri 4862 12326 4950 12414 sw
tri 4960 12326 5048 12414 ne
rect 5048 12410 5412 12414
rect 5048 12326 5190 12410
rect 4760 12290 4950 12326
rect 4586 12286 4950 12290
tri 4950 12286 4990 12326 sw
tri 5048 12286 5088 12326 ne
rect 5088 12290 5190 12326
rect 5310 12326 5412 12410
tri 5412 12326 5500 12414 sw
tri 5510 12326 5598 12414 ne
rect 5598 12410 5962 12414
rect 5598 12326 5740 12410
rect 5310 12290 5500 12326
rect 5088 12286 5500 12290
rect 4586 12238 4990 12286
rect 4086 12188 4488 12238
rect 3566 12158 3988 12188
rect 3074 12100 3468 12158
rect 2564 12060 2976 12100
tri 2976 12060 3016 12100 sw
tri 3074 12060 3114 12100 ne
rect 3114 12060 3468 12100
tri 3468 12060 3566 12158 sw
tri 3566 12060 3664 12158 ne
rect 3664 12100 3988 12158
tri 3988 12100 4076 12188 sw
tri 4086 12100 4174 12188 ne
rect 4174 12158 4488 12188
tri 4488 12158 4568 12238 sw
tri 4586 12158 4666 12238 ne
rect 4666 12188 4990 12238
tri 4990 12188 5088 12286 sw
tri 5088 12188 5186 12286 ne
rect 5186 12238 5500 12286
tri 5500 12238 5588 12326 sw
tri 5598 12238 5686 12326 ne
rect 5686 12290 5740 12326
rect 5860 12326 5962 12410
tri 5962 12326 6050 12414 sw
tri 6060 12326 6148 12414 ne
rect 6148 12410 6512 12414
rect 6148 12326 6290 12410
rect 5860 12290 6050 12326
rect 5686 12286 6050 12290
tri 6050 12286 6090 12326 sw
tri 6148 12286 6188 12326 ne
rect 6188 12290 6290 12326
rect 6410 12326 6512 12410
tri 6512 12326 6600 12414 sw
tri 6610 12326 6698 12414 ne
rect 6698 12410 7062 12414
rect 6698 12326 6840 12410
rect 6410 12290 6600 12326
rect 6188 12286 6600 12290
rect 5686 12238 6090 12286
rect 5186 12188 5588 12238
rect 4666 12158 5088 12188
rect 4174 12100 4568 12158
rect 3664 12060 4076 12100
tri 4076 12060 4116 12100 sw
tri 4174 12060 4214 12100 ne
rect 4214 12060 4568 12100
tri 4568 12060 4666 12158 sw
tri 4666 12060 4764 12158 ne
rect 4764 12100 5088 12158
tri 5088 12100 5176 12188 sw
tri 5186 12100 5274 12188 ne
rect 5274 12158 5588 12188
tri 5588 12158 5668 12238 sw
tri 5686 12158 5766 12238 ne
rect 5766 12188 6090 12238
tri 6090 12188 6188 12286 sw
tri 6188 12188 6286 12286 ne
rect 6286 12238 6600 12286
tri 6600 12238 6688 12326 sw
tri 6698 12238 6786 12326 ne
rect 6786 12290 6840 12326
rect 6960 12326 7062 12410
tri 7062 12326 7150 12414 sw
tri 7160 12326 7248 12414 ne
rect 7248 12410 7612 12414
rect 7248 12326 7390 12410
rect 6960 12290 7150 12326
rect 6786 12286 7150 12290
tri 7150 12286 7190 12326 sw
tri 7248 12286 7288 12326 ne
rect 7288 12290 7390 12326
rect 7510 12326 7612 12410
tri 7612 12326 7700 12414 sw
tri 7710 12326 7798 12414 ne
rect 7798 12410 8162 12414
rect 7798 12326 7940 12410
rect 7510 12290 7700 12326
rect 7288 12286 7700 12290
rect 6786 12238 7190 12286
rect 6286 12188 6688 12238
rect 5766 12158 6188 12188
rect 5274 12100 5668 12158
rect 4764 12060 5176 12100
tri 5176 12060 5216 12100 sw
tri 5274 12060 5314 12100 ne
rect 5314 12060 5668 12100
tri 5668 12060 5766 12158 sw
tri 5766 12060 5864 12158 ne
rect 5864 12100 6188 12158
tri 6188 12100 6276 12188 sw
tri 6286 12100 6374 12188 ne
rect 6374 12158 6688 12188
tri 6688 12158 6768 12238 sw
tri 6786 12158 6866 12238 ne
rect 6866 12188 7190 12238
tri 7190 12188 7288 12286 sw
tri 7288 12188 7386 12286 ne
rect 7386 12238 7700 12286
tri 7700 12238 7788 12326 sw
tri 7798 12238 7886 12326 ne
rect 7886 12290 7940 12326
rect 8060 12326 8162 12410
tri 8162 12326 8250 12414 sw
tri 8260 12326 8348 12414 ne
rect 8348 12410 8712 12414
rect 8348 12326 8490 12410
rect 8060 12290 8250 12326
rect 7886 12286 8250 12290
tri 8250 12286 8290 12326 sw
tri 8348 12286 8388 12326 ne
rect 8388 12290 8490 12326
rect 8610 12326 8712 12410
tri 8712 12326 8800 12414 sw
tri 8810 12326 8898 12414 ne
rect 8898 12410 9262 12414
rect 8898 12326 9040 12410
rect 8610 12290 8800 12326
rect 8388 12286 8800 12290
rect 7886 12238 8290 12286
rect 7386 12188 7788 12238
rect 6866 12158 7288 12188
rect 6374 12100 6768 12158
rect 5864 12060 6276 12100
tri 6276 12060 6316 12100 sw
tri 6374 12060 6414 12100 ne
rect 6414 12060 6768 12100
tri 6768 12060 6866 12158 sw
tri 6866 12060 6964 12158 ne
rect 6964 12100 7288 12158
tri 7288 12100 7376 12188 sw
tri 7386 12100 7474 12188 ne
rect 7474 12158 7788 12188
tri 7788 12158 7868 12238 sw
tri 7886 12158 7966 12238 ne
rect 7966 12188 8290 12238
tri 8290 12188 8388 12286 sw
tri 8388 12188 8486 12286 ne
rect 8486 12238 8800 12286
tri 8800 12238 8888 12326 sw
tri 8898 12238 8986 12326 ne
rect 8986 12290 9040 12326
rect 9160 12326 9262 12410
tri 9262 12326 9350 12414 sw
tri 9360 12326 9448 12414 ne
rect 9448 12410 9812 12414
rect 9448 12326 9590 12410
rect 9160 12290 9350 12326
rect 8986 12286 9350 12290
tri 9350 12286 9390 12326 sw
tri 9448 12286 9488 12326 ne
rect 9488 12290 9590 12326
rect 9710 12326 9812 12410
tri 9812 12326 9900 12414 sw
tri 9910 12326 9998 12414 ne
rect 9998 12410 10362 12414
rect 9998 12326 10140 12410
rect 9710 12290 9900 12326
rect 9488 12286 9900 12290
rect 8986 12238 9390 12286
rect 8486 12188 8888 12238
rect 7966 12158 8388 12188
rect 7474 12100 7868 12158
rect 6964 12060 7376 12100
tri 7376 12060 7416 12100 sw
tri 7474 12060 7514 12100 ne
rect 7514 12060 7868 12100
tri 7868 12060 7966 12158 sw
tri 7966 12060 8064 12158 ne
rect 8064 12100 8388 12158
tri 8388 12100 8476 12188 sw
tri 8486 12100 8574 12188 ne
rect 8574 12158 8888 12188
tri 8888 12158 8968 12238 sw
tri 8986 12158 9066 12238 ne
rect 9066 12188 9390 12238
tri 9390 12188 9488 12286 sw
tri 9488 12188 9586 12286 ne
rect 9586 12238 9900 12286
tri 9900 12238 9988 12326 sw
tri 9998 12238 10086 12326 ne
rect 10086 12290 10140 12326
rect 10260 12326 10362 12410
tri 10362 12326 10450 12414 sw
tri 10460 12326 10548 12414 ne
rect 10548 12410 10912 12414
rect 10548 12326 10690 12410
rect 10260 12290 10450 12326
rect 10086 12286 10450 12290
tri 10450 12286 10490 12326 sw
tri 10548 12286 10588 12326 ne
rect 10588 12290 10690 12326
rect 10810 12326 10912 12410
tri 10912 12326 11000 12414 sw
tri 11010 12326 11098 12414 ne
rect 11098 12410 11462 12414
rect 11098 12326 11240 12410
rect 10810 12290 11000 12326
rect 10588 12286 11000 12290
rect 10086 12238 10490 12286
rect 9586 12188 9988 12238
rect 9066 12158 9488 12188
rect 8574 12100 8968 12158
rect 8064 12060 8476 12100
tri 8476 12060 8516 12100 sw
tri 8574 12060 8614 12100 ne
rect 8614 12060 8968 12100
tri 8968 12060 9066 12158 sw
tri 9066 12060 9164 12158 ne
rect 9164 12100 9488 12158
tri 9488 12100 9576 12188 sw
tri 9586 12100 9674 12188 ne
rect 9674 12158 9988 12188
tri 9988 12158 10068 12238 sw
tri 10086 12158 10166 12238 ne
rect 10166 12188 10490 12238
tri 10490 12188 10588 12286 sw
tri 10588 12188 10686 12286 ne
rect 10686 12238 11000 12286
tri 11000 12238 11088 12326 sw
tri 11098 12238 11186 12326 ne
rect 11186 12290 11240 12326
rect 11360 12326 11462 12410
tri 11462 12326 11550 12414 sw
tri 11560 12326 11648 12414 ne
rect 11648 12410 12012 12414
rect 11648 12326 11790 12410
rect 11360 12290 11550 12326
rect 11186 12286 11550 12290
tri 11550 12286 11590 12326 sw
tri 11648 12286 11688 12326 ne
rect 11688 12290 11790 12326
rect 11910 12326 12012 12410
tri 12012 12326 12100 12414 sw
tri 12110 12326 12198 12414 ne
rect 12198 12410 12562 12414
rect 12198 12326 12340 12410
rect 11910 12290 12100 12326
rect 11688 12286 12100 12290
rect 11186 12238 11590 12286
rect 10686 12188 11088 12238
rect 10166 12158 10588 12188
rect 9674 12100 10068 12158
rect 9164 12060 9576 12100
tri 9576 12060 9616 12100 sw
tri 9674 12060 9714 12100 ne
rect 9714 12060 10068 12100
tri 10068 12060 10166 12158 sw
tri 10166 12060 10264 12158 ne
rect 10264 12100 10588 12158
tri 10588 12100 10676 12188 sw
tri 10686 12100 10774 12188 ne
rect 10774 12158 11088 12188
tri 11088 12158 11168 12238 sw
tri 11186 12158 11266 12238 ne
rect 11266 12188 11590 12238
tri 11590 12188 11688 12286 sw
tri 11688 12188 11786 12286 ne
rect 11786 12238 12100 12286
tri 12100 12238 12188 12326 sw
tri 12198 12238 12286 12326 ne
rect 12286 12290 12340 12326
rect 12460 12326 12562 12410
tri 12562 12326 12650 12414 sw
tri 12660 12326 12748 12414 ne
rect 12748 12410 13112 12414
rect 12748 12326 12890 12410
rect 12460 12290 12650 12326
rect 12286 12286 12650 12290
tri 12650 12286 12690 12326 sw
tri 12748 12286 12788 12326 ne
rect 12788 12290 12890 12326
rect 13010 12326 13112 12410
tri 13112 12326 13200 12414 sw
tri 13210 12326 13298 12414 ne
rect 13298 12410 15775 12414
rect 13298 12326 13440 12410
rect 13010 12290 13200 12326
rect 12788 12286 13200 12290
rect 12286 12238 12690 12286
rect 11786 12188 12188 12238
rect 11266 12158 11688 12188
rect 10774 12100 11168 12158
rect 10264 12060 10676 12100
tri 10676 12060 10716 12100 sw
tri 10774 12060 10814 12100 ne
rect 10814 12060 11168 12100
tri 11168 12060 11266 12158 sw
tri 11266 12060 11364 12158 ne
rect 11364 12100 11688 12158
tri 11688 12100 11776 12188 sw
tri 11786 12100 11874 12188 ne
rect 11874 12158 12188 12188
tri 12188 12158 12268 12238 sw
tri 12286 12158 12366 12238 ne
rect 12366 12188 12690 12238
tri 12690 12188 12788 12286 sw
tri 12788 12188 12886 12286 ne
rect 12886 12238 13200 12286
tri 13200 12238 13288 12326 sw
tri 13298 12238 13386 12326 ne
rect 13386 12290 13440 12326
rect 13560 12290 15775 12410
rect 13386 12238 15775 12290
rect 12886 12188 13288 12238
rect 12366 12158 12788 12188
rect 11874 12100 12268 12158
rect 11364 12060 11776 12100
tri 11776 12060 11816 12100 sw
tri 11874 12060 11914 12100 ne
rect 11914 12060 12268 12100
tri 12268 12060 12366 12158 sw
tri 12366 12060 12464 12158 ne
rect 12464 12100 12788 12158
tri 12788 12100 12876 12188 sw
tri 12886 12100 12974 12188 ne
rect 12974 12158 13288 12188
tri 13288 12158 13368 12238 sw
tri 13386 12158 13466 12238 ne
rect 13466 12158 14075 12238
rect 12974 12100 13368 12158
rect 12464 12060 12876 12100
tri 12876 12060 12916 12100 sw
tri 12974 12060 13014 12100 ne
rect 13014 12060 13368 12100
tri 13368 12060 13466 12158 sw
tri 13466 12060 13564 12158 ne
rect 13564 12138 14075 12158
rect 14175 12138 15775 12238
rect 13564 12060 15775 12138
rect -1025 12012 -284 12060
rect -1025 11912 -925 12012
rect -825 11962 -284 12012
tri -284 11962 -186 12060 sw
tri -186 11962 -88 12060 ne
rect -88 11962 266 12060
tri 266 11962 364 12060 sw
tri 364 11962 462 12060 ne
rect 462 11962 816 12060
tri 816 11962 914 12060 sw
tri 914 11962 1012 12060 ne
rect 1012 11962 1366 12060
tri 1366 11962 1464 12060 sw
tri 1464 11962 1562 12060 ne
rect 1562 11962 1916 12060
tri 1916 11962 2014 12060 sw
tri 2014 11962 2112 12060 ne
rect 2112 11962 2466 12060
tri 2466 11962 2564 12060 sw
tri 2564 11962 2662 12060 ne
rect 2662 11962 3016 12060
tri 3016 11962 3114 12060 sw
tri 3114 11962 3212 12060 ne
rect 3212 11962 3566 12060
tri 3566 11962 3664 12060 sw
tri 3664 11962 3762 12060 ne
rect 3762 11962 4116 12060
tri 4116 11962 4214 12060 sw
tri 4214 11962 4312 12060 ne
rect 4312 11962 4666 12060
tri 4666 11962 4764 12060 sw
tri 4764 11962 4862 12060 ne
rect 4862 11962 5216 12060
tri 5216 11962 5314 12060 sw
tri 5314 11962 5412 12060 ne
rect 5412 11962 5766 12060
tri 5766 11962 5864 12060 sw
tri 5864 11962 5962 12060 ne
rect 5962 11962 6316 12060
tri 6316 11962 6414 12060 sw
tri 6414 11962 6512 12060 ne
rect 6512 11962 6866 12060
tri 6866 11962 6964 12060 sw
tri 6964 11962 7062 12060 ne
rect 7062 11962 7416 12060
tri 7416 11962 7514 12060 sw
tri 7514 11962 7612 12060 ne
rect 7612 11962 7966 12060
tri 7966 11962 8064 12060 sw
tri 8064 11962 8162 12060 ne
rect 8162 11962 8516 12060
tri 8516 11962 8614 12060 sw
tri 8614 11962 8712 12060 ne
rect 8712 11962 9066 12060
tri 9066 11962 9164 12060 sw
tri 9164 11962 9262 12060 ne
rect 9262 11962 9616 12060
tri 9616 11962 9714 12060 sw
tri 9714 11962 9812 12060 ne
rect 9812 11962 10166 12060
tri 10166 11962 10264 12060 sw
tri 10264 11962 10362 12060 ne
rect 10362 11962 10716 12060
tri 10716 11962 10814 12060 sw
tri 10814 11962 10912 12060 ne
rect 10912 11962 11266 12060
tri 11266 11962 11364 12060 sw
tri 11364 11962 11462 12060 ne
rect 11462 11962 11816 12060
tri 11816 11962 11914 12060 sw
tri 11914 11962 12012 12060 ne
rect 12012 11962 12366 12060
tri 12366 11962 12464 12060 sw
tri 12464 11962 12562 12060 ne
rect 12562 11962 12916 12060
tri 12916 11962 13014 12060 sw
tri 13014 11962 13112 12060 ne
rect 13112 11962 13466 12060
tri 13466 11962 13564 12060 sw
tri 13564 11962 13662 12060 ne
rect 13662 11962 15775 12060
rect -825 11912 -186 11962
rect -1025 11864 -186 11912
tri -186 11864 -88 11962 sw
tri -88 11864 10 11962 ne
rect 10 11864 364 11962
tri 364 11864 462 11962 sw
tri 462 11864 560 11962 ne
rect 560 11864 914 11962
tri 914 11864 1012 11962 sw
tri 1012 11864 1110 11962 ne
rect 1110 11864 1464 11962
tri 1464 11864 1562 11962 sw
tri 1562 11864 1660 11962 ne
rect 1660 11864 2014 11962
tri 2014 11864 2112 11962 sw
tri 2112 11864 2210 11962 ne
rect 2210 11864 2564 11962
tri 2564 11864 2662 11962 sw
tri 2662 11864 2760 11962 ne
rect 2760 11864 3114 11962
tri 3114 11864 3212 11962 sw
tri 3212 11864 3310 11962 ne
rect 3310 11864 3664 11962
tri 3664 11864 3762 11962 sw
tri 3762 11864 3860 11962 ne
rect 3860 11864 4214 11962
tri 4214 11864 4312 11962 sw
tri 4312 11864 4410 11962 ne
rect 4410 11864 4764 11962
tri 4764 11864 4862 11962 sw
tri 4862 11864 4960 11962 ne
rect 4960 11864 5314 11962
tri 5314 11864 5412 11962 sw
tri 5412 11864 5510 11962 ne
rect 5510 11864 5864 11962
tri 5864 11864 5962 11962 sw
tri 5962 11864 6060 11962 ne
rect 6060 11864 6414 11962
tri 6414 11864 6512 11962 sw
tri 6512 11864 6610 11962 ne
rect 6610 11864 6964 11962
tri 6964 11864 7062 11962 sw
tri 7062 11864 7160 11962 ne
rect 7160 11864 7514 11962
tri 7514 11864 7612 11962 sw
tri 7612 11864 7710 11962 ne
rect 7710 11864 8064 11962
tri 8064 11864 8162 11962 sw
tri 8162 11864 8260 11962 ne
rect 8260 11864 8614 11962
tri 8614 11864 8712 11962 sw
tri 8712 11864 8810 11962 ne
rect 8810 11864 9164 11962
tri 9164 11864 9262 11962 sw
tri 9262 11864 9360 11962 ne
rect 9360 11864 9714 11962
tri 9714 11864 9812 11962 sw
tri 9812 11864 9910 11962 ne
rect 9910 11864 10264 11962
tri 10264 11864 10362 11962 sw
tri 10362 11864 10460 11962 ne
rect 10460 11864 10814 11962
tri 10814 11864 10912 11962 sw
tri 10912 11864 11010 11962 ne
rect 11010 11864 11364 11962
tri 11364 11864 11462 11962 sw
tri 11462 11864 11560 11962 ne
rect 11560 11864 11914 11962
tri 11914 11864 12012 11962 sw
tri 12012 11864 12110 11962 ne
rect 12110 11864 12464 11962
tri 12464 11864 12562 11962 sw
tri 12562 11864 12660 11962 ne
rect 12660 11864 13014 11962
tri 13014 11864 13112 11962 sw
tri 13112 11864 13210 11962 ne
rect 13210 11864 13564 11962
tri 13564 11864 13662 11962 sw
rect -1025 11860 -88 11864
rect -1025 11740 -310 11860
rect -190 11776 -88 11860
tri -88 11776 0 11864 sw
tri 10 11776 98 11864 ne
rect 98 11860 462 11864
rect 98 11776 240 11860
rect -190 11740 0 11776
rect -1025 11736 0 11740
tri 0 11736 40 11776 sw
tri 98 11736 138 11776 ne
rect 138 11740 240 11776
rect 360 11776 462 11860
tri 462 11776 550 11864 sw
tri 560 11776 648 11864 ne
rect 648 11860 1012 11864
rect 648 11776 790 11860
rect 360 11740 550 11776
rect 138 11736 550 11740
tri -412 11638 -314 11736 ne
rect -314 11638 40 11736
tri 40 11638 138 11736 sw
tri 138 11638 236 11736 ne
rect 236 11688 550 11736
tri 550 11688 638 11776 sw
tri 648 11688 736 11776 ne
rect 736 11740 790 11776
rect 910 11776 1012 11860
tri 1012 11776 1100 11864 sw
tri 1110 11776 1198 11864 ne
rect 1198 11860 1562 11864
rect 1198 11776 1340 11860
rect 910 11740 1100 11776
rect 736 11736 1100 11740
tri 1100 11736 1140 11776 sw
tri 1198 11736 1238 11776 ne
rect 1238 11740 1340 11776
rect 1460 11776 1562 11860
tri 1562 11776 1650 11864 sw
tri 1660 11776 1748 11864 ne
rect 1748 11860 2112 11864
rect 1748 11776 1890 11860
rect 1460 11740 1650 11776
rect 1238 11736 1650 11740
rect 736 11688 1140 11736
rect 236 11638 638 11688
rect -2525 11550 -412 11638
tri -412 11550 -324 11638 sw
tri -314 11550 -226 11638 ne
rect -226 11550 138 11638
tri 138 11550 226 11638 sw
tri 236 11550 324 11638 ne
rect 324 11608 638 11638
tri 638 11608 718 11688 sw
tri 736 11608 816 11688 ne
rect 816 11638 1140 11688
tri 1140 11638 1238 11736 sw
tri 1238 11638 1336 11736 ne
rect 1336 11688 1650 11736
tri 1650 11688 1738 11776 sw
tri 1748 11688 1836 11776 ne
rect 1836 11740 1890 11776
rect 2010 11776 2112 11860
tri 2112 11776 2200 11864 sw
tri 2210 11776 2298 11864 ne
rect 2298 11860 2662 11864
rect 2298 11776 2440 11860
rect 2010 11740 2200 11776
rect 1836 11736 2200 11740
tri 2200 11736 2240 11776 sw
tri 2298 11736 2338 11776 ne
rect 2338 11740 2440 11776
rect 2560 11776 2662 11860
tri 2662 11776 2750 11864 sw
tri 2760 11776 2848 11864 ne
rect 2848 11860 3212 11864
rect 2848 11776 2990 11860
rect 2560 11740 2750 11776
rect 2338 11736 2750 11740
rect 1836 11688 2240 11736
rect 1336 11638 1738 11688
rect 816 11608 1238 11638
rect 324 11550 718 11608
rect -2525 11510 -324 11550
tri -324 11510 -284 11550 sw
tri -226 11510 -186 11550 ne
rect -186 11510 226 11550
tri 226 11510 266 11550 sw
tri 324 11510 364 11550 ne
rect 364 11510 718 11550
tri 718 11510 816 11608 sw
tri 816 11510 914 11608 ne
rect 914 11550 1238 11608
tri 1238 11550 1326 11638 sw
tri 1336 11550 1424 11638 ne
rect 1424 11608 1738 11638
tri 1738 11608 1818 11688 sw
tri 1836 11608 1916 11688 ne
rect 1916 11638 2240 11688
tri 2240 11638 2338 11736 sw
tri 2338 11638 2436 11736 ne
rect 2436 11688 2750 11736
tri 2750 11688 2838 11776 sw
tri 2848 11688 2936 11776 ne
rect 2936 11740 2990 11776
rect 3110 11776 3212 11860
tri 3212 11776 3300 11864 sw
tri 3310 11776 3398 11864 ne
rect 3398 11860 3762 11864
rect 3398 11776 3540 11860
rect 3110 11740 3300 11776
rect 2936 11736 3300 11740
tri 3300 11736 3340 11776 sw
tri 3398 11736 3438 11776 ne
rect 3438 11740 3540 11776
rect 3660 11776 3762 11860
tri 3762 11776 3850 11864 sw
tri 3860 11776 3948 11864 ne
rect 3948 11860 4312 11864
rect 3948 11776 4090 11860
rect 3660 11740 3850 11776
rect 3438 11736 3850 11740
rect 2936 11688 3340 11736
rect 2436 11638 2838 11688
rect 1916 11608 2338 11638
rect 1424 11550 1818 11608
rect 914 11510 1326 11550
tri 1326 11510 1366 11550 sw
tri 1424 11510 1464 11550 ne
rect 1464 11510 1818 11550
tri 1818 11510 1916 11608 sw
tri 1916 11510 2014 11608 ne
rect 2014 11550 2338 11608
tri 2338 11550 2426 11638 sw
tri 2436 11550 2524 11638 ne
rect 2524 11608 2838 11638
tri 2838 11608 2918 11688 sw
tri 2936 11608 3016 11688 ne
rect 3016 11638 3340 11688
tri 3340 11638 3438 11736 sw
tri 3438 11638 3536 11736 ne
rect 3536 11688 3850 11736
tri 3850 11688 3938 11776 sw
tri 3948 11688 4036 11776 ne
rect 4036 11740 4090 11776
rect 4210 11776 4312 11860
tri 4312 11776 4400 11864 sw
tri 4410 11776 4498 11864 ne
rect 4498 11860 4862 11864
rect 4498 11776 4640 11860
rect 4210 11740 4400 11776
rect 4036 11736 4400 11740
tri 4400 11736 4440 11776 sw
tri 4498 11736 4538 11776 ne
rect 4538 11740 4640 11776
rect 4760 11776 4862 11860
tri 4862 11776 4950 11864 sw
tri 4960 11776 5048 11864 ne
rect 5048 11860 5412 11864
rect 5048 11776 5190 11860
rect 4760 11740 4950 11776
rect 4538 11736 4950 11740
rect 4036 11688 4440 11736
rect 3536 11638 3938 11688
rect 3016 11608 3438 11638
rect 2524 11550 2918 11608
rect 2014 11510 2426 11550
tri 2426 11510 2466 11550 sw
tri 2524 11510 2564 11550 ne
rect 2564 11510 2918 11550
tri 2918 11510 3016 11608 sw
tri 3016 11510 3114 11608 ne
rect 3114 11550 3438 11608
tri 3438 11550 3526 11638 sw
tri 3536 11550 3624 11638 ne
rect 3624 11608 3938 11638
tri 3938 11608 4018 11688 sw
tri 4036 11608 4116 11688 ne
rect 4116 11638 4440 11688
tri 4440 11638 4538 11736 sw
tri 4538 11638 4636 11736 ne
rect 4636 11688 4950 11736
tri 4950 11688 5038 11776 sw
tri 5048 11688 5136 11776 ne
rect 5136 11740 5190 11776
rect 5310 11776 5412 11860
tri 5412 11776 5500 11864 sw
tri 5510 11776 5598 11864 ne
rect 5598 11860 5962 11864
rect 5598 11776 5740 11860
rect 5310 11740 5500 11776
rect 5136 11736 5500 11740
tri 5500 11736 5540 11776 sw
tri 5598 11736 5638 11776 ne
rect 5638 11740 5740 11776
rect 5860 11776 5962 11860
tri 5962 11776 6050 11864 sw
tri 6060 11776 6148 11864 ne
rect 6148 11860 6512 11864
rect 6148 11776 6290 11860
rect 5860 11740 6050 11776
rect 5638 11736 6050 11740
rect 5136 11688 5540 11736
rect 4636 11638 5038 11688
rect 4116 11608 4538 11638
rect 3624 11550 4018 11608
rect 3114 11510 3526 11550
tri 3526 11510 3566 11550 sw
tri 3624 11510 3664 11550 ne
rect 3664 11510 4018 11550
tri 4018 11510 4116 11608 sw
tri 4116 11510 4214 11608 ne
rect 4214 11550 4538 11608
tri 4538 11550 4626 11638 sw
tri 4636 11550 4724 11638 ne
rect 4724 11608 5038 11638
tri 5038 11608 5118 11688 sw
tri 5136 11608 5216 11688 ne
rect 5216 11638 5540 11688
tri 5540 11638 5638 11736 sw
tri 5638 11638 5736 11736 ne
rect 5736 11688 6050 11736
tri 6050 11688 6138 11776 sw
tri 6148 11688 6236 11776 ne
rect 6236 11740 6290 11776
rect 6410 11776 6512 11860
tri 6512 11776 6600 11864 sw
tri 6610 11776 6698 11864 ne
rect 6698 11860 7062 11864
rect 6698 11776 6840 11860
rect 6410 11740 6600 11776
rect 6236 11736 6600 11740
tri 6600 11736 6640 11776 sw
tri 6698 11736 6738 11776 ne
rect 6738 11740 6840 11776
rect 6960 11776 7062 11860
tri 7062 11776 7150 11864 sw
tri 7160 11776 7248 11864 ne
rect 7248 11860 7612 11864
rect 7248 11776 7390 11860
rect 6960 11740 7150 11776
rect 6738 11736 7150 11740
rect 6236 11688 6640 11736
rect 5736 11638 6138 11688
rect 5216 11608 5638 11638
rect 4724 11550 5118 11608
rect 4214 11510 4626 11550
tri 4626 11510 4666 11550 sw
tri 4724 11510 4764 11550 ne
rect 4764 11510 5118 11550
tri 5118 11510 5216 11608 sw
tri 5216 11510 5314 11608 ne
rect 5314 11550 5638 11608
tri 5638 11550 5726 11638 sw
tri 5736 11550 5824 11638 ne
rect 5824 11608 6138 11638
tri 6138 11608 6218 11688 sw
tri 6236 11608 6316 11688 ne
rect 6316 11638 6640 11688
tri 6640 11638 6738 11736 sw
tri 6738 11638 6836 11736 ne
rect 6836 11688 7150 11736
tri 7150 11688 7238 11776 sw
tri 7248 11688 7336 11776 ne
rect 7336 11740 7390 11776
rect 7510 11776 7612 11860
tri 7612 11776 7700 11864 sw
tri 7710 11776 7798 11864 ne
rect 7798 11860 8162 11864
rect 7798 11776 7940 11860
rect 7510 11740 7700 11776
rect 7336 11736 7700 11740
tri 7700 11736 7740 11776 sw
tri 7798 11736 7838 11776 ne
rect 7838 11740 7940 11776
rect 8060 11776 8162 11860
tri 8162 11776 8250 11864 sw
tri 8260 11776 8348 11864 ne
rect 8348 11860 8712 11864
rect 8348 11776 8490 11860
rect 8060 11740 8250 11776
rect 7838 11736 8250 11740
rect 7336 11688 7740 11736
rect 6836 11638 7238 11688
rect 6316 11608 6738 11638
rect 5824 11550 6218 11608
rect 5314 11510 5726 11550
tri 5726 11510 5766 11550 sw
tri 5824 11510 5864 11550 ne
rect 5864 11510 6218 11550
tri 6218 11510 6316 11608 sw
tri 6316 11510 6414 11608 ne
rect 6414 11550 6738 11608
tri 6738 11550 6826 11638 sw
tri 6836 11550 6924 11638 ne
rect 6924 11608 7238 11638
tri 7238 11608 7318 11688 sw
tri 7336 11608 7416 11688 ne
rect 7416 11638 7740 11688
tri 7740 11638 7838 11736 sw
tri 7838 11638 7936 11736 ne
rect 7936 11688 8250 11736
tri 8250 11688 8338 11776 sw
tri 8348 11688 8436 11776 ne
rect 8436 11740 8490 11776
rect 8610 11776 8712 11860
tri 8712 11776 8800 11864 sw
tri 8810 11776 8898 11864 ne
rect 8898 11860 9262 11864
rect 8898 11776 9040 11860
rect 8610 11740 8800 11776
rect 8436 11736 8800 11740
tri 8800 11736 8840 11776 sw
tri 8898 11736 8938 11776 ne
rect 8938 11740 9040 11776
rect 9160 11776 9262 11860
tri 9262 11776 9350 11864 sw
tri 9360 11776 9448 11864 ne
rect 9448 11860 9812 11864
rect 9448 11776 9590 11860
rect 9160 11740 9350 11776
rect 8938 11736 9350 11740
rect 8436 11688 8840 11736
rect 7936 11638 8338 11688
rect 7416 11608 7838 11638
rect 6924 11550 7318 11608
rect 6414 11510 6826 11550
tri 6826 11510 6866 11550 sw
tri 6924 11510 6964 11550 ne
rect 6964 11510 7318 11550
tri 7318 11510 7416 11608 sw
tri 7416 11510 7514 11608 ne
rect 7514 11550 7838 11608
tri 7838 11550 7926 11638 sw
tri 7936 11550 8024 11638 ne
rect 8024 11608 8338 11638
tri 8338 11608 8418 11688 sw
tri 8436 11608 8516 11688 ne
rect 8516 11638 8840 11688
tri 8840 11638 8938 11736 sw
tri 8938 11638 9036 11736 ne
rect 9036 11688 9350 11736
tri 9350 11688 9438 11776 sw
tri 9448 11688 9536 11776 ne
rect 9536 11740 9590 11776
rect 9710 11776 9812 11860
tri 9812 11776 9900 11864 sw
tri 9910 11776 9998 11864 ne
rect 9998 11860 10362 11864
rect 9998 11776 10140 11860
rect 9710 11740 9900 11776
rect 9536 11736 9900 11740
tri 9900 11736 9940 11776 sw
tri 9998 11736 10038 11776 ne
rect 10038 11740 10140 11776
rect 10260 11776 10362 11860
tri 10362 11776 10450 11864 sw
tri 10460 11776 10548 11864 ne
rect 10548 11860 10912 11864
rect 10548 11776 10690 11860
rect 10260 11740 10450 11776
rect 10038 11736 10450 11740
rect 9536 11688 9940 11736
rect 9036 11638 9438 11688
rect 8516 11608 8938 11638
rect 8024 11550 8418 11608
rect 7514 11510 7926 11550
tri 7926 11510 7966 11550 sw
tri 8024 11510 8064 11550 ne
rect 8064 11510 8418 11550
tri 8418 11510 8516 11608 sw
tri 8516 11510 8614 11608 ne
rect 8614 11550 8938 11608
tri 8938 11550 9026 11638 sw
tri 9036 11550 9124 11638 ne
rect 9124 11608 9438 11638
tri 9438 11608 9518 11688 sw
tri 9536 11608 9616 11688 ne
rect 9616 11638 9940 11688
tri 9940 11638 10038 11736 sw
tri 10038 11638 10136 11736 ne
rect 10136 11688 10450 11736
tri 10450 11688 10538 11776 sw
tri 10548 11688 10636 11776 ne
rect 10636 11740 10690 11776
rect 10810 11776 10912 11860
tri 10912 11776 11000 11864 sw
tri 11010 11776 11098 11864 ne
rect 11098 11860 11462 11864
rect 11098 11776 11240 11860
rect 10810 11740 11000 11776
rect 10636 11736 11000 11740
tri 11000 11736 11040 11776 sw
tri 11098 11736 11138 11776 ne
rect 11138 11740 11240 11776
rect 11360 11776 11462 11860
tri 11462 11776 11550 11864 sw
tri 11560 11776 11648 11864 ne
rect 11648 11860 12012 11864
rect 11648 11776 11790 11860
rect 11360 11740 11550 11776
rect 11138 11736 11550 11740
rect 10636 11688 11040 11736
rect 10136 11638 10538 11688
rect 9616 11608 10038 11638
rect 9124 11550 9518 11608
rect 8614 11510 9026 11550
tri 9026 11510 9066 11550 sw
tri 9124 11510 9164 11550 ne
rect 9164 11510 9518 11550
tri 9518 11510 9616 11608 sw
tri 9616 11510 9714 11608 ne
rect 9714 11550 10038 11608
tri 10038 11550 10126 11638 sw
tri 10136 11550 10224 11638 ne
rect 10224 11608 10538 11638
tri 10538 11608 10618 11688 sw
tri 10636 11608 10716 11688 ne
rect 10716 11638 11040 11688
tri 11040 11638 11138 11736 sw
tri 11138 11638 11236 11736 ne
rect 11236 11688 11550 11736
tri 11550 11688 11638 11776 sw
tri 11648 11688 11736 11776 ne
rect 11736 11740 11790 11776
rect 11910 11776 12012 11860
tri 12012 11776 12100 11864 sw
tri 12110 11776 12198 11864 ne
rect 12198 11860 12562 11864
rect 12198 11776 12340 11860
rect 11910 11740 12100 11776
rect 11736 11736 12100 11740
tri 12100 11736 12140 11776 sw
tri 12198 11736 12238 11776 ne
rect 12238 11740 12340 11776
rect 12460 11776 12562 11860
tri 12562 11776 12650 11864 sw
tri 12660 11776 12748 11864 ne
rect 12748 11860 13112 11864
rect 12748 11776 12890 11860
rect 12460 11740 12650 11776
rect 12238 11736 12650 11740
rect 11736 11688 12140 11736
rect 11236 11638 11638 11688
rect 10716 11608 11138 11638
rect 10224 11550 10618 11608
rect 9714 11510 10126 11550
tri 10126 11510 10166 11550 sw
tri 10224 11510 10264 11550 ne
rect 10264 11510 10618 11550
tri 10618 11510 10716 11608 sw
tri 10716 11510 10814 11608 ne
rect 10814 11550 11138 11608
tri 11138 11550 11226 11638 sw
tri 11236 11550 11324 11638 ne
rect 11324 11608 11638 11638
tri 11638 11608 11718 11688 sw
tri 11736 11608 11816 11688 ne
rect 11816 11638 12140 11688
tri 12140 11638 12238 11736 sw
tri 12238 11638 12336 11736 ne
rect 12336 11688 12650 11736
tri 12650 11688 12738 11776 sw
tri 12748 11688 12836 11776 ne
rect 12836 11740 12890 11776
rect 13010 11776 13112 11860
tri 13112 11776 13200 11864 sw
tri 13210 11776 13298 11864 ne
rect 13298 11860 14275 11864
rect 13298 11776 13440 11860
rect 13010 11740 13200 11776
rect 12836 11736 13200 11740
tri 13200 11736 13240 11776 sw
tri 13298 11736 13338 11776 ne
rect 13338 11740 13440 11776
rect 13560 11740 14275 11860
rect 13338 11736 14275 11740
rect 12836 11688 13240 11736
rect 12336 11638 12738 11688
rect 11816 11608 12238 11638
rect 11324 11550 11718 11608
rect 10814 11510 11226 11550
tri 11226 11510 11266 11550 sw
tri 11324 11510 11364 11550 ne
rect 11364 11510 11718 11550
tri 11718 11510 11816 11608 sw
tri 11816 11510 11914 11608 ne
rect 11914 11550 12238 11608
tri 12238 11550 12326 11638 sw
tri 12336 11550 12424 11638 ne
rect 12424 11608 12738 11638
tri 12738 11608 12818 11688 sw
tri 12836 11608 12916 11688 ne
rect 12916 11638 13240 11688
tri 13240 11638 13338 11736 sw
tri 13338 11638 13436 11736 ne
rect 13436 11638 14275 11736
rect 12916 11608 13338 11638
rect 12424 11550 12818 11608
rect 11914 11510 12326 11550
tri 12326 11510 12366 11550 sw
tri 12424 11510 12464 11550 ne
rect 12464 11510 12818 11550
tri 12818 11510 12916 11608 sw
tri 12916 11510 13014 11608 ne
rect 13014 11550 13338 11608
tri 13338 11550 13426 11638 sw
tri 13436 11550 13524 11638 ne
rect 13524 11550 14275 11638
rect 13014 11510 13426 11550
tri 13426 11510 13466 11550 sw
tri 13524 11510 13564 11550 ne
rect 13564 11510 14275 11550
rect -2525 11412 -284 11510
tri -284 11412 -186 11510 sw
tri -186 11412 -88 11510 ne
rect -88 11412 266 11510
tri 266 11412 364 11510 sw
tri 364 11412 462 11510 ne
rect 462 11412 816 11510
tri 816 11412 914 11510 sw
tri 914 11412 1012 11510 ne
rect 1012 11412 1366 11510
tri 1366 11412 1464 11510 sw
tri 1464 11412 1562 11510 ne
rect 1562 11412 1916 11510
tri 1916 11412 2014 11510 sw
tri 2014 11412 2112 11510 ne
rect 2112 11412 2466 11510
tri 2466 11412 2564 11510 sw
tri 2564 11412 2662 11510 ne
rect 2662 11412 3016 11510
tri 3016 11412 3114 11510 sw
tri 3114 11412 3212 11510 ne
rect 3212 11412 3566 11510
tri 3566 11412 3664 11510 sw
tri 3664 11412 3762 11510 ne
rect 3762 11412 4116 11510
tri 4116 11412 4214 11510 sw
tri 4214 11412 4312 11510 ne
rect 4312 11412 4666 11510
tri 4666 11412 4764 11510 sw
tri 4764 11412 4862 11510 ne
rect 4862 11412 5216 11510
tri 5216 11412 5314 11510 sw
tri 5314 11412 5412 11510 ne
rect 5412 11412 5766 11510
tri 5766 11412 5864 11510 sw
tri 5864 11412 5962 11510 ne
rect 5962 11412 6316 11510
tri 6316 11412 6414 11510 sw
tri 6414 11412 6512 11510 ne
rect 6512 11412 6866 11510
tri 6866 11412 6964 11510 sw
tri 6964 11412 7062 11510 ne
rect 7062 11412 7416 11510
tri 7416 11412 7514 11510 sw
tri 7514 11412 7612 11510 ne
rect 7612 11412 7966 11510
tri 7966 11412 8064 11510 sw
tri 8064 11412 8162 11510 ne
rect 8162 11412 8516 11510
tri 8516 11412 8614 11510 sw
tri 8614 11412 8712 11510 ne
rect 8712 11412 9066 11510
tri 9066 11412 9164 11510 sw
tri 9164 11412 9262 11510 ne
rect 9262 11412 9616 11510
tri 9616 11412 9714 11510 sw
tri 9714 11412 9812 11510 ne
rect 9812 11412 10166 11510
tri 10166 11412 10264 11510 sw
tri 10264 11412 10362 11510 ne
rect 10362 11412 10716 11510
tri 10716 11412 10814 11510 sw
tri 10814 11412 10912 11510 ne
rect 10912 11412 11266 11510
tri 11266 11412 11364 11510 sw
tri 11364 11412 11462 11510 ne
rect 11462 11412 11816 11510
tri 11816 11412 11914 11510 sw
tri 11914 11412 12012 11510 ne
rect 12012 11412 12366 11510
tri 12366 11412 12464 11510 sw
tri 12464 11412 12562 11510 ne
rect 12562 11412 12916 11510
tri 12916 11412 13014 11510 sw
tri 13014 11412 13112 11510 ne
rect 13112 11412 13466 11510
tri 13466 11412 13564 11510 sw
tri 13564 11412 13662 11510 ne
rect 13662 11412 14275 11510
rect -2525 11314 -186 11412
tri -186 11314 -88 11412 sw
tri -88 11314 10 11412 ne
rect 10 11314 364 11412
tri 364 11314 462 11412 sw
tri 462 11314 560 11412 ne
rect 560 11314 914 11412
tri 914 11314 1012 11412 sw
tri 1012 11314 1110 11412 ne
rect 1110 11314 1464 11412
tri 1464 11314 1562 11412 sw
tri 1562 11314 1660 11412 ne
rect 1660 11314 2014 11412
tri 2014 11314 2112 11412 sw
tri 2112 11314 2210 11412 ne
rect 2210 11314 2564 11412
tri 2564 11314 2662 11412 sw
tri 2662 11314 2760 11412 ne
rect 2760 11314 3114 11412
tri 3114 11314 3212 11412 sw
tri 3212 11314 3310 11412 ne
rect 3310 11314 3664 11412
tri 3664 11314 3762 11412 sw
tri 3762 11314 3860 11412 ne
rect 3860 11314 4214 11412
tri 4214 11314 4312 11412 sw
tri 4312 11314 4410 11412 ne
rect 4410 11314 4764 11412
tri 4764 11314 4862 11412 sw
tri 4862 11314 4960 11412 ne
rect 4960 11314 5314 11412
tri 5314 11314 5412 11412 sw
tri 5412 11314 5510 11412 ne
rect 5510 11314 5864 11412
tri 5864 11314 5962 11412 sw
tri 5962 11314 6060 11412 ne
rect 6060 11314 6414 11412
tri 6414 11314 6512 11412 sw
tri 6512 11314 6610 11412 ne
rect 6610 11314 6964 11412
tri 6964 11314 7062 11412 sw
tri 7062 11314 7160 11412 ne
rect 7160 11314 7514 11412
tri 7514 11314 7612 11412 sw
tri 7612 11314 7710 11412 ne
rect 7710 11314 8064 11412
tri 8064 11314 8162 11412 sw
tri 8162 11314 8260 11412 ne
rect 8260 11314 8614 11412
tri 8614 11314 8712 11412 sw
tri 8712 11314 8810 11412 ne
rect 8810 11314 9164 11412
tri 9164 11314 9262 11412 sw
tri 9262 11314 9360 11412 ne
rect 9360 11314 9714 11412
tri 9714 11314 9812 11412 sw
tri 9812 11314 9910 11412 ne
rect 9910 11314 10264 11412
tri 10264 11314 10362 11412 sw
tri 10362 11314 10460 11412 ne
rect 10460 11314 10814 11412
tri 10814 11314 10912 11412 sw
tri 10912 11314 11010 11412 ne
rect 11010 11314 11364 11412
tri 11364 11314 11462 11412 sw
tri 11462 11314 11560 11412 ne
rect 11560 11314 11914 11412
tri 11914 11314 12012 11412 sw
tri 12012 11314 12110 11412 ne
rect 12110 11314 12464 11412
tri 12464 11314 12562 11412 sw
tri 12562 11314 12660 11412 ne
rect 12660 11314 13014 11412
tri 13014 11314 13112 11412 sw
tri 13112 11314 13210 11412 ne
rect 13210 11314 13564 11412
tri 13564 11314 13662 11412 sw
rect 14775 11314 15775 11962
rect -2525 11310 -88 11314
rect -2525 11190 -310 11310
rect -190 11226 -88 11310
tri -88 11226 0 11314 sw
tri 10 11226 98 11314 ne
rect 98 11310 462 11314
rect 98 11226 240 11310
rect -190 11190 0 11226
rect -2525 11186 0 11190
rect -2525 10538 -1525 11186
tri -412 11088 -314 11186 ne
rect -314 11138 0 11186
tri 0 11138 88 11226 sw
tri 98 11138 186 11226 ne
rect 186 11190 240 11226
rect 360 11226 462 11310
tri 462 11226 550 11314 sw
tri 560 11226 648 11314 ne
rect 648 11310 1012 11314
rect 648 11226 790 11310
rect 360 11190 550 11226
rect 186 11186 550 11190
tri 550 11186 590 11226 sw
tri 648 11186 688 11226 ne
rect 688 11190 790 11226
rect 910 11226 1012 11310
tri 1012 11226 1100 11314 sw
tri 1110 11226 1198 11314 ne
rect 1198 11310 1562 11314
rect 1198 11226 1340 11310
rect 910 11190 1100 11226
rect 688 11186 1100 11190
rect 186 11138 590 11186
rect -314 11088 88 11138
rect -1025 11000 -412 11088
tri -412 11000 -324 11088 sw
tri -314 11000 -226 11088 ne
rect -226 11058 88 11088
tri 88 11058 168 11138 sw
tri 186 11058 266 11138 ne
rect 266 11088 590 11138
tri 590 11088 688 11186 sw
tri 688 11088 786 11186 ne
rect 786 11138 1100 11186
tri 1100 11138 1188 11226 sw
tri 1198 11138 1286 11226 ne
rect 1286 11190 1340 11226
rect 1460 11226 1562 11310
tri 1562 11226 1650 11314 sw
tri 1660 11226 1748 11314 ne
rect 1748 11310 2112 11314
rect 1748 11226 1890 11310
rect 1460 11190 1650 11226
rect 1286 11186 1650 11190
tri 1650 11186 1690 11226 sw
tri 1748 11186 1788 11226 ne
rect 1788 11190 1890 11226
rect 2010 11226 2112 11310
tri 2112 11226 2200 11314 sw
tri 2210 11226 2298 11314 ne
rect 2298 11310 2662 11314
rect 2298 11226 2440 11310
rect 2010 11190 2200 11226
rect 1788 11186 2200 11190
rect 1286 11138 1690 11186
rect 786 11088 1188 11138
rect 266 11058 688 11088
rect -226 11000 168 11058
rect -1025 10960 -324 11000
tri -324 10960 -284 11000 sw
tri -226 10960 -186 11000 ne
rect -186 10960 168 11000
tri 168 10960 266 11058 sw
tri 266 10960 364 11058 ne
rect 364 11000 688 11058
tri 688 11000 776 11088 sw
tri 786 11000 874 11088 ne
rect 874 11058 1188 11088
tri 1188 11058 1268 11138 sw
tri 1286 11058 1366 11138 ne
rect 1366 11088 1690 11138
tri 1690 11088 1788 11186 sw
tri 1788 11088 1886 11186 ne
rect 1886 11138 2200 11186
tri 2200 11138 2288 11226 sw
tri 2298 11138 2386 11226 ne
rect 2386 11190 2440 11226
rect 2560 11226 2662 11310
tri 2662 11226 2750 11314 sw
tri 2760 11226 2848 11314 ne
rect 2848 11310 3212 11314
rect 2848 11226 2990 11310
rect 2560 11190 2750 11226
rect 2386 11186 2750 11190
tri 2750 11186 2790 11226 sw
tri 2848 11186 2888 11226 ne
rect 2888 11190 2990 11226
rect 3110 11226 3212 11310
tri 3212 11226 3300 11314 sw
tri 3310 11226 3398 11314 ne
rect 3398 11310 3762 11314
rect 3398 11226 3540 11310
rect 3110 11190 3300 11226
rect 2888 11186 3300 11190
rect 2386 11138 2790 11186
rect 1886 11088 2288 11138
rect 1366 11058 1788 11088
rect 874 11000 1268 11058
rect 364 10960 776 11000
tri 776 10960 816 11000 sw
tri 874 10960 914 11000 ne
rect 914 10960 1268 11000
tri 1268 10960 1366 11058 sw
tri 1366 10960 1464 11058 ne
rect 1464 11000 1788 11058
tri 1788 11000 1876 11088 sw
tri 1886 11000 1974 11088 ne
rect 1974 11058 2288 11088
tri 2288 11058 2368 11138 sw
tri 2386 11058 2466 11138 ne
rect 2466 11088 2790 11138
tri 2790 11088 2888 11186 sw
tri 2888 11088 2986 11186 ne
rect 2986 11138 3300 11186
tri 3300 11138 3388 11226 sw
tri 3398 11138 3486 11226 ne
rect 3486 11190 3540 11226
rect 3660 11226 3762 11310
tri 3762 11226 3850 11314 sw
tri 3860 11226 3948 11314 ne
rect 3948 11310 4312 11314
rect 3948 11226 4090 11310
rect 3660 11190 3850 11226
rect 3486 11186 3850 11190
tri 3850 11186 3890 11226 sw
tri 3948 11186 3988 11226 ne
rect 3988 11190 4090 11226
rect 4210 11226 4312 11310
tri 4312 11226 4400 11314 sw
tri 4410 11226 4498 11314 ne
rect 4498 11310 4862 11314
rect 4498 11226 4640 11310
rect 4210 11190 4400 11226
rect 3988 11186 4400 11190
rect 3486 11138 3890 11186
rect 2986 11088 3388 11138
rect 2466 11058 2888 11088
rect 1974 11000 2368 11058
rect 1464 10960 1876 11000
tri 1876 10960 1916 11000 sw
tri 1974 10960 2014 11000 ne
rect 2014 10960 2368 11000
tri 2368 10960 2466 11058 sw
tri 2466 10960 2564 11058 ne
rect 2564 11000 2888 11058
tri 2888 11000 2976 11088 sw
tri 2986 11000 3074 11088 ne
rect 3074 11058 3388 11088
tri 3388 11058 3468 11138 sw
tri 3486 11058 3566 11138 ne
rect 3566 11088 3890 11138
tri 3890 11088 3988 11186 sw
tri 3988 11088 4086 11186 ne
rect 4086 11138 4400 11186
tri 4400 11138 4488 11226 sw
tri 4498 11138 4586 11226 ne
rect 4586 11190 4640 11226
rect 4760 11226 4862 11310
tri 4862 11226 4950 11314 sw
tri 4960 11226 5048 11314 ne
rect 5048 11310 5412 11314
rect 5048 11226 5190 11310
rect 4760 11190 4950 11226
rect 4586 11186 4950 11190
tri 4950 11186 4990 11226 sw
tri 5048 11186 5088 11226 ne
rect 5088 11190 5190 11226
rect 5310 11226 5412 11310
tri 5412 11226 5500 11314 sw
tri 5510 11226 5598 11314 ne
rect 5598 11310 5962 11314
rect 5598 11226 5740 11310
rect 5310 11190 5500 11226
rect 5088 11186 5500 11190
rect 4586 11138 4990 11186
rect 4086 11088 4488 11138
rect 3566 11058 3988 11088
rect 3074 11000 3468 11058
rect 2564 10960 2976 11000
tri 2976 10960 3016 11000 sw
tri 3074 10960 3114 11000 ne
rect 3114 10960 3468 11000
tri 3468 10960 3566 11058 sw
tri 3566 10960 3664 11058 ne
rect 3664 11000 3988 11058
tri 3988 11000 4076 11088 sw
tri 4086 11000 4174 11088 ne
rect 4174 11058 4488 11088
tri 4488 11058 4568 11138 sw
tri 4586 11058 4666 11138 ne
rect 4666 11088 4990 11138
tri 4990 11088 5088 11186 sw
tri 5088 11088 5186 11186 ne
rect 5186 11138 5500 11186
tri 5500 11138 5588 11226 sw
tri 5598 11138 5686 11226 ne
rect 5686 11190 5740 11226
rect 5860 11226 5962 11310
tri 5962 11226 6050 11314 sw
tri 6060 11226 6148 11314 ne
rect 6148 11310 6512 11314
rect 6148 11226 6290 11310
rect 5860 11190 6050 11226
rect 5686 11186 6050 11190
tri 6050 11186 6090 11226 sw
tri 6148 11186 6188 11226 ne
rect 6188 11190 6290 11226
rect 6410 11226 6512 11310
tri 6512 11226 6600 11314 sw
tri 6610 11226 6698 11314 ne
rect 6698 11310 7062 11314
rect 6698 11226 6840 11310
rect 6410 11190 6600 11226
rect 6188 11186 6600 11190
rect 5686 11138 6090 11186
rect 5186 11088 5588 11138
rect 4666 11058 5088 11088
rect 4174 11000 4568 11058
rect 3664 10960 4076 11000
tri 4076 10960 4116 11000 sw
tri 4174 10960 4214 11000 ne
rect 4214 10960 4568 11000
tri 4568 10960 4666 11058 sw
tri 4666 10960 4764 11058 ne
rect 4764 11000 5088 11058
tri 5088 11000 5176 11088 sw
tri 5186 11000 5274 11088 ne
rect 5274 11058 5588 11088
tri 5588 11058 5668 11138 sw
tri 5686 11058 5766 11138 ne
rect 5766 11088 6090 11138
tri 6090 11088 6188 11186 sw
tri 6188 11088 6286 11186 ne
rect 6286 11138 6600 11186
tri 6600 11138 6688 11226 sw
tri 6698 11138 6786 11226 ne
rect 6786 11190 6840 11226
rect 6960 11226 7062 11310
tri 7062 11226 7150 11314 sw
tri 7160 11226 7248 11314 ne
rect 7248 11310 7612 11314
rect 7248 11226 7390 11310
rect 6960 11190 7150 11226
rect 6786 11186 7150 11190
tri 7150 11186 7190 11226 sw
tri 7248 11186 7288 11226 ne
rect 7288 11190 7390 11226
rect 7510 11226 7612 11310
tri 7612 11226 7700 11314 sw
tri 7710 11226 7798 11314 ne
rect 7798 11310 8162 11314
rect 7798 11226 7940 11310
rect 7510 11190 7700 11226
rect 7288 11186 7700 11190
rect 6786 11138 7190 11186
rect 6286 11088 6688 11138
rect 5766 11058 6188 11088
rect 5274 11000 5668 11058
rect 4764 10960 5176 11000
tri 5176 10960 5216 11000 sw
tri 5274 10960 5314 11000 ne
rect 5314 10960 5668 11000
tri 5668 10960 5766 11058 sw
tri 5766 10960 5864 11058 ne
rect 5864 11000 6188 11058
tri 6188 11000 6276 11088 sw
tri 6286 11000 6374 11088 ne
rect 6374 11058 6688 11088
tri 6688 11058 6768 11138 sw
tri 6786 11058 6866 11138 ne
rect 6866 11088 7190 11138
tri 7190 11088 7288 11186 sw
tri 7288 11088 7386 11186 ne
rect 7386 11138 7700 11186
tri 7700 11138 7788 11226 sw
tri 7798 11138 7886 11226 ne
rect 7886 11190 7940 11226
rect 8060 11226 8162 11310
tri 8162 11226 8250 11314 sw
tri 8260 11226 8348 11314 ne
rect 8348 11310 8712 11314
rect 8348 11226 8490 11310
rect 8060 11190 8250 11226
rect 7886 11186 8250 11190
tri 8250 11186 8290 11226 sw
tri 8348 11186 8388 11226 ne
rect 8388 11190 8490 11226
rect 8610 11226 8712 11310
tri 8712 11226 8800 11314 sw
tri 8810 11226 8898 11314 ne
rect 8898 11310 9262 11314
rect 8898 11226 9040 11310
rect 8610 11190 8800 11226
rect 8388 11186 8800 11190
rect 7886 11138 8290 11186
rect 7386 11088 7788 11138
rect 6866 11058 7288 11088
rect 6374 11000 6768 11058
rect 5864 10960 6276 11000
tri 6276 10960 6316 11000 sw
tri 6374 10960 6414 11000 ne
rect 6414 10960 6768 11000
tri 6768 10960 6866 11058 sw
tri 6866 10960 6964 11058 ne
rect 6964 11000 7288 11058
tri 7288 11000 7376 11088 sw
tri 7386 11000 7474 11088 ne
rect 7474 11058 7788 11088
tri 7788 11058 7868 11138 sw
tri 7886 11058 7966 11138 ne
rect 7966 11088 8290 11138
tri 8290 11088 8388 11186 sw
tri 8388 11088 8486 11186 ne
rect 8486 11138 8800 11186
tri 8800 11138 8888 11226 sw
tri 8898 11138 8986 11226 ne
rect 8986 11190 9040 11226
rect 9160 11226 9262 11310
tri 9262 11226 9350 11314 sw
tri 9360 11226 9448 11314 ne
rect 9448 11310 9812 11314
rect 9448 11226 9590 11310
rect 9160 11190 9350 11226
rect 8986 11186 9350 11190
tri 9350 11186 9390 11226 sw
tri 9448 11186 9488 11226 ne
rect 9488 11190 9590 11226
rect 9710 11226 9812 11310
tri 9812 11226 9900 11314 sw
tri 9910 11226 9998 11314 ne
rect 9998 11310 10362 11314
rect 9998 11226 10140 11310
rect 9710 11190 9900 11226
rect 9488 11186 9900 11190
rect 8986 11138 9390 11186
rect 8486 11088 8888 11138
rect 7966 11058 8388 11088
rect 7474 11000 7868 11058
rect 6964 10960 7376 11000
tri 7376 10960 7416 11000 sw
tri 7474 10960 7514 11000 ne
rect 7514 10960 7868 11000
tri 7868 10960 7966 11058 sw
tri 7966 10960 8064 11058 ne
rect 8064 11000 8388 11058
tri 8388 11000 8476 11088 sw
tri 8486 11000 8574 11088 ne
rect 8574 11058 8888 11088
tri 8888 11058 8968 11138 sw
tri 8986 11058 9066 11138 ne
rect 9066 11088 9390 11138
tri 9390 11088 9488 11186 sw
tri 9488 11088 9586 11186 ne
rect 9586 11138 9900 11186
tri 9900 11138 9988 11226 sw
tri 9998 11138 10086 11226 ne
rect 10086 11190 10140 11226
rect 10260 11226 10362 11310
tri 10362 11226 10450 11314 sw
tri 10460 11226 10548 11314 ne
rect 10548 11310 10912 11314
rect 10548 11226 10690 11310
rect 10260 11190 10450 11226
rect 10086 11186 10450 11190
tri 10450 11186 10490 11226 sw
tri 10548 11186 10588 11226 ne
rect 10588 11190 10690 11226
rect 10810 11226 10912 11310
tri 10912 11226 11000 11314 sw
tri 11010 11226 11098 11314 ne
rect 11098 11310 11462 11314
rect 11098 11226 11240 11310
rect 10810 11190 11000 11226
rect 10588 11186 11000 11190
rect 10086 11138 10490 11186
rect 9586 11088 9988 11138
rect 9066 11058 9488 11088
rect 8574 11000 8968 11058
rect 8064 10960 8476 11000
tri 8476 10960 8516 11000 sw
tri 8574 10960 8614 11000 ne
rect 8614 10960 8968 11000
tri 8968 10960 9066 11058 sw
tri 9066 10960 9164 11058 ne
rect 9164 11000 9488 11058
tri 9488 11000 9576 11088 sw
tri 9586 11000 9674 11088 ne
rect 9674 11058 9988 11088
tri 9988 11058 10068 11138 sw
tri 10086 11058 10166 11138 ne
rect 10166 11088 10490 11138
tri 10490 11088 10588 11186 sw
tri 10588 11088 10686 11186 ne
rect 10686 11138 11000 11186
tri 11000 11138 11088 11226 sw
tri 11098 11138 11186 11226 ne
rect 11186 11190 11240 11226
rect 11360 11226 11462 11310
tri 11462 11226 11550 11314 sw
tri 11560 11226 11648 11314 ne
rect 11648 11310 12012 11314
rect 11648 11226 11790 11310
rect 11360 11190 11550 11226
rect 11186 11186 11550 11190
tri 11550 11186 11590 11226 sw
tri 11648 11186 11688 11226 ne
rect 11688 11190 11790 11226
rect 11910 11226 12012 11310
tri 12012 11226 12100 11314 sw
tri 12110 11226 12198 11314 ne
rect 12198 11310 12562 11314
rect 12198 11226 12340 11310
rect 11910 11190 12100 11226
rect 11688 11186 12100 11190
rect 11186 11138 11590 11186
rect 10686 11088 11088 11138
rect 10166 11058 10588 11088
rect 9674 11000 10068 11058
rect 9164 10960 9576 11000
tri 9576 10960 9616 11000 sw
tri 9674 10960 9714 11000 ne
rect 9714 10960 10068 11000
tri 10068 10960 10166 11058 sw
tri 10166 10960 10264 11058 ne
rect 10264 11000 10588 11058
tri 10588 11000 10676 11088 sw
tri 10686 11000 10774 11088 ne
rect 10774 11058 11088 11088
tri 11088 11058 11168 11138 sw
tri 11186 11058 11266 11138 ne
rect 11266 11088 11590 11138
tri 11590 11088 11688 11186 sw
tri 11688 11088 11786 11186 ne
rect 11786 11138 12100 11186
tri 12100 11138 12188 11226 sw
tri 12198 11138 12286 11226 ne
rect 12286 11190 12340 11226
rect 12460 11226 12562 11310
tri 12562 11226 12650 11314 sw
tri 12660 11226 12748 11314 ne
rect 12748 11310 13112 11314
rect 12748 11226 12890 11310
rect 12460 11190 12650 11226
rect 12286 11186 12650 11190
tri 12650 11186 12690 11226 sw
tri 12748 11186 12788 11226 ne
rect 12788 11190 12890 11226
rect 13010 11226 13112 11310
tri 13112 11226 13200 11314 sw
tri 13210 11226 13298 11314 ne
rect 13298 11310 15775 11314
rect 13298 11226 13440 11310
rect 13010 11190 13200 11226
rect 12788 11186 13200 11190
rect 12286 11138 12690 11186
rect 11786 11088 12188 11138
rect 11266 11058 11688 11088
rect 10774 11000 11168 11058
rect 10264 10960 10676 11000
tri 10676 10960 10716 11000 sw
tri 10774 10960 10814 11000 ne
rect 10814 10960 11168 11000
tri 11168 10960 11266 11058 sw
tri 11266 10960 11364 11058 ne
rect 11364 11000 11688 11058
tri 11688 11000 11776 11088 sw
tri 11786 11000 11874 11088 ne
rect 11874 11058 12188 11088
tri 12188 11058 12268 11138 sw
tri 12286 11058 12366 11138 ne
rect 12366 11088 12690 11138
tri 12690 11088 12788 11186 sw
tri 12788 11088 12886 11186 ne
rect 12886 11138 13200 11186
tri 13200 11138 13288 11226 sw
tri 13298 11138 13386 11226 ne
rect 13386 11190 13440 11226
rect 13560 11190 15775 11310
rect 13386 11138 15775 11190
rect 12886 11088 13288 11138
rect 12366 11058 12788 11088
rect 11874 11000 12268 11058
rect 11364 10960 11776 11000
tri 11776 10960 11816 11000 sw
tri 11874 10960 11914 11000 ne
rect 11914 10960 12268 11000
tri 12268 10960 12366 11058 sw
tri 12366 10960 12464 11058 ne
rect 12464 11000 12788 11058
tri 12788 11000 12876 11088 sw
tri 12886 11000 12974 11088 ne
rect 12974 11058 13288 11088
tri 13288 11058 13368 11138 sw
tri 13386 11058 13466 11138 ne
rect 13466 11058 14075 11138
rect 12974 11000 13368 11058
rect 12464 10960 12876 11000
tri 12876 10960 12916 11000 sw
tri 12974 10960 13014 11000 ne
rect 13014 10960 13368 11000
tri 13368 10960 13466 11058 sw
tri 13466 10960 13564 11058 ne
rect 13564 11038 14075 11058
rect 14175 11038 15775 11138
rect 13564 10960 15775 11038
rect -1025 10912 -284 10960
rect -1025 10812 -925 10912
rect -825 10862 -284 10912
tri -284 10862 -186 10960 sw
tri -186 10862 -88 10960 ne
rect -88 10862 266 10960
tri 266 10862 364 10960 sw
tri 364 10862 462 10960 ne
rect 462 10862 816 10960
tri 816 10862 914 10960 sw
tri 914 10862 1012 10960 ne
rect 1012 10862 1366 10960
tri 1366 10862 1464 10960 sw
tri 1464 10862 1562 10960 ne
rect 1562 10862 1916 10960
tri 1916 10862 2014 10960 sw
tri 2014 10862 2112 10960 ne
rect 2112 10862 2466 10960
tri 2466 10862 2564 10960 sw
tri 2564 10862 2662 10960 ne
rect 2662 10862 3016 10960
tri 3016 10862 3114 10960 sw
tri 3114 10862 3212 10960 ne
rect 3212 10862 3566 10960
tri 3566 10862 3664 10960 sw
tri 3664 10862 3762 10960 ne
rect 3762 10862 4116 10960
tri 4116 10862 4214 10960 sw
tri 4214 10862 4312 10960 ne
rect 4312 10862 4666 10960
tri 4666 10862 4764 10960 sw
tri 4764 10862 4862 10960 ne
rect 4862 10862 5216 10960
tri 5216 10862 5314 10960 sw
tri 5314 10862 5412 10960 ne
rect 5412 10862 5766 10960
tri 5766 10862 5864 10960 sw
tri 5864 10862 5962 10960 ne
rect 5962 10862 6316 10960
tri 6316 10862 6414 10960 sw
tri 6414 10862 6512 10960 ne
rect 6512 10862 6866 10960
tri 6866 10862 6964 10960 sw
tri 6964 10862 7062 10960 ne
rect 7062 10862 7416 10960
tri 7416 10862 7514 10960 sw
tri 7514 10862 7612 10960 ne
rect 7612 10862 7966 10960
tri 7966 10862 8064 10960 sw
tri 8064 10862 8162 10960 ne
rect 8162 10862 8516 10960
tri 8516 10862 8614 10960 sw
tri 8614 10862 8712 10960 ne
rect 8712 10862 9066 10960
tri 9066 10862 9164 10960 sw
tri 9164 10862 9262 10960 ne
rect 9262 10862 9616 10960
tri 9616 10862 9714 10960 sw
tri 9714 10862 9812 10960 ne
rect 9812 10862 10166 10960
tri 10166 10862 10264 10960 sw
tri 10264 10862 10362 10960 ne
rect 10362 10862 10716 10960
tri 10716 10862 10814 10960 sw
tri 10814 10862 10912 10960 ne
rect 10912 10862 11266 10960
tri 11266 10862 11364 10960 sw
tri 11364 10862 11462 10960 ne
rect 11462 10862 11816 10960
tri 11816 10862 11914 10960 sw
tri 11914 10862 12012 10960 ne
rect 12012 10862 12366 10960
tri 12366 10862 12464 10960 sw
tri 12464 10862 12562 10960 ne
rect 12562 10862 12916 10960
tri 12916 10862 13014 10960 sw
tri 13014 10862 13112 10960 ne
rect 13112 10862 13466 10960
tri 13466 10862 13564 10960 sw
tri 13564 10862 13662 10960 ne
rect 13662 10862 15775 10960
rect -825 10812 -186 10862
rect -1025 10764 -186 10812
tri -186 10764 -88 10862 sw
tri -88 10764 10 10862 ne
rect 10 10764 364 10862
tri 364 10764 462 10862 sw
tri 462 10764 560 10862 ne
rect 560 10764 914 10862
tri 914 10764 1012 10862 sw
tri 1012 10764 1110 10862 ne
rect 1110 10764 1464 10862
tri 1464 10764 1562 10862 sw
tri 1562 10764 1660 10862 ne
rect 1660 10764 2014 10862
tri 2014 10764 2112 10862 sw
tri 2112 10764 2210 10862 ne
rect 2210 10764 2564 10862
tri 2564 10764 2662 10862 sw
tri 2662 10764 2760 10862 ne
rect 2760 10764 3114 10862
tri 3114 10764 3212 10862 sw
tri 3212 10764 3310 10862 ne
rect 3310 10764 3664 10862
tri 3664 10764 3762 10862 sw
tri 3762 10764 3860 10862 ne
rect 3860 10764 4214 10862
tri 4214 10764 4312 10862 sw
tri 4312 10764 4410 10862 ne
rect 4410 10764 4764 10862
tri 4764 10764 4862 10862 sw
tri 4862 10764 4960 10862 ne
rect 4960 10764 5314 10862
tri 5314 10764 5412 10862 sw
tri 5412 10764 5510 10862 ne
rect 5510 10764 5864 10862
tri 5864 10764 5962 10862 sw
tri 5962 10764 6060 10862 ne
rect 6060 10764 6414 10862
tri 6414 10764 6512 10862 sw
tri 6512 10764 6610 10862 ne
rect 6610 10764 6964 10862
tri 6964 10764 7062 10862 sw
tri 7062 10764 7160 10862 ne
rect 7160 10764 7514 10862
tri 7514 10764 7612 10862 sw
tri 7612 10764 7710 10862 ne
rect 7710 10764 8064 10862
tri 8064 10764 8162 10862 sw
tri 8162 10764 8260 10862 ne
rect 8260 10764 8614 10862
tri 8614 10764 8712 10862 sw
tri 8712 10764 8810 10862 ne
rect 8810 10764 9164 10862
tri 9164 10764 9262 10862 sw
tri 9262 10764 9360 10862 ne
rect 9360 10764 9714 10862
tri 9714 10764 9812 10862 sw
tri 9812 10764 9910 10862 ne
rect 9910 10764 10264 10862
tri 10264 10764 10362 10862 sw
tri 10362 10764 10460 10862 ne
rect 10460 10764 10814 10862
tri 10814 10764 10912 10862 sw
tri 10912 10764 11010 10862 ne
rect 11010 10764 11364 10862
tri 11364 10764 11462 10862 sw
tri 11462 10764 11560 10862 ne
rect 11560 10764 11914 10862
tri 11914 10764 12012 10862 sw
tri 12012 10764 12110 10862 ne
rect 12110 10764 12464 10862
tri 12464 10764 12562 10862 sw
tri 12562 10764 12660 10862 ne
rect 12660 10764 13014 10862
tri 13014 10764 13112 10862 sw
tri 13112 10764 13210 10862 ne
rect 13210 10764 13564 10862
tri 13564 10764 13662 10862 sw
rect -1025 10760 -88 10764
rect -1025 10640 -310 10760
rect -190 10676 -88 10760
tri -88 10676 0 10764 sw
tri 10 10676 98 10764 ne
rect 98 10760 462 10764
rect 98 10676 240 10760
rect -190 10640 0 10676
rect -1025 10636 0 10640
tri 0 10636 40 10676 sw
tri 98 10636 138 10676 ne
rect 138 10640 240 10676
rect 360 10676 462 10760
tri 462 10676 550 10764 sw
tri 560 10676 648 10764 ne
rect 648 10760 1012 10764
rect 648 10676 790 10760
rect 360 10640 550 10676
rect 138 10636 550 10640
tri -412 10538 -314 10636 ne
rect -314 10538 40 10636
tri 40 10538 138 10636 sw
tri 138 10538 236 10636 ne
rect 236 10588 550 10636
tri 550 10588 638 10676 sw
tri 648 10588 736 10676 ne
rect 736 10640 790 10676
rect 910 10676 1012 10760
tri 1012 10676 1100 10764 sw
tri 1110 10676 1198 10764 ne
rect 1198 10760 1562 10764
rect 1198 10676 1340 10760
rect 910 10640 1100 10676
rect 736 10636 1100 10640
tri 1100 10636 1140 10676 sw
tri 1198 10636 1238 10676 ne
rect 1238 10640 1340 10676
rect 1460 10676 1562 10760
tri 1562 10676 1650 10764 sw
tri 1660 10676 1748 10764 ne
rect 1748 10760 2112 10764
rect 1748 10676 1890 10760
rect 1460 10640 1650 10676
rect 1238 10636 1650 10640
rect 736 10588 1140 10636
rect 236 10538 638 10588
rect -2525 10450 -412 10538
tri -412 10450 -324 10538 sw
tri -314 10450 -226 10538 ne
rect -226 10450 138 10538
tri 138 10450 226 10538 sw
tri 236 10450 324 10538 ne
rect 324 10508 638 10538
tri 638 10508 718 10588 sw
tri 736 10508 816 10588 ne
rect 816 10538 1140 10588
tri 1140 10538 1238 10636 sw
tri 1238 10538 1336 10636 ne
rect 1336 10588 1650 10636
tri 1650 10588 1738 10676 sw
tri 1748 10588 1836 10676 ne
rect 1836 10640 1890 10676
rect 2010 10676 2112 10760
tri 2112 10676 2200 10764 sw
tri 2210 10676 2298 10764 ne
rect 2298 10760 2662 10764
rect 2298 10676 2440 10760
rect 2010 10640 2200 10676
rect 1836 10636 2200 10640
tri 2200 10636 2240 10676 sw
tri 2298 10636 2338 10676 ne
rect 2338 10640 2440 10676
rect 2560 10676 2662 10760
tri 2662 10676 2750 10764 sw
tri 2760 10676 2848 10764 ne
rect 2848 10760 3212 10764
rect 2848 10676 2990 10760
rect 2560 10640 2750 10676
rect 2338 10636 2750 10640
rect 1836 10588 2240 10636
rect 1336 10538 1738 10588
rect 816 10508 1238 10538
rect 324 10450 718 10508
rect -2525 10410 -324 10450
tri -324 10410 -284 10450 sw
tri -226 10410 -186 10450 ne
rect -186 10410 226 10450
tri 226 10410 266 10450 sw
tri 324 10410 364 10450 ne
rect 364 10410 718 10450
tri 718 10410 816 10508 sw
tri 816 10410 914 10508 ne
rect 914 10450 1238 10508
tri 1238 10450 1326 10538 sw
tri 1336 10450 1424 10538 ne
rect 1424 10508 1738 10538
tri 1738 10508 1818 10588 sw
tri 1836 10508 1916 10588 ne
rect 1916 10538 2240 10588
tri 2240 10538 2338 10636 sw
tri 2338 10538 2436 10636 ne
rect 2436 10588 2750 10636
tri 2750 10588 2838 10676 sw
tri 2848 10588 2936 10676 ne
rect 2936 10640 2990 10676
rect 3110 10676 3212 10760
tri 3212 10676 3300 10764 sw
tri 3310 10676 3398 10764 ne
rect 3398 10760 3762 10764
rect 3398 10676 3540 10760
rect 3110 10640 3300 10676
rect 2936 10636 3300 10640
tri 3300 10636 3340 10676 sw
tri 3398 10636 3438 10676 ne
rect 3438 10640 3540 10676
rect 3660 10676 3762 10760
tri 3762 10676 3850 10764 sw
tri 3860 10676 3948 10764 ne
rect 3948 10760 4312 10764
rect 3948 10676 4090 10760
rect 3660 10640 3850 10676
rect 3438 10636 3850 10640
rect 2936 10588 3340 10636
rect 2436 10538 2838 10588
rect 1916 10508 2338 10538
rect 1424 10450 1818 10508
rect 914 10410 1326 10450
tri 1326 10410 1366 10450 sw
tri 1424 10410 1464 10450 ne
rect 1464 10410 1818 10450
tri 1818 10410 1916 10508 sw
tri 1916 10410 2014 10508 ne
rect 2014 10450 2338 10508
tri 2338 10450 2426 10538 sw
tri 2436 10450 2524 10538 ne
rect 2524 10508 2838 10538
tri 2838 10508 2918 10588 sw
tri 2936 10508 3016 10588 ne
rect 3016 10538 3340 10588
tri 3340 10538 3438 10636 sw
tri 3438 10538 3536 10636 ne
rect 3536 10588 3850 10636
tri 3850 10588 3938 10676 sw
tri 3948 10588 4036 10676 ne
rect 4036 10640 4090 10676
rect 4210 10676 4312 10760
tri 4312 10676 4400 10764 sw
tri 4410 10676 4498 10764 ne
rect 4498 10760 4862 10764
rect 4498 10676 4640 10760
rect 4210 10640 4400 10676
rect 4036 10636 4400 10640
tri 4400 10636 4440 10676 sw
tri 4498 10636 4538 10676 ne
rect 4538 10640 4640 10676
rect 4760 10676 4862 10760
tri 4862 10676 4950 10764 sw
tri 4960 10676 5048 10764 ne
rect 5048 10760 5412 10764
rect 5048 10676 5190 10760
rect 4760 10640 4950 10676
rect 4538 10636 4950 10640
rect 4036 10588 4440 10636
rect 3536 10538 3938 10588
rect 3016 10508 3438 10538
rect 2524 10450 2918 10508
rect 2014 10410 2426 10450
tri 2426 10410 2466 10450 sw
tri 2524 10410 2564 10450 ne
rect 2564 10410 2918 10450
tri 2918 10410 3016 10508 sw
tri 3016 10410 3114 10508 ne
rect 3114 10450 3438 10508
tri 3438 10450 3526 10538 sw
tri 3536 10450 3624 10538 ne
rect 3624 10508 3938 10538
tri 3938 10508 4018 10588 sw
tri 4036 10508 4116 10588 ne
rect 4116 10538 4440 10588
tri 4440 10538 4538 10636 sw
tri 4538 10538 4636 10636 ne
rect 4636 10588 4950 10636
tri 4950 10588 5038 10676 sw
tri 5048 10588 5136 10676 ne
rect 5136 10640 5190 10676
rect 5310 10676 5412 10760
tri 5412 10676 5500 10764 sw
tri 5510 10676 5598 10764 ne
rect 5598 10760 5962 10764
rect 5598 10676 5740 10760
rect 5310 10640 5500 10676
rect 5136 10636 5500 10640
tri 5500 10636 5540 10676 sw
tri 5598 10636 5638 10676 ne
rect 5638 10640 5740 10676
rect 5860 10676 5962 10760
tri 5962 10676 6050 10764 sw
tri 6060 10676 6148 10764 ne
rect 6148 10760 6512 10764
rect 6148 10676 6290 10760
rect 5860 10640 6050 10676
rect 5638 10636 6050 10640
rect 5136 10588 5540 10636
rect 4636 10538 5038 10588
rect 4116 10508 4538 10538
rect 3624 10450 4018 10508
rect 3114 10410 3526 10450
tri 3526 10410 3566 10450 sw
tri 3624 10410 3664 10450 ne
rect 3664 10410 4018 10450
tri 4018 10410 4116 10508 sw
tri 4116 10410 4214 10508 ne
rect 4214 10450 4538 10508
tri 4538 10450 4626 10538 sw
tri 4636 10450 4724 10538 ne
rect 4724 10508 5038 10538
tri 5038 10508 5118 10588 sw
tri 5136 10508 5216 10588 ne
rect 5216 10538 5540 10588
tri 5540 10538 5638 10636 sw
tri 5638 10538 5736 10636 ne
rect 5736 10588 6050 10636
tri 6050 10588 6138 10676 sw
tri 6148 10588 6236 10676 ne
rect 6236 10640 6290 10676
rect 6410 10676 6512 10760
tri 6512 10676 6600 10764 sw
tri 6610 10676 6698 10764 ne
rect 6698 10760 7062 10764
rect 6698 10676 6840 10760
rect 6410 10640 6600 10676
rect 6236 10636 6600 10640
tri 6600 10636 6640 10676 sw
tri 6698 10636 6738 10676 ne
rect 6738 10640 6840 10676
rect 6960 10676 7062 10760
tri 7062 10676 7150 10764 sw
tri 7160 10676 7248 10764 ne
rect 7248 10760 7612 10764
rect 7248 10676 7390 10760
rect 6960 10640 7150 10676
rect 6738 10636 7150 10640
rect 6236 10588 6640 10636
rect 5736 10538 6138 10588
rect 5216 10508 5638 10538
rect 4724 10450 5118 10508
rect 4214 10410 4626 10450
tri 4626 10410 4666 10450 sw
tri 4724 10410 4764 10450 ne
rect 4764 10410 5118 10450
tri 5118 10410 5216 10508 sw
tri 5216 10410 5314 10508 ne
rect 5314 10450 5638 10508
tri 5638 10450 5726 10538 sw
tri 5736 10450 5824 10538 ne
rect 5824 10508 6138 10538
tri 6138 10508 6218 10588 sw
tri 6236 10508 6316 10588 ne
rect 6316 10538 6640 10588
tri 6640 10538 6738 10636 sw
tri 6738 10538 6836 10636 ne
rect 6836 10588 7150 10636
tri 7150 10588 7238 10676 sw
tri 7248 10588 7336 10676 ne
rect 7336 10640 7390 10676
rect 7510 10676 7612 10760
tri 7612 10676 7700 10764 sw
tri 7710 10676 7798 10764 ne
rect 7798 10760 8162 10764
rect 7798 10676 7940 10760
rect 7510 10640 7700 10676
rect 7336 10636 7700 10640
tri 7700 10636 7740 10676 sw
tri 7798 10636 7838 10676 ne
rect 7838 10640 7940 10676
rect 8060 10676 8162 10760
tri 8162 10676 8250 10764 sw
tri 8260 10676 8348 10764 ne
rect 8348 10760 8712 10764
rect 8348 10676 8490 10760
rect 8060 10640 8250 10676
rect 7838 10636 8250 10640
rect 7336 10588 7740 10636
rect 6836 10538 7238 10588
rect 6316 10508 6738 10538
rect 5824 10450 6218 10508
rect 5314 10410 5726 10450
tri 5726 10410 5766 10450 sw
tri 5824 10410 5864 10450 ne
rect 5864 10410 6218 10450
tri 6218 10410 6316 10508 sw
tri 6316 10410 6414 10508 ne
rect 6414 10450 6738 10508
tri 6738 10450 6826 10538 sw
tri 6836 10450 6924 10538 ne
rect 6924 10508 7238 10538
tri 7238 10508 7318 10588 sw
tri 7336 10508 7416 10588 ne
rect 7416 10538 7740 10588
tri 7740 10538 7838 10636 sw
tri 7838 10538 7936 10636 ne
rect 7936 10588 8250 10636
tri 8250 10588 8338 10676 sw
tri 8348 10588 8436 10676 ne
rect 8436 10640 8490 10676
rect 8610 10676 8712 10760
tri 8712 10676 8800 10764 sw
tri 8810 10676 8898 10764 ne
rect 8898 10760 9262 10764
rect 8898 10676 9040 10760
rect 8610 10640 8800 10676
rect 8436 10636 8800 10640
tri 8800 10636 8840 10676 sw
tri 8898 10636 8938 10676 ne
rect 8938 10640 9040 10676
rect 9160 10676 9262 10760
tri 9262 10676 9350 10764 sw
tri 9360 10676 9448 10764 ne
rect 9448 10760 9812 10764
rect 9448 10676 9590 10760
rect 9160 10640 9350 10676
rect 8938 10636 9350 10640
rect 8436 10588 8840 10636
rect 7936 10538 8338 10588
rect 7416 10508 7838 10538
rect 6924 10450 7318 10508
rect 6414 10410 6826 10450
tri 6826 10410 6866 10450 sw
tri 6924 10410 6964 10450 ne
rect 6964 10410 7318 10450
tri 7318 10410 7416 10508 sw
tri 7416 10410 7514 10508 ne
rect 7514 10450 7838 10508
tri 7838 10450 7926 10538 sw
tri 7936 10450 8024 10538 ne
rect 8024 10508 8338 10538
tri 8338 10508 8418 10588 sw
tri 8436 10508 8516 10588 ne
rect 8516 10538 8840 10588
tri 8840 10538 8938 10636 sw
tri 8938 10538 9036 10636 ne
rect 9036 10588 9350 10636
tri 9350 10588 9438 10676 sw
tri 9448 10588 9536 10676 ne
rect 9536 10640 9590 10676
rect 9710 10676 9812 10760
tri 9812 10676 9900 10764 sw
tri 9910 10676 9998 10764 ne
rect 9998 10760 10362 10764
rect 9998 10676 10140 10760
rect 9710 10640 9900 10676
rect 9536 10636 9900 10640
tri 9900 10636 9940 10676 sw
tri 9998 10636 10038 10676 ne
rect 10038 10640 10140 10676
rect 10260 10676 10362 10760
tri 10362 10676 10450 10764 sw
tri 10460 10676 10548 10764 ne
rect 10548 10760 10912 10764
rect 10548 10676 10690 10760
rect 10260 10640 10450 10676
rect 10038 10636 10450 10640
rect 9536 10588 9940 10636
rect 9036 10538 9438 10588
rect 8516 10508 8938 10538
rect 8024 10450 8418 10508
rect 7514 10410 7926 10450
tri 7926 10410 7966 10450 sw
tri 8024 10410 8064 10450 ne
rect 8064 10410 8418 10450
tri 8418 10410 8516 10508 sw
tri 8516 10410 8614 10508 ne
rect 8614 10450 8938 10508
tri 8938 10450 9026 10538 sw
tri 9036 10450 9124 10538 ne
rect 9124 10508 9438 10538
tri 9438 10508 9518 10588 sw
tri 9536 10508 9616 10588 ne
rect 9616 10538 9940 10588
tri 9940 10538 10038 10636 sw
tri 10038 10538 10136 10636 ne
rect 10136 10588 10450 10636
tri 10450 10588 10538 10676 sw
tri 10548 10588 10636 10676 ne
rect 10636 10640 10690 10676
rect 10810 10676 10912 10760
tri 10912 10676 11000 10764 sw
tri 11010 10676 11098 10764 ne
rect 11098 10760 11462 10764
rect 11098 10676 11240 10760
rect 10810 10640 11000 10676
rect 10636 10636 11000 10640
tri 11000 10636 11040 10676 sw
tri 11098 10636 11138 10676 ne
rect 11138 10640 11240 10676
rect 11360 10676 11462 10760
tri 11462 10676 11550 10764 sw
tri 11560 10676 11648 10764 ne
rect 11648 10760 12012 10764
rect 11648 10676 11790 10760
rect 11360 10640 11550 10676
rect 11138 10636 11550 10640
rect 10636 10588 11040 10636
rect 10136 10538 10538 10588
rect 9616 10508 10038 10538
rect 9124 10450 9518 10508
rect 8614 10410 9026 10450
tri 9026 10410 9066 10450 sw
tri 9124 10410 9164 10450 ne
rect 9164 10410 9518 10450
tri 9518 10410 9616 10508 sw
tri 9616 10410 9714 10508 ne
rect 9714 10450 10038 10508
tri 10038 10450 10126 10538 sw
tri 10136 10450 10224 10538 ne
rect 10224 10508 10538 10538
tri 10538 10508 10618 10588 sw
tri 10636 10508 10716 10588 ne
rect 10716 10538 11040 10588
tri 11040 10538 11138 10636 sw
tri 11138 10538 11236 10636 ne
rect 11236 10588 11550 10636
tri 11550 10588 11638 10676 sw
tri 11648 10588 11736 10676 ne
rect 11736 10640 11790 10676
rect 11910 10676 12012 10760
tri 12012 10676 12100 10764 sw
tri 12110 10676 12198 10764 ne
rect 12198 10760 12562 10764
rect 12198 10676 12340 10760
rect 11910 10640 12100 10676
rect 11736 10636 12100 10640
tri 12100 10636 12140 10676 sw
tri 12198 10636 12238 10676 ne
rect 12238 10640 12340 10676
rect 12460 10676 12562 10760
tri 12562 10676 12650 10764 sw
tri 12660 10676 12748 10764 ne
rect 12748 10760 13112 10764
rect 12748 10676 12890 10760
rect 12460 10640 12650 10676
rect 12238 10636 12650 10640
rect 11736 10588 12140 10636
rect 11236 10538 11638 10588
rect 10716 10508 11138 10538
rect 10224 10450 10618 10508
rect 9714 10410 10126 10450
tri 10126 10410 10166 10450 sw
tri 10224 10410 10264 10450 ne
rect 10264 10410 10618 10450
tri 10618 10410 10716 10508 sw
tri 10716 10410 10814 10508 ne
rect 10814 10450 11138 10508
tri 11138 10450 11226 10538 sw
tri 11236 10450 11324 10538 ne
rect 11324 10508 11638 10538
tri 11638 10508 11718 10588 sw
tri 11736 10508 11816 10588 ne
rect 11816 10538 12140 10588
tri 12140 10538 12238 10636 sw
tri 12238 10538 12336 10636 ne
rect 12336 10588 12650 10636
tri 12650 10588 12738 10676 sw
tri 12748 10588 12836 10676 ne
rect 12836 10640 12890 10676
rect 13010 10676 13112 10760
tri 13112 10676 13200 10764 sw
tri 13210 10676 13298 10764 ne
rect 13298 10760 14275 10764
rect 13298 10676 13440 10760
rect 13010 10640 13200 10676
rect 12836 10636 13200 10640
tri 13200 10636 13240 10676 sw
tri 13298 10636 13338 10676 ne
rect 13338 10640 13440 10676
rect 13560 10640 14275 10760
rect 13338 10636 14275 10640
rect 12836 10588 13240 10636
rect 12336 10538 12738 10588
rect 11816 10508 12238 10538
rect 11324 10450 11718 10508
rect 10814 10410 11226 10450
tri 11226 10410 11266 10450 sw
tri 11324 10410 11364 10450 ne
rect 11364 10410 11718 10450
tri 11718 10410 11816 10508 sw
tri 11816 10410 11914 10508 ne
rect 11914 10450 12238 10508
tri 12238 10450 12326 10538 sw
tri 12336 10450 12424 10538 ne
rect 12424 10508 12738 10538
tri 12738 10508 12818 10588 sw
tri 12836 10508 12916 10588 ne
rect 12916 10538 13240 10588
tri 13240 10538 13338 10636 sw
tri 13338 10538 13436 10636 ne
rect 13436 10538 14275 10636
rect 12916 10508 13338 10538
rect 12424 10450 12818 10508
rect 11914 10410 12326 10450
tri 12326 10410 12366 10450 sw
tri 12424 10410 12464 10450 ne
rect 12464 10410 12818 10450
tri 12818 10410 12916 10508 sw
tri 12916 10410 13014 10508 ne
rect 13014 10450 13338 10508
tri 13338 10450 13426 10538 sw
tri 13436 10450 13524 10538 ne
rect 13524 10450 14275 10538
rect 13014 10410 13426 10450
tri 13426 10410 13466 10450 sw
tri 13524 10410 13564 10450 ne
rect 13564 10410 14275 10450
rect -2525 10312 -284 10410
tri -284 10312 -186 10410 sw
tri -186 10312 -88 10410 ne
rect -88 10312 266 10410
tri 266 10312 364 10410 sw
tri 364 10312 462 10410 ne
rect 462 10312 816 10410
tri 816 10312 914 10410 sw
tri 914 10312 1012 10410 ne
rect 1012 10312 1366 10410
tri 1366 10312 1464 10410 sw
tri 1464 10312 1562 10410 ne
rect 1562 10312 1916 10410
tri 1916 10312 2014 10410 sw
tri 2014 10312 2112 10410 ne
rect 2112 10312 2466 10410
tri 2466 10312 2564 10410 sw
tri 2564 10312 2662 10410 ne
rect 2662 10312 3016 10410
tri 3016 10312 3114 10410 sw
tri 3114 10312 3212 10410 ne
rect 3212 10312 3566 10410
tri 3566 10312 3664 10410 sw
tri 3664 10312 3762 10410 ne
rect 3762 10312 4116 10410
tri 4116 10312 4214 10410 sw
tri 4214 10312 4312 10410 ne
rect 4312 10312 4666 10410
tri 4666 10312 4764 10410 sw
tri 4764 10312 4862 10410 ne
rect 4862 10312 5216 10410
tri 5216 10312 5314 10410 sw
tri 5314 10312 5412 10410 ne
rect 5412 10312 5766 10410
tri 5766 10312 5864 10410 sw
tri 5864 10312 5962 10410 ne
rect 5962 10312 6316 10410
tri 6316 10312 6414 10410 sw
tri 6414 10312 6512 10410 ne
rect 6512 10312 6866 10410
tri 6866 10312 6964 10410 sw
tri 6964 10312 7062 10410 ne
rect 7062 10312 7416 10410
tri 7416 10312 7514 10410 sw
tri 7514 10312 7612 10410 ne
rect 7612 10312 7966 10410
tri 7966 10312 8064 10410 sw
tri 8064 10312 8162 10410 ne
rect 8162 10312 8516 10410
tri 8516 10312 8614 10410 sw
tri 8614 10312 8712 10410 ne
rect 8712 10312 9066 10410
tri 9066 10312 9164 10410 sw
tri 9164 10312 9262 10410 ne
rect 9262 10312 9616 10410
tri 9616 10312 9714 10410 sw
tri 9714 10312 9812 10410 ne
rect 9812 10312 10166 10410
tri 10166 10312 10264 10410 sw
tri 10264 10312 10362 10410 ne
rect 10362 10312 10716 10410
tri 10716 10312 10814 10410 sw
tri 10814 10312 10912 10410 ne
rect 10912 10312 11266 10410
tri 11266 10312 11364 10410 sw
tri 11364 10312 11462 10410 ne
rect 11462 10312 11816 10410
tri 11816 10312 11914 10410 sw
tri 11914 10312 12012 10410 ne
rect 12012 10312 12366 10410
tri 12366 10312 12464 10410 sw
tri 12464 10312 12562 10410 ne
rect 12562 10312 12916 10410
tri 12916 10312 13014 10410 sw
tri 13014 10312 13112 10410 ne
rect 13112 10312 13466 10410
tri 13466 10312 13564 10410 sw
tri 13564 10312 13662 10410 ne
rect 13662 10312 14275 10410
rect -2525 10214 -186 10312
tri -186 10214 -88 10312 sw
tri -88 10214 10 10312 ne
rect 10 10214 364 10312
tri 364 10214 462 10312 sw
tri 462 10214 560 10312 ne
rect 560 10214 914 10312
tri 914 10214 1012 10312 sw
tri 1012 10214 1110 10312 ne
rect 1110 10214 1464 10312
tri 1464 10214 1562 10312 sw
tri 1562 10214 1660 10312 ne
rect 1660 10214 2014 10312
tri 2014 10214 2112 10312 sw
tri 2112 10214 2210 10312 ne
rect 2210 10214 2564 10312
tri 2564 10214 2662 10312 sw
tri 2662 10214 2760 10312 ne
rect 2760 10214 3114 10312
tri 3114 10214 3212 10312 sw
tri 3212 10214 3310 10312 ne
rect 3310 10214 3664 10312
tri 3664 10214 3762 10312 sw
tri 3762 10214 3860 10312 ne
rect 3860 10214 4214 10312
tri 4214 10214 4312 10312 sw
tri 4312 10214 4410 10312 ne
rect 4410 10214 4764 10312
tri 4764 10214 4862 10312 sw
tri 4862 10214 4960 10312 ne
rect 4960 10214 5314 10312
tri 5314 10214 5412 10312 sw
tri 5412 10214 5510 10312 ne
rect 5510 10214 5864 10312
tri 5864 10214 5962 10312 sw
tri 5962 10214 6060 10312 ne
rect 6060 10214 6414 10312
tri 6414 10214 6512 10312 sw
tri 6512 10214 6610 10312 ne
rect 6610 10214 6964 10312
tri 6964 10214 7062 10312 sw
tri 7062 10214 7160 10312 ne
rect 7160 10214 7514 10312
tri 7514 10214 7612 10312 sw
tri 7612 10214 7710 10312 ne
rect 7710 10214 8064 10312
tri 8064 10214 8162 10312 sw
tri 8162 10214 8260 10312 ne
rect 8260 10214 8614 10312
tri 8614 10214 8712 10312 sw
tri 8712 10214 8810 10312 ne
rect 8810 10214 9164 10312
tri 9164 10214 9262 10312 sw
tri 9262 10214 9360 10312 ne
rect 9360 10214 9714 10312
tri 9714 10214 9812 10312 sw
tri 9812 10214 9910 10312 ne
rect 9910 10214 10264 10312
tri 10264 10214 10362 10312 sw
tri 10362 10214 10460 10312 ne
rect 10460 10214 10814 10312
tri 10814 10214 10912 10312 sw
tri 10912 10214 11010 10312 ne
rect 11010 10214 11364 10312
tri 11364 10214 11462 10312 sw
tri 11462 10214 11560 10312 ne
rect 11560 10214 11914 10312
tri 11914 10214 12012 10312 sw
tri 12012 10214 12110 10312 ne
rect 12110 10214 12464 10312
tri 12464 10214 12562 10312 sw
tri 12562 10214 12660 10312 ne
rect 12660 10214 13014 10312
tri 13014 10214 13112 10312 sw
tri 13112 10214 13210 10312 ne
rect 13210 10214 13564 10312
tri 13564 10214 13662 10312 sw
rect 14775 10214 15775 10862
rect -2525 10210 -88 10214
rect -2525 10090 -310 10210
rect -190 10126 -88 10210
tri -88 10126 0 10214 sw
tri 10 10126 98 10214 ne
rect 98 10210 462 10214
rect 98 10126 240 10210
rect -190 10090 0 10126
rect -2525 10086 0 10090
rect -2525 9438 -1525 10086
tri -412 9988 -314 10086 ne
rect -314 10038 0 10086
tri 0 10038 88 10126 sw
tri 98 10038 186 10126 ne
rect 186 10090 240 10126
rect 360 10126 462 10210
tri 462 10126 550 10214 sw
tri 560 10126 648 10214 ne
rect 648 10210 1012 10214
rect 648 10126 790 10210
rect 360 10090 550 10126
rect 186 10086 550 10090
tri 550 10086 590 10126 sw
tri 648 10086 688 10126 ne
rect 688 10090 790 10126
rect 910 10126 1012 10210
tri 1012 10126 1100 10214 sw
tri 1110 10126 1198 10214 ne
rect 1198 10210 1562 10214
rect 1198 10126 1340 10210
rect 910 10090 1100 10126
rect 688 10086 1100 10090
rect 186 10038 590 10086
rect -314 9988 88 10038
rect -1025 9900 -412 9988
tri -412 9900 -324 9988 sw
tri -314 9900 -226 9988 ne
rect -226 9958 88 9988
tri 88 9958 168 10038 sw
tri 186 9958 266 10038 ne
rect 266 9988 590 10038
tri 590 9988 688 10086 sw
tri 688 9988 786 10086 ne
rect 786 10038 1100 10086
tri 1100 10038 1188 10126 sw
tri 1198 10038 1286 10126 ne
rect 1286 10090 1340 10126
rect 1460 10126 1562 10210
tri 1562 10126 1650 10214 sw
tri 1660 10126 1748 10214 ne
rect 1748 10210 2112 10214
rect 1748 10126 1890 10210
rect 1460 10090 1650 10126
rect 1286 10086 1650 10090
tri 1650 10086 1690 10126 sw
tri 1748 10086 1788 10126 ne
rect 1788 10090 1890 10126
rect 2010 10126 2112 10210
tri 2112 10126 2200 10214 sw
tri 2210 10126 2298 10214 ne
rect 2298 10210 2662 10214
rect 2298 10126 2440 10210
rect 2010 10090 2200 10126
rect 1788 10086 2200 10090
rect 1286 10038 1690 10086
rect 786 9988 1188 10038
rect 266 9958 688 9988
rect -226 9900 168 9958
rect -1025 9860 -324 9900
tri -324 9860 -284 9900 sw
tri -226 9860 -186 9900 ne
rect -186 9860 168 9900
tri 168 9860 266 9958 sw
tri 266 9860 364 9958 ne
rect 364 9900 688 9958
tri 688 9900 776 9988 sw
tri 786 9900 874 9988 ne
rect 874 9958 1188 9988
tri 1188 9958 1268 10038 sw
tri 1286 9958 1366 10038 ne
rect 1366 9988 1690 10038
tri 1690 9988 1788 10086 sw
tri 1788 9988 1886 10086 ne
rect 1886 10038 2200 10086
tri 2200 10038 2288 10126 sw
tri 2298 10038 2386 10126 ne
rect 2386 10090 2440 10126
rect 2560 10126 2662 10210
tri 2662 10126 2750 10214 sw
tri 2760 10126 2848 10214 ne
rect 2848 10210 3212 10214
rect 2848 10126 2990 10210
rect 2560 10090 2750 10126
rect 2386 10086 2750 10090
tri 2750 10086 2790 10126 sw
tri 2848 10086 2888 10126 ne
rect 2888 10090 2990 10126
rect 3110 10126 3212 10210
tri 3212 10126 3300 10214 sw
tri 3310 10126 3398 10214 ne
rect 3398 10210 3762 10214
rect 3398 10126 3540 10210
rect 3110 10090 3300 10126
rect 2888 10086 3300 10090
rect 2386 10038 2790 10086
rect 1886 9988 2288 10038
rect 1366 9958 1788 9988
rect 874 9900 1268 9958
rect 364 9860 776 9900
tri 776 9860 816 9900 sw
tri 874 9860 914 9900 ne
rect 914 9860 1268 9900
tri 1268 9860 1366 9958 sw
tri 1366 9860 1464 9958 ne
rect 1464 9900 1788 9958
tri 1788 9900 1876 9988 sw
tri 1886 9900 1974 9988 ne
rect 1974 9958 2288 9988
tri 2288 9958 2368 10038 sw
tri 2386 9958 2466 10038 ne
rect 2466 9988 2790 10038
tri 2790 9988 2888 10086 sw
tri 2888 9988 2986 10086 ne
rect 2986 10038 3300 10086
tri 3300 10038 3388 10126 sw
tri 3398 10038 3486 10126 ne
rect 3486 10090 3540 10126
rect 3660 10126 3762 10210
tri 3762 10126 3850 10214 sw
tri 3860 10126 3948 10214 ne
rect 3948 10210 4312 10214
rect 3948 10126 4090 10210
rect 3660 10090 3850 10126
rect 3486 10086 3850 10090
tri 3850 10086 3890 10126 sw
tri 3948 10086 3988 10126 ne
rect 3988 10090 4090 10126
rect 4210 10126 4312 10210
tri 4312 10126 4400 10214 sw
tri 4410 10126 4498 10214 ne
rect 4498 10210 4862 10214
rect 4498 10126 4640 10210
rect 4210 10090 4400 10126
rect 3988 10086 4400 10090
rect 3486 10038 3890 10086
rect 2986 9988 3388 10038
rect 2466 9958 2888 9988
rect 1974 9900 2368 9958
rect 1464 9860 1876 9900
tri 1876 9860 1916 9900 sw
tri 1974 9860 2014 9900 ne
rect 2014 9860 2368 9900
tri 2368 9860 2466 9958 sw
tri 2466 9860 2564 9958 ne
rect 2564 9900 2888 9958
tri 2888 9900 2976 9988 sw
tri 2986 9900 3074 9988 ne
rect 3074 9958 3388 9988
tri 3388 9958 3468 10038 sw
tri 3486 9958 3566 10038 ne
rect 3566 9988 3890 10038
tri 3890 9988 3988 10086 sw
tri 3988 9988 4086 10086 ne
rect 4086 10038 4400 10086
tri 4400 10038 4488 10126 sw
tri 4498 10038 4586 10126 ne
rect 4586 10090 4640 10126
rect 4760 10126 4862 10210
tri 4862 10126 4950 10214 sw
tri 4960 10126 5048 10214 ne
rect 5048 10210 5412 10214
rect 5048 10126 5190 10210
rect 4760 10090 4950 10126
rect 4586 10086 4950 10090
tri 4950 10086 4990 10126 sw
tri 5048 10086 5088 10126 ne
rect 5088 10090 5190 10126
rect 5310 10126 5412 10210
tri 5412 10126 5500 10214 sw
tri 5510 10126 5598 10214 ne
rect 5598 10210 5962 10214
rect 5598 10126 5740 10210
rect 5310 10090 5500 10126
rect 5088 10086 5500 10090
rect 4586 10038 4990 10086
rect 4086 9988 4488 10038
rect 3566 9958 3988 9988
rect 3074 9900 3468 9958
rect 2564 9860 2976 9900
tri 2976 9860 3016 9900 sw
tri 3074 9860 3114 9900 ne
rect 3114 9860 3468 9900
tri 3468 9860 3566 9958 sw
tri 3566 9860 3664 9958 ne
rect 3664 9900 3988 9958
tri 3988 9900 4076 9988 sw
tri 4086 9900 4174 9988 ne
rect 4174 9958 4488 9988
tri 4488 9958 4568 10038 sw
tri 4586 9958 4666 10038 ne
rect 4666 9988 4990 10038
tri 4990 9988 5088 10086 sw
tri 5088 9988 5186 10086 ne
rect 5186 10038 5500 10086
tri 5500 10038 5588 10126 sw
tri 5598 10038 5686 10126 ne
rect 5686 10090 5740 10126
rect 5860 10126 5962 10210
tri 5962 10126 6050 10214 sw
tri 6060 10126 6148 10214 ne
rect 6148 10210 6512 10214
rect 6148 10126 6290 10210
rect 5860 10090 6050 10126
rect 5686 10086 6050 10090
tri 6050 10086 6090 10126 sw
tri 6148 10086 6188 10126 ne
rect 6188 10090 6290 10126
rect 6410 10126 6512 10210
tri 6512 10126 6600 10214 sw
tri 6610 10126 6698 10214 ne
rect 6698 10210 7062 10214
rect 6698 10126 6840 10210
rect 6410 10090 6600 10126
rect 6188 10086 6600 10090
rect 5686 10038 6090 10086
rect 5186 9988 5588 10038
rect 4666 9958 5088 9988
rect 4174 9900 4568 9958
rect 3664 9860 4076 9900
tri 4076 9860 4116 9900 sw
tri 4174 9860 4214 9900 ne
rect 4214 9860 4568 9900
tri 4568 9860 4666 9958 sw
tri 4666 9860 4764 9958 ne
rect 4764 9900 5088 9958
tri 5088 9900 5176 9988 sw
tri 5186 9900 5274 9988 ne
rect 5274 9958 5588 9988
tri 5588 9958 5668 10038 sw
tri 5686 9958 5766 10038 ne
rect 5766 9988 6090 10038
tri 6090 9988 6188 10086 sw
tri 6188 9988 6286 10086 ne
rect 6286 10038 6600 10086
tri 6600 10038 6688 10126 sw
tri 6698 10038 6786 10126 ne
rect 6786 10090 6840 10126
rect 6960 10126 7062 10210
tri 7062 10126 7150 10214 sw
tri 7160 10126 7248 10214 ne
rect 7248 10210 7612 10214
rect 7248 10126 7390 10210
rect 6960 10090 7150 10126
rect 6786 10086 7150 10090
tri 7150 10086 7190 10126 sw
tri 7248 10086 7288 10126 ne
rect 7288 10090 7390 10126
rect 7510 10126 7612 10210
tri 7612 10126 7700 10214 sw
tri 7710 10126 7798 10214 ne
rect 7798 10210 8162 10214
rect 7798 10126 7940 10210
rect 7510 10090 7700 10126
rect 7288 10086 7700 10090
rect 6786 10038 7190 10086
rect 6286 9988 6688 10038
rect 5766 9958 6188 9988
rect 5274 9900 5668 9958
rect 4764 9860 5176 9900
tri 5176 9860 5216 9900 sw
tri 5274 9860 5314 9900 ne
rect 5314 9860 5668 9900
tri 5668 9860 5766 9958 sw
tri 5766 9860 5864 9958 ne
rect 5864 9900 6188 9958
tri 6188 9900 6276 9988 sw
tri 6286 9900 6374 9988 ne
rect 6374 9958 6688 9988
tri 6688 9958 6768 10038 sw
tri 6786 9958 6866 10038 ne
rect 6866 9988 7190 10038
tri 7190 9988 7288 10086 sw
tri 7288 9988 7386 10086 ne
rect 7386 10038 7700 10086
tri 7700 10038 7788 10126 sw
tri 7798 10038 7886 10126 ne
rect 7886 10090 7940 10126
rect 8060 10126 8162 10210
tri 8162 10126 8250 10214 sw
tri 8260 10126 8348 10214 ne
rect 8348 10210 8712 10214
rect 8348 10126 8490 10210
rect 8060 10090 8250 10126
rect 7886 10086 8250 10090
tri 8250 10086 8290 10126 sw
tri 8348 10086 8388 10126 ne
rect 8388 10090 8490 10126
rect 8610 10126 8712 10210
tri 8712 10126 8800 10214 sw
tri 8810 10126 8898 10214 ne
rect 8898 10210 9262 10214
rect 8898 10126 9040 10210
rect 8610 10090 8800 10126
rect 8388 10086 8800 10090
rect 7886 10038 8290 10086
rect 7386 9988 7788 10038
rect 6866 9958 7288 9988
rect 6374 9900 6768 9958
rect 5864 9860 6276 9900
tri 6276 9860 6316 9900 sw
tri 6374 9860 6414 9900 ne
rect 6414 9860 6768 9900
tri 6768 9860 6866 9958 sw
tri 6866 9860 6964 9958 ne
rect 6964 9900 7288 9958
tri 7288 9900 7376 9988 sw
tri 7386 9900 7474 9988 ne
rect 7474 9958 7788 9988
tri 7788 9958 7868 10038 sw
tri 7886 9958 7966 10038 ne
rect 7966 9988 8290 10038
tri 8290 9988 8388 10086 sw
tri 8388 9988 8486 10086 ne
rect 8486 10038 8800 10086
tri 8800 10038 8888 10126 sw
tri 8898 10038 8986 10126 ne
rect 8986 10090 9040 10126
rect 9160 10126 9262 10210
tri 9262 10126 9350 10214 sw
tri 9360 10126 9448 10214 ne
rect 9448 10210 9812 10214
rect 9448 10126 9590 10210
rect 9160 10090 9350 10126
rect 8986 10086 9350 10090
tri 9350 10086 9390 10126 sw
tri 9448 10086 9488 10126 ne
rect 9488 10090 9590 10126
rect 9710 10126 9812 10210
tri 9812 10126 9900 10214 sw
tri 9910 10126 9998 10214 ne
rect 9998 10210 10362 10214
rect 9998 10126 10140 10210
rect 9710 10090 9900 10126
rect 9488 10086 9900 10090
rect 8986 10038 9390 10086
rect 8486 9988 8888 10038
rect 7966 9958 8388 9988
rect 7474 9900 7868 9958
rect 6964 9860 7376 9900
tri 7376 9860 7416 9900 sw
tri 7474 9860 7514 9900 ne
rect 7514 9860 7868 9900
tri 7868 9860 7966 9958 sw
tri 7966 9860 8064 9958 ne
rect 8064 9900 8388 9958
tri 8388 9900 8476 9988 sw
tri 8486 9900 8574 9988 ne
rect 8574 9958 8888 9988
tri 8888 9958 8968 10038 sw
tri 8986 9958 9066 10038 ne
rect 9066 9988 9390 10038
tri 9390 9988 9488 10086 sw
tri 9488 9988 9586 10086 ne
rect 9586 10038 9900 10086
tri 9900 10038 9988 10126 sw
tri 9998 10038 10086 10126 ne
rect 10086 10090 10140 10126
rect 10260 10126 10362 10210
tri 10362 10126 10450 10214 sw
tri 10460 10126 10548 10214 ne
rect 10548 10210 10912 10214
rect 10548 10126 10690 10210
rect 10260 10090 10450 10126
rect 10086 10086 10450 10090
tri 10450 10086 10490 10126 sw
tri 10548 10086 10588 10126 ne
rect 10588 10090 10690 10126
rect 10810 10126 10912 10210
tri 10912 10126 11000 10214 sw
tri 11010 10126 11098 10214 ne
rect 11098 10210 11462 10214
rect 11098 10126 11240 10210
rect 10810 10090 11000 10126
rect 10588 10086 11000 10090
rect 10086 10038 10490 10086
rect 9586 9988 9988 10038
rect 9066 9958 9488 9988
rect 8574 9900 8968 9958
rect 8064 9860 8476 9900
tri 8476 9860 8516 9900 sw
tri 8574 9860 8614 9900 ne
rect 8614 9860 8968 9900
tri 8968 9860 9066 9958 sw
tri 9066 9860 9164 9958 ne
rect 9164 9900 9488 9958
tri 9488 9900 9576 9988 sw
tri 9586 9900 9674 9988 ne
rect 9674 9958 9988 9988
tri 9988 9958 10068 10038 sw
tri 10086 9958 10166 10038 ne
rect 10166 9988 10490 10038
tri 10490 9988 10588 10086 sw
tri 10588 9988 10686 10086 ne
rect 10686 10038 11000 10086
tri 11000 10038 11088 10126 sw
tri 11098 10038 11186 10126 ne
rect 11186 10090 11240 10126
rect 11360 10126 11462 10210
tri 11462 10126 11550 10214 sw
tri 11560 10126 11648 10214 ne
rect 11648 10210 12012 10214
rect 11648 10126 11790 10210
rect 11360 10090 11550 10126
rect 11186 10086 11550 10090
tri 11550 10086 11590 10126 sw
tri 11648 10086 11688 10126 ne
rect 11688 10090 11790 10126
rect 11910 10126 12012 10210
tri 12012 10126 12100 10214 sw
tri 12110 10126 12198 10214 ne
rect 12198 10210 12562 10214
rect 12198 10126 12340 10210
rect 11910 10090 12100 10126
rect 11688 10086 12100 10090
rect 11186 10038 11590 10086
rect 10686 9988 11088 10038
rect 10166 9958 10588 9988
rect 9674 9900 10068 9958
rect 9164 9860 9576 9900
tri 9576 9860 9616 9900 sw
tri 9674 9860 9714 9900 ne
rect 9714 9860 10068 9900
tri 10068 9860 10166 9958 sw
tri 10166 9860 10264 9958 ne
rect 10264 9900 10588 9958
tri 10588 9900 10676 9988 sw
tri 10686 9900 10774 9988 ne
rect 10774 9958 11088 9988
tri 11088 9958 11168 10038 sw
tri 11186 9958 11266 10038 ne
rect 11266 9988 11590 10038
tri 11590 9988 11688 10086 sw
tri 11688 9988 11786 10086 ne
rect 11786 10038 12100 10086
tri 12100 10038 12188 10126 sw
tri 12198 10038 12286 10126 ne
rect 12286 10090 12340 10126
rect 12460 10126 12562 10210
tri 12562 10126 12650 10214 sw
tri 12660 10126 12748 10214 ne
rect 12748 10210 13112 10214
rect 12748 10126 12890 10210
rect 12460 10090 12650 10126
rect 12286 10086 12650 10090
tri 12650 10086 12690 10126 sw
tri 12748 10086 12788 10126 ne
rect 12788 10090 12890 10126
rect 13010 10126 13112 10210
tri 13112 10126 13200 10214 sw
tri 13210 10126 13298 10214 ne
rect 13298 10210 15775 10214
rect 13298 10126 13440 10210
rect 13010 10090 13200 10126
rect 12788 10086 13200 10090
rect 12286 10038 12690 10086
rect 11786 9988 12188 10038
rect 11266 9958 11688 9988
rect 10774 9900 11168 9958
rect 10264 9860 10676 9900
tri 10676 9860 10716 9900 sw
tri 10774 9860 10814 9900 ne
rect 10814 9860 11168 9900
tri 11168 9860 11266 9958 sw
tri 11266 9860 11364 9958 ne
rect 11364 9900 11688 9958
tri 11688 9900 11776 9988 sw
tri 11786 9900 11874 9988 ne
rect 11874 9958 12188 9988
tri 12188 9958 12268 10038 sw
tri 12286 9958 12366 10038 ne
rect 12366 9988 12690 10038
tri 12690 9988 12788 10086 sw
tri 12788 9988 12886 10086 ne
rect 12886 10038 13200 10086
tri 13200 10038 13288 10126 sw
tri 13298 10038 13386 10126 ne
rect 13386 10090 13440 10126
rect 13560 10090 15775 10210
rect 13386 10038 15775 10090
rect 12886 9988 13288 10038
rect 12366 9958 12788 9988
rect 11874 9900 12268 9958
rect 11364 9860 11776 9900
tri 11776 9860 11816 9900 sw
tri 11874 9860 11914 9900 ne
rect 11914 9860 12268 9900
tri 12268 9860 12366 9958 sw
tri 12366 9860 12464 9958 ne
rect 12464 9900 12788 9958
tri 12788 9900 12876 9988 sw
tri 12886 9900 12974 9988 ne
rect 12974 9958 13288 9988
tri 13288 9958 13368 10038 sw
tri 13386 9958 13466 10038 ne
rect 13466 9958 14075 10038
rect 12974 9900 13368 9958
rect 12464 9860 12876 9900
tri 12876 9860 12916 9900 sw
tri 12974 9860 13014 9900 ne
rect 13014 9860 13368 9900
tri 13368 9860 13466 9958 sw
tri 13466 9860 13564 9958 ne
rect 13564 9938 14075 9958
rect 14175 9938 15775 10038
rect 13564 9860 15775 9938
rect -1025 9812 -284 9860
rect -1025 9712 -925 9812
rect -825 9762 -284 9812
tri -284 9762 -186 9860 sw
tri -186 9762 -88 9860 ne
rect -88 9762 266 9860
tri 266 9762 364 9860 sw
tri 364 9762 462 9860 ne
rect 462 9762 816 9860
tri 816 9762 914 9860 sw
tri 914 9762 1012 9860 ne
rect 1012 9762 1366 9860
tri 1366 9762 1464 9860 sw
tri 1464 9762 1562 9860 ne
rect 1562 9762 1916 9860
tri 1916 9762 2014 9860 sw
tri 2014 9762 2112 9860 ne
rect 2112 9762 2466 9860
tri 2466 9762 2564 9860 sw
tri 2564 9762 2662 9860 ne
rect 2662 9762 3016 9860
tri 3016 9762 3114 9860 sw
tri 3114 9762 3212 9860 ne
rect 3212 9762 3566 9860
tri 3566 9762 3664 9860 sw
tri 3664 9762 3762 9860 ne
rect 3762 9762 4116 9860
tri 4116 9762 4214 9860 sw
tri 4214 9762 4312 9860 ne
rect 4312 9762 4666 9860
tri 4666 9762 4764 9860 sw
tri 4764 9762 4862 9860 ne
rect 4862 9762 5216 9860
tri 5216 9762 5314 9860 sw
tri 5314 9762 5412 9860 ne
rect 5412 9762 5766 9860
tri 5766 9762 5864 9860 sw
tri 5864 9762 5962 9860 ne
rect 5962 9762 6316 9860
tri 6316 9762 6414 9860 sw
tri 6414 9762 6512 9860 ne
rect 6512 9762 6866 9860
tri 6866 9762 6964 9860 sw
tri 6964 9762 7062 9860 ne
rect 7062 9762 7416 9860
tri 7416 9762 7514 9860 sw
tri 7514 9762 7612 9860 ne
rect 7612 9762 7966 9860
tri 7966 9762 8064 9860 sw
tri 8064 9762 8162 9860 ne
rect 8162 9762 8516 9860
tri 8516 9762 8614 9860 sw
tri 8614 9762 8712 9860 ne
rect 8712 9762 9066 9860
tri 9066 9762 9164 9860 sw
tri 9164 9762 9262 9860 ne
rect 9262 9762 9616 9860
tri 9616 9762 9714 9860 sw
tri 9714 9762 9812 9860 ne
rect 9812 9762 10166 9860
tri 10166 9762 10264 9860 sw
tri 10264 9762 10362 9860 ne
rect 10362 9762 10716 9860
tri 10716 9762 10814 9860 sw
tri 10814 9762 10912 9860 ne
rect 10912 9762 11266 9860
tri 11266 9762 11364 9860 sw
tri 11364 9762 11462 9860 ne
rect 11462 9762 11816 9860
tri 11816 9762 11914 9860 sw
tri 11914 9762 12012 9860 ne
rect 12012 9762 12366 9860
tri 12366 9762 12464 9860 sw
tri 12464 9762 12562 9860 ne
rect 12562 9762 12916 9860
tri 12916 9762 13014 9860 sw
tri 13014 9762 13112 9860 ne
rect 13112 9762 13466 9860
tri 13466 9762 13564 9860 sw
tri 13564 9762 13662 9860 ne
rect 13662 9762 15775 9860
rect -825 9712 -186 9762
rect -1025 9664 -186 9712
tri -186 9664 -88 9762 sw
tri -88 9664 10 9762 ne
rect 10 9664 364 9762
tri 364 9664 462 9762 sw
tri 462 9664 560 9762 ne
rect 560 9664 914 9762
tri 914 9664 1012 9762 sw
tri 1012 9664 1110 9762 ne
rect 1110 9664 1464 9762
tri 1464 9664 1562 9762 sw
tri 1562 9664 1660 9762 ne
rect 1660 9664 2014 9762
tri 2014 9664 2112 9762 sw
tri 2112 9664 2210 9762 ne
rect 2210 9664 2564 9762
tri 2564 9664 2662 9762 sw
tri 2662 9664 2760 9762 ne
rect 2760 9664 3114 9762
tri 3114 9664 3212 9762 sw
tri 3212 9664 3310 9762 ne
rect 3310 9664 3664 9762
tri 3664 9664 3762 9762 sw
tri 3762 9664 3860 9762 ne
rect 3860 9664 4214 9762
tri 4214 9664 4312 9762 sw
tri 4312 9664 4410 9762 ne
rect 4410 9664 4764 9762
tri 4764 9664 4862 9762 sw
tri 4862 9664 4960 9762 ne
rect 4960 9664 5314 9762
tri 5314 9664 5412 9762 sw
tri 5412 9664 5510 9762 ne
rect 5510 9664 5864 9762
tri 5864 9664 5962 9762 sw
tri 5962 9664 6060 9762 ne
rect 6060 9664 6414 9762
tri 6414 9664 6512 9762 sw
tri 6512 9664 6610 9762 ne
rect 6610 9664 6964 9762
tri 6964 9664 7062 9762 sw
tri 7062 9664 7160 9762 ne
rect 7160 9664 7514 9762
tri 7514 9664 7612 9762 sw
tri 7612 9664 7710 9762 ne
rect 7710 9664 8064 9762
tri 8064 9664 8162 9762 sw
tri 8162 9664 8260 9762 ne
rect 8260 9664 8614 9762
tri 8614 9664 8712 9762 sw
tri 8712 9664 8810 9762 ne
rect 8810 9664 9164 9762
tri 9164 9664 9262 9762 sw
tri 9262 9664 9360 9762 ne
rect 9360 9664 9714 9762
tri 9714 9664 9812 9762 sw
tri 9812 9664 9910 9762 ne
rect 9910 9664 10264 9762
tri 10264 9664 10362 9762 sw
tri 10362 9664 10460 9762 ne
rect 10460 9664 10814 9762
tri 10814 9664 10912 9762 sw
tri 10912 9664 11010 9762 ne
rect 11010 9664 11364 9762
tri 11364 9664 11462 9762 sw
tri 11462 9664 11560 9762 ne
rect 11560 9664 11914 9762
tri 11914 9664 12012 9762 sw
tri 12012 9664 12110 9762 ne
rect 12110 9664 12464 9762
tri 12464 9664 12562 9762 sw
tri 12562 9664 12660 9762 ne
rect 12660 9664 13014 9762
tri 13014 9664 13112 9762 sw
tri 13112 9664 13210 9762 ne
rect 13210 9664 13564 9762
tri 13564 9664 13662 9762 sw
rect -1025 9660 -88 9664
rect -1025 9540 -310 9660
rect -190 9576 -88 9660
tri -88 9576 0 9664 sw
tri 10 9576 98 9664 ne
rect 98 9660 462 9664
rect 98 9576 240 9660
rect -190 9540 0 9576
rect -1025 9536 0 9540
tri 0 9536 40 9576 sw
tri 98 9536 138 9576 ne
rect 138 9540 240 9576
rect 360 9576 462 9660
tri 462 9576 550 9664 sw
tri 560 9576 648 9664 ne
rect 648 9660 1012 9664
rect 648 9576 790 9660
rect 360 9540 550 9576
rect 138 9536 550 9540
tri -412 9438 -314 9536 ne
rect -314 9438 40 9536
tri 40 9438 138 9536 sw
tri 138 9438 236 9536 ne
rect 236 9488 550 9536
tri 550 9488 638 9576 sw
tri 648 9488 736 9576 ne
rect 736 9540 790 9576
rect 910 9576 1012 9660
tri 1012 9576 1100 9664 sw
tri 1110 9576 1198 9664 ne
rect 1198 9660 1562 9664
rect 1198 9576 1340 9660
rect 910 9540 1100 9576
rect 736 9536 1100 9540
tri 1100 9536 1140 9576 sw
tri 1198 9536 1238 9576 ne
rect 1238 9540 1340 9576
rect 1460 9576 1562 9660
tri 1562 9576 1650 9664 sw
tri 1660 9576 1748 9664 ne
rect 1748 9660 2112 9664
rect 1748 9576 1890 9660
rect 1460 9540 1650 9576
rect 1238 9536 1650 9540
rect 736 9488 1140 9536
rect 236 9438 638 9488
rect -2525 9350 -412 9438
tri -412 9350 -324 9438 sw
tri -314 9350 -226 9438 ne
rect -226 9350 138 9438
tri 138 9350 226 9438 sw
tri 236 9350 324 9438 ne
rect 324 9408 638 9438
tri 638 9408 718 9488 sw
tri 736 9408 816 9488 ne
rect 816 9438 1140 9488
tri 1140 9438 1238 9536 sw
tri 1238 9438 1336 9536 ne
rect 1336 9488 1650 9536
tri 1650 9488 1738 9576 sw
tri 1748 9488 1836 9576 ne
rect 1836 9540 1890 9576
rect 2010 9576 2112 9660
tri 2112 9576 2200 9664 sw
tri 2210 9576 2298 9664 ne
rect 2298 9660 2662 9664
rect 2298 9576 2440 9660
rect 2010 9540 2200 9576
rect 1836 9536 2200 9540
tri 2200 9536 2240 9576 sw
tri 2298 9536 2338 9576 ne
rect 2338 9540 2440 9576
rect 2560 9576 2662 9660
tri 2662 9576 2750 9664 sw
tri 2760 9576 2848 9664 ne
rect 2848 9660 3212 9664
rect 2848 9576 2990 9660
rect 2560 9540 2750 9576
rect 2338 9536 2750 9540
rect 1836 9488 2240 9536
rect 1336 9438 1738 9488
rect 816 9408 1238 9438
rect 324 9350 718 9408
rect -2525 9310 -324 9350
tri -324 9310 -284 9350 sw
tri -226 9310 -186 9350 ne
rect -186 9310 226 9350
tri 226 9310 266 9350 sw
tri 324 9310 364 9350 ne
rect 364 9310 718 9350
tri 718 9310 816 9408 sw
tri 816 9310 914 9408 ne
rect 914 9350 1238 9408
tri 1238 9350 1326 9438 sw
tri 1336 9350 1424 9438 ne
rect 1424 9408 1738 9438
tri 1738 9408 1818 9488 sw
tri 1836 9408 1916 9488 ne
rect 1916 9438 2240 9488
tri 2240 9438 2338 9536 sw
tri 2338 9438 2436 9536 ne
rect 2436 9488 2750 9536
tri 2750 9488 2838 9576 sw
tri 2848 9488 2936 9576 ne
rect 2936 9540 2990 9576
rect 3110 9576 3212 9660
tri 3212 9576 3300 9664 sw
tri 3310 9576 3398 9664 ne
rect 3398 9660 3762 9664
rect 3398 9576 3540 9660
rect 3110 9540 3300 9576
rect 2936 9536 3300 9540
tri 3300 9536 3340 9576 sw
tri 3398 9536 3438 9576 ne
rect 3438 9540 3540 9576
rect 3660 9576 3762 9660
tri 3762 9576 3850 9664 sw
tri 3860 9576 3948 9664 ne
rect 3948 9660 4312 9664
rect 3948 9576 4090 9660
rect 3660 9540 3850 9576
rect 3438 9536 3850 9540
rect 2936 9488 3340 9536
rect 2436 9438 2838 9488
rect 1916 9408 2338 9438
rect 1424 9350 1818 9408
rect 914 9310 1326 9350
tri 1326 9310 1366 9350 sw
tri 1424 9310 1464 9350 ne
rect 1464 9310 1818 9350
tri 1818 9310 1916 9408 sw
tri 1916 9310 2014 9408 ne
rect 2014 9350 2338 9408
tri 2338 9350 2426 9438 sw
tri 2436 9350 2524 9438 ne
rect 2524 9408 2838 9438
tri 2838 9408 2918 9488 sw
tri 2936 9408 3016 9488 ne
rect 3016 9438 3340 9488
tri 3340 9438 3438 9536 sw
tri 3438 9438 3536 9536 ne
rect 3536 9488 3850 9536
tri 3850 9488 3938 9576 sw
tri 3948 9488 4036 9576 ne
rect 4036 9540 4090 9576
rect 4210 9576 4312 9660
tri 4312 9576 4400 9664 sw
tri 4410 9576 4498 9664 ne
rect 4498 9660 4862 9664
rect 4498 9576 4640 9660
rect 4210 9540 4400 9576
rect 4036 9536 4400 9540
tri 4400 9536 4440 9576 sw
tri 4498 9536 4538 9576 ne
rect 4538 9540 4640 9576
rect 4760 9576 4862 9660
tri 4862 9576 4950 9664 sw
tri 4960 9576 5048 9664 ne
rect 5048 9660 5412 9664
rect 5048 9576 5190 9660
rect 4760 9540 4950 9576
rect 4538 9536 4950 9540
rect 4036 9488 4440 9536
rect 3536 9438 3938 9488
rect 3016 9408 3438 9438
rect 2524 9350 2918 9408
rect 2014 9310 2426 9350
tri 2426 9310 2466 9350 sw
tri 2524 9310 2564 9350 ne
rect 2564 9310 2918 9350
tri 2918 9310 3016 9408 sw
tri 3016 9310 3114 9408 ne
rect 3114 9350 3438 9408
tri 3438 9350 3526 9438 sw
tri 3536 9350 3624 9438 ne
rect 3624 9408 3938 9438
tri 3938 9408 4018 9488 sw
tri 4036 9408 4116 9488 ne
rect 4116 9438 4440 9488
tri 4440 9438 4538 9536 sw
tri 4538 9438 4636 9536 ne
rect 4636 9488 4950 9536
tri 4950 9488 5038 9576 sw
tri 5048 9488 5136 9576 ne
rect 5136 9540 5190 9576
rect 5310 9576 5412 9660
tri 5412 9576 5500 9664 sw
tri 5510 9576 5598 9664 ne
rect 5598 9660 5962 9664
rect 5598 9576 5740 9660
rect 5310 9540 5500 9576
rect 5136 9536 5500 9540
tri 5500 9536 5540 9576 sw
tri 5598 9536 5638 9576 ne
rect 5638 9540 5740 9576
rect 5860 9576 5962 9660
tri 5962 9576 6050 9664 sw
tri 6060 9576 6148 9664 ne
rect 6148 9660 6512 9664
rect 6148 9576 6290 9660
rect 5860 9540 6050 9576
rect 5638 9536 6050 9540
rect 5136 9488 5540 9536
rect 4636 9438 5038 9488
rect 4116 9408 4538 9438
rect 3624 9350 4018 9408
rect 3114 9310 3526 9350
tri 3526 9310 3566 9350 sw
tri 3624 9310 3664 9350 ne
rect 3664 9310 4018 9350
tri 4018 9310 4116 9408 sw
tri 4116 9310 4214 9408 ne
rect 4214 9350 4538 9408
tri 4538 9350 4626 9438 sw
tri 4636 9350 4724 9438 ne
rect 4724 9408 5038 9438
tri 5038 9408 5118 9488 sw
tri 5136 9408 5216 9488 ne
rect 5216 9438 5540 9488
tri 5540 9438 5638 9536 sw
tri 5638 9438 5736 9536 ne
rect 5736 9488 6050 9536
tri 6050 9488 6138 9576 sw
tri 6148 9488 6236 9576 ne
rect 6236 9540 6290 9576
rect 6410 9576 6512 9660
tri 6512 9576 6600 9664 sw
tri 6610 9576 6698 9664 ne
rect 6698 9660 7062 9664
rect 6698 9576 6840 9660
rect 6410 9540 6600 9576
rect 6236 9536 6600 9540
tri 6600 9536 6640 9576 sw
tri 6698 9536 6738 9576 ne
rect 6738 9540 6840 9576
rect 6960 9576 7062 9660
tri 7062 9576 7150 9664 sw
tri 7160 9576 7248 9664 ne
rect 7248 9660 7612 9664
rect 7248 9576 7390 9660
rect 6960 9540 7150 9576
rect 6738 9536 7150 9540
rect 6236 9488 6640 9536
rect 5736 9438 6138 9488
rect 5216 9408 5638 9438
rect 4724 9350 5118 9408
rect 4214 9310 4626 9350
tri 4626 9310 4666 9350 sw
tri 4724 9310 4764 9350 ne
rect 4764 9310 5118 9350
tri 5118 9310 5216 9408 sw
tri 5216 9310 5314 9408 ne
rect 5314 9350 5638 9408
tri 5638 9350 5726 9438 sw
tri 5736 9350 5824 9438 ne
rect 5824 9408 6138 9438
tri 6138 9408 6218 9488 sw
tri 6236 9408 6316 9488 ne
rect 6316 9438 6640 9488
tri 6640 9438 6738 9536 sw
tri 6738 9438 6836 9536 ne
rect 6836 9488 7150 9536
tri 7150 9488 7238 9576 sw
tri 7248 9488 7336 9576 ne
rect 7336 9540 7390 9576
rect 7510 9576 7612 9660
tri 7612 9576 7700 9664 sw
tri 7710 9576 7798 9664 ne
rect 7798 9660 8162 9664
rect 7798 9576 7940 9660
rect 7510 9540 7700 9576
rect 7336 9536 7700 9540
tri 7700 9536 7740 9576 sw
tri 7798 9536 7838 9576 ne
rect 7838 9540 7940 9576
rect 8060 9576 8162 9660
tri 8162 9576 8250 9664 sw
tri 8260 9576 8348 9664 ne
rect 8348 9660 8712 9664
rect 8348 9576 8490 9660
rect 8060 9540 8250 9576
rect 7838 9536 8250 9540
rect 7336 9488 7740 9536
rect 6836 9438 7238 9488
rect 6316 9408 6738 9438
rect 5824 9350 6218 9408
rect 5314 9310 5726 9350
tri 5726 9310 5766 9350 sw
tri 5824 9310 5864 9350 ne
rect 5864 9310 6218 9350
tri 6218 9310 6316 9408 sw
tri 6316 9310 6414 9408 ne
rect 6414 9350 6738 9408
tri 6738 9350 6826 9438 sw
tri 6836 9350 6924 9438 ne
rect 6924 9408 7238 9438
tri 7238 9408 7318 9488 sw
tri 7336 9408 7416 9488 ne
rect 7416 9438 7740 9488
tri 7740 9438 7838 9536 sw
tri 7838 9438 7936 9536 ne
rect 7936 9488 8250 9536
tri 8250 9488 8338 9576 sw
tri 8348 9488 8436 9576 ne
rect 8436 9540 8490 9576
rect 8610 9576 8712 9660
tri 8712 9576 8800 9664 sw
tri 8810 9576 8898 9664 ne
rect 8898 9660 9262 9664
rect 8898 9576 9040 9660
rect 8610 9540 8800 9576
rect 8436 9536 8800 9540
tri 8800 9536 8840 9576 sw
tri 8898 9536 8938 9576 ne
rect 8938 9540 9040 9576
rect 9160 9576 9262 9660
tri 9262 9576 9350 9664 sw
tri 9360 9576 9448 9664 ne
rect 9448 9660 9812 9664
rect 9448 9576 9590 9660
rect 9160 9540 9350 9576
rect 8938 9536 9350 9540
rect 8436 9488 8840 9536
rect 7936 9438 8338 9488
rect 7416 9408 7838 9438
rect 6924 9350 7318 9408
rect 6414 9310 6826 9350
tri 6826 9310 6866 9350 sw
tri 6924 9310 6964 9350 ne
rect 6964 9310 7318 9350
tri 7318 9310 7416 9408 sw
tri 7416 9310 7514 9408 ne
rect 7514 9350 7838 9408
tri 7838 9350 7926 9438 sw
tri 7936 9350 8024 9438 ne
rect 8024 9408 8338 9438
tri 8338 9408 8418 9488 sw
tri 8436 9408 8516 9488 ne
rect 8516 9438 8840 9488
tri 8840 9438 8938 9536 sw
tri 8938 9438 9036 9536 ne
rect 9036 9488 9350 9536
tri 9350 9488 9438 9576 sw
tri 9448 9488 9536 9576 ne
rect 9536 9540 9590 9576
rect 9710 9576 9812 9660
tri 9812 9576 9900 9664 sw
tri 9910 9576 9998 9664 ne
rect 9998 9660 10362 9664
rect 9998 9576 10140 9660
rect 9710 9540 9900 9576
rect 9536 9536 9900 9540
tri 9900 9536 9940 9576 sw
tri 9998 9536 10038 9576 ne
rect 10038 9540 10140 9576
rect 10260 9576 10362 9660
tri 10362 9576 10450 9664 sw
tri 10460 9576 10548 9664 ne
rect 10548 9660 10912 9664
rect 10548 9576 10690 9660
rect 10260 9540 10450 9576
rect 10038 9536 10450 9540
rect 9536 9488 9940 9536
rect 9036 9438 9438 9488
rect 8516 9408 8938 9438
rect 8024 9350 8418 9408
rect 7514 9310 7926 9350
tri 7926 9310 7966 9350 sw
tri 8024 9310 8064 9350 ne
rect 8064 9310 8418 9350
tri 8418 9310 8516 9408 sw
tri 8516 9310 8614 9408 ne
rect 8614 9350 8938 9408
tri 8938 9350 9026 9438 sw
tri 9036 9350 9124 9438 ne
rect 9124 9408 9438 9438
tri 9438 9408 9518 9488 sw
tri 9536 9408 9616 9488 ne
rect 9616 9438 9940 9488
tri 9940 9438 10038 9536 sw
tri 10038 9438 10136 9536 ne
rect 10136 9488 10450 9536
tri 10450 9488 10538 9576 sw
tri 10548 9488 10636 9576 ne
rect 10636 9540 10690 9576
rect 10810 9576 10912 9660
tri 10912 9576 11000 9664 sw
tri 11010 9576 11098 9664 ne
rect 11098 9660 11462 9664
rect 11098 9576 11240 9660
rect 10810 9540 11000 9576
rect 10636 9536 11000 9540
tri 11000 9536 11040 9576 sw
tri 11098 9536 11138 9576 ne
rect 11138 9540 11240 9576
rect 11360 9576 11462 9660
tri 11462 9576 11550 9664 sw
tri 11560 9576 11648 9664 ne
rect 11648 9660 12012 9664
rect 11648 9576 11790 9660
rect 11360 9540 11550 9576
rect 11138 9536 11550 9540
rect 10636 9488 11040 9536
rect 10136 9438 10538 9488
rect 9616 9408 10038 9438
rect 9124 9350 9518 9408
rect 8614 9310 9026 9350
tri 9026 9310 9066 9350 sw
tri 9124 9310 9164 9350 ne
rect 9164 9310 9518 9350
tri 9518 9310 9616 9408 sw
tri 9616 9310 9714 9408 ne
rect 9714 9350 10038 9408
tri 10038 9350 10126 9438 sw
tri 10136 9350 10224 9438 ne
rect 10224 9408 10538 9438
tri 10538 9408 10618 9488 sw
tri 10636 9408 10716 9488 ne
rect 10716 9438 11040 9488
tri 11040 9438 11138 9536 sw
tri 11138 9438 11236 9536 ne
rect 11236 9488 11550 9536
tri 11550 9488 11638 9576 sw
tri 11648 9488 11736 9576 ne
rect 11736 9540 11790 9576
rect 11910 9576 12012 9660
tri 12012 9576 12100 9664 sw
tri 12110 9576 12198 9664 ne
rect 12198 9660 12562 9664
rect 12198 9576 12340 9660
rect 11910 9540 12100 9576
rect 11736 9536 12100 9540
tri 12100 9536 12140 9576 sw
tri 12198 9536 12238 9576 ne
rect 12238 9540 12340 9576
rect 12460 9576 12562 9660
tri 12562 9576 12650 9664 sw
tri 12660 9576 12748 9664 ne
rect 12748 9660 13112 9664
rect 12748 9576 12890 9660
rect 12460 9540 12650 9576
rect 12238 9536 12650 9540
rect 11736 9488 12140 9536
rect 11236 9438 11638 9488
rect 10716 9408 11138 9438
rect 10224 9350 10618 9408
rect 9714 9310 10126 9350
tri 10126 9310 10166 9350 sw
tri 10224 9310 10264 9350 ne
rect 10264 9310 10618 9350
tri 10618 9310 10716 9408 sw
tri 10716 9310 10814 9408 ne
rect 10814 9350 11138 9408
tri 11138 9350 11226 9438 sw
tri 11236 9350 11324 9438 ne
rect 11324 9408 11638 9438
tri 11638 9408 11718 9488 sw
tri 11736 9408 11816 9488 ne
rect 11816 9438 12140 9488
tri 12140 9438 12238 9536 sw
tri 12238 9438 12336 9536 ne
rect 12336 9488 12650 9536
tri 12650 9488 12738 9576 sw
tri 12748 9488 12836 9576 ne
rect 12836 9540 12890 9576
rect 13010 9576 13112 9660
tri 13112 9576 13200 9664 sw
tri 13210 9576 13298 9664 ne
rect 13298 9660 14275 9664
rect 13298 9576 13440 9660
rect 13010 9540 13200 9576
rect 12836 9536 13200 9540
tri 13200 9536 13240 9576 sw
tri 13298 9536 13338 9576 ne
rect 13338 9540 13440 9576
rect 13560 9540 14275 9660
rect 13338 9536 14275 9540
rect 12836 9488 13240 9536
rect 12336 9438 12738 9488
rect 11816 9408 12238 9438
rect 11324 9350 11718 9408
rect 10814 9310 11226 9350
tri 11226 9310 11266 9350 sw
tri 11324 9310 11364 9350 ne
rect 11364 9310 11718 9350
tri 11718 9310 11816 9408 sw
tri 11816 9310 11914 9408 ne
rect 11914 9350 12238 9408
tri 12238 9350 12326 9438 sw
tri 12336 9350 12424 9438 ne
rect 12424 9408 12738 9438
tri 12738 9408 12818 9488 sw
tri 12836 9408 12916 9488 ne
rect 12916 9438 13240 9488
tri 13240 9438 13338 9536 sw
tri 13338 9438 13436 9536 ne
rect 13436 9438 14275 9536
rect 12916 9408 13338 9438
rect 12424 9350 12818 9408
rect 11914 9310 12326 9350
tri 12326 9310 12366 9350 sw
tri 12424 9310 12464 9350 ne
rect 12464 9310 12818 9350
tri 12818 9310 12916 9408 sw
tri 12916 9310 13014 9408 ne
rect 13014 9350 13338 9408
tri 13338 9350 13426 9438 sw
tri 13436 9350 13524 9438 ne
rect 13524 9350 14275 9438
rect 13014 9310 13426 9350
tri 13426 9310 13466 9350 sw
tri 13524 9310 13564 9350 ne
rect 13564 9310 14275 9350
rect -2525 9212 -284 9310
tri -284 9212 -186 9310 sw
tri -186 9212 -88 9310 ne
rect -88 9212 266 9310
tri 266 9212 364 9310 sw
tri 364 9212 462 9310 ne
rect 462 9212 816 9310
tri 816 9212 914 9310 sw
tri 914 9212 1012 9310 ne
rect 1012 9212 1366 9310
tri 1366 9212 1464 9310 sw
tri 1464 9212 1562 9310 ne
rect 1562 9212 1916 9310
tri 1916 9212 2014 9310 sw
tri 2014 9212 2112 9310 ne
rect 2112 9212 2466 9310
tri 2466 9212 2564 9310 sw
tri 2564 9212 2662 9310 ne
rect 2662 9212 3016 9310
tri 3016 9212 3114 9310 sw
tri 3114 9212 3212 9310 ne
rect 3212 9212 3566 9310
tri 3566 9212 3664 9310 sw
tri 3664 9212 3762 9310 ne
rect 3762 9212 4116 9310
tri 4116 9212 4214 9310 sw
tri 4214 9212 4312 9310 ne
rect 4312 9212 4666 9310
tri 4666 9212 4764 9310 sw
tri 4764 9212 4862 9310 ne
rect 4862 9212 5216 9310
tri 5216 9212 5314 9310 sw
tri 5314 9212 5412 9310 ne
rect 5412 9212 5766 9310
tri 5766 9212 5864 9310 sw
tri 5864 9212 5962 9310 ne
rect 5962 9212 6316 9310
tri 6316 9212 6414 9310 sw
tri 6414 9212 6512 9310 ne
rect 6512 9212 6866 9310
tri 6866 9212 6964 9310 sw
tri 6964 9212 7062 9310 ne
rect 7062 9212 7416 9310
tri 7416 9212 7514 9310 sw
tri 7514 9212 7612 9310 ne
rect 7612 9212 7966 9310
tri 7966 9212 8064 9310 sw
tri 8064 9212 8162 9310 ne
rect 8162 9212 8516 9310
tri 8516 9212 8614 9310 sw
tri 8614 9212 8712 9310 ne
rect 8712 9212 9066 9310
tri 9066 9212 9164 9310 sw
tri 9164 9212 9262 9310 ne
rect 9262 9212 9616 9310
tri 9616 9212 9714 9310 sw
tri 9714 9212 9812 9310 ne
rect 9812 9212 10166 9310
tri 10166 9212 10264 9310 sw
tri 10264 9212 10362 9310 ne
rect 10362 9212 10716 9310
tri 10716 9212 10814 9310 sw
tri 10814 9212 10912 9310 ne
rect 10912 9212 11266 9310
tri 11266 9212 11364 9310 sw
tri 11364 9212 11462 9310 ne
rect 11462 9212 11816 9310
tri 11816 9212 11914 9310 sw
tri 11914 9212 12012 9310 ne
rect 12012 9212 12366 9310
tri 12366 9212 12464 9310 sw
tri 12464 9212 12562 9310 ne
rect 12562 9212 12916 9310
tri 12916 9212 13014 9310 sw
tri 13014 9212 13112 9310 ne
rect 13112 9212 13466 9310
tri 13466 9212 13564 9310 sw
tri 13564 9212 13662 9310 ne
rect 13662 9212 14275 9310
rect -2525 9114 -186 9212
tri -186 9114 -88 9212 sw
tri -88 9114 10 9212 ne
rect 10 9114 364 9212
tri 364 9114 462 9212 sw
tri 462 9114 560 9212 ne
rect 560 9114 914 9212
tri 914 9114 1012 9212 sw
tri 1012 9114 1110 9212 ne
rect 1110 9114 1464 9212
tri 1464 9114 1562 9212 sw
tri 1562 9114 1660 9212 ne
rect 1660 9114 2014 9212
tri 2014 9114 2112 9212 sw
tri 2112 9114 2210 9212 ne
rect 2210 9114 2564 9212
tri 2564 9114 2662 9212 sw
tri 2662 9114 2760 9212 ne
rect 2760 9114 3114 9212
tri 3114 9114 3212 9212 sw
tri 3212 9114 3310 9212 ne
rect 3310 9114 3664 9212
tri 3664 9114 3762 9212 sw
tri 3762 9114 3860 9212 ne
rect 3860 9114 4214 9212
tri 4214 9114 4312 9212 sw
tri 4312 9114 4410 9212 ne
rect 4410 9114 4764 9212
tri 4764 9114 4862 9212 sw
tri 4862 9114 4960 9212 ne
rect 4960 9114 5314 9212
tri 5314 9114 5412 9212 sw
tri 5412 9114 5510 9212 ne
rect 5510 9114 5864 9212
tri 5864 9114 5962 9212 sw
tri 5962 9114 6060 9212 ne
rect 6060 9114 6414 9212
tri 6414 9114 6512 9212 sw
tri 6512 9114 6610 9212 ne
rect 6610 9114 6964 9212
tri 6964 9114 7062 9212 sw
tri 7062 9114 7160 9212 ne
rect 7160 9114 7514 9212
tri 7514 9114 7612 9212 sw
tri 7612 9114 7710 9212 ne
rect 7710 9114 8064 9212
tri 8064 9114 8162 9212 sw
tri 8162 9114 8260 9212 ne
rect 8260 9114 8614 9212
tri 8614 9114 8712 9212 sw
tri 8712 9114 8810 9212 ne
rect 8810 9114 9164 9212
tri 9164 9114 9262 9212 sw
tri 9262 9114 9360 9212 ne
rect 9360 9114 9714 9212
tri 9714 9114 9812 9212 sw
tri 9812 9114 9910 9212 ne
rect 9910 9114 10264 9212
tri 10264 9114 10362 9212 sw
tri 10362 9114 10460 9212 ne
rect 10460 9114 10814 9212
tri 10814 9114 10912 9212 sw
tri 10912 9114 11010 9212 ne
rect 11010 9114 11364 9212
tri 11364 9114 11462 9212 sw
tri 11462 9114 11560 9212 ne
rect 11560 9114 11914 9212
tri 11914 9114 12012 9212 sw
tri 12012 9114 12110 9212 ne
rect 12110 9114 12464 9212
tri 12464 9114 12562 9212 sw
tri 12562 9114 12660 9212 ne
rect 12660 9114 13014 9212
tri 13014 9114 13112 9212 sw
tri 13112 9114 13210 9212 ne
rect 13210 9114 13564 9212
tri 13564 9114 13662 9212 sw
rect 14775 9114 15775 9762
rect -2525 9110 -88 9114
rect -2525 8990 -310 9110
rect -190 9026 -88 9110
tri -88 9026 0 9114 sw
tri 10 9026 98 9114 ne
rect 98 9110 462 9114
rect 98 9026 240 9110
rect -190 8990 0 9026
rect -2525 8986 0 8990
rect -2525 8338 -1525 8986
tri -412 8888 -314 8986 ne
rect -314 8938 0 8986
tri 0 8938 88 9026 sw
tri 98 8938 186 9026 ne
rect 186 8990 240 9026
rect 360 9026 462 9110
tri 462 9026 550 9114 sw
tri 560 9026 648 9114 ne
rect 648 9110 1012 9114
rect 648 9026 790 9110
rect 360 8990 550 9026
rect 186 8986 550 8990
tri 550 8986 590 9026 sw
tri 648 8986 688 9026 ne
rect 688 8990 790 9026
rect 910 9026 1012 9110
tri 1012 9026 1100 9114 sw
tri 1110 9026 1198 9114 ne
rect 1198 9110 1562 9114
rect 1198 9026 1340 9110
rect 910 8990 1100 9026
rect 688 8986 1100 8990
rect 186 8938 590 8986
rect -314 8888 88 8938
rect -1025 8800 -412 8888
tri -412 8800 -324 8888 sw
tri -314 8800 -226 8888 ne
rect -226 8858 88 8888
tri 88 8858 168 8938 sw
tri 186 8858 266 8938 ne
rect 266 8888 590 8938
tri 590 8888 688 8986 sw
tri 688 8888 786 8986 ne
rect 786 8938 1100 8986
tri 1100 8938 1188 9026 sw
tri 1198 8938 1286 9026 ne
rect 1286 8990 1340 9026
rect 1460 9026 1562 9110
tri 1562 9026 1650 9114 sw
tri 1660 9026 1748 9114 ne
rect 1748 9110 2112 9114
rect 1748 9026 1890 9110
rect 1460 8990 1650 9026
rect 1286 8986 1650 8990
tri 1650 8986 1690 9026 sw
tri 1748 8986 1788 9026 ne
rect 1788 8990 1890 9026
rect 2010 9026 2112 9110
tri 2112 9026 2200 9114 sw
tri 2210 9026 2298 9114 ne
rect 2298 9110 2662 9114
rect 2298 9026 2440 9110
rect 2010 8990 2200 9026
rect 1788 8986 2200 8990
rect 1286 8938 1690 8986
rect 786 8888 1188 8938
rect 266 8858 688 8888
rect -226 8800 168 8858
rect -1025 8760 -324 8800
tri -324 8760 -284 8800 sw
tri -226 8760 -186 8800 ne
rect -186 8760 168 8800
tri 168 8760 266 8858 sw
tri 266 8760 364 8858 ne
rect 364 8800 688 8858
tri 688 8800 776 8888 sw
tri 786 8800 874 8888 ne
rect 874 8858 1188 8888
tri 1188 8858 1268 8938 sw
tri 1286 8858 1366 8938 ne
rect 1366 8888 1690 8938
tri 1690 8888 1788 8986 sw
tri 1788 8888 1886 8986 ne
rect 1886 8938 2200 8986
tri 2200 8938 2288 9026 sw
tri 2298 8938 2386 9026 ne
rect 2386 8990 2440 9026
rect 2560 9026 2662 9110
tri 2662 9026 2750 9114 sw
tri 2760 9026 2848 9114 ne
rect 2848 9110 3212 9114
rect 2848 9026 2990 9110
rect 2560 8990 2750 9026
rect 2386 8986 2750 8990
tri 2750 8986 2790 9026 sw
tri 2848 8986 2888 9026 ne
rect 2888 8990 2990 9026
rect 3110 9026 3212 9110
tri 3212 9026 3300 9114 sw
tri 3310 9026 3398 9114 ne
rect 3398 9110 3762 9114
rect 3398 9026 3540 9110
rect 3110 8990 3300 9026
rect 2888 8986 3300 8990
rect 2386 8938 2790 8986
rect 1886 8888 2288 8938
rect 1366 8858 1788 8888
rect 874 8800 1268 8858
rect 364 8760 776 8800
tri 776 8760 816 8800 sw
tri 874 8760 914 8800 ne
rect 914 8760 1268 8800
tri 1268 8760 1366 8858 sw
tri 1366 8760 1464 8858 ne
rect 1464 8800 1788 8858
tri 1788 8800 1876 8888 sw
tri 1886 8800 1974 8888 ne
rect 1974 8858 2288 8888
tri 2288 8858 2368 8938 sw
tri 2386 8858 2466 8938 ne
rect 2466 8888 2790 8938
tri 2790 8888 2888 8986 sw
tri 2888 8888 2986 8986 ne
rect 2986 8938 3300 8986
tri 3300 8938 3388 9026 sw
tri 3398 8938 3486 9026 ne
rect 3486 8990 3540 9026
rect 3660 9026 3762 9110
tri 3762 9026 3850 9114 sw
tri 3860 9026 3948 9114 ne
rect 3948 9110 4312 9114
rect 3948 9026 4090 9110
rect 3660 8990 3850 9026
rect 3486 8986 3850 8990
tri 3850 8986 3890 9026 sw
tri 3948 8986 3988 9026 ne
rect 3988 8990 4090 9026
rect 4210 9026 4312 9110
tri 4312 9026 4400 9114 sw
tri 4410 9026 4498 9114 ne
rect 4498 9110 4862 9114
rect 4498 9026 4640 9110
rect 4210 8990 4400 9026
rect 3988 8986 4400 8990
rect 3486 8938 3890 8986
rect 2986 8888 3388 8938
rect 2466 8858 2888 8888
rect 1974 8800 2368 8858
rect 1464 8760 1876 8800
tri 1876 8760 1916 8800 sw
tri 1974 8760 2014 8800 ne
rect 2014 8760 2368 8800
tri 2368 8760 2466 8858 sw
tri 2466 8760 2564 8858 ne
rect 2564 8800 2888 8858
tri 2888 8800 2976 8888 sw
tri 2986 8800 3074 8888 ne
rect 3074 8858 3388 8888
tri 3388 8858 3468 8938 sw
tri 3486 8858 3566 8938 ne
rect 3566 8888 3890 8938
tri 3890 8888 3988 8986 sw
tri 3988 8888 4086 8986 ne
rect 4086 8938 4400 8986
tri 4400 8938 4488 9026 sw
tri 4498 8938 4586 9026 ne
rect 4586 8990 4640 9026
rect 4760 9026 4862 9110
tri 4862 9026 4950 9114 sw
tri 4960 9026 5048 9114 ne
rect 5048 9110 5412 9114
rect 5048 9026 5190 9110
rect 4760 8990 4950 9026
rect 4586 8986 4950 8990
tri 4950 8986 4990 9026 sw
tri 5048 8986 5088 9026 ne
rect 5088 8990 5190 9026
rect 5310 9026 5412 9110
tri 5412 9026 5500 9114 sw
tri 5510 9026 5598 9114 ne
rect 5598 9110 5962 9114
rect 5598 9026 5740 9110
rect 5310 8990 5500 9026
rect 5088 8986 5500 8990
rect 4586 8938 4990 8986
rect 4086 8888 4488 8938
rect 3566 8858 3988 8888
rect 3074 8800 3468 8858
rect 2564 8760 2976 8800
tri 2976 8760 3016 8800 sw
tri 3074 8760 3114 8800 ne
rect 3114 8760 3468 8800
tri 3468 8760 3566 8858 sw
tri 3566 8760 3664 8858 ne
rect 3664 8800 3988 8858
tri 3988 8800 4076 8888 sw
tri 4086 8800 4174 8888 ne
rect 4174 8858 4488 8888
tri 4488 8858 4568 8938 sw
tri 4586 8858 4666 8938 ne
rect 4666 8888 4990 8938
tri 4990 8888 5088 8986 sw
tri 5088 8888 5186 8986 ne
rect 5186 8938 5500 8986
tri 5500 8938 5588 9026 sw
tri 5598 8938 5686 9026 ne
rect 5686 8990 5740 9026
rect 5860 9026 5962 9110
tri 5962 9026 6050 9114 sw
tri 6060 9026 6148 9114 ne
rect 6148 9110 6512 9114
rect 6148 9026 6290 9110
rect 5860 8990 6050 9026
rect 5686 8986 6050 8990
tri 6050 8986 6090 9026 sw
tri 6148 8986 6188 9026 ne
rect 6188 8990 6290 9026
rect 6410 9026 6512 9110
tri 6512 9026 6600 9114 sw
tri 6610 9026 6698 9114 ne
rect 6698 9110 7062 9114
rect 6698 9026 6840 9110
rect 6410 8990 6600 9026
rect 6188 8986 6600 8990
rect 5686 8938 6090 8986
rect 5186 8888 5588 8938
rect 4666 8858 5088 8888
rect 4174 8800 4568 8858
rect 3664 8760 4076 8800
tri 4076 8760 4116 8800 sw
tri 4174 8760 4214 8800 ne
rect 4214 8760 4568 8800
tri 4568 8760 4666 8858 sw
tri 4666 8760 4764 8858 ne
rect 4764 8800 5088 8858
tri 5088 8800 5176 8888 sw
tri 5186 8800 5274 8888 ne
rect 5274 8858 5588 8888
tri 5588 8858 5668 8938 sw
tri 5686 8858 5766 8938 ne
rect 5766 8888 6090 8938
tri 6090 8888 6188 8986 sw
tri 6188 8888 6286 8986 ne
rect 6286 8938 6600 8986
tri 6600 8938 6688 9026 sw
tri 6698 8938 6786 9026 ne
rect 6786 8990 6840 9026
rect 6960 9026 7062 9110
tri 7062 9026 7150 9114 sw
tri 7160 9026 7248 9114 ne
rect 7248 9110 7612 9114
rect 7248 9026 7390 9110
rect 6960 8990 7150 9026
rect 6786 8986 7150 8990
tri 7150 8986 7190 9026 sw
tri 7248 8986 7288 9026 ne
rect 7288 8990 7390 9026
rect 7510 9026 7612 9110
tri 7612 9026 7700 9114 sw
tri 7710 9026 7798 9114 ne
rect 7798 9110 8162 9114
rect 7798 9026 7940 9110
rect 7510 8990 7700 9026
rect 7288 8986 7700 8990
rect 6786 8938 7190 8986
rect 6286 8888 6688 8938
rect 5766 8858 6188 8888
rect 5274 8800 5668 8858
rect 4764 8760 5176 8800
tri 5176 8760 5216 8800 sw
tri 5274 8760 5314 8800 ne
rect 5314 8760 5668 8800
tri 5668 8760 5766 8858 sw
tri 5766 8760 5864 8858 ne
rect 5864 8800 6188 8858
tri 6188 8800 6276 8888 sw
tri 6286 8800 6374 8888 ne
rect 6374 8858 6688 8888
tri 6688 8858 6768 8938 sw
tri 6786 8858 6866 8938 ne
rect 6866 8888 7190 8938
tri 7190 8888 7288 8986 sw
tri 7288 8888 7386 8986 ne
rect 7386 8938 7700 8986
tri 7700 8938 7788 9026 sw
tri 7798 8938 7886 9026 ne
rect 7886 8990 7940 9026
rect 8060 9026 8162 9110
tri 8162 9026 8250 9114 sw
tri 8260 9026 8348 9114 ne
rect 8348 9110 8712 9114
rect 8348 9026 8490 9110
rect 8060 8990 8250 9026
rect 7886 8986 8250 8990
tri 8250 8986 8290 9026 sw
tri 8348 8986 8388 9026 ne
rect 8388 8990 8490 9026
rect 8610 9026 8712 9110
tri 8712 9026 8800 9114 sw
tri 8810 9026 8898 9114 ne
rect 8898 9110 9262 9114
rect 8898 9026 9040 9110
rect 8610 8990 8800 9026
rect 8388 8986 8800 8990
rect 7886 8938 8290 8986
rect 7386 8888 7788 8938
rect 6866 8858 7288 8888
rect 6374 8800 6768 8858
rect 5864 8760 6276 8800
tri 6276 8760 6316 8800 sw
tri 6374 8760 6414 8800 ne
rect 6414 8760 6768 8800
tri 6768 8760 6866 8858 sw
tri 6866 8760 6964 8858 ne
rect 6964 8800 7288 8858
tri 7288 8800 7376 8888 sw
tri 7386 8800 7474 8888 ne
rect 7474 8858 7788 8888
tri 7788 8858 7868 8938 sw
tri 7886 8858 7966 8938 ne
rect 7966 8888 8290 8938
tri 8290 8888 8388 8986 sw
tri 8388 8888 8486 8986 ne
rect 8486 8938 8800 8986
tri 8800 8938 8888 9026 sw
tri 8898 8938 8986 9026 ne
rect 8986 8990 9040 9026
rect 9160 9026 9262 9110
tri 9262 9026 9350 9114 sw
tri 9360 9026 9448 9114 ne
rect 9448 9110 9812 9114
rect 9448 9026 9590 9110
rect 9160 8990 9350 9026
rect 8986 8986 9350 8990
tri 9350 8986 9390 9026 sw
tri 9448 8986 9488 9026 ne
rect 9488 8990 9590 9026
rect 9710 9026 9812 9110
tri 9812 9026 9900 9114 sw
tri 9910 9026 9998 9114 ne
rect 9998 9110 10362 9114
rect 9998 9026 10140 9110
rect 9710 8990 9900 9026
rect 9488 8986 9900 8990
rect 8986 8938 9390 8986
rect 8486 8888 8888 8938
rect 7966 8858 8388 8888
rect 7474 8800 7868 8858
rect 6964 8760 7376 8800
tri 7376 8760 7416 8800 sw
tri 7474 8760 7514 8800 ne
rect 7514 8760 7868 8800
tri 7868 8760 7966 8858 sw
tri 7966 8760 8064 8858 ne
rect 8064 8800 8388 8858
tri 8388 8800 8476 8888 sw
tri 8486 8800 8574 8888 ne
rect 8574 8858 8888 8888
tri 8888 8858 8968 8938 sw
tri 8986 8858 9066 8938 ne
rect 9066 8888 9390 8938
tri 9390 8888 9488 8986 sw
tri 9488 8888 9586 8986 ne
rect 9586 8938 9900 8986
tri 9900 8938 9988 9026 sw
tri 9998 8938 10086 9026 ne
rect 10086 8990 10140 9026
rect 10260 9026 10362 9110
tri 10362 9026 10450 9114 sw
tri 10460 9026 10548 9114 ne
rect 10548 9110 10912 9114
rect 10548 9026 10690 9110
rect 10260 8990 10450 9026
rect 10086 8986 10450 8990
tri 10450 8986 10490 9026 sw
tri 10548 8986 10588 9026 ne
rect 10588 8990 10690 9026
rect 10810 9026 10912 9110
tri 10912 9026 11000 9114 sw
tri 11010 9026 11098 9114 ne
rect 11098 9110 11462 9114
rect 11098 9026 11240 9110
rect 10810 8990 11000 9026
rect 10588 8986 11000 8990
rect 10086 8938 10490 8986
rect 9586 8888 9988 8938
rect 9066 8858 9488 8888
rect 8574 8800 8968 8858
rect 8064 8760 8476 8800
tri 8476 8760 8516 8800 sw
tri 8574 8760 8614 8800 ne
rect 8614 8760 8968 8800
tri 8968 8760 9066 8858 sw
tri 9066 8760 9164 8858 ne
rect 9164 8800 9488 8858
tri 9488 8800 9576 8888 sw
tri 9586 8800 9674 8888 ne
rect 9674 8858 9988 8888
tri 9988 8858 10068 8938 sw
tri 10086 8858 10166 8938 ne
rect 10166 8888 10490 8938
tri 10490 8888 10588 8986 sw
tri 10588 8888 10686 8986 ne
rect 10686 8938 11000 8986
tri 11000 8938 11088 9026 sw
tri 11098 8938 11186 9026 ne
rect 11186 8990 11240 9026
rect 11360 9026 11462 9110
tri 11462 9026 11550 9114 sw
tri 11560 9026 11648 9114 ne
rect 11648 9110 12012 9114
rect 11648 9026 11790 9110
rect 11360 8990 11550 9026
rect 11186 8986 11550 8990
tri 11550 8986 11590 9026 sw
tri 11648 8986 11688 9026 ne
rect 11688 8990 11790 9026
rect 11910 9026 12012 9110
tri 12012 9026 12100 9114 sw
tri 12110 9026 12198 9114 ne
rect 12198 9110 12562 9114
rect 12198 9026 12340 9110
rect 11910 8990 12100 9026
rect 11688 8986 12100 8990
rect 11186 8938 11590 8986
rect 10686 8888 11088 8938
rect 10166 8858 10588 8888
rect 9674 8800 10068 8858
rect 9164 8760 9576 8800
tri 9576 8760 9616 8800 sw
tri 9674 8760 9714 8800 ne
rect 9714 8760 10068 8800
tri 10068 8760 10166 8858 sw
tri 10166 8760 10264 8858 ne
rect 10264 8800 10588 8858
tri 10588 8800 10676 8888 sw
tri 10686 8800 10774 8888 ne
rect 10774 8858 11088 8888
tri 11088 8858 11168 8938 sw
tri 11186 8858 11266 8938 ne
rect 11266 8888 11590 8938
tri 11590 8888 11688 8986 sw
tri 11688 8888 11786 8986 ne
rect 11786 8938 12100 8986
tri 12100 8938 12188 9026 sw
tri 12198 8938 12286 9026 ne
rect 12286 8990 12340 9026
rect 12460 9026 12562 9110
tri 12562 9026 12650 9114 sw
tri 12660 9026 12748 9114 ne
rect 12748 9110 13112 9114
rect 12748 9026 12890 9110
rect 12460 8990 12650 9026
rect 12286 8986 12650 8990
tri 12650 8986 12690 9026 sw
tri 12748 8986 12788 9026 ne
rect 12788 8990 12890 9026
rect 13010 9026 13112 9110
tri 13112 9026 13200 9114 sw
tri 13210 9026 13298 9114 ne
rect 13298 9110 15775 9114
rect 13298 9026 13440 9110
rect 13010 8990 13200 9026
rect 12788 8986 13200 8990
rect 12286 8938 12690 8986
rect 11786 8888 12188 8938
rect 11266 8858 11688 8888
rect 10774 8800 11168 8858
rect 10264 8760 10676 8800
tri 10676 8760 10716 8800 sw
tri 10774 8760 10814 8800 ne
rect 10814 8760 11168 8800
tri 11168 8760 11266 8858 sw
tri 11266 8760 11364 8858 ne
rect 11364 8800 11688 8858
tri 11688 8800 11776 8888 sw
tri 11786 8800 11874 8888 ne
rect 11874 8858 12188 8888
tri 12188 8858 12268 8938 sw
tri 12286 8858 12366 8938 ne
rect 12366 8888 12690 8938
tri 12690 8888 12788 8986 sw
tri 12788 8888 12886 8986 ne
rect 12886 8938 13200 8986
tri 13200 8938 13288 9026 sw
tri 13298 8938 13386 9026 ne
rect 13386 8990 13440 9026
rect 13560 8990 15775 9110
rect 13386 8938 15775 8990
rect 12886 8888 13288 8938
rect 12366 8858 12788 8888
rect 11874 8800 12268 8858
rect 11364 8760 11776 8800
tri 11776 8760 11816 8800 sw
tri 11874 8760 11914 8800 ne
rect 11914 8760 12268 8800
tri 12268 8760 12366 8858 sw
tri 12366 8760 12464 8858 ne
rect 12464 8800 12788 8858
tri 12788 8800 12876 8888 sw
tri 12886 8800 12974 8888 ne
rect 12974 8858 13288 8888
tri 13288 8858 13368 8938 sw
tri 13386 8858 13466 8938 ne
rect 13466 8858 14075 8938
rect 12974 8800 13368 8858
rect 12464 8760 12876 8800
tri 12876 8760 12916 8800 sw
tri 12974 8760 13014 8800 ne
rect 13014 8760 13368 8800
tri 13368 8760 13466 8858 sw
tri 13466 8760 13564 8858 ne
rect 13564 8838 14075 8858
rect 14175 8838 15775 8938
rect 13564 8760 15775 8838
rect -1025 8712 -284 8760
rect -1025 8612 -925 8712
rect -825 8662 -284 8712
tri -284 8662 -186 8760 sw
tri -186 8662 -88 8760 ne
rect -88 8662 266 8760
tri 266 8662 364 8760 sw
tri 364 8662 462 8760 ne
rect 462 8662 816 8760
tri 816 8662 914 8760 sw
tri 914 8662 1012 8760 ne
rect 1012 8662 1366 8760
tri 1366 8662 1464 8760 sw
tri 1464 8662 1562 8760 ne
rect 1562 8662 1916 8760
tri 1916 8662 2014 8760 sw
tri 2014 8662 2112 8760 ne
rect 2112 8662 2466 8760
tri 2466 8662 2564 8760 sw
tri 2564 8662 2662 8760 ne
rect 2662 8662 3016 8760
tri 3016 8662 3114 8760 sw
tri 3114 8662 3212 8760 ne
rect 3212 8662 3566 8760
tri 3566 8662 3664 8760 sw
tri 3664 8662 3762 8760 ne
rect 3762 8662 4116 8760
tri 4116 8662 4214 8760 sw
tri 4214 8662 4312 8760 ne
rect 4312 8662 4666 8760
tri 4666 8662 4764 8760 sw
tri 4764 8662 4862 8760 ne
rect 4862 8662 5216 8760
tri 5216 8662 5314 8760 sw
tri 5314 8662 5412 8760 ne
rect 5412 8662 5766 8760
tri 5766 8662 5864 8760 sw
tri 5864 8662 5962 8760 ne
rect 5962 8662 6316 8760
tri 6316 8662 6414 8760 sw
tri 6414 8662 6512 8760 ne
rect 6512 8662 6866 8760
tri 6866 8662 6964 8760 sw
tri 6964 8662 7062 8760 ne
rect 7062 8662 7416 8760
tri 7416 8662 7514 8760 sw
tri 7514 8662 7612 8760 ne
rect 7612 8662 7966 8760
tri 7966 8662 8064 8760 sw
tri 8064 8662 8162 8760 ne
rect 8162 8662 8516 8760
tri 8516 8662 8614 8760 sw
tri 8614 8662 8712 8760 ne
rect 8712 8662 9066 8760
tri 9066 8662 9164 8760 sw
tri 9164 8662 9262 8760 ne
rect 9262 8662 9616 8760
tri 9616 8662 9714 8760 sw
tri 9714 8662 9812 8760 ne
rect 9812 8662 10166 8760
tri 10166 8662 10264 8760 sw
tri 10264 8662 10362 8760 ne
rect 10362 8662 10716 8760
tri 10716 8662 10814 8760 sw
tri 10814 8662 10912 8760 ne
rect 10912 8662 11266 8760
tri 11266 8662 11364 8760 sw
tri 11364 8662 11462 8760 ne
rect 11462 8662 11816 8760
tri 11816 8662 11914 8760 sw
tri 11914 8662 12012 8760 ne
rect 12012 8662 12366 8760
tri 12366 8662 12464 8760 sw
tri 12464 8662 12562 8760 ne
rect 12562 8662 12916 8760
tri 12916 8662 13014 8760 sw
tri 13014 8662 13112 8760 ne
rect 13112 8662 13466 8760
tri 13466 8662 13564 8760 sw
tri 13564 8662 13662 8760 ne
rect 13662 8662 15775 8760
rect -825 8612 -186 8662
rect -1025 8564 -186 8612
tri -186 8564 -88 8662 sw
tri -88 8564 10 8662 ne
rect 10 8564 364 8662
tri 364 8564 462 8662 sw
tri 462 8564 560 8662 ne
rect 560 8564 914 8662
tri 914 8564 1012 8662 sw
tri 1012 8564 1110 8662 ne
rect 1110 8564 1464 8662
tri 1464 8564 1562 8662 sw
tri 1562 8564 1660 8662 ne
rect 1660 8564 2014 8662
tri 2014 8564 2112 8662 sw
tri 2112 8564 2210 8662 ne
rect 2210 8564 2564 8662
tri 2564 8564 2662 8662 sw
tri 2662 8564 2760 8662 ne
rect 2760 8564 3114 8662
tri 3114 8564 3212 8662 sw
tri 3212 8564 3310 8662 ne
rect 3310 8564 3664 8662
tri 3664 8564 3762 8662 sw
tri 3762 8564 3860 8662 ne
rect 3860 8564 4214 8662
tri 4214 8564 4312 8662 sw
tri 4312 8564 4410 8662 ne
rect 4410 8564 4764 8662
tri 4764 8564 4862 8662 sw
tri 4862 8564 4960 8662 ne
rect 4960 8564 5314 8662
tri 5314 8564 5412 8662 sw
tri 5412 8564 5510 8662 ne
rect 5510 8564 5864 8662
tri 5864 8564 5962 8662 sw
tri 5962 8564 6060 8662 ne
rect 6060 8564 6414 8662
tri 6414 8564 6512 8662 sw
tri 6512 8564 6610 8662 ne
rect 6610 8564 6964 8662
tri 6964 8564 7062 8662 sw
tri 7062 8564 7160 8662 ne
rect 7160 8564 7514 8662
tri 7514 8564 7612 8662 sw
tri 7612 8564 7710 8662 ne
rect 7710 8564 8064 8662
tri 8064 8564 8162 8662 sw
tri 8162 8564 8260 8662 ne
rect 8260 8564 8614 8662
tri 8614 8564 8712 8662 sw
tri 8712 8564 8810 8662 ne
rect 8810 8564 9164 8662
tri 9164 8564 9262 8662 sw
tri 9262 8564 9360 8662 ne
rect 9360 8564 9714 8662
tri 9714 8564 9812 8662 sw
tri 9812 8564 9910 8662 ne
rect 9910 8564 10264 8662
tri 10264 8564 10362 8662 sw
tri 10362 8564 10460 8662 ne
rect 10460 8564 10814 8662
tri 10814 8564 10912 8662 sw
tri 10912 8564 11010 8662 ne
rect 11010 8564 11364 8662
tri 11364 8564 11462 8662 sw
tri 11462 8564 11560 8662 ne
rect 11560 8564 11914 8662
tri 11914 8564 12012 8662 sw
tri 12012 8564 12110 8662 ne
rect 12110 8564 12464 8662
tri 12464 8564 12562 8662 sw
tri 12562 8564 12660 8662 ne
rect 12660 8564 13014 8662
tri 13014 8564 13112 8662 sw
tri 13112 8564 13210 8662 ne
rect 13210 8564 13564 8662
tri 13564 8564 13662 8662 sw
rect -1025 8560 -88 8564
rect -1025 8440 -310 8560
rect -190 8476 -88 8560
tri -88 8476 0 8564 sw
tri 10 8476 98 8564 ne
rect 98 8560 462 8564
rect 98 8476 240 8560
rect -190 8440 0 8476
rect -1025 8436 0 8440
tri 0 8436 40 8476 sw
tri 98 8436 138 8476 ne
rect 138 8440 240 8476
rect 360 8476 462 8560
tri 462 8476 550 8564 sw
tri 560 8476 648 8564 ne
rect 648 8560 1012 8564
rect 648 8476 790 8560
rect 360 8440 550 8476
rect 138 8436 550 8440
tri -412 8338 -314 8436 ne
rect -314 8338 40 8436
tri 40 8338 138 8436 sw
tri 138 8338 236 8436 ne
rect 236 8388 550 8436
tri 550 8388 638 8476 sw
tri 648 8388 736 8476 ne
rect 736 8440 790 8476
rect 910 8476 1012 8560
tri 1012 8476 1100 8564 sw
tri 1110 8476 1198 8564 ne
rect 1198 8560 1562 8564
rect 1198 8476 1340 8560
rect 910 8440 1100 8476
rect 736 8436 1100 8440
tri 1100 8436 1140 8476 sw
tri 1198 8436 1238 8476 ne
rect 1238 8440 1340 8476
rect 1460 8476 1562 8560
tri 1562 8476 1650 8564 sw
tri 1660 8476 1748 8564 ne
rect 1748 8560 2112 8564
rect 1748 8476 1890 8560
rect 1460 8440 1650 8476
rect 1238 8436 1650 8440
rect 736 8388 1140 8436
rect 236 8338 638 8388
rect -2525 8250 -412 8338
tri -412 8250 -324 8338 sw
tri -314 8250 -226 8338 ne
rect -226 8250 138 8338
tri 138 8250 226 8338 sw
tri 236 8250 324 8338 ne
rect 324 8308 638 8338
tri 638 8308 718 8388 sw
tri 736 8308 816 8388 ne
rect 816 8338 1140 8388
tri 1140 8338 1238 8436 sw
tri 1238 8338 1336 8436 ne
rect 1336 8388 1650 8436
tri 1650 8388 1738 8476 sw
tri 1748 8388 1836 8476 ne
rect 1836 8440 1890 8476
rect 2010 8476 2112 8560
tri 2112 8476 2200 8564 sw
tri 2210 8476 2298 8564 ne
rect 2298 8560 2662 8564
rect 2298 8476 2440 8560
rect 2010 8440 2200 8476
rect 1836 8436 2200 8440
tri 2200 8436 2240 8476 sw
tri 2298 8436 2338 8476 ne
rect 2338 8440 2440 8476
rect 2560 8476 2662 8560
tri 2662 8476 2750 8564 sw
tri 2760 8476 2848 8564 ne
rect 2848 8560 3212 8564
rect 2848 8476 2990 8560
rect 2560 8440 2750 8476
rect 2338 8436 2750 8440
rect 1836 8388 2240 8436
rect 1336 8338 1738 8388
rect 816 8308 1238 8338
rect 324 8250 718 8308
rect -2525 8210 -324 8250
tri -324 8210 -284 8250 sw
tri -226 8210 -186 8250 ne
rect -186 8210 226 8250
tri 226 8210 266 8250 sw
tri 324 8210 364 8250 ne
rect 364 8210 718 8250
tri 718 8210 816 8308 sw
tri 816 8210 914 8308 ne
rect 914 8250 1238 8308
tri 1238 8250 1326 8338 sw
tri 1336 8250 1424 8338 ne
rect 1424 8308 1738 8338
tri 1738 8308 1818 8388 sw
tri 1836 8308 1916 8388 ne
rect 1916 8338 2240 8388
tri 2240 8338 2338 8436 sw
tri 2338 8338 2436 8436 ne
rect 2436 8388 2750 8436
tri 2750 8388 2838 8476 sw
tri 2848 8388 2936 8476 ne
rect 2936 8440 2990 8476
rect 3110 8476 3212 8560
tri 3212 8476 3300 8564 sw
tri 3310 8476 3398 8564 ne
rect 3398 8560 3762 8564
rect 3398 8476 3540 8560
rect 3110 8440 3300 8476
rect 2936 8436 3300 8440
tri 3300 8436 3340 8476 sw
tri 3398 8436 3438 8476 ne
rect 3438 8440 3540 8476
rect 3660 8476 3762 8560
tri 3762 8476 3850 8564 sw
tri 3860 8476 3948 8564 ne
rect 3948 8560 4312 8564
rect 3948 8476 4090 8560
rect 3660 8440 3850 8476
rect 3438 8436 3850 8440
rect 2936 8388 3340 8436
rect 2436 8338 2838 8388
rect 1916 8308 2338 8338
rect 1424 8250 1818 8308
rect 914 8210 1326 8250
tri 1326 8210 1366 8250 sw
tri 1424 8210 1464 8250 ne
rect 1464 8210 1818 8250
tri 1818 8210 1916 8308 sw
tri 1916 8210 2014 8308 ne
rect 2014 8250 2338 8308
tri 2338 8250 2426 8338 sw
tri 2436 8250 2524 8338 ne
rect 2524 8308 2838 8338
tri 2838 8308 2918 8388 sw
tri 2936 8308 3016 8388 ne
rect 3016 8338 3340 8388
tri 3340 8338 3438 8436 sw
tri 3438 8338 3536 8436 ne
rect 3536 8388 3850 8436
tri 3850 8388 3938 8476 sw
tri 3948 8388 4036 8476 ne
rect 4036 8440 4090 8476
rect 4210 8476 4312 8560
tri 4312 8476 4400 8564 sw
tri 4410 8476 4498 8564 ne
rect 4498 8560 4862 8564
rect 4498 8476 4640 8560
rect 4210 8440 4400 8476
rect 4036 8436 4400 8440
tri 4400 8436 4440 8476 sw
tri 4498 8436 4538 8476 ne
rect 4538 8440 4640 8476
rect 4760 8476 4862 8560
tri 4862 8476 4950 8564 sw
tri 4960 8476 5048 8564 ne
rect 5048 8560 5412 8564
rect 5048 8476 5190 8560
rect 4760 8440 4950 8476
rect 4538 8436 4950 8440
rect 4036 8388 4440 8436
rect 3536 8338 3938 8388
rect 3016 8308 3438 8338
rect 2524 8250 2918 8308
rect 2014 8210 2426 8250
tri 2426 8210 2466 8250 sw
tri 2524 8210 2564 8250 ne
rect 2564 8210 2918 8250
tri 2918 8210 3016 8308 sw
tri 3016 8210 3114 8308 ne
rect 3114 8250 3438 8308
tri 3438 8250 3526 8338 sw
tri 3536 8250 3624 8338 ne
rect 3624 8308 3938 8338
tri 3938 8308 4018 8388 sw
tri 4036 8308 4116 8388 ne
rect 4116 8338 4440 8388
tri 4440 8338 4538 8436 sw
tri 4538 8338 4636 8436 ne
rect 4636 8388 4950 8436
tri 4950 8388 5038 8476 sw
tri 5048 8388 5136 8476 ne
rect 5136 8440 5190 8476
rect 5310 8476 5412 8560
tri 5412 8476 5500 8564 sw
tri 5510 8476 5598 8564 ne
rect 5598 8560 5962 8564
rect 5598 8476 5740 8560
rect 5310 8440 5500 8476
rect 5136 8436 5500 8440
tri 5500 8436 5540 8476 sw
tri 5598 8436 5638 8476 ne
rect 5638 8440 5740 8476
rect 5860 8476 5962 8560
tri 5962 8476 6050 8564 sw
tri 6060 8476 6148 8564 ne
rect 6148 8560 6512 8564
rect 6148 8476 6290 8560
rect 5860 8440 6050 8476
rect 5638 8436 6050 8440
rect 5136 8388 5540 8436
rect 4636 8338 5038 8388
rect 4116 8308 4538 8338
rect 3624 8250 4018 8308
rect 3114 8210 3526 8250
tri 3526 8210 3566 8250 sw
tri 3624 8210 3664 8250 ne
rect 3664 8210 4018 8250
tri 4018 8210 4116 8308 sw
tri 4116 8210 4214 8308 ne
rect 4214 8250 4538 8308
tri 4538 8250 4626 8338 sw
tri 4636 8250 4724 8338 ne
rect 4724 8308 5038 8338
tri 5038 8308 5118 8388 sw
tri 5136 8308 5216 8388 ne
rect 5216 8338 5540 8388
tri 5540 8338 5638 8436 sw
tri 5638 8338 5736 8436 ne
rect 5736 8388 6050 8436
tri 6050 8388 6138 8476 sw
tri 6148 8388 6236 8476 ne
rect 6236 8440 6290 8476
rect 6410 8476 6512 8560
tri 6512 8476 6600 8564 sw
tri 6610 8476 6698 8564 ne
rect 6698 8560 7062 8564
rect 6698 8476 6840 8560
rect 6410 8440 6600 8476
rect 6236 8436 6600 8440
tri 6600 8436 6640 8476 sw
tri 6698 8436 6738 8476 ne
rect 6738 8440 6840 8476
rect 6960 8476 7062 8560
tri 7062 8476 7150 8564 sw
tri 7160 8476 7248 8564 ne
rect 7248 8560 7612 8564
rect 7248 8476 7390 8560
rect 6960 8440 7150 8476
rect 6738 8436 7150 8440
rect 6236 8388 6640 8436
rect 5736 8338 6138 8388
rect 5216 8308 5638 8338
rect 4724 8250 5118 8308
rect 4214 8210 4626 8250
tri 4626 8210 4666 8250 sw
tri 4724 8210 4764 8250 ne
rect 4764 8210 5118 8250
tri 5118 8210 5216 8308 sw
tri 5216 8210 5314 8308 ne
rect 5314 8250 5638 8308
tri 5638 8250 5726 8338 sw
tri 5736 8250 5824 8338 ne
rect 5824 8308 6138 8338
tri 6138 8308 6218 8388 sw
tri 6236 8308 6316 8388 ne
rect 6316 8338 6640 8388
tri 6640 8338 6738 8436 sw
tri 6738 8338 6836 8436 ne
rect 6836 8388 7150 8436
tri 7150 8388 7238 8476 sw
tri 7248 8388 7336 8476 ne
rect 7336 8440 7390 8476
rect 7510 8476 7612 8560
tri 7612 8476 7700 8564 sw
tri 7710 8476 7798 8564 ne
rect 7798 8560 8162 8564
rect 7798 8476 7940 8560
rect 7510 8440 7700 8476
rect 7336 8436 7700 8440
tri 7700 8436 7740 8476 sw
tri 7798 8436 7838 8476 ne
rect 7838 8440 7940 8476
rect 8060 8476 8162 8560
tri 8162 8476 8250 8564 sw
tri 8260 8476 8348 8564 ne
rect 8348 8560 8712 8564
rect 8348 8476 8490 8560
rect 8060 8440 8250 8476
rect 7838 8436 8250 8440
rect 7336 8388 7740 8436
rect 6836 8338 7238 8388
rect 6316 8308 6738 8338
rect 5824 8250 6218 8308
rect 5314 8210 5726 8250
tri 5726 8210 5766 8250 sw
tri 5824 8210 5864 8250 ne
rect 5864 8210 6218 8250
tri 6218 8210 6316 8308 sw
tri 6316 8210 6414 8308 ne
rect 6414 8250 6738 8308
tri 6738 8250 6826 8338 sw
tri 6836 8250 6924 8338 ne
rect 6924 8308 7238 8338
tri 7238 8308 7318 8388 sw
tri 7336 8308 7416 8388 ne
rect 7416 8338 7740 8388
tri 7740 8338 7838 8436 sw
tri 7838 8338 7936 8436 ne
rect 7936 8388 8250 8436
tri 8250 8388 8338 8476 sw
tri 8348 8388 8436 8476 ne
rect 8436 8440 8490 8476
rect 8610 8476 8712 8560
tri 8712 8476 8800 8564 sw
tri 8810 8476 8898 8564 ne
rect 8898 8560 9262 8564
rect 8898 8476 9040 8560
rect 8610 8440 8800 8476
rect 8436 8436 8800 8440
tri 8800 8436 8840 8476 sw
tri 8898 8436 8938 8476 ne
rect 8938 8440 9040 8476
rect 9160 8476 9262 8560
tri 9262 8476 9350 8564 sw
tri 9360 8476 9448 8564 ne
rect 9448 8560 9812 8564
rect 9448 8476 9590 8560
rect 9160 8440 9350 8476
rect 8938 8436 9350 8440
rect 8436 8388 8840 8436
rect 7936 8338 8338 8388
rect 7416 8308 7838 8338
rect 6924 8250 7318 8308
rect 6414 8210 6826 8250
tri 6826 8210 6866 8250 sw
tri 6924 8210 6964 8250 ne
rect 6964 8210 7318 8250
tri 7318 8210 7416 8308 sw
tri 7416 8210 7514 8308 ne
rect 7514 8250 7838 8308
tri 7838 8250 7926 8338 sw
tri 7936 8250 8024 8338 ne
rect 8024 8308 8338 8338
tri 8338 8308 8418 8388 sw
tri 8436 8308 8516 8388 ne
rect 8516 8338 8840 8388
tri 8840 8338 8938 8436 sw
tri 8938 8338 9036 8436 ne
rect 9036 8388 9350 8436
tri 9350 8388 9438 8476 sw
tri 9448 8388 9536 8476 ne
rect 9536 8440 9590 8476
rect 9710 8476 9812 8560
tri 9812 8476 9900 8564 sw
tri 9910 8476 9998 8564 ne
rect 9998 8560 10362 8564
rect 9998 8476 10140 8560
rect 9710 8440 9900 8476
rect 9536 8436 9900 8440
tri 9900 8436 9940 8476 sw
tri 9998 8436 10038 8476 ne
rect 10038 8440 10140 8476
rect 10260 8476 10362 8560
tri 10362 8476 10450 8564 sw
tri 10460 8476 10548 8564 ne
rect 10548 8560 10912 8564
rect 10548 8476 10690 8560
rect 10260 8440 10450 8476
rect 10038 8436 10450 8440
rect 9536 8388 9940 8436
rect 9036 8338 9438 8388
rect 8516 8308 8938 8338
rect 8024 8250 8418 8308
rect 7514 8210 7926 8250
tri 7926 8210 7966 8250 sw
tri 8024 8210 8064 8250 ne
rect 8064 8210 8418 8250
tri 8418 8210 8516 8308 sw
tri 8516 8210 8614 8308 ne
rect 8614 8250 8938 8308
tri 8938 8250 9026 8338 sw
tri 9036 8250 9124 8338 ne
rect 9124 8308 9438 8338
tri 9438 8308 9518 8388 sw
tri 9536 8308 9616 8388 ne
rect 9616 8338 9940 8388
tri 9940 8338 10038 8436 sw
tri 10038 8338 10136 8436 ne
rect 10136 8388 10450 8436
tri 10450 8388 10538 8476 sw
tri 10548 8388 10636 8476 ne
rect 10636 8440 10690 8476
rect 10810 8476 10912 8560
tri 10912 8476 11000 8564 sw
tri 11010 8476 11098 8564 ne
rect 11098 8560 11462 8564
rect 11098 8476 11240 8560
rect 10810 8440 11000 8476
rect 10636 8436 11000 8440
tri 11000 8436 11040 8476 sw
tri 11098 8436 11138 8476 ne
rect 11138 8440 11240 8476
rect 11360 8476 11462 8560
tri 11462 8476 11550 8564 sw
tri 11560 8476 11648 8564 ne
rect 11648 8560 12012 8564
rect 11648 8476 11790 8560
rect 11360 8440 11550 8476
rect 11138 8436 11550 8440
rect 10636 8388 11040 8436
rect 10136 8338 10538 8388
rect 9616 8308 10038 8338
rect 9124 8250 9518 8308
rect 8614 8210 9026 8250
tri 9026 8210 9066 8250 sw
tri 9124 8210 9164 8250 ne
rect 9164 8210 9518 8250
tri 9518 8210 9616 8308 sw
tri 9616 8210 9714 8308 ne
rect 9714 8250 10038 8308
tri 10038 8250 10126 8338 sw
tri 10136 8250 10224 8338 ne
rect 10224 8308 10538 8338
tri 10538 8308 10618 8388 sw
tri 10636 8308 10716 8388 ne
rect 10716 8338 11040 8388
tri 11040 8338 11138 8436 sw
tri 11138 8338 11236 8436 ne
rect 11236 8388 11550 8436
tri 11550 8388 11638 8476 sw
tri 11648 8388 11736 8476 ne
rect 11736 8440 11790 8476
rect 11910 8476 12012 8560
tri 12012 8476 12100 8564 sw
tri 12110 8476 12198 8564 ne
rect 12198 8560 12562 8564
rect 12198 8476 12340 8560
rect 11910 8440 12100 8476
rect 11736 8436 12100 8440
tri 12100 8436 12140 8476 sw
tri 12198 8436 12238 8476 ne
rect 12238 8440 12340 8476
rect 12460 8476 12562 8560
tri 12562 8476 12650 8564 sw
tri 12660 8476 12748 8564 ne
rect 12748 8560 13112 8564
rect 12748 8476 12890 8560
rect 12460 8440 12650 8476
rect 12238 8436 12650 8440
rect 11736 8388 12140 8436
rect 11236 8338 11638 8388
rect 10716 8308 11138 8338
rect 10224 8250 10618 8308
rect 9714 8210 10126 8250
tri 10126 8210 10166 8250 sw
tri 10224 8210 10264 8250 ne
rect 10264 8210 10618 8250
tri 10618 8210 10716 8308 sw
tri 10716 8210 10814 8308 ne
rect 10814 8250 11138 8308
tri 11138 8250 11226 8338 sw
tri 11236 8250 11324 8338 ne
rect 11324 8308 11638 8338
tri 11638 8308 11718 8388 sw
tri 11736 8308 11816 8388 ne
rect 11816 8338 12140 8388
tri 12140 8338 12238 8436 sw
tri 12238 8338 12336 8436 ne
rect 12336 8388 12650 8436
tri 12650 8388 12738 8476 sw
tri 12748 8388 12836 8476 ne
rect 12836 8440 12890 8476
rect 13010 8476 13112 8560
tri 13112 8476 13200 8564 sw
tri 13210 8476 13298 8564 ne
rect 13298 8560 14275 8564
rect 13298 8476 13440 8560
rect 13010 8440 13200 8476
rect 12836 8436 13200 8440
tri 13200 8436 13240 8476 sw
tri 13298 8436 13338 8476 ne
rect 13338 8440 13440 8476
rect 13560 8440 14275 8560
rect 13338 8436 14275 8440
rect 12836 8388 13240 8436
rect 12336 8338 12738 8388
rect 11816 8308 12238 8338
rect 11324 8250 11718 8308
rect 10814 8210 11226 8250
tri 11226 8210 11266 8250 sw
tri 11324 8210 11364 8250 ne
rect 11364 8210 11718 8250
tri 11718 8210 11816 8308 sw
tri 11816 8210 11914 8308 ne
rect 11914 8250 12238 8308
tri 12238 8250 12326 8338 sw
tri 12336 8250 12424 8338 ne
rect 12424 8308 12738 8338
tri 12738 8308 12818 8388 sw
tri 12836 8308 12916 8388 ne
rect 12916 8338 13240 8388
tri 13240 8338 13338 8436 sw
tri 13338 8338 13436 8436 ne
rect 13436 8338 14275 8436
rect 12916 8308 13338 8338
rect 12424 8250 12818 8308
rect 11914 8210 12326 8250
tri 12326 8210 12366 8250 sw
tri 12424 8210 12464 8250 ne
rect 12464 8210 12818 8250
tri 12818 8210 12916 8308 sw
tri 12916 8210 13014 8308 ne
rect 13014 8250 13338 8308
tri 13338 8250 13426 8338 sw
tri 13436 8250 13524 8338 ne
rect 13524 8250 14275 8338
rect 13014 8210 13426 8250
tri 13426 8210 13466 8250 sw
tri 13524 8210 13564 8250 ne
rect 13564 8210 14275 8250
rect -2525 8112 -284 8210
tri -284 8112 -186 8210 sw
tri -186 8112 -88 8210 ne
rect -88 8112 266 8210
tri 266 8112 364 8210 sw
tri 364 8112 462 8210 ne
rect 462 8112 816 8210
tri 816 8112 914 8210 sw
tri 914 8112 1012 8210 ne
rect 1012 8112 1366 8210
tri 1366 8112 1464 8210 sw
tri 1464 8112 1562 8210 ne
rect 1562 8112 1916 8210
tri 1916 8112 2014 8210 sw
tri 2014 8112 2112 8210 ne
rect 2112 8112 2466 8210
tri 2466 8112 2564 8210 sw
tri 2564 8112 2662 8210 ne
rect 2662 8112 3016 8210
tri 3016 8112 3114 8210 sw
tri 3114 8112 3212 8210 ne
rect 3212 8112 3566 8210
tri 3566 8112 3664 8210 sw
tri 3664 8112 3762 8210 ne
rect 3762 8112 4116 8210
tri 4116 8112 4214 8210 sw
tri 4214 8112 4312 8210 ne
rect 4312 8112 4666 8210
tri 4666 8112 4764 8210 sw
tri 4764 8112 4862 8210 ne
rect 4862 8112 5216 8210
tri 5216 8112 5314 8210 sw
tri 5314 8112 5412 8210 ne
rect 5412 8112 5766 8210
tri 5766 8112 5864 8210 sw
tri 5864 8112 5962 8210 ne
rect 5962 8112 6316 8210
tri 6316 8112 6414 8210 sw
tri 6414 8112 6512 8210 ne
rect 6512 8112 6866 8210
tri 6866 8112 6964 8210 sw
tri 6964 8112 7062 8210 ne
rect 7062 8112 7416 8210
tri 7416 8112 7514 8210 sw
tri 7514 8112 7612 8210 ne
rect 7612 8112 7966 8210
tri 7966 8112 8064 8210 sw
tri 8064 8112 8162 8210 ne
rect 8162 8112 8516 8210
tri 8516 8112 8614 8210 sw
tri 8614 8112 8712 8210 ne
rect 8712 8112 9066 8210
tri 9066 8112 9164 8210 sw
tri 9164 8112 9262 8210 ne
rect 9262 8112 9616 8210
tri 9616 8112 9714 8210 sw
tri 9714 8112 9812 8210 ne
rect 9812 8112 10166 8210
tri 10166 8112 10264 8210 sw
tri 10264 8112 10362 8210 ne
rect 10362 8112 10716 8210
tri 10716 8112 10814 8210 sw
tri 10814 8112 10912 8210 ne
rect 10912 8112 11266 8210
tri 11266 8112 11364 8210 sw
tri 11364 8112 11462 8210 ne
rect 11462 8112 11816 8210
tri 11816 8112 11914 8210 sw
tri 11914 8112 12012 8210 ne
rect 12012 8112 12366 8210
tri 12366 8112 12464 8210 sw
tri 12464 8112 12562 8210 ne
rect 12562 8112 12916 8210
tri 12916 8112 13014 8210 sw
tri 13014 8112 13112 8210 ne
rect 13112 8112 13466 8210
tri 13466 8112 13564 8210 sw
tri 13564 8112 13662 8210 ne
rect 13662 8112 14275 8210
rect -2525 8014 -186 8112
tri -186 8014 -88 8112 sw
tri -88 8014 10 8112 ne
rect 10 8014 364 8112
tri 364 8014 462 8112 sw
tri 462 8014 560 8112 ne
rect 560 8014 914 8112
tri 914 8014 1012 8112 sw
tri 1012 8014 1110 8112 ne
rect 1110 8014 1464 8112
tri 1464 8014 1562 8112 sw
tri 1562 8014 1660 8112 ne
rect 1660 8014 2014 8112
tri 2014 8014 2112 8112 sw
tri 2112 8014 2210 8112 ne
rect 2210 8014 2564 8112
tri 2564 8014 2662 8112 sw
tri 2662 8014 2760 8112 ne
rect 2760 8014 3114 8112
tri 3114 8014 3212 8112 sw
tri 3212 8014 3310 8112 ne
rect 3310 8014 3664 8112
tri 3664 8014 3762 8112 sw
tri 3762 8014 3860 8112 ne
rect 3860 8014 4214 8112
tri 4214 8014 4312 8112 sw
tri 4312 8014 4410 8112 ne
rect 4410 8014 4764 8112
tri 4764 8014 4862 8112 sw
tri 4862 8014 4960 8112 ne
rect 4960 8014 5314 8112
tri 5314 8014 5412 8112 sw
tri 5412 8014 5510 8112 ne
rect 5510 8014 5864 8112
tri 5864 8014 5962 8112 sw
tri 5962 8014 6060 8112 ne
rect 6060 8014 6414 8112
tri 6414 8014 6512 8112 sw
tri 6512 8014 6610 8112 ne
rect 6610 8014 6964 8112
tri 6964 8014 7062 8112 sw
tri 7062 8014 7160 8112 ne
rect 7160 8014 7514 8112
tri 7514 8014 7612 8112 sw
tri 7612 8014 7710 8112 ne
rect 7710 8014 8064 8112
tri 8064 8014 8162 8112 sw
tri 8162 8014 8260 8112 ne
rect 8260 8014 8614 8112
tri 8614 8014 8712 8112 sw
tri 8712 8014 8810 8112 ne
rect 8810 8014 9164 8112
tri 9164 8014 9262 8112 sw
tri 9262 8014 9360 8112 ne
rect 9360 8014 9714 8112
tri 9714 8014 9812 8112 sw
tri 9812 8014 9910 8112 ne
rect 9910 8014 10264 8112
tri 10264 8014 10362 8112 sw
tri 10362 8014 10460 8112 ne
rect 10460 8014 10814 8112
tri 10814 8014 10912 8112 sw
tri 10912 8014 11010 8112 ne
rect 11010 8014 11364 8112
tri 11364 8014 11462 8112 sw
tri 11462 8014 11560 8112 ne
rect 11560 8014 11914 8112
tri 11914 8014 12012 8112 sw
tri 12012 8014 12110 8112 ne
rect 12110 8014 12464 8112
tri 12464 8014 12562 8112 sw
tri 12562 8014 12660 8112 ne
rect 12660 8014 13014 8112
tri 13014 8014 13112 8112 sw
tri 13112 8014 13210 8112 ne
rect 13210 8014 13564 8112
tri 13564 8014 13662 8112 sw
rect 14775 8014 15775 8662
rect -2525 8010 -88 8014
rect -2525 7890 -310 8010
rect -190 7926 -88 8010
tri -88 7926 0 8014 sw
tri 10 7926 98 8014 ne
rect 98 8010 462 8014
rect 98 7926 240 8010
rect -190 7890 0 7926
rect -2525 7886 0 7890
rect -2525 7238 -1525 7886
tri -412 7788 -314 7886 ne
rect -314 7838 0 7886
tri 0 7838 88 7926 sw
tri 98 7838 186 7926 ne
rect 186 7890 240 7926
rect 360 7926 462 8010
tri 462 7926 550 8014 sw
tri 560 7926 648 8014 ne
rect 648 8010 1012 8014
rect 648 7926 790 8010
rect 360 7890 550 7926
rect 186 7886 550 7890
tri 550 7886 590 7926 sw
tri 648 7886 688 7926 ne
rect 688 7890 790 7926
rect 910 7926 1012 8010
tri 1012 7926 1100 8014 sw
tri 1110 7926 1198 8014 ne
rect 1198 8010 1562 8014
rect 1198 7926 1340 8010
rect 910 7890 1100 7926
rect 688 7886 1100 7890
rect 186 7838 590 7886
rect -314 7788 88 7838
rect -1025 7700 -412 7788
tri -412 7700 -324 7788 sw
tri -314 7700 -226 7788 ne
rect -226 7758 88 7788
tri 88 7758 168 7838 sw
tri 186 7758 266 7838 ne
rect 266 7788 590 7838
tri 590 7788 688 7886 sw
tri 688 7788 786 7886 ne
rect 786 7838 1100 7886
tri 1100 7838 1188 7926 sw
tri 1198 7838 1286 7926 ne
rect 1286 7890 1340 7926
rect 1460 7926 1562 8010
tri 1562 7926 1650 8014 sw
tri 1660 7926 1748 8014 ne
rect 1748 8010 2112 8014
rect 1748 7926 1890 8010
rect 1460 7890 1650 7926
rect 1286 7886 1650 7890
tri 1650 7886 1690 7926 sw
tri 1748 7886 1788 7926 ne
rect 1788 7890 1890 7926
rect 2010 7926 2112 8010
tri 2112 7926 2200 8014 sw
tri 2210 7926 2298 8014 ne
rect 2298 8010 2662 8014
rect 2298 7926 2440 8010
rect 2010 7890 2200 7926
rect 1788 7886 2200 7890
rect 1286 7838 1690 7886
rect 786 7788 1188 7838
rect 266 7758 688 7788
rect -226 7700 168 7758
rect -1025 7660 -324 7700
tri -324 7660 -284 7700 sw
tri -226 7660 -186 7700 ne
rect -186 7660 168 7700
tri 168 7660 266 7758 sw
tri 266 7660 364 7758 ne
rect 364 7700 688 7758
tri 688 7700 776 7788 sw
tri 786 7700 874 7788 ne
rect 874 7758 1188 7788
tri 1188 7758 1268 7838 sw
tri 1286 7758 1366 7838 ne
rect 1366 7788 1690 7838
tri 1690 7788 1788 7886 sw
tri 1788 7788 1886 7886 ne
rect 1886 7838 2200 7886
tri 2200 7838 2288 7926 sw
tri 2298 7838 2386 7926 ne
rect 2386 7890 2440 7926
rect 2560 7926 2662 8010
tri 2662 7926 2750 8014 sw
tri 2760 7926 2848 8014 ne
rect 2848 8010 3212 8014
rect 2848 7926 2990 8010
rect 2560 7890 2750 7926
rect 2386 7886 2750 7890
tri 2750 7886 2790 7926 sw
tri 2848 7886 2888 7926 ne
rect 2888 7890 2990 7926
rect 3110 7926 3212 8010
tri 3212 7926 3300 8014 sw
tri 3310 7926 3398 8014 ne
rect 3398 8010 3762 8014
rect 3398 7926 3540 8010
rect 3110 7890 3300 7926
rect 2888 7886 3300 7890
rect 2386 7838 2790 7886
rect 1886 7788 2288 7838
rect 1366 7758 1788 7788
rect 874 7700 1268 7758
rect 364 7660 776 7700
tri 776 7660 816 7700 sw
tri 874 7660 914 7700 ne
rect 914 7660 1268 7700
tri 1268 7660 1366 7758 sw
tri 1366 7660 1464 7758 ne
rect 1464 7700 1788 7758
tri 1788 7700 1876 7788 sw
tri 1886 7700 1974 7788 ne
rect 1974 7758 2288 7788
tri 2288 7758 2368 7838 sw
tri 2386 7758 2466 7838 ne
rect 2466 7788 2790 7838
tri 2790 7788 2888 7886 sw
tri 2888 7788 2986 7886 ne
rect 2986 7838 3300 7886
tri 3300 7838 3388 7926 sw
tri 3398 7838 3486 7926 ne
rect 3486 7890 3540 7926
rect 3660 7926 3762 8010
tri 3762 7926 3850 8014 sw
tri 3860 7926 3948 8014 ne
rect 3948 8010 4312 8014
rect 3948 7926 4090 8010
rect 3660 7890 3850 7926
rect 3486 7886 3850 7890
tri 3850 7886 3890 7926 sw
tri 3948 7886 3988 7926 ne
rect 3988 7890 4090 7926
rect 4210 7926 4312 8010
tri 4312 7926 4400 8014 sw
tri 4410 7926 4498 8014 ne
rect 4498 8010 4862 8014
rect 4498 7926 4640 8010
rect 4210 7890 4400 7926
rect 3988 7886 4400 7890
rect 3486 7838 3890 7886
rect 2986 7788 3388 7838
rect 2466 7758 2888 7788
rect 1974 7700 2368 7758
rect 1464 7660 1876 7700
tri 1876 7660 1916 7700 sw
tri 1974 7660 2014 7700 ne
rect 2014 7660 2368 7700
tri 2368 7660 2466 7758 sw
tri 2466 7660 2564 7758 ne
rect 2564 7700 2888 7758
tri 2888 7700 2976 7788 sw
tri 2986 7700 3074 7788 ne
rect 3074 7758 3388 7788
tri 3388 7758 3468 7838 sw
tri 3486 7758 3566 7838 ne
rect 3566 7788 3890 7838
tri 3890 7788 3988 7886 sw
tri 3988 7788 4086 7886 ne
rect 4086 7838 4400 7886
tri 4400 7838 4488 7926 sw
tri 4498 7838 4586 7926 ne
rect 4586 7890 4640 7926
rect 4760 7926 4862 8010
tri 4862 7926 4950 8014 sw
tri 4960 7926 5048 8014 ne
rect 5048 8010 5412 8014
rect 5048 7926 5190 8010
rect 4760 7890 4950 7926
rect 4586 7886 4950 7890
tri 4950 7886 4990 7926 sw
tri 5048 7886 5088 7926 ne
rect 5088 7890 5190 7926
rect 5310 7926 5412 8010
tri 5412 7926 5500 8014 sw
tri 5510 7926 5598 8014 ne
rect 5598 8010 5962 8014
rect 5598 7926 5740 8010
rect 5310 7890 5500 7926
rect 5088 7886 5500 7890
rect 4586 7838 4990 7886
rect 4086 7788 4488 7838
rect 3566 7758 3988 7788
rect 3074 7700 3468 7758
rect 2564 7660 2976 7700
tri 2976 7660 3016 7700 sw
tri 3074 7660 3114 7700 ne
rect 3114 7660 3468 7700
tri 3468 7660 3566 7758 sw
tri 3566 7660 3664 7758 ne
rect 3664 7700 3988 7758
tri 3988 7700 4076 7788 sw
tri 4086 7700 4174 7788 ne
rect 4174 7758 4488 7788
tri 4488 7758 4568 7838 sw
tri 4586 7758 4666 7838 ne
rect 4666 7788 4990 7838
tri 4990 7788 5088 7886 sw
tri 5088 7788 5186 7886 ne
rect 5186 7838 5500 7886
tri 5500 7838 5588 7926 sw
tri 5598 7838 5686 7926 ne
rect 5686 7890 5740 7926
rect 5860 7926 5962 8010
tri 5962 7926 6050 8014 sw
tri 6060 7926 6148 8014 ne
rect 6148 8010 6512 8014
rect 6148 7926 6290 8010
rect 5860 7890 6050 7926
rect 5686 7886 6050 7890
tri 6050 7886 6090 7926 sw
tri 6148 7886 6188 7926 ne
rect 6188 7890 6290 7926
rect 6410 7926 6512 8010
tri 6512 7926 6600 8014 sw
tri 6610 7926 6698 8014 ne
rect 6698 8010 7062 8014
rect 6698 7926 6840 8010
rect 6410 7890 6600 7926
rect 6188 7886 6600 7890
rect 5686 7838 6090 7886
rect 5186 7788 5588 7838
rect 4666 7758 5088 7788
rect 4174 7700 4568 7758
rect 3664 7660 4076 7700
tri 4076 7660 4116 7700 sw
tri 4174 7660 4214 7700 ne
rect 4214 7660 4568 7700
tri 4568 7660 4666 7758 sw
tri 4666 7660 4764 7758 ne
rect 4764 7700 5088 7758
tri 5088 7700 5176 7788 sw
tri 5186 7700 5274 7788 ne
rect 5274 7758 5588 7788
tri 5588 7758 5668 7838 sw
tri 5686 7758 5766 7838 ne
rect 5766 7788 6090 7838
tri 6090 7788 6188 7886 sw
tri 6188 7788 6286 7886 ne
rect 6286 7838 6600 7886
tri 6600 7838 6688 7926 sw
tri 6698 7838 6786 7926 ne
rect 6786 7890 6840 7926
rect 6960 7926 7062 8010
tri 7062 7926 7150 8014 sw
tri 7160 7926 7248 8014 ne
rect 7248 8010 7612 8014
rect 7248 7926 7390 8010
rect 6960 7890 7150 7926
rect 6786 7886 7150 7890
tri 7150 7886 7190 7926 sw
tri 7248 7886 7288 7926 ne
rect 7288 7890 7390 7926
rect 7510 7926 7612 8010
tri 7612 7926 7700 8014 sw
tri 7710 7926 7798 8014 ne
rect 7798 8010 8162 8014
rect 7798 7926 7940 8010
rect 7510 7890 7700 7926
rect 7288 7886 7700 7890
rect 6786 7838 7190 7886
rect 6286 7788 6688 7838
rect 5766 7758 6188 7788
rect 5274 7700 5668 7758
rect 4764 7660 5176 7700
tri 5176 7660 5216 7700 sw
tri 5274 7660 5314 7700 ne
rect 5314 7660 5668 7700
tri 5668 7660 5766 7758 sw
tri 5766 7660 5864 7758 ne
rect 5864 7700 6188 7758
tri 6188 7700 6276 7788 sw
tri 6286 7700 6374 7788 ne
rect 6374 7758 6688 7788
tri 6688 7758 6768 7838 sw
tri 6786 7758 6866 7838 ne
rect 6866 7788 7190 7838
tri 7190 7788 7288 7886 sw
tri 7288 7788 7386 7886 ne
rect 7386 7838 7700 7886
tri 7700 7838 7788 7926 sw
tri 7798 7838 7886 7926 ne
rect 7886 7890 7940 7926
rect 8060 7926 8162 8010
tri 8162 7926 8250 8014 sw
tri 8260 7926 8348 8014 ne
rect 8348 8010 8712 8014
rect 8348 7926 8490 8010
rect 8060 7890 8250 7926
rect 7886 7886 8250 7890
tri 8250 7886 8290 7926 sw
tri 8348 7886 8388 7926 ne
rect 8388 7890 8490 7926
rect 8610 7926 8712 8010
tri 8712 7926 8800 8014 sw
tri 8810 7926 8898 8014 ne
rect 8898 8010 9262 8014
rect 8898 7926 9040 8010
rect 8610 7890 8800 7926
rect 8388 7886 8800 7890
rect 7886 7838 8290 7886
rect 7386 7788 7788 7838
rect 6866 7758 7288 7788
rect 6374 7700 6768 7758
rect 5864 7660 6276 7700
tri 6276 7660 6316 7700 sw
tri 6374 7660 6414 7700 ne
rect 6414 7660 6768 7700
tri 6768 7660 6866 7758 sw
tri 6866 7660 6964 7758 ne
rect 6964 7700 7288 7758
tri 7288 7700 7376 7788 sw
tri 7386 7700 7474 7788 ne
rect 7474 7758 7788 7788
tri 7788 7758 7868 7838 sw
tri 7886 7758 7966 7838 ne
rect 7966 7788 8290 7838
tri 8290 7788 8388 7886 sw
tri 8388 7788 8486 7886 ne
rect 8486 7838 8800 7886
tri 8800 7838 8888 7926 sw
tri 8898 7838 8986 7926 ne
rect 8986 7890 9040 7926
rect 9160 7926 9262 8010
tri 9262 7926 9350 8014 sw
tri 9360 7926 9448 8014 ne
rect 9448 8010 9812 8014
rect 9448 7926 9590 8010
rect 9160 7890 9350 7926
rect 8986 7886 9350 7890
tri 9350 7886 9390 7926 sw
tri 9448 7886 9488 7926 ne
rect 9488 7890 9590 7926
rect 9710 7926 9812 8010
tri 9812 7926 9900 8014 sw
tri 9910 7926 9998 8014 ne
rect 9998 8010 10362 8014
rect 9998 7926 10140 8010
rect 9710 7890 9900 7926
rect 9488 7886 9900 7890
rect 8986 7838 9390 7886
rect 8486 7788 8888 7838
rect 7966 7758 8388 7788
rect 7474 7700 7868 7758
rect 6964 7660 7376 7700
tri 7376 7660 7416 7700 sw
tri 7474 7660 7514 7700 ne
rect 7514 7660 7868 7700
tri 7868 7660 7966 7758 sw
tri 7966 7660 8064 7758 ne
rect 8064 7700 8388 7758
tri 8388 7700 8476 7788 sw
tri 8486 7700 8574 7788 ne
rect 8574 7758 8888 7788
tri 8888 7758 8968 7838 sw
tri 8986 7758 9066 7838 ne
rect 9066 7788 9390 7838
tri 9390 7788 9488 7886 sw
tri 9488 7788 9586 7886 ne
rect 9586 7838 9900 7886
tri 9900 7838 9988 7926 sw
tri 9998 7838 10086 7926 ne
rect 10086 7890 10140 7926
rect 10260 7926 10362 8010
tri 10362 7926 10450 8014 sw
tri 10460 7926 10548 8014 ne
rect 10548 8010 10912 8014
rect 10548 7926 10690 8010
rect 10260 7890 10450 7926
rect 10086 7886 10450 7890
tri 10450 7886 10490 7926 sw
tri 10548 7886 10588 7926 ne
rect 10588 7890 10690 7926
rect 10810 7926 10912 8010
tri 10912 7926 11000 8014 sw
tri 11010 7926 11098 8014 ne
rect 11098 8010 11462 8014
rect 11098 7926 11240 8010
rect 10810 7890 11000 7926
rect 10588 7886 11000 7890
rect 10086 7838 10490 7886
rect 9586 7788 9988 7838
rect 9066 7758 9488 7788
rect 8574 7700 8968 7758
rect 8064 7660 8476 7700
tri 8476 7660 8516 7700 sw
tri 8574 7660 8614 7700 ne
rect 8614 7660 8968 7700
tri 8968 7660 9066 7758 sw
tri 9066 7660 9164 7758 ne
rect 9164 7700 9488 7758
tri 9488 7700 9576 7788 sw
tri 9586 7700 9674 7788 ne
rect 9674 7758 9988 7788
tri 9988 7758 10068 7838 sw
tri 10086 7758 10166 7838 ne
rect 10166 7788 10490 7838
tri 10490 7788 10588 7886 sw
tri 10588 7788 10686 7886 ne
rect 10686 7838 11000 7886
tri 11000 7838 11088 7926 sw
tri 11098 7838 11186 7926 ne
rect 11186 7890 11240 7926
rect 11360 7926 11462 8010
tri 11462 7926 11550 8014 sw
tri 11560 7926 11648 8014 ne
rect 11648 8010 12012 8014
rect 11648 7926 11790 8010
rect 11360 7890 11550 7926
rect 11186 7886 11550 7890
tri 11550 7886 11590 7926 sw
tri 11648 7886 11688 7926 ne
rect 11688 7890 11790 7926
rect 11910 7926 12012 8010
tri 12012 7926 12100 8014 sw
tri 12110 7926 12198 8014 ne
rect 12198 8010 12562 8014
rect 12198 7926 12340 8010
rect 11910 7890 12100 7926
rect 11688 7886 12100 7890
rect 11186 7838 11590 7886
rect 10686 7788 11088 7838
rect 10166 7758 10588 7788
rect 9674 7700 10068 7758
rect 9164 7660 9576 7700
tri 9576 7660 9616 7700 sw
tri 9674 7660 9714 7700 ne
rect 9714 7660 10068 7700
tri 10068 7660 10166 7758 sw
tri 10166 7660 10264 7758 ne
rect 10264 7700 10588 7758
tri 10588 7700 10676 7788 sw
tri 10686 7700 10774 7788 ne
rect 10774 7758 11088 7788
tri 11088 7758 11168 7838 sw
tri 11186 7758 11266 7838 ne
rect 11266 7788 11590 7838
tri 11590 7788 11688 7886 sw
tri 11688 7788 11786 7886 ne
rect 11786 7838 12100 7886
tri 12100 7838 12188 7926 sw
tri 12198 7838 12286 7926 ne
rect 12286 7890 12340 7926
rect 12460 7926 12562 8010
tri 12562 7926 12650 8014 sw
tri 12660 7926 12748 8014 ne
rect 12748 8010 13112 8014
rect 12748 7926 12890 8010
rect 12460 7890 12650 7926
rect 12286 7886 12650 7890
tri 12650 7886 12690 7926 sw
tri 12748 7886 12788 7926 ne
rect 12788 7890 12890 7926
rect 13010 7926 13112 8010
tri 13112 7926 13200 8014 sw
tri 13210 7926 13298 8014 ne
rect 13298 8010 15775 8014
rect 13298 7926 13440 8010
rect 13010 7890 13200 7926
rect 12788 7886 13200 7890
rect 12286 7838 12690 7886
rect 11786 7788 12188 7838
rect 11266 7758 11688 7788
rect 10774 7700 11168 7758
rect 10264 7660 10676 7700
tri 10676 7660 10716 7700 sw
tri 10774 7660 10814 7700 ne
rect 10814 7660 11168 7700
tri 11168 7660 11266 7758 sw
tri 11266 7660 11364 7758 ne
rect 11364 7700 11688 7758
tri 11688 7700 11776 7788 sw
tri 11786 7700 11874 7788 ne
rect 11874 7758 12188 7788
tri 12188 7758 12268 7838 sw
tri 12286 7758 12366 7838 ne
rect 12366 7788 12690 7838
tri 12690 7788 12788 7886 sw
tri 12788 7788 12886 7886 ne
rect 12886 7838 13200 7886
tri 13200 7838 13288 7926 sw
tri 13298 7838 13386 7926 ne
rect 13386 7890 13440 7926
rect 13560 7890 15775 8010
rect 13386 7838 15775 7890
rect 12886 7788 13288 7838
rect 12366 7758 12788 7788
rect 11874 7700 12268 7758
rect 11364 7660 11776 7700
tri 11776 7660 11816 7700 sw
tri 11874 7660 11914 7700 ne
rect 11914 7660 12268 7700
tri 12268 7660 12366 7758 sw
tri 12366 7660 12464 7758 ne
rect 12464 7700 12788 7758
tri 12788 7700 12876 7788 sw
tri 12886 7700 12974 7788 ne
rect 12974 7758 13288 7788
tri 13288 7758 13368 7838 sw
tri 13386 7758 13466 7838 ne
rect 13466 7758 14075 7838
rect 12974 7700 13368 7758
rect 12464 7660 12876 7700
tri 12876 7660 12916 7700 sw
tri 12974 7660 13014 7700 ne
rect 13014 7660 13368 7700
tri 13368 7660 13466 7758 sw
tri 13466 7660 13564 7758 ne
rect 13564 7738 14075 7758
rect 14175 7738 15775 7838
rect 13564 7660 15775 7738
rect -1025 7612 -284 7660
rect -1025 7512 -925 7612
rect -825 7562 -284 7612
tri -284 7562 -186 7660 sw
tri -186 7562 -88 7660 ne
rect -88 7562 266 7660
tri 266 7562 364 7660 sw
tri 364 7562 462 7660 ne
rect 462 7562 816 7660
tri 816 7562 914 7660 sw
tri 914 7562 1012 7660 ne
rect 1012 7562 1366 7660
tri 1366 7562 1464 7660 sw
tri 1464 7562 1562 7660 ne
rect 1562 7562 1916 7660
tri 1916 7562 2014 7660 sw
tri 2014 7562 2112 7660 ne
rect 2112 7562 2466 7660
tri 2466 7562 2564 7660 sw
tri 2564 7562 2662 7660 ne
rect 2662 7562 3016 7660
tri 3016 7562 3114 7660 sw
tri 3114 7562 3212 7660 ne
rect 3212 7562 3566 7660
tri 3566 7562 3664 7660 sw
tri 3664 7562 3762 7660 ne
rect 3762 7562 4116 7660
tri 4116 7562 4214 7660 sw
tri 4214 7562 4312 7660 ne
rect 4312 7562 4666 7660
tri 4666 7562 4764 7660 sw
tri 4764 7562 4862 7660 ne
rect 4862 7562 5216 7660
tri 5216 7562 5314 7660 sw
tri 5314 7562 5412 7660 ne
rect 5412 7562 5766 7660
tri 5766 7562 5864 7660 sw
tri 5864 7562 5962 7660 ne
rect 5962 7562 6316 7660
tri 6316 7562 6414 7660 sw
tri 6414 7562 6512 7660 ne
rect 6512 7562 6866 7660
tri 6866 7562 6964 7660 sw
tri 6964 7562 7062 7660 ne
rect 7062 7562 7416 7660
tri 7416 7562 7514 7660 sw
tri 7514 7562 7612 7660 ne
rect 7612 7562 7966 7660
tri 7966 7562 8064 7660 sw
tri 8064 7562 8162 7660 ne
rect 8162 7562 8516 7660
tri 8516 7562 8614 7660 sw
tri 8614 7562 8712 7660 ne
rect 8712 7562 9066 7660
tri 9066 7562 9164 7660 sw
tri 9164 7562 9262 7660 ne
rect 9262 7562 9616 7660
tri 9616 7562 9714 7660 sw
tri 9714 7562 9812 7660 ne
rect 9812 7562 10166 7660
tri 10166 7562 10264 7660 sw
tri 10264 7562 10362 7660 ne
rect 10362 7562 10716 7660
tri 10716 7562 10814 7660 sw
tri 10814 7562 10912 7660 ne
rect 10912 7562 11266 7660
tri 11266 7562 11364 7660 sw
tri 11364 7562 11462 7660 ne
rect 11462 7562 11816 7660
tri 11816 7562 11914 7660 sw
tri 11914 7562 12012 7660 ne
rect 12012 7562 12366 7660
tri 12366 7562 12464 7660 sw
tri 12464 7562 12562 7660 ne
rect 12562 7562 12916 7660
tri 12916 7562 13014 7660 sw
tri 13014 7562 13112 7660 ne
rect 13112 7562 13466 7660
tri 13466 7562 13564 7660 sw
tri 13564 7562 13662 7660 ne
rect 13662 7562 15775 7660
rect -825 7512 -186 7562
rect -1025 7464 -186 7512
tri -186 7464 -88 7562 sw
tri -88 7464 10 7562 ne
rect 10 7464 364 7562
tri 364 7464 462 7562 sw
tri 462 7464 560 7562 ne
rect 560 7464 914 7562
tri 914 7464 1012 7562 sw
tri 1012 7464 1110 7562 ne
rect 1110 7464 1464 7562
tri 1464 7464 1562 7562 sw
tri 1562 7464 1660 7562 ne
rect 1660 7464 2014 7562
tri 2014 7464 2112 7562 sw
tri 2112 7464 2210 7562 ne
rect 2210 7464 2564 7562
tri 2564 7464 2662 7562 sw
tri 2662 7464 2760 7562 ne
rect 2760 7464 3114 7562
tri 3114 7464 3212 7562 sw
tri 3212 7464 3310 7562 ne
rect 3310 7464 3664 7562
tri 3664 7464 3762 7562 sw
tri 3762 7464 3860 7562 ne
rect 3860 7464 4214 7562
tri 4214 7464 4312 7562 sw
tri 4312 7464 4410 7562 ne
rect 4410 7464 4764 7562
tri 4764 7464 4862 7562 sw
tri 4862 7464 4960 7562 ne
rect 4960 7464 5314 7562
tri 5314 7464 5412 7562 sw
tri 5412 7464 5510 7562 ne
rect 5510 7464 5864 7562
tri 5864 7464 5962 7562 sw
tri 5962 7464 6060 7562 ne
rect 6060 7464 6414 7562
tri 6414 7464 6512 7562 sw
tri 6512 7464 6610 7562 ne
rect 6610 7464 6964 7562
tri 6964 7464 7062 7562 sw
tri 7062 7464 7160 7562 ne
rect 7160 7464 7514 7562
tri 7514 7464 7612 7562 sw
tri 7612 7464 7710 7562 ne
rect 7710 7464 8064 7562
tri 8064 7464 8162 7562 sw
tri 8162 7464 8260 7562 ne
rect 8260 7464 8614 7562
tri 8614 7464 8712 7562 sw
tri 8712 7464 8810 7562 ne
rect 8810 7464 9164 7562
tri 9164 7464 9262 7562 sw
tri 9262 7464 9360 7562 ne
rect 9360 7464 9714 7562
tri 9714 7464 9812 7562 sw
tri 9812 7464 9910 7562 ne
rect 9910 7464 10264 7562
tri 10264 7464 10362 7562 sw
tri 10362 7464 10460 7562 ne
rect 10460 7464 10814 7562
tri 10814 7464 10912 7562 sw
tri 10912 7464 11010 7562 ne
rect 11010 7464 11364 7562
tri 11364 7464 11462 7562 sw
tri 11462 7464 11560 7562 ne
rect 11560 7464 11914 7562
tri 11914 7464 12012 7562 sw
tri 12012 7464 12110 7562 ne
rect 12110 7464 12464 7562
tri 12464 7464 12562 7562 sw
tri 12562 7464 12660 7562 ne
rect 12660 7464 13014 7562
tri 13014 7464 13112 7562 sw
tri 13112 7464 13210 7562 ne
rect 13210 7464 13564 7562
tri 13564 7464 13662 7562 sw
rect -1025 7460 -88 7464
rect -1025 7340 -310 7460
rect -190 7376 -88 7460
tri -88 7376 0 7464 sw
tri 10 7376 98 7464 ne
rect 98 7460 462 7464
rect 98 7376 240 7460
rect -190 7340 0 7376
rect -1025 7336 0 7340
tri 0 7336 40 7376 sw
tri 98 7336 138 7376 ne
rect 138 7340 240 7376
rect 360 7376 462 7460
tri 462 7376 550 7464 sw
tri 560 7376 648 7464 ne
rect 648 7460 1012 7464
rect 648 7376 790 7460
rect 360 7340 550 7376
rect 138 7336 550 7340
tri -412 7238 -314 7336 ne
rect -314 7238 40 7336
tri 40 7238 138 7336 sw
tri 138 7238 236 7336 ne
rect 236 7288 550 7336
tri 550 7288 638 7376 sw
tri 648 7288 736 7376 ne
rect 736 7340 790 7376
rect 910 7376 1012 7460
tri 1012 7376 1100 7464 sw
tri 1110 7376 1198 7464 ne
rect 1198 7460 1562 7464
rect 1198 7376 1340 7460
rect 910 7340 1100 7376
rect 736 7336 1100 7340
tri 1100 7336 1140 7376 sw
tri 1198 7336 1238 7376 ne
rect 1238 7340 1340 7376
rect 1460 7376 1562 7460
tri 1562 7376 1650 7464 sw
tri 1660 7376 1748 7464 ne
rect 1748 7460 2112 7464
rect 1748 7376 1890 7460
rect 1460 7340 1650 7376
rect 1238 7336 1650 7340
rect 736 7288 1140 7336
rect 236 7238 638 7288
rect -2525 7150 -412 7238
tri -412 7150 -324 7238 sw
tri -314 7150 -226 7238 ne
rect -226 7150 138 7238
tri 138 7150 226 7238 sw
tri 236 7150 324 7238 ne
rect 324 7208 638 7238
tri 638 7208 718 7288 sw
tri 736 7208 816 7288 ne
rect 816 7238 1140 7288
tri 1140 7238 1238 7336 sw
tri 1238 7238 1336 7336 ne
rect 1336 7288 1650 7336
tri 1650 7288 1738 7376 sw
tri 1748 7288 1836 7376 ne
rect 1836 7340 1890 7376
rect 2010 7376 2112 7460
tri 2112 7376 2200 7464 sw
tri 2210 7376 2298 7464 ne
rect 2298 7460 2662 7464
rect 2298 7376 2440 7460
rect 2010 7340 2200 7376
rect 1836 7336 2200 7340
tri 2200 7336 2240 7376 sw
tri 2298 7336 2338 7376 ne
rect 2338 7340 2440 7376
rect 2560 7376 2662 7460
tri 2662 7376 2750 7464 sw
tri 2760 7376 2848 7464 ne
rect 2848 7460 3212 7464
rect 2848 7376 2990 7460
rect 2560 7340 2750 7376
rect 2338 7336 2750 7340
rect 1836 7288 2240 7336
rect 1336 7238 1738 7288
rect 816 7208 1238 7238
rect 324 7150 718 7208
rect -2525 7110 -324 7150
tri -324 7110 -284 7150 sw
tri -226 7110 -186 7150 ne
rect -186 7110 226 7150
tri 226 7110 266 7150 sw
tri 324 7110 364 7150 ne
rect 364 7110 718 7150
tri 718 7110 816 7208 sw
tri 816 7110 914 7208 ne
rect 914 7150 1238 7208
tri 1238 7150 1326 7238 sw
tri 1336 7150 1424 7238 ne
rect 1424 7208 1738 7238
tri 1738 7208 1818 7288 sw
tri 1836 7208 1916 7288 ne
rect 1916 7238 2240 7288
tri 2240 7238 2338 7336 sw
tri 2338 7238 2436 7336 ne
rect 2436 7288 2750 7336
tri 2750 7288 2838 7376 sw
tri 2848 7288 2936 7376 ne
rect 2936 7340 2990 7376
rect 3110 7376 3212 7460
tri 3212 7376 3300 7464 sw
tri 3310 7376 3398 7464 ne
rect 3398 7460 3762 7464
rect 3398 7376 3540 7460
rect 3110 7340 3300 7376
rect 2936 7336 3300 7340
tri 3300 7336 3340 7376 sw
tri 3398 7336 3438 7376 ne
rect 3438 7340 3540 7376
rect 3660 7376 3762 7460
tri 3762 7376 3850 7464 sw
tri 3860 7376 3948 7464 ne
rect 3948 7460 4312 7464
rect 3948 7376 4090 7460
rect 3660 7340 3850 7376
rect 3438 7336 3850 7340
rect 2936 7288 3340 7336
rect 2436 7238 2838 7288
rect 1916 7208 2338 7238
rect 1424 7150 1818 7208
rect 914 7110 1326 7150
tri 1326 7110 1366 7150 sw
tri 1424 7110 1464 7150 ne
rect 1464 7110 1818 7150
tri 1818 7110 1916 7208 sw
tri 1916 7110 2014 7208 ne
rect 2014 7150 2338 7208
tri 2338 7150 2426 7238 sw
tri 2436 7150 2524 7238 ne
rect 2524 7208 2838 7238
tri 2838 7208 2918 7288 sw
tri 2936 7208 3016 7288 ne
rect 3016 7238 3340 7288
tri 3340 7238 3438 7336 sw
tri 3438 7238 3536 7336 ne
rect 3536 7288 3850 7336
tri 3850 7288 3938 7376 sw
tri 3948 7288 4036 7376 ne
rect 4036 7340 4090 7376
rect 4210 7376 4312 7460
tri 4312 7376 4400 7464 sw
tri 4410 7376 4498 7464 ne
rect 4498 7460 4862 7464
rect 4498 7376 4640 7460
rect 4210 7340 4400 7376
rect 4036 7336 4400 7340
tri 4400 7336 4440 7376 sw
tri 4498 7336 4538 7376 ne
rect 4538 7340 4640 7376
rect 4760 7376 4862 7460
tri 4862 7376 4950 7464 sw
tri 4960 7376 5048 7464 ne
rect 5048 7460 5412 7464
rect 5048 7376 5190 7460
rect 4760 7340 4950 7376
rect 4538 7336 4950 7340
rect 4036 7288 4440 7336
rect 3536 7238 3938 7288
rect 3016 7208 3438 7238
rect 2524 7150 2918 7208
rect 2014 7110 2426 7150
tri 2426 7110 2466 7150 sw
tri 2524 7110 2564 7150 ne
rect 2564 7110 2918 7150
tri 2918 7110 3016 7208 sw
tri 3016 7110 3114 7208 ne
rect 3114 7150 3438 7208
tri 3438 7150 3526 7238 sw
tri 3536 7150 3624 7238 ne
rect 3624 7208 3938 7238
tri 3938 7208 4018 7288 sw
tri 4036 7208 4116 7288 ne
rect 4116 7238 4440 7288
tri 4440 7238 4538 7336 sw
tri 4538 7238 4636 7336 ne
rect 4636 7288 4950 7336
tri 4950 7288 5038 7376 sw
tri 5048 7288 5136 7376 ne
rect 5136 7340 5190 7376
rect 5310 7376 5412 7460
tri 5412 7376 5500 7464 sw
tri 5510 7376 5598 7464 ne
rect 5598 7460 5962 7464
rect 5598 7376 5740 7460
rect 5310 7340 5500 7376
rect 5136 7336 5500 7340
tri 5500 7336 5540 7376 sw
tri 5598 7336 5638 7376 ne
rect 5638 7340 5740 7376
rect 5860 7376 5962 7460
tri 5962 7376 6050 7464 sw
tri 6060 7376 6148 7464 ne
rect 6148 7460 6512 7464
rect 6148 7376 6290 7460
rect 5860 7340 6050 7376
rect 5638 7336 6050 7340
rect 5136 7288 5540 7336
rect 4636 7238 5038 7288
rect 4116 7208 4538 7238
rect 3624 7150 4018 7208
rect 3114 7110 3526 7150
tri 3526 7110 3566 7150 sw
tri 3624 7110 3664 7150 ne
rect 3664 7110 4018 7150
tri 4018 7110 4116 7208 sw
tri 4116 7110 4214 7208 ne
rect 4214 7150 4538 7208
tri 4538 7150 4626 7238 sw
tri 4636 7150 4724 7238 ne
rect 4724 7208 5038 7238
tri 5038 7208 5118 7288 sw
tri 5136 7208 5216 7288 ne
rect 5216 7238 5540 7288
tri 5540 7238 5638 7336 sw
tri 5638 7238 5736 7336 ne
rect 5736 7288 6050 7336
tri 6050 7288 6138 7376 sw
tri 6148 7288 6236 7376 ne
rect 6236 7340 6290 7376
rect 6410 7376 6512 7460
tri 6512 7376 6600 7464 sw
tri 6610 7376 6698 7464 ne
rect 6698 7460 7062 7464
rect 6698 7376 6840 7460
rect 6410 7340 6600 7376
rect 6236 7336 6600 7340
tri 6600 7336 6640 7376 sw
tri 6698 7336 6738 7376 ne
rect 6738 7340 6840 7376
rect 6960 7376 7062 7460
tri 7062 7376 7150 7464 sw
tri 7160 7376 7248 7464 ne
rect 7248 7460 7612 7464
rect 7248 7376 7390 7460
rect 6960 7340 7150 7376
rect 6738 7336 7150 7340
rect 6236 7288 6640 7336
rect 5736 7238 6138 7288
rect 5216 7208 5638 7238
rect 4724 7150 5118 7208
rect 4214 7110 4626 7150
tri 4626 7110 4666 7150 sw
tri 4724 7110 4764 7150 ne
rect 4764 7110 5118 7150
tri 5118 7110 5216 7208 sw
tri 5216 7110 5314 7208 ne
rect 5314 7150 5638 7208
tri 5638 7150 5726 7238 sw
tri 5736 7150 5824 7238 ne
rect 5824 7208 6138 7238
tri 6138 7208 6218 7288 sw
tri 6236 7208 6316 7288 ne
rect 6316 7238 6640 7288
tri 6640 7238 6738 7336 sw
tri 6738 7238 6836 7336 ne
rect 6836 7288 7150 7336
tri 7150 7288 7238 7376 sw
tri 7248 7288 7336 7376 ne
rect 7336 7340 7390 7376
rect 7510 7376 7612 7460
tri 7612 7376 7700 7464 sw
tri 7710 7376 7798 7464 ne
rect 7798 7460 8162 7464
rect 7798 7376 7940 7460
rect 7510 7340 7700 7376
rect 7336 7336 7700 7340
tri 7700 7336 7740 7376 sw
tri 7798 7336 7838 7376 ne
rect 7838 7340 7940 7376
rect 8060 7376 8162 7460
tri 8162 7376 8250 7464 sw
tri 8260 7376 8348 7464 ne
rect 8348 7460 8712 7464
rect 8348 7376 8490 7460
rect 8060 7340 8250 7376
rect 7838 7336 8250 7340
rect 7336 7288 7740 7336
rect 6836 7238 7238 7288
rect 6316 7208 6738 7238
rect 5824 7150 6218 7208
rect 5314 7110 5726 7150
tri 5726 7110 5766 7150 sw
tri 5824 7110 5864 7150 ne
rect 5864 7110 6218 7150
tri 6218 7110 6316 7208 sw
tri 6316 7110 6414 7208 ne
rect 6414 7150 6738 7208
tri 6738 7150 6826 7238 sw
tri 6836 7150 6924 7238 ne
rect 6924 7208 7238 7238
tri 7238 7208 7318 7288 sw
tri 7336 7208 7416 7288 ne
rect 7416 7238 7740 7288
tri 7740 7238 7838 7336 sw
tri 7838 7238 7936 7336 ne
rect 7936 7288 8250 7336
tri 8250 7288 8338 7376 sw
tri 8348 7288 8436 7376 ne
rect 8436 7340 8490 7376
rect 8610 7376 8712 7460
tri 8712 7376 8800 7464 sw
tri 8810 7376 8898 7464 ne
rect 8898 7460 9262 7464
rect 8898 7376 9040 7460
rect 8610 7340 8800 7376
rect 8436 7336 8800 7340
tri 8800 7336 8840 7376 sw
tri 8898 7336 8938 7376 ne
rect 8938 7340 9040 7376
rect 9160 7376 9262 7460
tri 9262 7376 9350 7464 sw
tri 9360 7376 9448 7464 ne
rect 9448 7460 9812 7464
rect 9448 7376 9590 7460
rect 9160 7340 9350 7376
rect 8938 7336 9350 7340
rect 8436 7288 8840 7336
rect 7936 7238 8338 7288
rect 7416 7208 7838 7238
rect 6924 7150 7318 7208
rect 6414 7110 6826 7150
tri 6826 7110 6866 7150 sw
tri 6924 7110 6964 7150 ne
rect 6964 7110 7318 7150
tri 7318 7110 7416 7208 sw
tri 7416 7110 7514 7208 ne
rect 7514 7150 7838 7208
tri 7838 7150 7926 7238 sw
tri 7936 7150 8024 7238 ne
rect 8024 7208 8338 7238
tri 8338 7208 8418 7288 sw
tri 8436 7208 8516 7288 ne
rect 8516 7238 8840 7288
tri 8840 7238 8938 7336 sw
tri 8938 7238 9036 7336 ne
rect 9036 7288 9350 7336
tri 9350 7288 9438 7376 sw
tri 9448 7288 9536 7376 ne
rect 9536 7340 9590 7376
rect 9710 7376 9812 7460
tri 9812 7376 9900 7464 sw
tri 9910 7376 9998 7464 ne
rect 9998 7460 10362 7464
rect 9998 7376 10140 7460
rect 9710 7340 9900 7376
rect 9536 7336 9900 7340
tri 9900 7336 9940 7376 sw
tri 9998 7336 10038 7376 ne
rect 10038 7340 10140 7376
rect 10260 7376 10362 7460
tri 10362 7376 10450 7464 sw
tri 10460 7376 10548 7464 ne
rect 10548 7460 10912 7464
rect 10548 7376 10690 7460
rect 10260 7340 10450 7376
rect 10038 7336 10450 7340
rect 9536 7288 9940 7336
rect 9036 7238 9438 7288
rect 8516 7208 8938 7238
rect 8024 7150 8418 7208
rect 7514 7110 7926 7150
tri 7926 7110 7966 7150 sw
tri 8024 7110 8064 7150 ne
rect 8064 7110 8418 7150
tri 8418 7110 8516 7208 sw
tri 8516 7110 8614 7208 ne
rect 8614 7150 8938 7208
tri 8938 7150 9026 7238 sw
tri 9036 7150 9124 7238 ne
rect 9124 7208 9438 7238
tri 9438 7208 9518 7288 sw
tri 9536 7208 9616 7288 ne
rect 9616 7238 9940 7288
tri 9940 7238 10038 7336 sw
tri 10038 7238 10136 7336 ne
rect 10136 7288 10450 7336
tri 10450 7288 10538 7376 sw
tri 10548 7288 10636 7376 ne
rect 10636 7340 10690 7376
rect 10810 7376 10912 7460
tri 10912 7376 11000 7464 sw
tri 11010 7376 11098 7464 ne
rect 11098 7460 11462 7464
rect 11098 7376 11240 7460
rect 10810 7340 11000 7376
rect 10636 7336 11000 7340
tri 11000 7336 11040 7376 sw
tri 11098 7336 11138 7376 ne
rect 11138 7340 11240 7376
rect 11360 7376 11462 7460
tri 11462 7376 11550 7464 sw
tri 11560 7376 11648 7464 ne
rect 11648 7460 12012 7464
rect 11648 7376 11790 7460
rect 11360 7340 11550 7376
rect 11138 7336 11550 7340
rect 10636 7288 11040 7336
rect 10136 7238 10538 7288
rect 9616 7208 10038 7238
rect 9124 7150 9518 7208
rect 8614 7110 9026 7150
tri 9026 7110 9066 7150 sw
tri 9124 7110 9164 7150 ne
rect 9164 7110 9518 7150
tri 9518 7110 9616 7208 sw
tri 9616 7110 9714 7208 ne
rect 9714 7150 10038 7208
tri 10038 7150 10126 7238 sw
tri 10136 7150 10224 7238 ne
rect 10224 7208 10538 7238
tri 10538 7208 10618 7288 sw
tri 10636 7208 10716 7288 ne
rect 10716 7238 11040 7288
tri 11040 7238 11138 7336 sw
tri 11138 7238 11236 7336 ne
rect 11236 7288 11550 7336
tri 11550 7288 11638 7376 sw
tri 11648 7288 11736 7376 ne
rect 11736 7340 11790 7376
rect 11910 7376 12012 7460
tri 12012 7376 12100 7464 sw
tri 12110 7376 12198 7464 ne
rect 12198 7460 12562 7464
rect 12198 7376 12340 7460
rect 11910 7340 12100 7376
rect 11736 7336 12100 7340
tri 12100 7336 12140 7376 sw
tri 12198 7336 12238 7376 ne
rect 12238 7340 12340 7376
rect 12460 7376 12562 7460
tri 12562 7376 12650 7464 sw
tri 12660 7376 12748 7464 ne
rect 12748 7460 13112 7464
rect 12748 7376 12890 7460
rect 12460 7340 12650 7376
rect 12238 7336 12650 7340
rect 11736 7288 12140 7336
rect 11236 7238 11638 7288
rect 10716 7208 11138 7238
rect 10224 7150 10618 7208
rect 9714 7110 10126 7150
tri 10126 7110 10166 7150 sw
tri 10224 7110 10264 7150 ne
rect 10264 7110 10618 7150
tri 10618 7110 10716 7208 sw
tri 10716 7110 10814 7208 ne
rect 10814 7150 11138 7208
tri 11138 7150 11226 7238 sw
tri 11236 7150 11324 7238 ne
rect 11324 7208 11638 7238
tri 11638 7208 11718 7288 sw
tri 11736 7208 11816 7288 ne
rect 11816 7238 12140 7288
tri 12140 7238 12238 7336 sw
tri 12238 7238 12336 7336 ne
rect 12336 7288 12650 7336
tri 12650 7288 12738 7376 sw
tri 12748 7288 12836 7376 ne
rect 12836 7340 12890 7376
rect 13010 7376 13112 7460
tri 13112 7376 13200 7464 sw
tri 13210 7376 13298 7464 ne
rect 13298 7460 14275 7464
rect 13298 7376 13440 7460
rect 13010 7340 13200 7376
rect 12836 7336 13200 7340
tri 13200 7336 13240 7376 sw
tri 13298 7336 13338 7376 ne
rect 13338 7340 13440 7376
rect 13560 7340 14275 7460
rect 13338 7336 14275 7340
rect 12836 7288 13240 7336
rect 12336 7238 12738 7288
rect 11816 7208 12238 7238
rect 11324 7150 11718 7208
rect 10814 7110 11226 7150
tri 11226 7110 11266 7150 sw
tri 11324 7110 11364 7150 ne
rect 11364 7110 11718 7150
tri 11718 7110 11816 7208 sw
tri 11816 7110 11914 7208 ne
rect 11914 7150 12238 7208
tri 12238 7150 12326 7238 sw
tri 12336 7150 12424 7238 ne
rect 12424 7208 12738 7238
tri 12738 7208 12818 7288 sw
tri 12836 7208 12916 7288 ne
rect 12916 7238 13240 7288
tri 13240 7238 13338 7336 sw
tri 13338 7238 13436 7336 ne
rect 13436 7238 14275 7336
rect 12916 7208 13338 7238
rect 12424 7150 12818 7208
rect 11914 7110 12326 7150
tri 12326 7110 12366 7150 sw
tri 12424 7110 12464 7150 ne
rect 12464 7110 12818 7150
tri 12818 7110 12916 7208 sw
tri 12916 7110 13014 7208 ne
rect 13014 7150 13338 7208
tri 13338 7150 13426 7238 sw
tri 13436 7150 13524 7238 ne
rect 13524 7150 14275 7238
rect 13014 7110 13426 7150
tri 13426 7110 13466 7150 sw
tri 13524 7110 13564 7150 ne
rect 13564 7110 14275 7150
rect -2525 7012 -284 7110
tri -284 7012 -186 7110 sw
tri -186 7012 -88 7110 ne
rect -88 7012 266 7110
tri 266 7012 364 7110 sw
tri 364 7012 462 7110 ne
rect 462 7012 816 7110
tri 816 7012 914 7110 sw
tri 914 7012 1012 7110 ne
rect 1012 7012 1366 7110
tri 1366 7012 1464 7110 sw
tri 1464 7012 1562 7110 ne
rect 1562 7012 1916 7110
tri 1916 7012 2014 7110 sw
tri 2014 7012 2112 7110 ne
rect 2112 7012 2466 7110
tri 2466 7012 2564 7110 sw
tri 2564 7012 2662 7110 ne
rect 2662 7012 3016 7110
tri 3016 7012 3114 7110 sw
tri 3114 7012 3212 7110 ne
rect 3212 7012 3566 7110
tri 3566 7012 3664 7110 sw
tri 3664 7012 3762 7110 ne
rect 3762 7012 4116 7110
tri 4116 7012 4214 7110 sw
tri 4214 7012 4312 7110 ne
rect 4312 7012 4666 7110
tri 4666 7012 4764 7110 sw
tri 4764 7012 4862 7110 ne
rect 4862 7012 5216 7110
tri 5216 7012 5314 7110 sw
tri 5314 7012 5412 7110 ne
rect 5412 7012 5766 7110
tri 5766 7012 5864 7110 sw
tri 5864 7012 5962 7110 ne
rect 5962 7012 6316 7110
tri 6316 7012 6414 7110 sw
tri 6414 7012 6512 7110 ne
rect 6512 7012 6866 7110
tri 6866 7012 6964 7110 sw
tri 6964 7012 7062 7110 ne
rect 7062 7012 7416 7110
tri 7416 7012 7514 7110 sw
tri 7514 7012 7612 7110 ne
rect 7612 7012 7966 7110
tri 7966 7012 8064 7110 sw
tri 8064 7012 8162 7110 ne
rect 8162 7012 8516 7110
tri 8516 7012 8614 7110 sw
tri 8614 7012 8712 7110 ne
rect 8712 7012 9066 7110
tri 9066 7012 9164 7110 sw
tri 9164 7012 9262 7110 ne
rect 9262 7012 9616 7110
tri 9616 7012 9714 7110 sw
tri 9714 7012 9812 7110 ne
rect 9812 7012 10166 7110
tri 10166 7012 10264 7110 sw
tri 10264 7012 10362 7110 ne
rect 10362 7012 10716 7110
tri 10716 7012 10814 7110 sw
tri 10814 7012 10912 7110 ne
rect 10912 7012 11266 7110
tri 11266 7012 11364 7110 sw
tri 11364 7012 11462 7110 ne
rect 11462 7012 11816 7110
tri 11816 7012 11914 7110 sw
tri 11914 7012 12012 7110 ne
rect 12012 7012 12366 7110
tri 12366 7012 12464 7110 sw
tri 12464 7012 12562 7110 ne
rect 12562 7012 12916 7110
tri 12916 7012 13014 7110 sw
tri 13014 7012 13112 7110 ne
rect 13112 7012 13466 7110
tri 13466 7012 13564 7110 sw
tri 13564 7012 13662 7110 ne
rect 13662 7012 14275 7110
rect -2525 6914 -186 7012
tri -186 6914 -88 7012 sw
tri -88 6914 10 7012 ne
rect 10 6914 364 7012
tri 364 6914 462 7012 sw
tri 462 6914 560 7012 ne
rect 560 6914 914 7012
tri 914 6914 1012 7012 sw
tri 1012 6914 1110 7012 ne
rect 1110 6914 1464 7012
tri 1464 6914 1562 7012 sw
tri 1562 6914 1660 7012 ne
rect 1660 6914 2014 7012
tri 2014 6914 2112 7012 sw
tri 2112 6914 2210 7012 ne
rect 2210 6914 2564 7012
tri 2564 6914 2662 7012 sw
tri 2662 6914 2760 7012 ne
rect 2760 6914 3114 7012
tri 3114 6914 3212 7012 sw
tri 3212 6914 3310 7012 ne
rect 3310 6914 3664 7012
tri 3664 6914 3762 7012 sw
tri 3762 6914 3860 7012 ne
rect 3860 6914 4214 7012
tri 4214 6914 4312 7012 sw
tri 4312 6914 4410 7012 ne
rect 4410 6914 4764 7012
tri 4764 6914 4862 7012 sw
tri 4862 6914 4960 7012 ne
rect 4960 6914 5314 7012
tri 5314 6914 5412 7012 sw
tri 5412 6914 5510 7012 ne
rect 5510 6914 5864 7012
tri 5864 6914 5962 7012 sw
tri 5962 6914 6060 7012 ne
rect 6060 6914 6414 7012
tri 6414 6914 6512 7012 sw
tri 6512 6914 6610 7012 ne
rect 6610 6914 6964 7012
tri 6964 6914 7062 7012 sw
tri 7062 6914 7160 7012 ne
rect 7160 6914 7514 7012
tri 7514 6914 7612 7012 sw
tri 7612 6914 7710 7012 ne
rect 7710 6914 8064 7012
tri 8064 6914 8162 7012 sw
tri 8162 6914 8260 7012 ne
rect 8260 6914 8614 7012
tri 8614 6914 8712 7012 sw
tri 8712 6914 8810 7012 ne
rect 8810 6914 9164 7012
tri 9164 6914 9262 7012 sw
tri 9262 6914 9360 7012 ne
rect 9360 6914 9714 7012
tri 9714 6914 9812 7012 sw
tri 9812 6914 9910 7012 ne
rect 9910 6914 10264 7012
tri 10264 6914 10362 7012 sw
tri 10362 6914 10460 7012 ne
rect 10460 6914 10814 7012
tri 10814 6914 10912 7012 sw
tri 10912 6914 11010 7012 ne
rect 11010 6914 11364 7012
tri 11364 6914 11462 7012 sw
tri 11462 6914 11560 7012 ne
rect 11560 6914 11914 7012
tri 11914 6914 12012 7012 sw
tri 12012 6914 12110 7012 ne
rect 12110 6914 12464 7012
tri 12464 6914 12562 7012 sw
tri 12562 6914 12660 7012 ne
rect 12660 6914 13014 7012
tri 13014 6914 13112 7012 sw
tri 13112 6914 13210 7012 ne
rect 13210 6914 13564 7012
tri 13564 6914 13662 7012 sw
rect 14775 6914 15775 7562
rect -2525 6910 -88 6914
rect -2525 6790 -310 6910
rect -190 6826 -88 6910
tri -88 6826 0 6914 sw
tri 10 6826 98 6914 ne
rect 98 6910 462 6914
rect 98 6826 240 6910
rect -190 6790 0 6826
rect -2525 6786 0 6790
rect -2525 6138 -1525 6786
tri -412 6688 -314 6786 ne
rect -314 6738 0 6786
tri 0 6738 88 6826 sw
tri 98 6738 186 6826 ne
rect 186 6790 240 6826
rect 360 6826 462 6910
tri 462 6826 550 6914 sw
tri 560 6826 648 6914 ne
rect 648 6910 1012 6914
rect 648 6826 790 6910
rect 360 6790 550 6826
rect 186 6786 550 6790
tri 550 6786 590 6826 sw
tri 648 6786 688 6826 ne
rect 688 6790 790 6826
rect 910 6826 1012 6910
tri 1012 6826 1100 6914 sw
tri 1110 6826 1198 6914 ne
rect 1198 6910 1562 6914
rect 1198 6826 1340 6910
rect 910 6790 1100 6826
rect 688 6786 1100 6790
rect 186 6738 590 6786
rect -314 6688 88 6738
rect -1025 6600 -412 6688
tri -412 6600 -324 6688 sw
tri -314 6600 -226 6688 ne
rect -226 6658 88 6688
tri 88 6658 168 6738 sw
tri 186 6658 266 6738 ne
rect 266 6688 590 6738
tri 590 6688 688 6786 sw
tri 688 6688 786 6786 ne
rect 786 6738 1100 6786
tri 1100 6738 1188 6826 sw
tri 1198 6738 1286 6826 ne
rect 1286 6790 1340 6826
rect 1460 6826 1562 6910
tri 1562 6826 1650 6914 sw
tri 1660 6826 1748 6914 ne
rect 1748 6910 2112 6914
rect 1748 6826 1890 6910
rect 1460 6790 1650 6826
rect 1286 6786 1650 6790
tri 1650 6786 1690 6826 sw
tri 1748 6786 1788 6826 ne
rect 1788 6790 1890 6826
rect 2010 6826 2112 6910
tri 2112 6826 2200 6914 sw
tri 2210 6826 2298 6914 ne
rect 2298 6910 2662 6914
rect 2298 6826 2440 6910
rect 2010 6790 2200 6826
rect 1788 6786 2200 6790
rect 1286 6738 1690 6786
rect 786 6688 1188 6738
rect 266 6658 688 6688
rect -226 6600 168 6658
rect -1025 6560 -324 6600
tri -324 6560 -284 6600 sw
tri -226 6560 -186 6600 ne
rect -186 6560 168 6600
tri 168 6560 266 6658 sw
tri 266 6560 364 6658 ne
rect 364 6600 688 6658
tri 688 6600 776 6688 sw
tri 786 6600 874 6688 ne
rect 874 6658 1188 6688
tri 1188 6658 1268 6738 sw
tri 1286 6658 1366 6738 ne
rect 1366 6688 1690 6738
tri 1690 6688 1788 6786 sw
tri 1788 6688 1886 6786 ne
rect 1886 6738 2200 6786
tri 2200 6738 2288 6826 sw
tri 2298 6738 2386 6826 ne
rect 2386 6790 2440 6826
rect 2560 6826 2662 6910
tri 2662 6826 2750 6914 sw
tri 2760 6826 2848 6914 ne
rect 2848 6910 3212 6914
rect 2848 6826 2990 6910
rect 2560 6790 2750 6826
rect 2386 6786 2750 6790
tri 2750 6786 2790 6826 sw
tri 2848 6786 2888 6826 ne
rect 2888 6790 2990 6826
rect 3110 6826 3212 6910
tri 3212 6826 3300 6914 sw
tri 3310 6826 3398 6914 ne
rect 3398 6910 3762 6914
rect 3398 6826 3540 6910
rect 3110 6790 3300 6826
rect 2888 6786 3300 6790
rect 2386 6738 2790 6786
rect 1886 6688 2288 6738
rect 1366 6658 1788 6688
rect 874 6600 1268 6658
rect 364 6560 776 6600
tri 776 6560 816 6600 sw
tri 874 6560 914 6600 ne
rect 914 6560 1268 6600
tri 1268 6560 1366 6658 sw
tri 1366 6560 1464 6658 ne
rect 1464 6600 1788 6658
tri 1788 6600 1876 6688 sw
tri 1886 6600 1974 6688 ne
rect 1974 6658 2288 6688
tri 2288 6658 2368 6738 sw
tri 2386 6658 2466 6738 ne
rect 2466 6688 2790 6738
tri 2790 6688 2888 6786 sw
tri 2888 6688 2986 6786 ne
rect 2986 6738 3300 6786
tri 3300 6738 3388 6826 sw
tri 3398 6738 3486 6826 ne
rect 3486 6790 3540 6826
rect 3660 6826 3762 6910
tri 3762 6826 3850 6914 sw
tri 3860 6826 3948 6914 ne
rect 3948 6910 4312 6914
rect 3948 6826 4090 6910
rect 3660 6790 3850 6826
rect 3486 6786 3850 6790
tri 3850 6786 3890 6826 sw
tri 3948 6786 3988 6826 ne
rect 3988 6790 4090 6826
rect 4210 6826 4312 6910
tri 4312 6826 4400 6914 sw
tri 4410 6826 4498 6914 ne
rect 4498 6910 4862 6914
rect 4498 6826 4640 6910
rect 4210 6790 4400 6826
rect 3988 6786 4400 6790
rect 3486 6738 3890 6786
rect 2986 6688 3388 6738
rect 2466 6658 2888 6688
rect 1974 6600 2368 6658
rect 1464 6560 1876 6600
tri 1876 6560 1916 6600 sw
tri 1974 6560 2014 6600 ne
rect 2014 6560 2368 6600
tri 2368 6560 2466 6658 sw
tri 2466 6560 2564 6658 ne
rect 2564 6600 2888 6658
tri 2888 6600 2976 6688 sw
tri 2986 6600 3074 6688 ne
rect 3074 6658 3388 6688
tri 3388 6658 3468 6738 sw
tri 3486 6658 3566 6738 ne
rect 3566 6688 3890 6738
tri 3890 6688 3988 6786 sw
tri 3988 6688 4086 6786 ne
rect 4086 6738 4400 6786
tri 4400 6738 4488 6826 sw
tri 4498 6738 4586 6826 ne
rect 4586 6790 4640 6826
rect 4760 6826 4862 6910
tri 4862 6826 4950 6914 sw
tri 4960 6826 5048 6914 ne
rect 5048 6910 5412 6914
rect 5048 6826 5190 6910
rect 4760 6790 4950 6826
rect 4586 6786 4950 6790
tri 4950 6786 4990 6826 sw
tri 5048 6786 5088 6826 ne
rect 5088 6790 5190 6826
rect 5310 6826 5412 6910
tri 5412 6826 5500 6914 sw
tri 5510 6826 5598 6914 ne
rect 5598 6910 5962 6914
rect 5598 6826 5740 6910
rect 5310 6790 5500 6826
rect 5088 6786 5500 6790
rect 4586 6738 4990 6786
rect 4086 6688 4488 6738
rect 3566 6658 3988 6688
rect 3074 6600 3468 6658
rect 2564 6560 2976 6600
tri 2976 6560 3016 6600 sw
tri 3074 6560 3114 6600 ne
rect 3114 6560 3468 6600
tri 3468 6560 3566 6658 sw
tri 3566 6560 3664 6658 ne
rect 3664 6600 3988 6658
tri 3988 6600 4076 6688 sw
tri 4086 6600 4174 6688 ne
rect 4174 6658 4488 6688
tri 4488 6658 4568 6738 sw
tri 4586 6658 4666 6738 ne
rect 4666 6688 4990 6738
tri 4990 6688 5088 6786 sw
tri 5088 6688 5186 6786 ne
rect 5186 6738 5500 6786
tri 5500 6738 5588 6826 sw
tri 5598 6738 5686 6826 ne
rect 5686 6790 5740 6826
rect 5860 6826 5962 6910
tri 5962 6826 6050 6914 sw
tri 6060 6826 6148 6914 ne
rect 6148 6910 6512 6914
rect 6148 6826 6290 6910
rect 5860 6790 6050 6826
rect 5686 6786 6050 6790
tri 6050 6786 6090 6826 sw
tri 6148 6786 6188 6826 ne
rect 6188 6790 6290 6826
rect 6410 6826 6512 6910
tri 6512 6826 6600 6914 sw
tri 6610 6826 6698 6914 ne
rect 6698 6910 7062 6914
rect 6698 6826 6840 6910
rect 6410 6790 6600 6826
rect 6188 6786 6600 6790
rect 5686 6738 6090 6786
rect 5186 6688 5588 6738
rect 4666 6658 5088 6688
rect 4174 6600 4568 6658
rect 3664 6560 4076 6600
tri 4076 6560 4116 6600 sw
tri 4174 6560 4214 6600 ne
rect 4214 6560 4568 6600
tri 4568 6560 4666 6658 sw
tri 4666 6560 4764 6658 ne
rect 4764 6600 5088 6658
tri 5088 6600 5176 6688 sw
tri 5186 6600 5274 6688 ne
rect 5274 6658 5588 6688
tri 5588 6658 5668 6738 sw
tri 5686 6658 5766 6738 ne
rect 5766 6688 6090 6738
tri 6090 6688 6188 6786 sw
tri 6188 6688 6286 6786 ne
rect 6286 6738 6600 6786
tri 6600 6738 6688 6826 sw
tri 6698 6738 6786 6826 ne
rect 6786 6790 6840 6826
rect 6960 6826 7062 6910
tri 7062 6826 7150 6914 sw
tri 7160 6826 7248 6914 ne
rect 7248 6910 7612 6914
rect 7248 6826 7390 6910
rect 6960 6790 7150 6826
rect 6786 6786 7150 6790
tri 7150 6786 7190 6826 sw
tri 7248 6786 7288 6826 ne
rect 7288 6790 7390 6826
rect 7510 6826 7612 6910
tri 7612 6826 7700 6914 sw
tri 7710 6826 7798 6914 ne
rect 7798 6910 8162 6914
rect 7798 6826 7940 6910
rect 7510 6790 7700 6826
rect 7288 6786 7700 6790
rect 6786 6738 7190 6786
rect 6286 6688 6688 6738
rect 5766 6658 6188 6688
rect 5274 6600 5668 6658
rect 4764 6560 5176 6600
tri 5176 6560 5216 6600 sw
tri 5274 6560 5314 6600 ne
rect 5314 6560 5668 6600
tri 5668 6560 5766 6658 sw
tri 5766 6560 5864 6658 ne
rect 5864 6600 6188 6658
tri 6188 6600 6276 6688 sw
tri 6286 6600 6374 6688 ne
rect 6374 6658 6688 6688
tri 6688 6658 6768 6738 sw
tri 6786 6658 6866 6738 ne
rect 6866 6688 7190 6738
tri 7190 6688 7288 6786 sw
tri 7288 6688 7386 6786 ne
rect 7386 6738 7700 6786
tri 7700 6738 7788 6826 sw
tri 7798 6738 7886 6826 ne
rect 7886 6790 7940 6826
rect 8060 6826 8162 6910
tri 8162 6826 8250 6914 sw
tri 8260 6826 8348 6914 ne
rect 8348 6910 8712 6914
rect 8348 6826 8490 6910
rect 8060 6790 8250 6826
rect 7886 6786 8250 6790
tri 8250 6786 8290 6826 sw
tri 8348 6786 8388 6826 ne
rect 8388 6790 8490 6826
rect 8610 6826 8712 6910
tri 8712 6826 8800 6914 sw
tri 8810 6826 8898 6914 ne
rect 8898 6910 9262 6914
rect 8898 6826 9040 6910
rect 8610 6790 8800 6826
rect 8388 6786 8800 6790
rect 7886 6738 8290 6786
rect 7386 6688 7788 6738
rect 6866 6658 7288 6688
rect 6374 6600 6768 6658
rect 5864 6560 6276 6600
tri 6276 6560 6316 6600 sw
tri 6374 6560 6414 6600 ne
rect 6414 6560 6768 6600
tri 6768 6560 6866 6658 sw
tri 6866 6560 6964 6658 ne
rect 6964 6600 7288 6658
tri 7288 6600 7376 6688 sw
tri 7386 6600 7474 6688 ne
rect 7474 6658 7788 6688
tri 7788 6658 7868 6738 sw
tri 7886 6658 7966 6738 ne
rect 7966 6688 8290 6738
tri 8290 6688 8388 6786 sw
tri 8388 6688 8486 6786 ne
rect 8486 6738 8800 6786
tri 8800 6738 8888 6826 sw
tri 8898 6738 8986 6826 ne
rect 8986 6790 9040 6826
rect 9160 6826 9262 6910
tri 9262 6826 9350 6914 sw
tri 9360 6826 9448 6914 ne
rect 9448 6910 9812 6914
rect 9448 6826 9590 6910
rect 9160 6790 9350 6826
rect 8986 6786 9350 6790
tri 9350 6786 9390 6826 sw
tri 9448 6786 9488 6826 ne
rect 9488 6790 9590 6826
rect 9710 6826 9812 6910
tri 9812 6826 9900 6914 sw
tri 9910 6826 9998 6914 ne
rect 9998 6910 10362 6914
rect 9998 6826 10140 6910
rect 9710 6790 9900 6826
rect 9488 6786 9900 6790
rect 8986 6738 9390 6786
rect 8486 6688 8888 6738
rect 7966 6658 8388 6688
rect 7474 6600 7868 6658
rect 6964 6560 7376 6600
tri 7376 6560 7416 6600 sw
tri 7474 6560 7514 6600 ne
rect 7514 6560 7868 6600
tri 7868 6560 7966 6658 sw
tri 7966 6560 8064 6658 ne
rect 8064 6600 8388 6658
tri 8388 6600 8476 6688 sw
tri 8486 6600 8574 6688 ne
rect 8574 6658 8888 6688
tri 8888 6658 8968 6738 sw
tri 8986 6658 9066 6738 ne
rect 9066 6688 9390 6738
tri 9390 6688 9488 6786 sw
tri 9488 6688 9586 6786 ne
rect 9586 6738 9900 6786
tri 9900 6738 9988 6826 sw
tri 9998 6738 10086 6826 ne
rect 10086 6790 10140 6826
rect 10260 6826 10362 6910
tri 10362 6826 10450 6914 sw
tri 10460 6826 10548 6914 ne
rect 10548 6910 10912 6914
rect 10548 6826 10690 6910
rect 10260 6790 10450 6826
rect 10086 6786 10450 6790
tri 10450 6786 10490 6826 sw
tri 10548 6786 10588 6826 ne
rect 10588 6790 10690 6826
rect 10810 6826 10912 6910
tri 10912 6826 11000 6914 sw
tri 11010 6826 11098 6914 ne
rect 11098 6910 11462 6914
rect 11098 6826 11240 6910
rect 10810 6790 11000 6826
rect 10588 6786 11000 6790
rect 10086 6738 10490 6786
rect 9586 6688 9988 6738
rect 9066 6658 9488 6688
rect 8574 6600 8968 6658
rect 8064 6560 8476 6600
tri 8476 6560 8516 6600 sw
tri 8574 6560 8614 6600 ne
rect 8614 6560 8968 6600
tri 8968 6560 9066 6658 sw
tri 9066 6560 9164 6658 ne
rect 9164 6600 9488 6658
tri 9488 6600 9576 6688 sw
tri 9586 6600 9674 6688 ne
rect 9674 6658 9988 6688
tri 9988 6658 10068 6738 sw
tri 10086 6658 10166 6738 ne
rect 10166 6688 10490 6738
tri 10490 6688 10588 6786 sw
tri 10588 6688 10686 6786 ne
rect 10686 6738 11000 6786
tri 11000 6738 11088 6826 sw
tri 11098 6738 11186 6826 ne
rect 11186 6790 11240 6826
rect 11360 6826 11462 6910
tri 11462 6826 11550 6914 sw
tri 11560 6826 11648 6914 ne
rect 11648 6910 12012 6914
rect 11648 6826 11790 6910
rect 11360 6790 11550 6826
rect 11186 6786 11550 6790
tri 11550 6786 11590 6826 sw
tri 11648 6786 11688 6826 ne
rect 11688 6790 11790 6826
rect 11910 6826 12012 6910
tri 12012 6826 12100 6914 sw
tri 12110 6826 12198 6914 ne
rect 12198 6910 12562 6914
rect 12198 6826 12340 6910
rect 11910 6790 12100 6826
rect 11688 6786 12100 6790
rect 11186 6738 11590 6786
rect 10686 6688 11088 6738
rect 10166 6658 10588 6688
rect 9674 6600 10068 6658
rect 9164 6560 9576 6600
tri 9576 6560 9616 6600 sw
tri 9674 6560 9714 6600 ne
rect 9714 6560 10068 6600
tri 10068 6560 10166 6658 sw
tri 10166 6560 10264 6658 ne
rect 10264 6600 10588 6658
tri 10588 6600 10676 6688 sw
tri 10686 6600 10774 6688 ne
rect 10774 6658 11088 6688
tri 11088 6658 11168 6738 sw
tri 11186 6658 11266 6738 ne
rect 11266 6688 11590 6738
tri 11590 6688 11688 6786 sw
tri 11688 6688 11786 6786 ne
rect 11786 6738 12100 6786
tri 12100 6738 12188 6826 sw
tri 12198 6738 12286 6826 ne
rect 12286 6790 12340 6826
rect 12460 6826 12562 6910
tri 12562 6826 12650 6914 sw
tri 12660 6826 12748 6914 ne
rect 12748 6910 13112 6914
rect 12748 6826 12890 6910
rect 12460 6790 12650 6826
rect 12286 6786 12650 6790
tri 12650 6786 12690 6826 sw
tri 12748 6786 12788 6826 ne
rect 12788 6790 12890 6826
rect 13010 6826 13112 6910
tri 13112 6826 13200 6914 sw
tri 13210 6826 13298 6914 ne
rect 13298 6910 15775 6914
rect 13298 6826 13440 6910
rect 13010 6790 13200 6826
rect 12788 6786 13200 6790
rect 12286 6738 12690 6786
rect 11786 6688 12188 6738
rect 11266 6658 11688 6688
rect 10774 6600 11168 6658
rect 10264 6560 10676 6600
tri 10676 6560 10716 6600 sw
tri 10774 6560 10814 6600 ne
rect 10814 6560 11168 6600
tri 11168 6560 11266 6658 sw
tri 11266 6560 11364 6658 ne
rect 11364 6600 11688 6658
tri 11688 6600 11776 6688 sw
tri 11786 6600 11874 6688 ne
rect 11874 6658 12188 6688
tri 12188 6658 12268 6738 sw
tri 12286 6658 12366 6738 ne
rect 12366 6688 12690 6738
tri 12690 6688 12788 6786 sw
tri 12788 6688 12886 6786 ne
rect 12886 6738 13200 6786
tri 13200 6738 13288 6826 sw
tri 13298 6738 13386 6826 ne
rect 13386 6790 13440 6826
rect 13560 6790 15775 6910
rect 13386 6738 15775 6790
rect 12886 6688 13288 6738
rect 12366 6658 12788 6688
rect 11874 6600 12268 6658
rect 11364 6560 11776 6600
tri 11776 6560 11816 6600 sw
tri 11874 6560 11914 6600 ne
rect 11914 6560 12268 6600
tri 12268 6560 12366 6658 sw
tri 12366 6560 12464 6658 ne
rect 12464 6600 12788 6658
tri 12788 6600 12876 6688 sw
tri 12886 6600 12974 6688 ne
rect 12974 6658 13288 6688
tri 13288 6658 13368 6738 sw
tri 13386 6658 13466 6738 ne
rect 13466 6658 14075 6738
rect 12974 6600 13368 6658
rect 12464 6560 12876 6600
tri 12876 6560 12916 6600 sw
tri 12974 6560 13014 6600 ne
rect 13014 6560 13368 6600
tri 13368 6560 13466 6658 sw
tri 13466 6560 13564 6658 ne
rect 13564 6638 14075 6658
rect 14175 6638 15775 6738
rect 13564 6560 15775 6638
rect -1025 6512 -284 6560
rect -1025 6412 -925 6512
rect -825 6462 -284 6512
tri -284 6462 -186 6560 sw
tri -186 6462 -88 6560 ne
rect -88 6462 266 6560
tri 266 6462 364 6560 sw
tri 364 6462 462 6560 ne
rect 462 6462 816 6560
tri 816 6462 914 6560 sw
tri 914 6462 1012 6560 ne
rect 1012 6462 1366 6560
tri 1366 6462 1464 6560 sw
tri 1464 6462 1562 6560 ne
rect 1562 6462 1916 6560
tri 1916 6462 2014 6560 sw
tri 2014 6462 2112 6560 ne
rect 2112 6462 2466 6560
tri 2466 6462 2564 6560 sw
tri 2564 6462 2662 6560 ne
rect 2662 6462 3016 6560
tri 3016 6462 3114 6560 sw
tri 3114 6462 3212 6560 ne
rect 3212 6462 3566 6560
tri 3566 6462 3664 6560 sw
tri 3664 6462 3762 6560 ne
rect 3762 6462 4116 6560
tri 4116 6462 4214 6560 sw
tri 4214 6462 4312 6560 ne
rect 4312 6462 4666 6560
tri 4666 6462 4764 6560 sw
tri 4764 6462 4862 6560 ne
rect 4862 6462 5216 6560
tri 5216 6462 5314 6560 sw
tri 5314 6462 5412 6560 ne
rect 5412 6462 5766 6560
tri 5766 6462 5864 6560 sw
tri 5864 6462 5962 6560 ne
rect 5962 6462 6316 6560
tri 6316 6462 6414 6560 sw
tri 6414 6462 6512 6560 ne
rect 6512 6462 6866 6560
tri 6866 6462 6964 6560 sw
tri 6964 6462 7062 6560 ne
rect 7062 6462 7416 6560
tri 7416 6462 7514 6560 sw
tri 7514 6462 7612 6560 ne
rect 7612 6462 7966 6560
tri 7966 6462 8064 6560 sw
tri 8064 6462 8162 6560 ne
rect 8162 6462 8516 6560
tri 8516 6462 8614 6560 sw
tri 8614 6462 8712 6560 ne
rect 8712 6462 9066 6560
tri 9066 6462 9164 6560 sw
tri 9164 6462 9262 6560 ne
rect 9262 6462 9616 6560
tri 9616 6462 9714 6560 sw
tri 9714 6462 9812 6560 ne
rect 9812 6462 10166 6560
tri 10166 6462 10264 6560 sw
tri 10264 6462 10362 6560 ne
rect 10362 6462 10716 6560
tri 10716 6462 10814 6560 sw
tri 10814 6462 10912 6560 ne
rect 10912 6462 11266 6560
tri 11266 6462 11364 6560 sw
tri 11364 6462 11462 6560 ne
rect 11462 6462 11816 6560
tri 11816 6462 11914 6560 sw
tri 11914 6462 12012 6560 ne
rect 12012 6462 12366 6560
tri 12366 6462 12464 6560 sw
tri 12464 6462 12562 6560 ne
rect 12562 6462 12916 6560
tri 12916 6462 13014 6560 sw
tri 13014 6462 13112 6560 ne
rect 13112 6462 13466 6560
tri 13466 6462 13564 6560 sw
tri 13564 6462 13662 6560 ne
rect 13662 6462 15775 6560
rect -825 6412 -186 6462
rect -1025 6364 -186 6412
tri -186 6364 -88 6462 sw
tri -88 6364 10 6462 ne
rect 10 6364 364 6462
tri 364 6364 462 6462 sw
tri 462 6364 560 6462 ne
rect 560 6364 914 6462
tri 914 6364 1012 6462 sw
tri 1012 6364 1110 6462 ne
rect 1110 6364 1464 6462
tri 1464 6364 1562 6462 sw
tri 1562 6364 1660 6462 ne
rect 1660 6364 2014 6462
tri 2014 6364 2112 6462 sw
tri 2112 6364 2210 6462 ne
rect 2210 6364 2564 6462
tri 2564 6364 2662 6462 sw
tri 2662 6364 2760 6462 ne
rect 2760 6364 3114 6462
tri 3114 6364 3212 6462 sw
tri 3212 6364 3310 6462 ne
rect 3310 6364 3664 6462
tri 3664 6364 3762 6462 sw
tri 3762 6364 3860 6462 ne
rect 3860 6364 4214 6462
tri 4214 6364 4312 6462 sw
tri 4312 6364 4410 6462 ne
rect 4410 6364 4764 6462
tri 4764 6364 4862 6462 sw
tri 4862 6364 4960 6462 ne
rect 4960 6364 5314 6462
tri 5314 6364 5412 6462 sw
tri 5412 6364 5510 6462 ne
rect 5510 6364 5864 6462
tri 5864 6364 5962 6462 sw
tri 5962 6364 6060 6462 ne
rect 6060 6364 6414 6462
tri 6414 6364 6512 6462 sw
tri 6512 6364 6610 6462 ne
rect 6610 6364 6964 6462
tri 6964 6364 7062 6462 sw
tri 7062 6364 7160 6462 ne
rect 7160 6364 7514 6462
tri 7514 6364 7612 6462 sw
tri 7612 6364 7710 6462 ne
rect 7710 6364 8064 6462
tri 8064 6364 8162 6462 sw
tri 8162 6364 8260 6462 ne
rect 8260 6364 8614 6462
tri 8614 6364 8712 6462 sw
tri 8712 6364 8810 6462 ne
rect 8810 6364 9164 6462
tri 9164 6364 9262 6462 sw
tri 9262 6364 9360 6462 ne
rect 9360 6364 9714 6462
tri 9714 6364 9812 6462 sw
tri 9812 6364 9910 6462 ne
rect 9910 6364 10264 6462
tri 10264 6364 10362 6462 sw
tri 10362 6364 10460 6462 ne
rect 10460 6364 10814 6462
tri 10814 6364 10912 6462 sw
tri 10912 6364 11010 6462 ne
rect 11010 6364 11364 6462
tri 11364 6364 11462 6462 sw
tri 11462 6364 11560 6462 ne
rect 11560 6364 11914 6462
tri 11914 6364 12012 6462 sw
tri 12012 6364 12110 6462 ne
rect 12110 6364 12464 6462
tri 12464 6364 12562 6462 sw
tri 12562 6364 12660 6462 ne
rect 12660 6364 13014 6462
tri 13014 6364 13112 6462 sw
tri 13112 6364 13210 6462 ne
rect 13210 6364 13564 6462
tri 13564 6364 13662 6462 sw
rect -1025 6360 -88 6364
rect -1025 6240 -310 6360
rect -190 6276 -88 6360
tri -88 6276 0 6364 sw
tri 10 6276 98 6364 ne
rect 98 6360 462 6364
rect 98 6276 240 6360
rect -190 6240 0 6276
rect -1025 6236 0 6240
tri 0 6236 40 6276 sw
tri 98 6236 138 6276 ne
rect 138 6240 240 6276
rect 360 6276 462 6360
tri 462 6276 550 6364 sw
tri 560 6276 648 6364 ne
rect 648 6360 1012 6364
rect 648 6276 790 6360
rect 360 6240 550 6276
rect 138 6236 550 6240
tri -412 6138 -314 6236 ne
rect -314 6138 40 6236
tri 40 6138 138 6236 sw
tri 138 6138 236 6236 ne
rect 236 6188 550 6236
tri 550 6188 638 6276 sw
tri 648 6188 736 6276 ne
rect 736 6240 790 6276
rect 910 6276 1012 6360
tri 1012 6276 1100 6364 sw
tri 1110 6276 1198 6364 ne
rect 1198 6360 1562 6364
rect 1198 6276 1340 6360
rect 910 6240 1100 6276
rect 736 6236 1100 6240
tri 1100 6236 1140 6276 sw
tri 1198 6236 1238 6276 ne
rect 1238 6240 1340 6276
rect 1460 6276 1562 6360
tri 1562 6276 1650 6364 sw
tri 1660 6276 1748 6364 ne
rect 1748 6360 2112 6364
rect 1748 6276 1890 6360
rect 1460 6240 1650 6276
rect 1238 6236 1650 6240
rect 736 6188 1140 6236
rect 236 6138 638 6188
rect -2525 6050 -412 6138
tri -412 6050 -324 6138 sw
tri -314 6050 -226 6138 ne
rect -226 6050 138 6138
tri 138 6050 226 6138 sw
tri 236 6050 324 6138 ne
rect 324 6108 638 6138
tri 638 6108 718 6188 sw
tri 736 6108 816 6188 ne
rect 816 6138 1140 6188
tri 1140 6138 1238 6236 sw
tri 1238 6138 1336 6236 ne
rect 1336 6188 1650 6236
tri 1650 6188 1738 6276 sw
tri 1748 6188 1836 6276 ne
rect 1836 6240 1890 6276
rect 2010 6276 2112 6360
tri 2112 6276 2200 6364 sw
tri 2210 6276 2298 6364 ne
rect 2298 6360 2662 6364
rect 2298 6276 2440 6360
rect 2010 6240 2200 6276
rect 1836 6236 2200 6240
tri 2200 6236 2240 6276 sw
tri 2298 6236 2338 6276 ne
rect 2338 6240 2440 6276
rect 2560 6276 2662 6360
tri 2662 6276 2750 6364 sw
tri 2760 6276 2848 6364 ne
rect 2848 6360 3212 6364
rect 2848 6276 2990 6360
rect 2560 6240 2750 6276
rect 2338 6236 2750 6240
rect 1836 6188 2240 6236
rect 1336 6138 1738 6188
rect 816 6108 1238 6138
rect 324 6050 718 6108
rect -2525 6010 -324 6050
tri -324 6010 -284 6050 sw
tri -226 6010 -186 6050 ne
rect -186 6010 226 6050
tri 226 6010 266 6050 sw
tri 324 6010 364 6050 ne
rect 364 6010 718 6050
tri 718 6010 816 6108 sw
tri 816 6010 914 6108 ne
rect 914 6050 1238 6108
tri 1238 6050 1326 6138 sw
tri 1336 6050 1424 6138 ne
rect 1424 6108 1738 6138
tri 1738 6108 1818 6188 sw
tri 1836 6108 1916 6188 ne
rect 1916 6138 2240 6188
tri 2240 6138 2338 6236 sw
tri 2338 6138 2436 6236 ne
rect 2436 6188 2750 6236
tri 2750 6188 2838 6276 sw
tri 2848 6188 2936 6276 ne
rect 2936 6240 2990 6276
rect 3110 6276 3212 6360
tri 3212 6276 3300 6364 sw
tri 3310 6276 3398 6364 ne
rect 3398 6360 3762 6364
rect 3398 6276 3540 6360
rect 3110 6240 3300 6276
rect 2936 6236 3300 6240
tri 3300 6236 3340 6276 sw
tri 3398 6236 3438 6276 ne
rect 3438 6240 3540 6276
rect 3660 6276 3762 6360
tri 3762 6276 3850 6364 sw
tri 3860 6276 3948 6364 ne
rect 3948 6360 4312 6364
rect 3948 6276 4090 6360
rect 3660 6240 3850 6276
rect 3438 6236 3850 6240
rect 2936 6188 3340 6236
rect 2436 6138 2838 6188
rect 1916 6108 2338 6138
rect 1424 6050 1818 6108
rect 914 6010 1326 6050
tri 1326 6010 1366 6050 sw
tri 1424 6010 1464 6050 ne
rect 1464 6010 1818 6050
tri 1818 6010 1916 6108 sw
tri 1916 6010 2014 6108 ne
rect 2014 6050 2338 6108
tri 2338 6050 2426 6138 sw
tri 2436 6050 2524 6138 ne
rect 2524 6108 2838 6138
tri 2838 6108 2918 6188 sw
tri 2936 6108 3016 6188 ne
rect 3016 6138 3340 6188
tri 3340 6138 3438 6236 sw
tri 3438 6138 3536 6236 ne
rect 3536 6188 3850 6236
tri 3850 6188 3938 6276 sw
tri 3948 6188 4036 6276 ne
rect 4036 6240 4090 6276
rect 4210 6276 4312 6360
tri 4312 6276 4400 6364 sw
tri 4410 6276 4498 6364 ne
rect 4498 6360 4862 6364
rect 4498 6276 4640 6360
rect 4210 6240 4400 6276
rect 4036 6236 4400 6240
tri 4400 6236 4440 6276 sw
tri 4498 6236 4538 6276 ne
rect 4538 6240 4640 6276
rect 4760 6276 4862 6360
tri 4862 6276 4950 6364 sw
tri 4960 6276 5048 6364 ne
rect 5048 6360 5412 6364
rect 5048 6276 5190 6360
rect 4760 6240 4950 6276
rect 4538 6236 4950 6240
rect 4036 6188 4440 6236
rect 3536 6138 3938 6188
rect 3016 6108 3438 6138
rect 2524 6050 2918 6108
rect 2014 6010 2426 6050
tri 2426 6010 2466 6050 sw
tri 2524 6010 2564 6050 ne
rect 2564 6010 2918 6050
tri 2918 6010 3016 6108 sw
tri 3016 6010 3114 6108 ne
rect 3114 6050 3438 6108
tri 3438 6050 3526 6138 sw
tri 3536 6050 3624 6138 ne
rect 3624 6108 3938 6138
tri 3938 6108 4018 6188 sw
tri 4036 6108 4116 6188 ne
rect 4116 6138 4440 6188
tri 4440 6138 4538 6236 sw
tri 4538 6138 4636 6236 ne
rect 4636 6188 4950 6236
tri 4950 6188 5038 6276 sw
tri 5048 6188 5136 6276 ne
rect 5136 6240 5190 6276
rect 5310 6276 5412 6360
tri 5412 6276 5500 6364 sw
tri 5510 6276 5598 6364 ne
rect 5598 6360 5962 6364
rect 5598 6276 5740 6360
rect 5310 6240 5500 6276
rect 5136 6236 5500 6240
tri 5500 6236 5540 6276 sw
tri 5598 6236 5638 6276 ne
rect 5638 6240 5740 6276
rect 5860 6276 5962 6360
tri 5962 6276 6050 6364 sw
tri 6060 6276 6148 6364 ne
rect 6148 6360 6512 6364
rect 6148 6276 6290 6360
rect 5860 6240 6050 6276
rect 5638 6236 6050 6240
rect 5136 6188 5540 6236
rect 4636 6138 5038 6188
rect 4116 6108 4538 6138
rect 3624 6050 4018 6108
rect 3114 6010 3526 6050
tri 3526 6010 3566 6050 sw
tri 3624 6010 3664 6050 ne
rect 3664 6010 4018 6050
tri 4018 6010 4116 6108 sw
tri 4116 6010 4214 6108 ne
rect 4214 6050 4538 6108
tri 4538 6050 4626 6138 sw
tri 4636 6050 4724 6138 ne
rect 4724 6108 5038 6138
tri 5038 6108 5118 6188 sw
tri 5136 6108 5216 6188 ne
rect 5216 6138 5540 6188
tri 5540 6138 5638 6236 sw
tri 5638 6138 5736 6236 ne
rect 5736 6188 6050 6236
tri 6050 6188 6138 6276 sw
tri 6148 6188 6236 6276 ne
rect 6236 6240 6290 6276
rect 6410 6276 6512 6360
tri 6512 6276 6600 6364 sw
tri 6610 6276 6698 6364 ne
rect 6698 6360 7062 6364
rect 6698 6276 6840 6360
rect 6410 6240 6600 6276
rect 6236 6236 6600 6240
tri 6600 6236 6640 6276 sw
tri 6698 6236 6738 6276 ne
rect 6738 6240 6840 6276
rect 6960 6276 7062 6360
tri 7062 6276 7150 6364 sw
tri 7160 6276 7248 6364 ne
rect 7248 6360 7612 6364
rect 7248 6276 7390 6360
rect 6960 6240 7150 6276
rect 6738 6236 7150 6240
rect 6236 6188 6640 6236
rect 5736 6138 6138 6188
rect 5216 6108 5638 6138
rect 4724 6050 5118 6108
rect 4214 6010 4626 6050
tri 4626 6010 4666 6050 sw
tri 4724 6010 4764 6050 ne
rect 4764 6010 5118 6050
tri 5118 6010 5216 6108 sw
tri 5216 6010 5314 6108 ne
rect 5314 6050 5638 6108
tri 5638 6050 5726 6138 sw
tri 5736 6050 5824 6138 ne
rect 5824 6108 6138 6138
tri 6138 6108 6218 6188 sw
tri 6236 6108 6316 6188 ne
rect 6316 6138 6640 6188
tri 6640 6138 6738 6236 sw
tri 6738 6138 6836 6236 ne
rect 6836 6188 7150 6236
tri 7150 6188 7238 6276 sw
tri 7248 6188 7336 6276 ne
rect 7336 6240 7390 6276
rect 7510 6276 7612 6360
tri 7612 6276 7700 6364 sw
tri 7710 6276 7798 6364 ne
rect 7798 6360 8162 6364
rect 7798 6276 7940 6360
rect 7510 6240 7700 6276
rect 7336 6236 7700 6240
tri 7700 6236 7740 6276 sw
tri 7798 6236 7838 6276 ne
rect 7838 6240 7940 6276
rect 8060 6276 8162 6360
tri 8162 6276 8250 6364 sw
tri 8260 6276 8348 6364 ne
rect 8348 6360 8712 6364
rect 8348 6276 8490 6360
rect 8060 6240 8250 6276
rect 7838 6236 8250 6240
rect 7336 6188 7740 6236
rect 6836 6138 7238 6188
rect 6316 6108 6738 6138
rect 5824 6050 6218 6108
rect 5314 6010 5726 6050
tri 5726 6010 5766 6050 sw
tri 5824 6010 5864 6050 ne
rect 5864 6010 6218 6050
tri 6218 6010 6316 6108 sw
tri 6316 6010 6414 6108 ne
rect 6414 6050 6738 6108
tri 6738 6050 6826 6138 sw
tri 6836 6050 6924 6138 ne
rect 6924 6108 7238 6138
tri 7238 6108 7318 6188 sw
tri 7336 6108 7416 6188 ne
rect 7416 6138 7740 6188
tri 7740 6138 7838 6236 sw
tri 7838 6138 7936 6236 ne
rect 7936 6188 8250 6236
tri 8250 6188 8338 6276 sw
tri 8348 6188 8436 6276 ne
rect 8436 6240 8490 6276
rect 8610 6276 8712 6360
tri 8712 6276 8800 6364 sw
tri 8810 6276 8898 6364 ne
rect 8898 6360 9262 6364
rect 8898 6276 9040 6360
rect 8610 6240 8800 6276
rect 8436 6236 8800 6240
tri 8800 6236 8840 6276 sw
tri 8898 6236 8938 6276 ne
rect 8938 6240 9040 6276
rect 9160 6276 9262 6360
tri 9262 6276 9350 6364 sw
tri 9360 6276 9448 6364 ne
rect 9448 6360 9812 6364
rect 9448 6276 9590 6360
rect 9160 6240 9350 6276
rect 8938 6236 9350 6240
rect 8436 6188 8840 6236
rect 7936 6138 8338 6188
rect 7416 6108 7838 6138
rect 6924 6050 7318 6108
rect 6414 6010 6826 6050
tri 6826 6010 6866 6050 sw
tri 6924 6010 6964 6050 ne
rect 6964 6010 7318 6050
tri 7318 6010 7416 6108 sw
tri 7416 6010 7514 6108 ne
rect 7514 6050 7838 6108
tri 7838 6050 7926 6138 sw
tri 7936 6050 8024 6138 ne
rect 8024 6108 8338 6138
tri 8338 6108 8418 6188 sw
tri 8436 6108 8516 6188 ne
rect 8516 6138 8840 6188
tri 8840 6138 8938 6236 sw
tri 8938 6138 9036 6236 ne
rect 9036 6188 9350 6236
tri 9350 6188 9438 6276 sw
tri 9448 6188 9536 6276 ne
rect 9536 6240 9590 6276
rect 9710 6276 9812 6360
tri 9812 6276 9900 6364 sw
tri 9910 6276 9998 6364 ne
rect 9998 6360 10362 6364
rect 9998 6276 10140 6360
rect 9710 6240 9900 6276
rect 9536 6236 9900 6240
tri 9900 6236 9940 6276 sw
tri 9998 6236 10038 6276 ne
rect 10038 6240 10140 6276
rect 10260 6276 10362 6360
tri 10362 6276 10450 6364 sw
tri 10460 6276 10548 6364 ne
rect 10548 6360 10912 6364
rect 10548 6276 10690 6360
rect 10260 6240 10450 6276
rect 10038 6236 10450 6240
rect 9536 6188 9940 6236
rect 9036 6138 9438 6188
rect 8516 6108 8938 6138
rect 8024 6050 8418 6108
rect 7514 6010 7926 6050
tri 7926 6010 7966 6050 sw
tri 8024 6010 8064 6050 ne
rect 8064 6010 8418 6050
tri 8418 6010 8516 6108 sw
tri 8516 6010 8614 6108 ne
rect 8614 6050 8938 6108
tri 8938 6050 9026 6138 sw
tri 9036 6050 9124 6138 ne
rect 9124 6108 9438 6138
tri 9438 6108 9518 6188 sw
tri 9536 6108 9616 6188 ne
rect 9616 6138 9940 6188
tri 9940 6138 10038 6236 sw
tri 10038 6138 10136 6236 ne
rect 10136 6188 10450 6236
tri 10450 6188 10538 6276 sw
tri 10548 6188 10636 6276 ne
rect 10636 6240 10690 6276
rect 10810 6276 10912 6360
tri 10912 6276 11000 6364 sw
tri 11010 6276 11098 6364 ne
rect 11098 6360 11462 6364
rect 11098 6276 11240 6360
rect 10810 6240 11000 6276
rect 10636 6236 11000 6240
tri 11000 6236 11040 6276 sw
tri 11098 6236 11138 6276 ne
rect 11138 6240 11240 6276
rect 11360 6276 11462 6360
tri 11462 6276 11550 6364 sw
tri 11560 6276 11648 6364 ne
rect 11648 6360 12012 6364
rect 11648 6276 11790 6360
rect 11360 6240 11550 6276
rect 11138 6236 11550 6240
rect 10636 6188 11040 6236
rect 10136 6138 10538 6188
rect 9616 6108 10038 6138
rect 9124 6050 9518 6108
rect 8614 6010 9026 6050
tri 9026 6010 9066 6050 sw
tri 9124 6010 9164 6050 ne
rect 9164 6010 9518 6050
tri 9518 6010 9616 6108 sw
tri 9616 6010 9714 6108 ne
rect 9714 6050 10038 6108
tri 10038 6050 10126 6138 sw
tri 10136 6050 10224 6138 ne
rect 10224 6108 10538 6138
tri 10538 6108 10618 6188 sw
tri 10636 6108 10716 6188 ne
rect 10716 6138 11040 6188
tri 11040 6138 11138 6236 sw
tri 11138 6138 11236 6236 ne
rect 11236 6188 11550 6236
tri 11550 6188 11638 6276 sw
tri 11648 6188 11736 6276 ne
rect 11736 6240 11790 6276
rect 11910 6276 12012 6360
tri 12012 6276 12100 6364 sw
tri 12110 6276 12198 6364 ne
rect 12198 6360 12562 6364
rect 12198 6276 12340 6360
rect 11910 6240 12100 6276
rect 11736 6236 12100 6240
tri 12100 6236 12140 6276 sw
tri 12198 6236 12238 6276 ne
rect 12238 6240 12340 6276
rect 12460 6276 12562 6360
tri 12562 6276 12650 6364 sw
tri 12660 6276 12748 6364 ne
rect 12748 6360 13112 6364
rect 12748 6276 12890 6360
rect 12460 6240 12650 6276
rect 12238 6236 12650 6240
rect 11736 6188 12140 6236
rect 11236 6138 11638 6188
rect 10716 6108 11138 6138
rect 10224 6050 10618 6108
rect 9714 6010 10126 6050
tri 10126 6010 10166 6050 sw
tri 10224 6010 10264 6050 ne
rect 10264 6010 10618 6050
tri 10618 6010 10716 6108 sw
tri 10716 6010 10814 6108 ne
rect 10814 6050 11138 6108
tri 11138 6050 11226 6138 sw
tri 11236 6050 11324 6138 ne
rect 11324 6108 11638 6138
tri 11638 6108 11718 6188 sw
tri 11736 6108 11816 6188 ne
rect 11816 6138 12140 6188
tri 12140 6138 12238 6236 sw
tri 12238 6138 12336 6236 ne
rect 12336 6188 12650 6236
tri 12650 6188 12738 6276 sw
tri 12748 6188 12836 6276 ne
rect 12836 6240 12890 6276
rect 13010 6276 13112 6360
tri 13112 6276 13200 6364 sw
tri 13210 6276 13298 6364 ne
rect 13298 6360 14275 6364
rect 13298 6276 13440 6360
rect 13010 6240 13200 6276
rect 12836 6236 13200 6240
tri 13200 6236 13240 6276 sw
tri 13298 6236 13338 6276 ne
rect 13338 6240 13440 6276
rect 13560 6240 14275 6360
rect 13338 6236 14275 6240
rect 12836 6188 13240 6236
rect 12336 6138 12738 6188
rect 11816 6108 12238 6138
rect 11324 6050 11718 6108
rect 10814 6010 11226 6050
tri 11226 6010 11266 6050 sw
tri 11324 6010 11364 6050 ne
rect 11364 6010 11718 6050
tri 11718 6010 11816 6108 sw
tri 11816 6010 11914 6108 ne
rect 11914 6050 12238 6108
tri 12238 6050 12326 6138 sw
tri 12336 6050 12424 6138 ne
rect 12424 6108 12738 6138
tri 12738 6108 12818 6188 sw
tri 12836 6108 12916 6188 ne
rect 12916 6138 13240 6188
tri 13240 6138 13338 6236 sw
tri 13338 6138 13436 6236 ne
rect 13436 6138 14275 6236
rect 12916 6108 13338 6138
rect 12424 6050 12818 6108
rect 11914 6010 12326 6050
tri 12326 6010 12366 6050 sw
tri 12424 6010 12464 6050 ne
rect 12464 6010 12818 6050
tri 12818 6010 12916 6108 sw
tri 12916 6010 13014 6108 ne
rect 13014 6050 13338 6108
tri 13338 6050 13426 6138 sw
tri 13436 6050 13524 6138 ne
rect 13524 6050 14275 6138
rect 13014 6010 13426 6050
tri 13426 6010 13466 6050 sw
tri 13524 6010 13564 6050 ne
rect 13564 6010 14275 6050
rect -2525 5912 -284 6010
tri -284 5912 -186 6010 sw
tri -186 5912 -88 6010 ne
rect -88 5912 266 6010
tri 266 5912 364 6010 sw
tri 364 5912 462 6010 ne
rect 462 5912 816 6010
tri 816 5912 914 6010 sw
tri 914 5912 1012 6010 ne
rect 1012 5912 1366 6010
tri 1366 5912 1464 6010 sw
tri 1464 5912 1562 6010 ne
rect 1562 5912 1916 6010
tri 1916 5912 2014 6010 sw
tri 2014 5912 2112 6010 ne
rect 2112 5912 2466 6010
tri 2466 5912 2564 6010 sw
tri 2564 5912 2662 6010 ne
rect 2662 5912 3016 6010
tri 3016 5912 3114 6010 sw
tri 3114 5912 3212 6010 ne
rect 3212 5912 3566 6010
tri 3566 5912 3664 6010 sw
tri 3664 5912 3762 6010 ne
rect 3762 5912 4116 6010
tri 4116 5912 4214 6010 sw
tri 4214 5912 4312 6010 ne
rect 4312 5912 4666 6010
tri 4666 5912 4764 6010 sw
tri 4764 5912 4862 6010 ne
rect 4862 5912 5216 6010
tri 5216 5912 5314 6010 sw
tri 5314 5912 5412 6010 ne
rect 5412 5912 5766 6010
tri 5766 5912 5864 6010 sw
tri 5864 5912 5962 6010 ne
rect 5962 5912 6316 6010
tri 6316 5912 6414 6010 sw
tri 6414 5912 6512 6010 ne
rect 6512 5912 6866 6010
tri 6866 5912 6964 6010 sw
tri 6964 5912 7062 6010 ne
rect 7062 5912 7416 6010
tri 7416 5912 7514 6010 sw
tri 7514 5912 7612 6010 ne
rect 7612 5912 7966 6010
tri 7966 5912 8064 6010 sw
tri 8064 5912 8162 6010 ne
rect 8162 5912 8516 6010
tri 8516 5912 8614 6010 sw
tri 8614 5912 8712 6010 ne
rect 8712 5912 9066 6010
tri 9066 5912 9164 6010 sw
tri 9164 5912 9262 6010 ne
rect 9262 5912 9616 6010
tri 9616 5912 9714 6010 sw
tri 9714 5912 9812 6010 ne
rect 9812 5912 10166 6010
tri 10166 5912 10264 6010 sw
tri 10264 5912 10362 6010 ne
rect 10362 5912 10716 6010
tri 10716 5912 10814 6010 sw
tri 10814 5912 10912 6010 ne
rect 10912 5912 11266 6010
tri 11266 5912 11364 6010 sw
tri 11364 5912 11462 6010 ne
rect 11462 5912 11816 6010
tri 11816 5912 11914 6010 sw
tri 11914 5912 12012 6010 ne
rect 12012 5912 12366 6010
tri 12366 5912 12464 6010 sw
tri 12464 5912 12562 6010 ne
rect 12562 5912 12916 6010
tri 12916 5912 13014 6010 sw
tri 13014 5912 13112 6010 ne
rect 13112 5912 13466 6010
tri 13466 5912 13564 6010 sw
tri 13564 5912 13662 6010 ne
rect 13662 5912 14275 6010
rect -2525 5814 -186 5912
tri -186 5814 -88 5912 sw
tri -88 5814 10 5912 ne
rect 10 5814 364 5912
tri 364 5814 462 5912 sw
tri 462 5814 560 5912 ne
rect 560 5814 914 5912
tri 914 5814 1012 5912 sw
tri 1012 5814 1110 5912 ne
rect 1110 5814 1464 5912
tri 1464 5814 1562 5912 sw
tri 1562 5814 1660 5912 ne
rect 1660 5814 2014 5912
tri 2014 5814 2112 5912 sw
tri 2112 5814 2210 5912 ne
rect 2210 5814 2564 5912
tri 2564 5814 2662 5912 sw
tri 2662 5814 2760 5912 ne
rect 2760 5814 3114 5912
tri 3114 5814 3212 5912 sw
tri 3212 5814 3310 5912 ne
rect 3310 5814 3664 5912
tri 3664 5814 3762 5912 sw
tri 3762 5814 3860 5912 ne
rect 3860 5814 4214 5912
tri 4214 5814 4312 5912 sw
tri 4312 5814 4410 5912 ne
rect 4410 5814 4764 5912
tri 4764 5814 4862 5912 sw
tri 4862 5814 4960 5912 ne
rect 4960 5814 5314 5912
tri 5314 5814 5412 5912 sw
tri 5412 5814 5510 5912 ne
rect 5510 5814 5864 5912
tri 5864 5814 5962 5912 sw
tri 5962 5814 6060 5912 ne
rect 6060 5814 6414 5912
tri 6414 5814 6512 5912 sw
tri 6512 5814 6610 5912 ne
rect 6610 5814 6964 5912
tri 6964 5814 7062 5912 sw
tri 7062 5814 7160 5912 ne
rect 7160 5814 7514 5912
tri 7514 5814 7612 5912 sw
tri 7612 5814 7710 5912 ne
rect 7710 5814 8064 5912
tri 8064 5814 8162 5912 sw
tri 8162 5814 8260 5912 ne
rect 8260 5814 8614 5912
tri 8614 5814 8712 5912 sw
tri 8712 5814 8810 5912 ne
rect 8810 5814 9164 5912
tri 9164 5814 9262 5912 sw
tri 9262 5814 9360 5912 ne
rect 9360 5814 9714 5912
tri 9714 5814 9812 5912 sw
tri 9812 5814 9910 5912 ne
rect 9910 5814 10264 5912
tri 10264 5814 10362 5912 sw
tri 10362 5814 10460 5912 ne
rect 10460 5814 10814 5912
tri 10814 5814 10912 5912 sw
tri 10912 5814 11010 5912 ne
rect 11010 5814 11364 5912
tri 11364 5814 11462 5912 sw
tri 11462 5814 11560 5912 ne
rect 11560 5814 11914 5912
tri 11914 5814 12012 5912 sw
tri 12012 5814 12110 5912 ne
rect 12110 5814 12464 5912
tri 12464 5814 12562 5912 sw
tri 12562 5814 12660 5912 ne
rect 12660 5814 13014 5912
tri 13014 5814 13112 5912 sw
tri 13112 5814 13210 5912 ne
rect 13210 5814 13564 5912
tri 13564 5814 13662 5912 sw
rect 14775 5814 15775 6462
rect -2525 5810 -88 5814
rect -2525 5690 -310 5810
rect -190 5726 -88 5810
tri -88 5726 0 5814 sw
tri 10 5726 98 5814 ne
rect 98 5810 462 5814
rect 98 5726 240 5810
rect -190 5690 0 5726
rect -2525 5686 0 5690
rect -2525 5038 -1525 5686
tri -412 5588 -314 5686 ne
rect -314 5638 0 5686
tri 0 5638 88 5726 sw
tri 98 5638 186 5726 ne
rect 186 5690 240 5726
rect 360 5726 462 5810
tri 462 5726 550 5814 sw
tri 560 5726 648 5814 ne
rect 648 5810 1012 5814
rect 648 5726 790 5810
rect 360 5690 550 5726
rect 186 5686 550 5690
tri 550 5686 590 5726 sw
tri 648 5686 688 5726 ne
rect 688 5690 790 5726
rect 910 5726 1012 5810
tri 1012 5726 1100 5814 sw
tri 1110 5726 1198 5814 ne
rect 1198 5810 1562 5814
rect 1198 5726 1340 5810
rect 910 5690 1100 5726
rect 688 5686 1100 5690
rect 186 5638 590 5686
rect -314 5588 88 5638
rect -1025 5500 -412 5588
tri -412 5500 -324 5588 sw
tri -314 5500 -226 5588 ne
rect -226 5558 88 5588
tri 88 5558 168 5638 sw
tri 186 5558 266 5638 ne
rect 266 5588 590 5638
tri 590 5588 688 5686 sw
tri 688 5588 786 5686 ne
rect 786 5638 1100 5686
tri 1100 5638 1188 5726 sw
tri 1198 5638 1286 5726 ne
rect 1286 5690 1340 5726
rect 1460 5726 1562 5810
tri 1562 5726 1650 5814 sw
tri 1660 5726 1748 5814 ne
rect 1748 5810 2112 5814
rect 1748 5726 1890 5810
rect 1460 5690 1650 5726
rect 1286 5686 1650 5690
tri 1650 5686 1690 5726 sw
tri 1748 5686 1788 5726 ne
rect 1788 5690 1890 5726
rect 2010 5726 2112 5810
tri 2112 5726 2200 5814 sw
tri 2210 5726 2298 5814 ne
rect 2298 5810 2662 5814
rect 2298 5726 2440 5810
rect 2010 5690 2200 5726
rect 1788 5686 2200 5690
rect 1286 5638 1690 5686
rect 786 5588 1188 5638
rect 266 5558 688 5588
rect -226 5500 168 5558
rect -1025 5460 -324 5500
tri -324 5460 -284 5500 sw
tri -226 5460 -186 5500 ne
rect -186 5460 168 5500
tri 168 5460 266 5558 sw
tri 266 5460 364 5558 ne
rect 364 5500 688 5558
tri 688 5500 776 5588 sw
tri 786 5500 874 5588 ne
rect 874 5558 1188 5588
tri 1188 5558 1268 5638 sw
tri 1286 5558 1366 5638 ne
rect 1366 5588 1690 5638
tri 1690 5588 1788 5686 sw
tri 1788 5588 1886 5686 ne
rect 1886 5638 2200 5686
tri 2200 5638 2288 5726 sw
tri 2298 5638 2386 5726 ne
rect 2386 5690 2440 5726
rect 2560 5726 2662 5810
tri 2662 5726 2750 5814 sw
tri 2760 5726 2848 5814 ne
rect 2848 5810 3212 5814
rect 2848 5726 2990 5810
rect 2560 5690 2750 5726
rect 2386 5686 2750 5690
tri 2750 5686 2790 5726 sw
tri 2848 5686 2888 5726 ne
rect 2888 5690 2990 5726
rect 3110 5726 3212 5810
tri 3212 5726 3300 5814 sw
tri 3310 5726 3398 5814 ne
rect 3398 5810 3762 5814
rect 3398 5726 3540 5810
rect 3110 5690 3300 5726
rect 2888 5686 3300 5690
rect 2386 5638 2790 5686
rect 1886 5588 2288 5638
rect 1366 5558 1788 5588
rect 874 5500 1268 5558
rect 364 5460 776 5500
tri 776 5460 816 5500 sw
tri 874 5460 914 5500 ne
rect 914 5460 1268 5500
tri 1268 5460 1366 5558 sw
tri 1366 5460 1464 5558 ne
rect 1464 5500 1788 5558
tri 1788 5500 1876 5588 sw
tri 1886 5500 1974 5588 ne
rect 1974 5558 2288 5588
tri 2288 5558 2368 5638 sw
tri 2386 5558 2466 5638 ne
rect 2466 5588 2790 5638
tri 2790 5588 2888 5686 sw
tri 2888 5588 2986 5686 ne
rect 2986 5638 3300 5686
tri 3300 5638 3388 5726 sw
tri 3398 5638 3486 5726 ne
rect 3486 5690 3540 5726
rect 3660 5726 3762 5810
tri 3762 5726 3850 5814 sw
tri 3860 5726 3948 5814 ne
rect 3948 5810 4312 5814
rect 3948 5726 4090 5810
rect 3660 5690 3850 5726
rect 3486 5686 3850 5690
tri 3850 5686 3890 5726 sw
tri 3948 5686 3988 5726 ne
rect 3988 5690 4090 5726
rect 4210 5726 4312 5810
tri 4312 5726 4400 5814 sw
tri 4410 5726 4498 5814 ne
rect 4498 5810 4862 5814
rect 4498 5726 4640 5810
rect 4210 5690 4400 5726
rect 3988 5686 4400 5690
rect 3486 5638 3890 5686
rect 2986 5588 3388 5638
rect 2466 5558 2888 5588
rect 1974 5500 2368 5558
rect 1464 5460 1876 5500
tri 1876 5460 1916 5500 sw
tri 1974 5460 2014 5500 ne
rect 2014 5460 2368 5500
tri 2368 5460 2466 5558 sw
tri 2466 5460 2564 5558 ne
rect 2564 5500 2888 5558
tri 2888 5500 2976 5588 sw
tri 2986 5500 3074 5588 ne
rect 3074 5558 3388 5588
tri 3388 5558 3468 5638 sw
tri 3486 5558 3566 5638 ne
rect 3566 5588 3890 5638
tri 3890 5588 3988 5686 sw
tri 3988 5588 4086 5686 ne
rect 4086 5638 4400 5686
tri 4400 5638 4488 5726 sw
tri 4498 5638 4586 5726 ne
rect 4586 5690 4640 5726
rect 4760 5726 4862 5810
tri 4862 5726 4950 5814 sw
tri 4960 5726 5048 5814 ne
rect 5048 5810 5412 5814
rect 5048 5726 5190 5810
rect 4760 5690 4950 5726
rect 4586 5686 4950 5690
tri 4950 5686 4990 5726 sw
tri 5048 5686 5088 5726 ne
rect 5088 5690 5190 5726
rect 5310 5726 5412 5810
tri 5412 5726 5500 5814 sw
tri 5510 5726 5598 5814 ne
rect 5598 5810 5962 5814
rect 5598 5726 5740 5810
rect 5310 5690 5500 5726
rect 5088 5686 5500 5690
rect 4586 5638 4990 5686
rect 4086 5588 4488 5638
rect 3566 5558 3988 5588
rect 3074 5500 3468 5558
rect 2564 5460 2976 5500
tri 2976 5460 3016 5500 sw
tri 3074 5460 3114 5500 ne
rect 3114 5460 3468 5500
tri 3468 5460 3566 5558 sw
tri 3566 5460 3664 5558 ne
rect 3664 5500 3988 5558
tri 3988 5500 4076 5588 sw
tri 4086 5500 4174 5588 ne
rect 4174 5558 4488 5588
tri 4488 5558 4568 5638 sw
tri 4586 5558 4666 5638 ne
rect 4666 5588 4990 5638
tri 4990 5588 5088 5686 sw
tri 5088 5588 5186 5686 ne
rect 5186 5638 5500 5686
tri 5500 5638 5588 5726 sw
tri 5598 5638 5686 5726 ne
rect 5686 5690 5740 5726
rect 5860 5726 5962 5810
tri 5962 5726 6050 5814 sw
tri 6060 5726 6148 5814 ne
rect 6148 5810 6512 5814
rect 6148 5726 6290 5810
rect 5860 5690 6050 5726
rect 5686 5686 6050 5690
tri 6050 5686 6090 5726 sw
tri 6148 5686 6188 5726 ne
rect 6188 5690 6290 5726
rect 6410 5726 6512 5810
tri 6512 5726 6600 5814 sw
tri 6610 5726 6698 5814 ne
rect 6698 5810 7062 5814
rect 6698 5726 6840 5810
rect 6410 5690 6600 5726
rect 6188 5686 6600 5690
rect 5686 5638 6090 5686
rect 5186 5588 5588 5638
rect 4666 5558 5088 5588
rect 4174 5500 4568 5558
rect 3664 5460 4076 5500
tri 4076 5460 4116 5500 sw
tri 4174 5460 4214 5500 ne
rect 4214 5460 4568 5500
tri 4568 5460 4666 5558 sw
tri 4666 5460 4764 5558 ne
rect 4764 5500 5088 5558
tri 5088 5500 5176 5588 sw
tri 5186 5500 5274 5588 ne
rect 5274 5558 5588 5588
tri 5588 5558 5668 5638 sw
tri 5686 5558 5766 5638 ne
rect 5766 5588 6090 5638
tri 6090 5588 6188 5686 sw
tri 6188 5588 6286 5686 ne
rect 6286 5638 6600 5686
tri 6600 5638 6688 5726 sw
tri 6698 5638 6786 5726 ne
rect 6786 5690 6840 5726
rect 6960 5726 7062 5810
tri 7062 5726 7150 5814 sw
tri 7160 5726 7248 5814 ne
rect 7248 5810 7612 5814
rect 7248 5726 7390 5810
rect 6960 5690 7150 5726
rect 6786 5686 7150 5690
tri 7150 5686 7190 5726 sw
tri 7248 5686 7288 5726 ne
rect 7288 5690 7390 5726
rect 7510 5726 7612 5810
tri 7612 5726 7700 5814 sw
tri 7710 5726 7798 5814 ne
rect 7798 5810 8162 5814
rect 7798 5726 7940 5810
rect 7510 5690 7700 5726
rect 7288 5686 7700 5690
rect 6786 5638 7190 5686
rect 6286 5588 6688 5638
rect 5766 5558 6188 5588
rect 5274 5500 5668 5558
rect 4764 5460 5176 5500
tri 5176 5460 5216 5500 sw
tri 5274 5460 5314 5500 ne
rect 5314 5460 5668 5500
tri 5668 5460 5766 5558 sw
tri 5766 5460 5864 5558 ne
rect 5864 5500 6188 5558
tri 6188 5500 6276 5588 sw
tri 6286 5500 6374 5588 ne
rect 6374 5558 6688 5588
tri 6688 5558 6768 5638 sw
tri 6786 5558 6866 5638 ne
rect 6866 5588 7190 5638
tri 7190 5588 7288 5686 sw
tri 7288 5588 7386 5686 ne
rect 7386 5638 7700 5686
tri 7700 5638 7788 5726 sw
tri 7798 5638 7886 5726 ne
rect 7886 5690 7940 5726
rect 8060 5726 8162 5810
tri 8162 5726 8250 5814 sw
tri 8260 5726 8348 5814 ne
rect 8348 5810 8712 5814
rect 8348 5726 8490 5810
rect 8060 5690 8250 5726
rect 7886 5686 8250 5690
tri 8250 5686 8290 5726 sw
tri 8348 5686 8388 5726 ne
rect 8388 5690 8490 5726
rect 8610 5726 8712 5810
tri 8712 5726 8800 5814 sw
tri 8810 5726 8898 5814 ne
rect 8898 5810 9262 5814
rect 8898 5726 9040 5810
rect 8610 5690 8800 5726
rect 8388 5686 8800 5690
rect 7886 5638 8290 5686
rect 7386 5588 7788 5638
rect 6866 5558 7288 5588
rect 6374 5500 6768 5558
rect 5864 5460 6276 5500
tri 6276 5460 6316 5500 sw
tri 6374 5460 6414 5500 ne
rect 6414 5460 6768 5500
tri 6768 5460 6866 5558 sw
tri 6866 5460 6964 5558 ne
rect 6964 5500 7288 5558
tri 7288 5500 7376 5588 sw
tri 7386 5500 7474 5588 ne
rect 7474 5558 7788 5588
tri 7788 5558 7868 5638 sw
tri 7886 5558 7966 5638 ne
rect 7966 5588 8290 5638
tri 8290 5588 8388 5686 sw
tri 8388 5588 8486 5686 ne
rect 8486 5638 8800 5686
tri 8800 5638 8888 5726 sw
tri 8898 5638 8986 5726 ne
rect 8986 5690 9040 5726
rect 9160 5726 9262 5810
tri 9262 5726 9350 5814 sw
tri 9360 5726 9448 5814 ne
rect 9448 5810 9812 5814
rect 9448 5726 9590 5810
rect 9160 5690 9350 5726
rect 8986 5686 9350 5690
tri 9350 5686 9390 5726 sw
tri 9448 5686 9488 5726 ne
rect 9488 5690 9590 5726
rect 9710 5726 9812 5810
tri 9812 5726 9900 5814 sw
tri 9910 5726 9998 5814 ne
rect 9998 5810 10362 5814
rect 9998 5726 10140 5810
rect 9710 5690 9900 5726
rect 9488 5686 9900 5690
rect 8986 5638 9390 5686
rect 8486 5588 8888 5638
rect 7966 5558 8388 5588
rect 7474 5500 7868 5558
rect 6964 5460 7376 5500
tri 7376 5460 7416 5500 sw
tri 7474 5460 7514 5500 ne
rect 7514 5460 7868 5500
tri 7868 5460 7966 5558 sw
tri 7966 5460 8064 5558 ne
rect 8064 5500 8388 5558
tri 8388 5500 8476 5588 sw
tri 8486 5500 8574 5588 ne
rect 8574 5558 8888 5588
tri 8888 5558 8968 5638 sw
tri 8986 5558 9066 5638 ne
rect 9066 5588 9390 5638
tri 9390 5588 9488 5686 sw
tri 9488 5588 9586 5686 ne
rect 9586 5638 9900 5686
tri 9900 5638 9988 5726 sw
tri 9998 5638 10086 5726 ne
rect 10086 5690 10140 5726
rect 10260 5726 10362 5810
tri 10362 5726 10450 5814 sw
tri 10460 5726 10548 5814 ne
rect 10548 5810 10912 5814
rect 10548 5726 10690 5810
rect 10260 5690 10450 5726
rect 10086 5686 10450 5690
tri 10450 5686 10490 5726 sw
tri 10548 5686 10588 5726 ne
rect 10588 5690 10690 5726
rect 10810 5726 10912 5810
tri 10912 5726 11000 5814 sw
tri 11010 5726 11098 5814 ne
rect 11098 5810 11462 5814
rect 11098 5726 11240 5810
rect 10810 5690 11000 5726
rect 10588 5686 11000 5690
rect 10086 5638 10490 5686
rect 9586 5588 9988 5638
rect 9066 5558 9488 5588
rect 8574 5500 8968 5558
rect 8064 5460 8476 5500
tri 8476 5460 8516 5500 sw
tri 8574 5460 8614 5500 ne
rect 8614 5460 8968 5500
tri 8968 5460 9066 5558 sw
tri 9066 5460 9164 5558 ne
rect 9164 5500 9488 5558
tri 9488 5500 9576 5588 sw
tri 9586 5500 9674 5588 ne
rect 9674 5558 9988 5588
tri 9988 5558 10068 5638 sw
tri 10086 5558 10166 5638 ne
rect 10166 5588 10490 5638
tri 10490 5588 10588 5686 sw
tri 10588 5588 10686 5686 ne
rect 10686 5638 11000 5686
tri 11000 5638 11088 5726 sw
tri 11098 5638 11186 5726 ne
rect 11186 5690 11240 5726
rect 11360 5726 11462 5810
tri 11462 5726 11550 5814 sw
tri 11560 5726 11648 5814 ne
rect 11648 5810 12012 5814
rect 11648 5726 11790 5810
rect 11360 5690 11550 5726
rect 11186 5686 11550 5690
tri 11550 5686 11590 5726 sw
tri 11648 5686 11688 5726 ne
rect 11688 5690 11790 5726
rect 11910 5726 12012 5810
tri 12012 5726 12100 5814 sw
tri 12110 5726 12198 5814 ne
rect 12198 5810 12562 5814
rect 12198 5726 12340 5810
rect 11910 5690 12100 5726
rect 11688 5686 12100 5690
rect 11186 5638 11590 5686
rect 10686 5588 11088 5638
rect 10166 5558 10588 5588
rect 9674 5500 10068 5558
rect 9164 5460 9576 5500
tri 9576 5460 9616 5500 sw
tri 9674 5460 9714 5500 ne
rect 9714 5460 10068 5500
tri 10068 5460 10166 5558 sw
tri 10166 5460 10264 5558 ne
rect 10264 5500 10588 5558
tri 10588 5500 10676 5588 sw
tri 10686 5500 10774 5588 ne
rect 10774 5558 11088 5588
tri 11088 5558 11168 5638 sw
tri 11186 5558 11266 5638 ne
rect 11266 5588 11590 5638
tri 11590 5588 11688 5686 sw
tri 11688 5588 11786 5686 ne
rect 11786 5638 12100 5686
tri 12100 5638 12188 5726 sw
tri 12198 5638 12286 5726 ne
rect 12286 5690 12340 5726
rect 12460 5726 12562 5810
tri 12562 5726 12650 5814 sw
tri 12660 5726 12748 5814 ne
rect 12748 5810 13112 5814
rect 12748 5726 12890 5810
rect 12460 5690 12650 5726
rect 12286 5686 12650 5690
tri 12650 5686 12690 5726 sw
tri 12748 5686 12788 5726 ne
rect 12788 5690 12890 5726
rect 13010 5726 13112 5810
tri 13112 5726 13200 5814 sw
tri 13210 5726 13298 5814 ne
rect 13298 5810 15775 5814
rect 13298 5726 13440 5810
rect 13010 5690 13200 5726
rect 12788 5686 13200 5690
rect 12286 5638 12690 5686
rect 11786 5588 12188 5638
rect 11266 5558 11688 5588
rect 10774 5500 11168 5558
rect 10264 5460 10676 5500
tri 10676 5460 10716 5500 sw
tri 10774 5460 10814 5500 ne
rect 10814 5460 11168 5500
tri 11168 5460 11266 5558 sw
tri 11266 5460 11364 5558 ne
rect 11364 5500 11688 5558
tri 11688 5500 11776 5588 sw
tri 11786 5500 11874 5588 ne
rect 11874 5558 12188 5588
tri 12188 5558 12268 5638 sw
tri 12286 5558 12366 5638 ne
rect 12366 5588 12690 5638
tri 12690 5588 12788 5686 sw
tri 12788 5588 12886 5686 ne
rect 12886 5638 13200 5686
tri 13200 5638 13288 5726 sw
tri 13298 5638 13386 5726 ne
rect 13386 5690 13440 5726
rect 13560 5690 15775 5810
rect 13386 5638 15775 5690
rect 12886 5588 13288 5638
rect 12366 5558 12788 5588
rect 11874 5500 12268 5558
rect 11364 5460 11776 5500
tri 11776 5460 11816 5500 sw
tri 11874 5460 11914 5500 ne
rect 11914 5460 12268 5500
tri 12268 5460 12366 5558 sw
tri 12366 5460 12464 5558 ne
rect 12464 5500 12788 5558
tri 12788 5500 12876 5588 sw
tri 12886 5500 12974 5588 ne
rect 12974 5558 13288 5588
tri 13288 5558 13368 5638 sw
tri 13386 5558 13466 5638 ne
rect 13466 5558 14075 5638
rect 12974 5500 13368 5558
rect 12464 5460 12876 5500
tri 12876 5460 12916 5500 sw
tri 12974 5460 13014 5500 ne
rect 13014 5460 13368 5500
tri 13368 5460 13466 5558 sw
tri 13466 5460 13564 5558 ne
rect 13564 5538 14075 5558
rect 14175 5538 15775 5638
rect 13564 5460 15775 5538
rect -1025 5412 -284 5460
rect -1025 5312 -925 5412
rect -825 5362 -284 5412
tri -284 5362 -186 5460 sw
tri -186 5362 -88 5460 ne
rect -88 5362 266 5460
tri 266 5362 364 5460 sw
tri 364 5362 462 5460 ne
rect 462 5362 816 5460
tri 816 5362 914 5460 sw
tri 914 5362 1012 5460 ne
rect 1012 5362 1366 5460
tri 1366 5362 1464 5460 sw
tri 1464 5362 1562 5460 ne
rect 1562 5362 1916 5460
tri 1916 5362 2014 5460 sw
tri 2014 5362 2112 5460 ne
rect 2112 5362 2466 5460
tri 2466 5362 2564 5460 sw
tri 2564 5362 2662 5460 ne
rect 2662 5362 3016 5460
tri 3016 5362 3114 5460 sw
tri 3114 5362 3212 5460 ne
rect 3212 5362 3566 5460
tri 3566 5362 3664 5460 sw
tri 3664 5362 3762 5460 ne
rect 3762 5362 4116 5460
tri 4116 5362 4214 5460 sw
tri 4214 5362 4312 5460 ne
rect 4312 5362 4666 5460
tri 4666 5362 4764 5460 sw
tri 4764 5362 4862 5460 ne
rect 4862 5362 5216 5460
tri 5216 5362 5314 5460 sw
tri 5314 5362 5412 5460 ne
rect 5412 5362 5766 5460
tri 5766 5362 5864 5460 sw
tri 5864 5362 5962 5460 ne
rect 5962 5362 6316 5460
tri 6316 5362 6414 5460 sw
tri 6414 5362 6512 5460 ne
rect 6512 5362 6866 5460
tri 6866 5362 6964 5460 sw
tri 6964 5362 7062 5460 ne
rect 7062 5362 7416 5460
tri 7416 5362 7514 5460 sw
tri 7514 5362 7612 5460 ne
rect 7612 5362 7966 5460
tri 7966 5362 8064 5460 sw
tri 8064 5362 8162 5460 ne
rect 8162 5362 8516 5460
tri 8516 5362 8614 5460 sw
tri 8614 5362 8712 5460 ne
rect 8712 5362 9066 5460
tri 9066 5362 9164 5460 sw
tri 9164 5362 9262 5460 ne
rect 9262 5362 9616 5460
tri 9616 5362 9714 5460 sw
tri 9714 5362 9812 5460 ne
rect 9812 5362 10166 5460
tri 10166 5362 10264 5460 sw
tri 10264 5362 10362 5460 ne
rect 10362 5362 10716 5460
tri 10716 5362 10814 5460 sw
tri 10814 5362 10912 5460 ne
rect 10912 5362 11266 5460
tri 11266 5362 11364 5460 sw
tri 11364 5362 11462 5460 ne
rect 11462 5362 11816 5460
tri 11816 5362 11914 5460 sw
tri 11914 5362 12012 5460 ne
rect 12012 5362 12366 5460
tri 12366 5362 12464 5460 sw
tri 12464 5362 12562 5460 ne
rect 12562 5362 12916 5460
tri 12916 5362 13014 5460 sw
tri 13014 5362 13112 5460 ne
rect 13112 5362 13466 5460
tri 13466 5362 13564 5460 sw
tri 13564 5362 13662 5460 ne
rect 13662 5362 15775 5460
rect -825 5312 -186 5362
rect -1025 5264 -186 5312
tri -186 5264 -88 5362 sw
tri -88 5264 10 5362 ne
rect 10 5264 364 5362
tri 364 5264 462 5362 sw
tri 462 5264 560 5362 ne
rect 560 5264 914 5362
tri 914 5264 1012 5362 sw
tri 1012 5264 1110 5362 ne
rect 1110 5264 1464 5362
tri 1464 5264 1562 5362 sw
tri 1562 5264 1660 5362 ne
rect 1660 5264 2014 5362
tri 2014 5264 2112 5362 sw
tri 2112 5264 2210 5362 ne
rect 2210 5264 2564 5362
tri 2564 5264 2662 5362 sw
tri 2662 5264 2760 5362 ne
rect 2760 5264 3114 5362
tri 3114 5264 3212 5362 sw
tri 3212 5264 3310 5362 ne
rect 3310 5264 3664 5362
tri 3664 5264 3762 5362 sw
tri 3762 5264 3860 5362 ne
rect 3860 5264 4214 5362
tri 4214 5264 4312 5362 sw
tri 4312 5264 4410 5362 ne
rect 4410 5264 4764 5362
tri 4764 5264 4862 5362 sw
tri 4862 5264 4960 5362 ne
rect 4960 5264 5314 5362
tri 5314 5264 5412 5362 sw
tri 5412 5264 5510 5362 ne
rect 5510 5264 5864 5362
tri 5864 5264 5962 5362 sw
tri 5962 5264 6060 5362 ne
rect 6060 5264 6414 5362
tri 6414 5264 6512 5362 sw
tri 6512 5264 6610 5362 ne
rect 6610 5264 6964 5362
tri 6964 5264 7062 5362 sw
tri 7062 5264 7160 5362 ne
rect 7160 5264 7514 5362
tri 7514 5264 7612 5362 sw
tri 7612 5264 7710 5362 ne
rect 7710 5264 8064 5362
tri 8064 5264 8162 5362 sw
tri 8162 5264 8260 5362 ne
rect 8260 5264 8614 5362
tri 8614 5264 8712 5362 sw
tri 8712 5264 8810 5362 ne
rect 8810 5264 9164 5362
tri 9164 5264 9262 5362 sw
tri 9262 5264 9360 5362 ne
rect 9360 5264 9714 5362
tri 9714 5264 9812 5362 sw
tri 9812 5264 9910 5362 ne
rect 9910 5264 10264 5362
tri 10264 5264 10362 5362 sw
tri 10362 5264 10460 5362 ne
rect 10460 5264 10814 5362
tri 10814 5264 10912 5362 sw
tri 10912 5264 11010 5362 ne
rect 11010 5264 11364 5362
tri 11364 5264 11462 5362 sw
tri 11462 5264 11560 5362 ne
rect 11560 5264 11914 5362
tri 11914 5264 12012 5362 sw
tri 12012 5264 12110 5362 ne
rect 12110 5264 12464 5362
tri 12464 5264 12562 5362 sw
tri 12562 5264 12660 5362 ne
rect 12660 5264 13014 5362
tri 13014 5264 13112 5362 sw
tri 13112 5264 13210 5362 ne
rect 13210 5264 13564 5362
tri 13564 5264 13662 5362 sw
rect -1025 5260 -88 5264
rect -1025 5140 -310 5260
rect -190 5176 -88 5260
tri -88 5176 0 5264 sw
tri 10 5176 98 5264 ne
rect 98 5260 462 5264
rect 98 5176 240 5260
rect -190 5140 0 5176
rect -1025 5136 0 5140
tri 0 5136 40 5176 sw
tri 98 5136 138 5176 ne
rect 138 5140 240 5176
rect 360 5176 462 5260
tri 462 5176 550 5264 sw
tri 560 5176 648 5264 ne
rect 648 5260 1012 5264
rect 648 5176 790 5260
rect 360 5140 550 5176
rect 138 5136 550 5140
tri -412 5038 -314 5136 ne
rect -314 5038 40 5136
tri 40 5038 138 5136 sw
tri 138 5038 236 5136 ne
rect 236 5088 550 5136
tri 550 5088 638 5176 sw
tri 648 5088 736 5176 ne
rect 736 5140 790 5176
rect 910 5176 1012 5260
tri 1012 5176 1100 5264 sw
tri 1110 5176 1198 5264 ne
rect 1198 5260 1562 5264
rect 1198 5176 1340 5260
rect 910 5140 1100 5176
rect 736 5136 1100 5140
tri 1100 5136 1140 5176 sw
tri 1198 5136 1238 5176 ne
rect 1238 5140 1340 5176
rect 1460 5176 1562 5260
tri 1562 5176 1650 5264 sw
tri 1660 5176 1748 5264 ne
rect 1748 5260 2112 5264
rect 1748 5176 1890 5260
rect 1460 5140 1650 5176
rect 1238 5136 1650 5140
rect 736 5088 1140 5136
rect 236 5038 638 5088
rect -2525 4950 -412 5038
tri -412 4950 -324 5038 sw
tri -314 4950 -226 5038 ne
rect -226 4950 138 5038
tri 138 4950 226 5038 sw
tri 236 4950 324 5038 ne
rect 324 5008 638 5038
tri 638 5008 718 5088 sw
tri 736 5008 816 5088 ne
rect 816 5038 1140 5088
tri 1140 5038 1238 5136 sw
tri 1238 5038 1336 5136 ne
rect 1336 5088 1650 5136
tri 1650 5088 1738 5176 sw
tri 1748 5088 1836 5176 ne
rect 1836 5140 1890 5176
rect 2010 5176 2112 5260
tri 2112 5176 2200 5264 sw
tri 2210 5176 2298 5264 ne
rect 2298 5260 2662 5264
rect 2298 5176 2440 5260
rect 2010 5140 2200 5176
rect 1836 5136 2200 5140
tri 2200 5136 2240 5176 sw
tri 2298 5136 2338 5176 ne
rect 2338 5140 2440 5176
rect 2560 5176 2662 5260
tri 2662 5176 2750 5264 sw
tri 2760 5176 2848 5264 ne
rect 2848 5260 3212 5264
rect 2848 5176 2990 5260
rect 2560 5140 2750 5176
rect 2338 5136 2750 5140
rect 1836 5088 2240 5136
rect 1336 5038 1738 5088
rect 816 5008 1238 5038
rect 324 4950 718 5008
rect -2525 4910 -324 4950
tri -324 4910 -284 4950 sw
tri -226 4910 -186 4950 ne
rect -186 4910 226 4950
tri 226 4910 266 4950 sw
tri 324 4910 364 4950 ne
rect 364 4910 718 4950
tri 718 4910 816 5008 sw
tri 816 4910 914 5008 ne
rect 914 4950 1238 5008
tri 1238 4950 1326 5038 sw
tri 1336 4950 1424 5038 ne
rect 1424 5008 1738 5038
tri 1738 5008 1818 5088 sw
tri 1836 5008 1916 5088 ne
rect 1916 5038 2240 5088
tri 2240 5038 2338 5136 sw
tri 2338 5038 2436 5136 ne
rect 2436 5088 2750 5136
tri 2750 5088 2838 5176 sw
tri 2848 5088 2936 5176 ne
rect 2936 5140 2990 5176
rect 3110 5176 3212 5260
tri 3212 5176 3300 5264 sw
tri 3310 5176 3398 5264 ne
rect 3398 5260 3762 5264
rect 3398 5176 3540 5260
rect 3110 5140 3300 5176
rect 2936 5136 3300 5140
tri 3300 5136 3340 5176 sw
tri 3398 5136 3438 5176 ne
rect 3438 5140 3540 5176
rect 3660 5176 3762 5260
tri 3762 5176 3850 5264 sw
tri 3860 5176 3948 5264 ne
rect 3948 5260 4312 5264
rect 3948 5176 4090 5260
rect 3660 5140 3850 5176
rect 3438 5136 3850 5140
rect 2936 5088 3340 5136
rect 2436 5038 2838 5088
rect 1916 5008 2338 5038
rect 1424 4950 1818 5008
rect 914 4910 1326 4950
tri 1326 4910 1366 4950 sw
tri 1424 4910 1464 4950 ne
rect 1464 4910 1818 4950
tri 1818 4910 1916 5008 sw
tri 1916 4910 2014 5008 ne
rect 2014 4950 2338 5008
tri 2338 4950 2426 5038 sw
tri 2436 4950 2524 5038 ne
rect 2524 5008 2838 5038
tri 2838 5008 2918 5088 sw
tri 2936 5008 3016 5088 ne
rect 3016 5038 3340 5088
tri 3340 5038 3438 5136 sw
tri 3438 5038 3536 5136 ne
rect 3536 5088 3850 5136
tri 3850 5088 3938 5176 sw
tri 3948 5088 4036 5176 ne
rect 4036 5140 4090 5176
rect 4210 5176 4312 5260
tri 4312 5176 4400 5264 sw
tri 4410 5176 4498 5264 ne
rect 4498 5260 4862 5264
rect 4498 5176 4640 5260
rect 4210 5140 4400 5176
rect 4036 5136 4400 5140
tri 4400 5136 4440 5176 sw
tri 4498 5136 4538 5176 ne
rect 4538 5140 4640 5176
rect 4760 5176 4862 5260
tri 4862 5176 4950 5264 sw
tri 4960 5176 5048 5264 ne
rect 5048 5260 5412 5264
rect 5048 5176 5190 5260
rect 4760 5140 4950 5176
rect 4538 5136 4950 5140
rect 4036 5088 4440 5136
rect 3536 5038 3938 5088
rect 3016 5008 3438 5038
rect 2524 4950 2918 5008
rect 2014 4910 2426 4950
tri 2426 4910 2466 4950 sw
tri 2524 4910 2564 4950 ne
rect 2564 4910 2918 4950
tri 2918 4910 3016 5008 sw
tri 3016 4910 3114 5008 ne
rect 3114 4950 3438 5008
tri 3438 4950 3526 5038 sw
tri 3536 4950 3624 5038 ne
rect 3624 5008 3938 5038
tri 3938 5008 4018 5088 sw
tri 4036 5008 4116 5088 ne
rect 4116 5038 4440 5088
tri 4440 5038 4538 5136 sw
tri 4538 5038 4636 5136 ne
rect 4636 5088 4950 5136
tri 4950 5088 5038 5176 sw
tri 5048 5088 5136 5176 ne
rect 5136 5140 5190 5176
rect 5310 5176 5412 5260
tri 5412 5176 5500 5264 sw
tri 5510 5176 5598 5264 ne
rect 5598 5260 5962 5264
rect 5598 5176 5740 5260
rect 5310 5140 5500 5176
rect 5136 5136 5500 5140
tri 5500 5136 5540 5176 sw
tri 5598 5136 5638 5176 ne
rect 5638 5140 5740 5176
rect 5860 5176 5962 5260
tri 5962 5176 6050 5264 sw
tri 6060 5176 6148 5264 ne
rect 6148 5260 6512 5264
rect 6148 5176 6290 5260
rect 5860 5140 6050 5176
rect 5638 5136 6050 5140
rect 5136 5088 5540 5136
rect 4636 5038 5038 5088
rect 4116 5008 4538 5038
rect 3624 4950 4018 5008
rect 3114 4910 3526 4950
tri 3526 4910 3566 4950 sw
tri 3624 4910 3664 4950 ne
rect 3664 4910 4018 4950
tri 4018 4910 4116 5008 sw
tri 4116 4910 4214 5008 ne
rect 4214 4950 4538 5008
tri 4538 4950 4626 5038 sw
tri 4636 4950 4724 5038 ne
rect 4724 5008 5038 5038
tri 5038 5008 5118 5088 sw
tri 5136 5008 5216 5088 ne
rect 5216 5038 5540 5088
tri 5540 5038 5638 5136 sw
tri 5638 5038 5736 5136 ne
rect 5736 5088 6050 5136
tri 6050 5088 6138 5176 sw
tri 6148 5088 6236 5176 ne
rect 6236 5140 6290 5176
rect 6410 5176 6512 5260
tri 6512 5176 6600 5264 sw
tri 6610 5176 6698 5264 ne
rect 6698 5260 7062 5264
rect 6698 5176 6840 5260
rect 6410 5140 6600 5176
rect 6236 5136 6600 5140
tri 6600 5136 6640 5176 sw
tri 6698 5136 6738 5176 ne
rect 6738 5140 6840 5176
rect 6960 5176 7062 5260
tri 7062 5176 7150 5264 sw
tri 7160 5176 7248 5264 ne
rect 7248 5260 7612 5264
rect 7248 5176 7390 5260
rect 6960 5140 7150 5176
rect 6738 5136 7150 5140
rect 6236 5088 6640 5136
rect 5736 5038 6138 5088
rect 5216 5008 5638 5038
rect 4724 4950 5118 5008
rect 4214 4910 4626 4950
tri 4626 4910 4666 4950 sw
tri 4724 4910 4764 4950 ne
rect 4764 4910 5118 4950
tri 5118 4910 5216 5008 sw
tri 5216 4910 5314 5008 ne
rect 5314 4950 5638 5008
tri 5638 4950 5726 5038 sw
tri 5736 4950 5824 5038 ne
rect 5824 5008 6138 5038
tri 6138 5008 6218 5088 sw
tri 6236 5008 6316 5088 ne
rect 6316 5038 6640 5088
tri 6640 5038 6738 5136 sw
tri 6738 5038 6836 5136 ne
rect 6836 5088 7150 5136
tri 7150 5088 7238 5176 sw
tri 7248 5088 7336 5176 ne
rect 7336 5140 7390 5176
rect 7510 5176 7612 5260
tri 7612 5176 7700 5264 sw
tri 7710 5176 7798 5264 ne
rect 7798 5260 8162 5264
rect 7798 5176 7940 5260
rect 7510 5140 7700 5176
rect 7336 5136 7700 5140
tri 7700 5136 7740 5176 sw
tri 7798 5136 7838 5176 ne
rect 7838 5140 7940 5176
rect 8060 5176 8162 5260
tri 8162 5176 8250 5264 sw
tri 8260 5176 8348 5264 ne
rect 8348 5260 8712 5264
rect 8348 5176 8490 5260
rect 8060 5140 8250 5176
rect 7838 5136 8250 5140
rect 7336 5088 7740 5136
rect 6836 5038 7238 5088
rect 6316 5008 6738 5038
rect 5824 4950 6218 5008
rect 5314 4910 5726 4950
tri 5726 4910 5766 4950 sw
tri 5824 4910 5864 4950 ne
rect 5864 4910 6218 4950
tri 6218 4910 6316 5008 sw
tri 6316 4910 6414 5008 ne
rect 6414 4950 6738 5008
tri 6738 4950 6826 5038 sw
tri 6836 4950 6924 5038 ne
rect 6924 5008 7238 5038
tri 7238 5008 7318 5088 sw
tri 7336 5008 7416 5088 ne
rect 7416 5038 7740 5088
tri 7740 5038 7838 5136 sw
tri 7838 5038 7936 5136 ne
rect 7936 5088 8250 5136
tri 8250 5088 8338 5176 sw
tri 8348 5088 8436 5176 ne
rect 8436 5140 8490 5176
rect 8610 5176 8712 5260
tri 8712 5176 8800 5264 sw
tri 8810 5176 8898 5264 ne
rect 8898 5260 9262 5264
rect 8898 5176 9040 5260
rect 8610 5140 8800 5176
rect 8436 5136 8800 5140
tri 8800 5136 8840 5176 sw
tri 8898 5136 8938 5176 ne
rect 8938 5140 9040 5176
rect 9160 5176 9262 5260
tri 9262 5176 9350 5264 sw
tri 9360 5176 9448 5264 ne
rect 9448 5260 9812 5264
rect 9448 5176 9590 5260
rect 9160 5140 9350 5176
rect 8938 5136 9350 5140
rect 8436 5088 8840 5136
rect 7936 5038 8338 5088
rect 7416 5008 7838 5038
rect 6924 4950 7318 5008
rect 6414 4910 6826 4950
tri 6826 4910 6866 4950 sw
tri 6924 4910 6964 4950 ne
rect 6964 4910 7318 4950
tri 7318 4910 7416 5008 sw
tri 7416 4910 7514 5008 ne
rect 7514 4950 7838 5008
tri 7838 4950 7926 5038 sw
tri 7936 4950 8024 5038 ne
rect 8024 5008 8338 5038
tri 8338 5008 8418 5088 sw
tri 8436 5008 8516 5088 ne
rect 8516 5038 8840 5088
tri 8840 5038 8938 5136 sw
tri 8938 5038 9036 5136 ne
rect 9036 5088 9350 5136
tri 9350 5088 9438 5176 sw
tri 9448 5088 9536 5176 ne
rect 9536 5140 9590 5176
rect 9710 5176 9812 5260
tri 9812 5176 9900 5264 sw
tri 9910 5176 9998 5264 ne
rect 9998 5260 10362 5264
rect 9998 5176 10140 5260
rect 9710 5140 9900 5176
rect 9536 5136 9900 5140
tri 9900 5136 9940 5176 sw
tri 9998 5136 10038 5176 ne
rect 10038 5140 10140 5176
rect 10260 5176 10362 5260
tri 10362 5176 10450 5264 sw
tri 10460 5176 10548 5264 ne
rect 10548 5260 10912 5264
rect 10548 5176 10690 5260
rect 10260 5140 10450 5176
rect 10038 5136 10450 5140
rect 9536 5088 9940 5136
rect 9036 5038 9438 5088
rect 8516 5008 8938 5038
rect 8024 4950 8418 5008
rect 7514 4910 7926 4950
tri 7926 4910 7966 4950 sw
tri 8024 4910 8064 4950 ne
rect 8064 4910 8418 4950
tri 8418 4910 8516 5008 sw
tri 8516 4910 8614 5008 ne
rect 8614 4950 8938 5008
tri 8938 4950 9026 5038 sw
tri 9036 4950 9124 5038 ne
rect 9124 5008 9438 5038
tri 9438 5008 9518 5088 sw
tri 9536 5008 9616 5088 ne
rect 9616 5038 9940 5088
tri 9940 5038 10038 5136 sw
tri 10038 5038 10136 5136 ne
rect 10136 5088 10450 5136
tri 10450 5088 10538 5176 sw
tri 10548 5088 10636 5176 ne
rect 10636 5140 10690 5176
rect 10810 5176 10912 5260
tri 10912 5176 11000 5264 sw
tri 11010 5176 11098 5264 ne
rect 11098 5260 11462 5264
rect 11098 5176 11240 5260
rect 10810 5140 11000 5176
rect 10636 5136 11000 5140
tri 11000 5136 11040 5176 sw
tri 11098 5136 11138 5176 ne
rect 11138 5140 11240 5176
rect 11360 5176 11462 5260
tri 11462 5176 11550 5264 sw
tri 11560 5176 11648 5264 ne
rect 11648 5260 12012 5264
rect 11648 5176 11790 5260
rect 11360 5140 11550 5176
rect 11138 5136 11550 5140
rect 10636 5088 11040 5136
rect 10136 5038 10538 5088
rect 9616 5008 10038 5038
rect 9124 4950 9518 5008
rect 8614 4910 9026 4950
tri 9026 4910 9066 4950 sw
tri 9124 4910 9164 4950 ne
rect 9164 4910 9518 4950
tri 9518 4910 9616 5008 sw
tri 9616 4910 9714 5008 ne
rect 9714 4950 10038 5008
tri 10038 4950 10126 5038 sw
tri 10136 4950 10224 5038 ne
rect 10224 5008 10538 5038
tri 10538 5008 10618 5088 sw
tri 10636 5008 10716 5088 ne
rect 10716 5038 11040 5088
tri 11040 5038 11138 5136 sw
tri 11138 5038 11236 5136 ne
rect 11236 5088 11550 5136
tri 11550 5088 11638 5176 sw
tri 11648 5088 11736 5176 ne
rect 11736 5140 11790 5176
rect 11910 5176 12012 5260
tri 12012 5176 12100 5264 sw
tri 12110 5176 12198 5264 ne
rect 12198 5260 12562 5264
rect 12198 5176 12340 5260
rect 11910 5140 12100 5176
rect 11736 5136 12100 5140
tri 12100 5136 12140 5176 sw
tri 12198 5136 12238 5176 ne
rect 12238 5140 12340 5176
rect 12460 5176 12562 5260
tri 12562 5176 12650 5264 sw
tri 12660 5176 12748 5264 ne
rect 12748 5260 13112 5264
rect 12748 5176 12890 5260
rect 12460 5140 12650 5176
rect 12238 5136 12650 5140
rect 11736 5088 12140 5136
rect 11236 5038 11638 5088
rect 10716 5008 11138 5038
rect 10224 4950 10618 5008
rect 9714 4910 10126 4950
tri 10126 4910 10166 4950 sw
tri 10224 4910 10264 4950 ne
rect 10264 4910 10618 4950
tri 10618 4910 10716 5008 sw
tri 10716 4910 10814 5008 ne
rect 10814 4950 11138 5008
tri 11138 4950 11226 5038 sw
tri 11236 4950 11324 5038 ne
rect 11324 5008 11638 5038
tri 11638 5008 11718 5088 sw
tri 11736 5008 11816 5088 ne
rect 11816 5038 12140 5088
tri 12140 5038 12238 5136 sw
tri 12238 5038 12336 5136 ne
rect 12336 5088 12650 5136
tri 12650 5088 12738 5176 sw
tri 12748 5088 12836 5176 ne
rect 12836 5140 12890 5176
rect 13010 5176 13112 5260
tri 13112 5176 13200 5264 sw
tri 13210 5176 13298 5264 ne
rect 13298 5260 14275 5264
rect 13298 5176 13440 5260
rect 13010 5140 13200 5176
rect 12836 5136 13200 5140
tri 13200 5136 13240 5176 sw
tri 13298 5136 13338 5176 ne
rect 13338 5140 13440 5176
rect 13560 5140 14275 5260
rect 13338 5136 14275 5140
rect 12836 5088 13240 5136
rect 12336 5038 12738 5088
rect 11816 5008 12238 5038
rect 11324 4950 11718 5008
rect 10814 4910 11226 4950
tri 11226 4910 11266 4950 sw
tri 11324 4910 11364 4950 ne
rect 11364 4910 11718 4950
tri 11718 4910 11816 5008 sw
tri 11816 4910 11914 5008 ne
rect 11914 4950 12238 5008
tri 12238 4950 12326 5038 sw
tri 12336 4950 12424 5038 ne
rect 12424 5008 12738 5038
tri 12738 5008 12818 5088 sw
tri 12836 5008 12916 5088 ne
rect 12916 5038 13240 5088
tri 13240 5038 13338 5136 sw
tri 13338 5038 13436 5136 ne
rect 13436 5038 14275 5136
rect 12916 5008 13338 5038
rect 12424 4950 12818 5008
rect 11914 4910 12326 4950
tri 12326 4910 12366 4950 sw
tri 12424 4910 12464 4950 ne
rect 12464 4910 12818 4950
tri 12818 4910 12916 5008 sw
tri 12916 4910 13014 5008 ne
rect 13014 4950 13338 5008
tri 13338 4950 13426 5038 sw
tri 13436 4950 13524 5038 ne
rect 13524 4950 14275 5038
rect 13014 4910 13426 4950
tri 13426 4910 13466 4950 sw
tri 13524 4910 13564 4950 ne
rect 13564 4910 14275 4950
rect -2525 4812 -284 4910
tri -284 4812 -186 4910 sw
tri -186 4812 -88 4910 ne
rect -88 4812 266 4910
tri 266 4812 364 4910 sw
tri 364 4812 462 4910 ne
rect 462 4812 816 4910
tri 816 4812 914 4910 sw
tri 914 4812 1012 4910 ne
rect 1012 4812 1366 4910
tri 1366 4812 1464 4910 sw
tri 1464 4812 1562 4910 ne
rect 1562 4812 1916 4910
tri 1916 4812 2014 4910 sw
tri 2014 4812 2112 4910 ne
rect 2112 4812 2466 4910
tri 2466 4812 2564 4910 sw
tri 2564 4812 2662 4910 ne
rect 2662 4812 3016 4910
tri 3016 4812 3114 4910 sw
tri 3114 4812 3212 4910 ne
rect 3212 4812 3566 4910
tri 3566 4812 3664 4910 sw
tri 3664 4812 3762 4910 ne
rect 3762 4812 4116 4910
tri 4116 4812 4214 4910 sw
tri 4214 4812 4312 4910 ne
rect 4312 4812 4666 4910
tri 4666 4812 4764 4910 sw
tri 4764 4812 4862 4910 ne
rect 4862 4812 5216 4910
tri 5216 4812 5314 4910 sw
tri 5314 4812 5412 4910 ne
rect 5412 4812 5766 4910
tri 5766 4812 5864 4910 sw
tri 5864 4812 5962 4910 ne
rect 5962 4812 6316 4910
tri 6316 4812 6414 4910 sw
tri 6414 4812 6512 4910 ne
rect 6512 4812 6866 4910
tri 6866 4812 6964 4910 sw
tri 6964 4812 7062 4910 ne
rect 7062 4812 7416 4910
tri 7416 4812 7514 4910 sw
tri 7514 4812 7612 4910 ne
rect 7612 4812 7966 4910
tri 7966 4812 8064 4910 sw
tri 8064 4812 8162 4910 ne
rect 8162 4812 8516 4910
tri 8516 4812 8614 4910 sw
tri 8614 4812 8712 4910 ne
rect 8712 4812 9066 4910
tri 9066 4812 9164 4910 sw
tri 9164 4812 9262 4910 ne
rect 9262 4812 9616 4910
tri 9616 4812 9714 4910 sw
tri 9714 4812 9812 4910 ne
rect 9812 4812 10166 4910
tri 10166 4812 10264 4910 sw
tri 10264 4812 10362 4910 ne
rect 10362 4812 10716 4910
tri 10716 4812 10814 4910 sw
tri 10814 4812 10912 4910 ne
rect 10912 4812 11266 4910
tri 11266 4812 11364 4910 sw
tri 11364 4812 11462 4910 ne
rect 11462 4812 11816 4910
tri 11816 4812 11914 4910 sw
tri 11914 4812 12012 4910 ne
rect 12012 4812 12366 4910
tri 12366 4812 12464 4910 sw
tri 12464 4812 12562 4910 ne
rect 12562 4812 12916 4910
tri 12916 4812 13014 4910 sw
tri 13014 4812 13112 4910 ne
rect 13112 4812 13466 4910
tri 13466 4812 13564 4910 sw
tri 13564 4812 13662 4910 ne
rect 13662 4812 14275 4910
rect -2525 4714 -186 4812
tri -186 4714 -88 4812 sw
tri -88 4714 10 4812 ne
rect 10 4714 364 4812
tri 364 4714 462 4812 sw
tri 462 4714 560 4812 ne
rect 560 4714 914 4812
tri 914 4714 1012 4812 sw
tri 1012 4714 1110 4812 ne
rect 1110 4714 1464 4812
tri 1464 4714 1562 4812 sw
tri 1562 4714 1660 4812 ne
rect 1660 4714 2014 4812
tri 2014 4714 2112 4812 sw
tri 2112 4714 2210 4812 ne
rect 2210 4714 2564 4812
tri 2564 4714 2662 4812 sw
tri 2662 4714 2760 4812 ne
rect 2760 4714 3114 4812
tri 3114 4714 3212 4812 sw
tri 3212 4714 3310 4812 ne
rect 3310 4714 3664 4812
tri 3664 4714 3762 4812 sw
tri 3762 4714 3860 4812 ne
rect 3860 4714 4214 4812
tri 4214 4714 4312 4812 sw
tri 4312 4714 4410 4812 ne
rect 4410 4714 4764 4812
tri 4764 4714 4862 4812 sw
tri 4862 4714 4960 4812 ne
rect 4960 4714 5314 4812
tri 5314 4714 5412 4812 sw
tri 5412 4714 5510 4812 ne
rect 5510 4714 5864 4812
tri 5864 4714 5962 4812 sw
tri 5962 4714 6060 4812 ne
rect 6060 4714 6414 4812
tri 6414 4714 6512 4812 sw
tri 6512 4714 6610 4812 ne
rect 6610 4714 6964 4812
tri 6964 4714 7062 4812 sw
tri 7062 4714 7160 4812 ne
rect 7160 4714 7514 4812
tri 7514 4714 7612 4812 sw
tri 7612 4714 7710 4812 ne
rect 7710 4714 8064 4812
tri 8064 4714 8162 4812 sw
tri 8162 4714 8260 4812 ne
rect 8260 4714 8614 4812
tri 8614 4714 8712 4812 sw
tri 8712 4714 8810 4812 ne
rect 8810 4714 9164 4812
tri 9164 4714 9262 4812 sw
tri 9262 4714 9360 4812 ne
rect 9360 4714 9714 4812
tri 9714 4714 9812 4812 sw
tri 9812 4714 9910 4812 ne
rect 9910 4714 10264 4812
tri 10264 4714 10362 4812 sw
tri 10362 4714 10460 4812 ne
rect 10460 4714 10814 4812
tri 10814 4714 10912 4812 sw
tri 10912 4714 11010 4812 ne
rect 11010 4714 11364 4812
tri 11364 4714 11462 4812 sw
tri 11462 4714 11560 4812 ne
rect 11560 4714 11914 4812
tri 11914 4714 12012 4812 sw
tri 12012 4714 12110 4812 ne
rect 12110 4714 12464 4812
tri 12464 4714 12562 4812 sw
tri 12562 4714 12660 4812 ne
rect 12660 4714 13014 4812
tri 13014 4714 13112 4812 sw
tri 13112 4714 13210 4812 ne
rect 13210 4714 13564 4812
tri 13564 4714 13662 4812 sw
rect 14775 4714 15775 5362
rect -2525 4710 -88 4714
rect -2525 4590 -310 4710
rect -190 4626 -88 4710
tri -88 4626 0 4714 sw
tri 10 4626 98 4714 ne
rect 98 4710 462 4714
rect 98 4626 240 4710
rect -190 4590 0 4626
rect -2525 4586 0 4590
rect -2525 3938 -1525 4586
tri -412 4488 -314 4586 ne
rect -314 4538 0 4586
tri 0 4538 88 4626 sw
tri 98 4538 186 4626 ne
rect 186 4590 240 4626
rect 360 4626 462 4710
tri 462 4626 550 4714 sw
tri 560 4626 648 4714 ne
rect 648 4710 1012 4714
rect 648 4626 790 4710
rect 360 4590 550 4626
rect 186 4586 550 4590
tri 550 4586 590 4626 sw
tri 648 4586 688 4626 ne
rect 688 4590 790 4626
rect 910 4626 1012 4710
tri 1012 4626 1100 4714 sw
tri 1110 4626 1198 4714 ne
rect 1198 4710 1562 4714
rect 1198 4626 1340 4710
rect 910 4590 1100 4626
rect 688 4586 1100 4590
rect 186 4538 590 4586
rect -314 4488 88 4538
rect -1025 4400 -412 4488
tri -412 4400 -324 4488 sw
tri -314 4400 -226 4488 ne
rect -226 4458 88 4488
tri 88 4458 168 4538 sw
tri 186 4458 266 4538 ne
rect 266 4488 590 4538
tri 590 4488 688 4586 sw
tri 688 4488 786 4586 ne
rect 786 4538 1100 4586
tri 1100 4538 1188 4626 sw
tri 1198 4538 1286 4626 ne
rect 1286 4590 1340 4626
rect 1460 4626 1562 4710
tri 1562 4626 1650 4714 sw
tri 1660 4626 1748 4714 ne
rect 1748 4710 2112 4714
rect 1748 4626 1890 4710
rect 1460 4590 1650 4626
rect 1286 4586 1650 4590
tri 1650 4586 1690 4626 sw
tri 1748 4586 1788 4626 ne
rect 1788 4590 1890 4626
rect 2010 4626 2112 4710
tri 2112 4626 2200 4714 sw
tri 2210 4626 2298 4714 ne
rect 2298 4710 2662 4714
rect 2298 4626 2440 4710
rect 2010 4590 2200 4626
rect 1788 4586 2200 4590
rect 1286 4538 1690 4586
rect 786 4488 1188 4538
rect 266 4458 688 4488
rect -226 4400 168 4458
rect -1025 4360 -324 4400
tri -324 4360 -284 4400 sw
tri -226 4360 -186 4400 ne
rect -186 4360 168 4400
tri 168 4360 266 4458 sw
tri 266 4360 364 4458 ne
rect 364 4400 688 4458
tri 688 4400 776 4488 sw
tri 786 4400 874 4488 ne
rect 874 4458 1188 4488
tri 1188 4458 1268 4538 sw
tri 1286 4458 1366 4538 ne
rect 1366 4488 1690 4538
tri 1690 4488 1788 4586 sw
tri 1788 4488 1886 4586 ne
rect 1886 4538 2200 4586
tri 2200 4538 2288 4626 sw
tri 2298 4538 2386 4626 ne
rect 2386 4590 2440 4626
rect 2560 4626 2662 4710
tri 2662 4626 2750 4714 sw
tri 2760 4626 2848 4714 ne
rect 2848 4710 3212 4714
rect 2848 4626 2990 4710
rect 2560 4590 2750 4626
rect 2386 4586 2750 4590
tri 2750 4586 2790 4626 sw
tri 2848 4586 2888 4626 ne
rect 2888 4590 2990 4626
rect 3110 4626 3212 4710
tri 3212 4626 3300 4714 sw
tri 3310 4626 3398 4714 ne
rect 3398 4710 3762 4714
rect 3398 4626 3540 4710
rect 3110 4590 3300 4626
rect 2888 4586 3300 4590
rect 2386 4538 2790 4586
rect 1886 4488 2288 4538
rect 1366 4458 1788 4488
rect 874 4400 1268 4458
rect 364 4360 776 4400
tri 776 4360 816 4400 sw
tri 874 4360 914 4400 ne
rect 914 4360 1268 4400
tri 1268 4360 1366 4458 sw
tri 1366 4360 1464 4458 ne
rect 1464 4400 1788 4458
tri 1788 4400 1876 4488 sw
tri 1886 4400 1974 4488 ne
rect 1974 4458 2288 4488
tri 2288 4458 2368 4538 sw
tri 2386 4458 2466 4538 ne
rect 2466 4488 2790 4538
tri 2790 4488 2888 4586 sw
tri 2888 4488 2986 4586 ne
rect 2986 4538 3300 4586
tri 3300 4538 3388 4626 sw
tri 3398 4538 3486 4626 ne
rect 3486 4590 3540 4626
rect 3660 4626 3762 4710
tri 3762 4626 3850 4714 sw
tri 3860 4626 3948 4714 ne
rect 3948 4710 4312 4714
rect 3948 4626 4090 4710
rect 3660 4590 3850 4626
rect 3486 4586 3850 4590
tri 3850 4586 3890 4626 sw
tri 3948 4586 3988 4626 ne
rect 3988 4590 4090 4626
rect 4210 4626 4312 4710
tri 4312 4626 4400 4714 sw
tri 4410 4626 4498 4714 ne
rect 4498 4710 4862 4714
rect 4498 4626 4640 4710
rect 4210 4590 4400 4626
rect 3988 4586 4400 4590
rect 3486 4538 3890 4586
rect 2986 4488 3388 4538
rect 2466 4458 2888 4488
rect 1974 4400 2368 4458
rect 1464 4360 1876 4400
tri 1876 4360 1916 4400 sw
tri 1974 4360 2014 4400 ne
rect 2014 4360 2368 4400
tri 2368 4360 2466 4458 sw
tri 2466 4360 2564 4458 ne
rect 2564 4400 2888 4458
tri 2888 4400 2976 4488 sw
tri 2986 4400 3074 4488 ne
rect 3074 4458 3388 4488
tri 3388 4458 3468 4538 sw
tri 3486 4458 3566 4538 ne
rect 3566 4488 3890 4538
tri 3890 4488 3988 4586 sw
tri 3988 4488 4086 4586 ne
rect 4086 4538 4400 4586
tri 4400 4538 4488 4626 sw
tri 4498 4538 4586 4626 ne
rect 4586 4590 4640 4626
rect 4760 4626 4862 4710
tri 4862 4626 4950 4714 sw
tri 4960 4626 5048 4714 ne
rect 5048 4710 5412 4714
rect 5048 4626 5190 4710
rect 4760 4590 4950 4626
rect 4586 4586 4950 4590
tri 4950 4586 4990 4626 sw
tri 5048 4586 5088 4626 ne
rect 5088 4590 5190 4626
rect 5310 4626 5412 4710
tri 5412 4626 5500 4714 sw
tri 5510 4626 5598 4714 ne
rect 5598 4710 5962 4714
rect 5598 4626 5740 4710
rect 5310 4590 5500 4626
rect 5088 4586 5500 4590
rect 4586 4538 4990 4586
rect 4086 4488 4488 4538
rect 3566 4458 3988 4488
rect 3074 4400 3468 4458
rect 2564 4360 2976 4400
tri 2976 4360 3016 4400 sw
tri 3074 4360 3114 4400 ne
rect 3114 4360 3468 4400
tri 3468 4360 3566 4458 sw
tri 3566 4360 3664 4458 ne
rect 3664 4400 3988 4458
tri 3988 4400 4076 4488 sw
tri 4086 4400 4174 4488 ne
rect 4174 4458 4488 4488
tri 4488 4458 4568 4538 sw
tri 4586 4458 4666 4538 ne
rect 4666 4488 4990 4538
tri 4990 4488 5088 4586 sw
tri 5088 4488 5186 4586 ne
rect 5186 4538 5500 4586
tri 5500 4538 5588 4626 sw
tri 5598 4538 5686 4626 ne
rect 5686 4590 5740 4626
rect 5860 4626 5962 4710
tri 5962 4626 6050 4714 sw
tri 6060 4626 6148 4714 ne
rect 6148 4710 6512 4714
rect 6148 4626 6290 4710
rect 5860 4590 6050 4626
rect 5686 4586 6050 4590
tri 6050 4586 6090 4626 sw
tri 6148 4586 6188 4626 ne
rect 6188 4590 6290 4626
rect 6410 4626 6512 4710
tri 6512 4626 6600 4714 sw
tri 6610 4626 6698 4714 ne
rect 6698 4710 7062 4714
rect 6698 4626 6840 4710
rect 6410 4590 6600 4626
rect 6188 4586 6600 4590
rect 5686 4538 6090 4586
rect 5186 4488 5588 4538
rect 4666 4458 5088 4488
rect 4174 4400 4568 4458
rect 3664 4360 4076 4400
tri 4076 4360 4116 4400 sw
tri 4174 4360 4214 4400 ne
rect 4214 4360 4568 4400
tri 4568 4360 4666 4458 sw
tri 4666 4360 4764 4458 ne
rect 4764 4400 5088 4458
tri 5088 4400 5176 4488 sw
tri 5186 4400 5274 4488 ne
rect 5274 4458 5588 4488
tri 5588 4458 5668 4538 sw
tri 5686 4458 5766 4538 ne
rect 5766 4488 6090 4538
tri 6090 4488 6188 4586 sw
tri 6188 4488 6286 4586 ne
rect 6286 4538 6600 4586
tri 6600 4538 6688 4626 sw
tri 6698 4538 6786 4626 ne
rect 6786 4590 6840 4626
rect 6960 4626 7062 4710
tri 7062 4626 7150 4714 sw
tri 7160 4626 7248 4714 ne
rect 7248 4710 7612 4714
rect 7248 4626 7390 4710
rect 6960 4590 7150 4626
rect 6786 4586 7150 4590
tri 7150 4586 7190 4626 sw
tri 7248 4586 7288 4626 ne
rect 7288 4590 7390 4626
rect 7510 4626 7612 4710
tri 7612 4626 7700 4714 sw
tri 7710 4626 7798 4714 ne
rect 7798 4710 8162 4714
rect 7798 4626 7940 4710
rect 7510 4590 7700 4626
rect 7288 4586 7700 4590
rect 6786 4538 7190 4586
rect 6286 4488 6688 4538
rect 5766 4458 6188 4488
rect 5274 4400 5668 4458
rect 4764 4360 5176 4400
tri 5176 4360 5216 4400 sw
tri 5274 4360 5314 4400 ne
rect 5314 4360 5668 4400
tri 5668 4360 5766 4458 sw
tri 5766 4360 5864 4458 ne
rect 5864 4400 6188 4458
tri 6188 4400 6276 4488 sw
tri 6286 4400 6374 4488 ne
rect 6374 4458 6688 4488
tri 6688 4458 6768 4538 sw
tri 6786 4458 6866 4538 ne
rect 6866 4488 7190 4538
tri 7190 4488 7288 4586 sw
tri 7288 4488 7386 4586 ne
rect 7386 4538 7700 4586
tri 7700 4538 7788 4626 sw
tri 7798 4538 7886 4626 ne
rect 7886 4590 7940 4626
rect 8060 4626 8162 4710
tri 8162 4626 8250 4714 sw
tri 8260 4626 8348 4714 ne
rect 8348 4710 8712 4714
rect 8348 4626 8490 4710
rect 8060 4590 8250 4626
rect 7886 4586 8250 4590
tri 8250 4586 8290 4626 sw
tri 8348 4586 8388 4626 ne
rect 8388 4590 8490 4626
rect 8610 4626 8712 4710
tri 8712 4626 8800 4714 sw
tri 8810 4626 8898 4714 ne
rect 8898 4710 9262 4714
rect 8898 4626 9040 4710
rect 8610 4590 8800 4626
rect 8388 4586 8800 4590
rect 7886 4538 8290 4586
rect 7386 4488 7788 4538
rect 6866 4458 7288 4488
rect 6374 4400 6768 4458
rect 5864 4360 6276 4400
tri 6276 4360 6316 4400 sw
tri 6374 4360 6414 4400 ne
rect 6414 4360 6768 4400
tri 6768 4360 6866 4458 sw
tri 6866 4360 6964 4458 ne
rect 6964 4400 7288 4458
tri 7288 4400 7376 4488 sw
tri 7386 4400 7474 4488 ne
rect 7474 4458 7788 4488
tri 7788 4458 7868 4538 sw
tri 7886 4458 7966 4538 ne
rect 7966 4488 8290 4538
tri 8290 4488 8388 4586 sw
tri 8388 4488 8486 4586 ne
rect 8486 4538 8800 4586
tri 8800 4538 8888 4626 sw
tri 8898 4538 8986 4626 ne
rect 8986 4590 9040 4626
rect 9160 4626 9262 4710
tri 9262 4626 9350 4714 sw
tri 9360 4626 9448 4714 ne
rect 9448 4710 9812 4714
rect 9448 4626 9590 4710
rect 9160 4590 9350 4626
rect 8986 4586 9350 4590
tri 9350 4586 9390 4626 sw
tri 9448 4586 9488 4626 ne
rect 9488 4590 9590 4626
rect 9710 4626 9812 4710
tri 9812 4626 9900 4714 sw
tri 9910 4626 9998 4714 ne
rect 9998 4710 10362 4714
rect 9998 4626 10140 4710
rect 9710 4590 9900 4626
rect 9488 4586 9900 4590
rect 8986 4538 9390 4586
rect 8486 4488 8888 4538
rect 7966 4458 8388 4488
rect 7474 4400 7868 4458
rect 6964 4360 7376 4400
tri 7376 4360 7416 4400 sw
tri 7474 4360 7514 4400 ne
rect 7514 4360 7868 4400
tri 7868 4360 7966 4458 sw
tri 7966 4360 8064 4458 ne
rect 8064 4400 8388 4458
tri 8388 4400 8476 4488 sw
tri 8486 4400 8574 4488 ne
rect 8574 4458 8888 4488
tri 8888 4458 8968 4538 sw
tri 8986 4458 9066 4538 ne
rect 9066 4488 9390 4538
tri 9390 4488 9488 4586 sw
tri 9488 4488 9586 4586 ne
rect 9586 4538 9900 4586
tri 9900 4538 9988 4626 sw
tri 9998 4538 10086 4626 ne
rect 10086 4590 10140 4626
rect 10260 4626 10362 4710
tri 10362 4626 10450 4714 sw
tri 10460 4626 10548 4714 ne
rect 10548 4710 10912 4714
rect 10548 4626 10690 4710
rect 10260 4590 10450 4626
rect 10086 4586 10450 4590
tri 10450 4586 10490 4626 sw
tri 10548 4586 10588 4626 ne
rect 10588 4590 10690 4626
rect 10810 4626 10912 4710
tri 10912 4626 11000 4714 sw
tri 11010 4626 11098 4714 ne
rect 11098 4710 11462 4714
rect 11098 4626 11240 4710
rect 10810 4590 11000 4626
rect 10588 4586 11000 4590
rect 10086 4538 10490 4586
rect 9586 4488 9988 4538
rect 9066 4458 9488 4488
rect 8574 4400 8968 4458
rect 8064 4360 8476 4400
tri 8476 4360 8516 4400 sw
tri 8574 4360 8614 4400 ne
rect 8614 4360 8968 4400
tri 8968 4360 9066 4458 sw
tri 9066 4360 9164 4458 ne
rect 9164 4400 9488 4458
tri 9488 4400 9576 4488 sw
tri 9586 4400 9674 4488 ne
rect 9674 4458 9988 4488
tri 9988 4458 10068 4538 sw
tri 10086 4458 10166 4538 ne
rect 10166 4488 10490 4538
tri 10490 4488 10588 4586 sw
tri 10588 4488 10686 4586 ne
rect 10686 4538 11000 4586
tri 11000 4538 11088 4626 sw
tri 11098 4538 11186 4626 ne
rect 11186 4590 11240 4626
rect 11360 4626 11462 4710
tri 11462 4626 11550 4714 sw
tri 11560 4626 11648 4714 ne
rect 11648 4710 12012 4714
rect 11648 4626 11790 4710
rect 11360 4590 11550 4626
rect 11186 4586 11550 4590
tri 11550 4586 11590 4626 sw
tri 11648 4586 11688 4626 ne
rect 11688 4590 11790 4626
rect 11910 4626 12012 4710
tri 12012 4626 12100 4714 sw
tri 12110 4626 12198 4714 ne
rect 12198 4710 12562 4714
rect 12198 4626 12340 4710
rect 11910 4590 12100 4626
rect 11688 4586 12100 4590
rect 11186 4538 11590 4586
rect 10686 4488 11088 4538
rect 10166 4458 10588 4488
rect 9674 4400 10068 4458
rect 9164 4360 9576 4400
tri 9576 4360 9616 4400 sw
tri 9674 4360 9714 4400 ne
rect 9714 4360 10068 4400
tri 10068 4360 10166 4458 sw
tri 10166 4360 10264 4458 ne
rect 10264 4400 10588 4458
tri 10588 4400 10676 4488 sw
tri 10686 4400 10774 4488 ne
rect 10774 4458 11088 4488
tri 11088 4458 11168 4538 sw
tri 11186 4458 11266 4538 ne
rect 11266 4488 11590 4538
tri 11590 4488 11688 4586 sw
tri 11688 4488 11786 4586 ne
rect 11786 4538 12100 4586
tri 12100 4538 12188 4626 sw
tri 12198 4538 12286 4626 ne
rect 12286 4590 12340 4626
rect 12460 4626 12562 4710
tri 12562 4626 12650 4714 sw
tri 12660 4626 12748 4714 ne
rect 12748 4710 13112 4714
rect 12748 4626 12890 4710
rect 12460 4590 12650 4626
rect 12286 4586 12650 4590
tri 12650 4586 12690 4626 sw
tri 12748 4586 12788 4626 ne
rect 12788 4590 12890 4626
rect 13010 4626 13112 4710
tri 13112 4626 13200 4714 sw
tri 13210 4626 13298 4714 ne
rect 13298 4710 15775 4714
rect 13298 4626 13440 4710
rect 13010 4590 13200 4626
rect 12788 4586 13200 4590
rect 12286 4538 12690 4586
rect 11786 4488 12188 4538
rect 11266 4458 11688 4488
rect 10774 4400 11168 4458
rect 10264 4360 10676 4400
tri 10676 4360 10716 4400 sw
tri 10774 4360 10814 4400 ne
rect 10814 4360 11168 4400
tri 11168 4360 11266 4458 sw
tri 11266 4360 11364 4458 ne
rect 11364 4400 11688 4458
tri 11688 4400 11776 4488 sw
tri 11786 4400 11874 4488 ne
rect 11874 4458 12188 4488
tri 12188 4458 12268 4538 sw
tri 12286 4458 12366 4538 ne
rect 12366 4488 12690 4538
tri 12690 4488 12788 4586 sw
tri 12788 4488 12886 4586 ne
rect 12886 4538 13200 4586
tri 13200 4538 13288 4626 sw
tri 13298 4538 13386 4626 ne
rect 13386 4590 13440 4626
rect 13560 4590 15775 4710
rect 13386 4538 15775 4590
rect 12886 4488 13288 4538
rect 12366 4458 12788 4488
rect 11874 4400 12268 4458
rect 11364 4360 11776 4400
tri 11776 4360 11816 4400 sw
tri 11874 4360 11914 4400 ne
rect 11914 4360 12268 4400
tri 12268 4360 12366 4458 sw
tri 12366 4360 12464 4458 ne
rect 12464 4400 12788 4458
tri 12788 4400 12876 4488 sw
tri 12886 4400 12974 4488 ne
rect 12974 4458 13288 4488
tri 13288 4458 13368 4538 sw
tri 13386 4458 13466 4538 ne
rect 13466 4458 14075 4538
rect 12974 4400 13368 4458
rect 12464 4360 12876 4400
tri 12876 4360 12916 4400 sw
tri 12974 4360 13014 4400 ne
rect 13014 4360 13368 4400
tri 13368 4360 13466 4458 sw
tri 13466 4360 13564 4458 ne
rect 13564 4438 14075 4458
rect 14175 4438 15775 4538
rect 13564 4360 15775 4438
rect -1025 4312 -284 4360
rect -1025 4212 -925 4312
rect -825 4262 -284 4312
tri -284 4262 -186 4360 sw
tri -186 4262 -88 4360 ne
rect -88 4262 266 4360
tri 266 4262 364 4360 sw
tri 364 4262 462 4360 ne
rect 462 4262 816 4360
tri 816 4262 914 4360 sw
tri 914 4262 1012 4360 ne
rect 1012 4262 1366 4360
tri 1366 4262 1464 4360 sw
tri 1464 4262 1562 4360 ne
rect 1562 4262 1916 4360
tri 1916 4262 2014 4360 sw
tri 2014 4262 2112 4360 ne
rect 2112 4262 2466 4360
tri 2466 4262 2564 4360 sw
tri 2564 4262 2662 4360 ne
rect 2662 4262 3016 4360
tri 3016 4262 3114 4360 sw
tri 3114 4262 3212 4360 ne
rect 3212 4262 3566 4360
tri 3566 4262 3664 4360 sw
tri 3664 4262 3762 4360 ne
rect 3762 4262 4116 4360
tri 4116 4262 4214 4360 sw
tri 4214 4262 4312 4360 ne
rect 4312 4262 4666 4360
tri 4666 4262 4764 4360 sw
tri 4764 4262 4862 4360 ne
rect 4862 4262 5216 4360
tri 5216 4262 5314 4360 sw
tri 5314 4262 5412 4360 ne
rect 5412 4262 5766 4360
tri 5766 4262 5864 4360 sw
tri 5864 4262 5962 4360 ne
rect 5962 4262 6316 4360
tri 6316 4262 6414 4360 sw
tri 6414 4262 6512 4360 ne
rect 6512 4262 6866 4360
tri 6866 4262 6964 4360 sw
tri 6964 4262 7062 4360 ne
rect 7062 4262 7416 4360
tri 7416 4262 7514 4360 sw
tri 7514 4262 7612 4360 ne
rect 7612 4262 7966 4360
tri 7966 4262 8064 4360 sw
tri 8064 4262 8162 4360 ne
rect 8162 4262 8516 4360
tri 8516 4262 8614 4360 sw
tri 8614 4262 8712 4360 ne
rect 8712 4262 9066 4360
tri 9066 4262 9164 4360 sw
tri 9164 4262 9262 4360 ne
rect 9262 4262 9616 4360
tri 9616 4262 9714 4360 sw
tri 9714 4262 9812 4360 ne
rect 9812 4262 10166 4360
tri 10166 4262 10264 4360 sw
tri 10264 4262 10362 4360 ne
rect 10362 4262 10716 4360
tri 10716 4262 10814 4360 sw
tri 10814 4262 10912 4360 ne
rect 10912 4262 11266 4360
tri 11266 4262 11364 4360 sw
tri 11364 4262 11462 4360 ne
rect 11462 4262 11816 4360
tri 11816 4262 11914 4360 sw
tri 11914 4262 12012 4360 ne
rect 12012 4262 12366 4360
tri 12366 4262 12464 4360 sw
tri 12464 4262 12562 4360 ne
rect 12562 4262 12916 4360
tri 12916 4262 13014 4360 sw
tri 13014 4262 13112 4360 ne
rect 13112 4262 13466 4360
tri 13466 4262 13564 4360 sw
tri 13564 4262 13662 4360 ne
rect 13662 4262 15775 4360
rect -825 4212 -186 4262
rect -1025 4164 -186 4212
tri -186 4164 -88 4262 sw
tri -88 4164 10 4262 ne
rect 10 4164 364 4262
tri 364 4164 462 4262 sw
tri 462 4164 560 4262 ne
rect 560 4164 914 4262
tri 914 4164 1012 4262 sw
tri 1012 4164 1110 4262 ne
rect 1110 4164 1464 4262
tri 1464 4164 1562 4262 sw
tri 1562 4164 1660 4262 ne
rect 1660 4164 2014 4262
tri 2014 4164 2112 4262 sw
tri 2112 4164 2210 4262 ne
rect 2210 4164 2564 4262
tri 2564 4164 2662 4262 sw
tri 2662 4164 2760 4262 ne
rect 2760 4164 3114 4262
tri 3114 4164 3212 4262 sw
tri 3212 4164 3310 4262 ne
rect 3310 4164 3664 4262
tri 3664 4164 3762 4262 sw
tri 3762 4164 3860 4262 ne
rect 3860 4164 4214 4262
tri 4214 4164 4312 4262 sw
tri 4312 4164 4410 4262 ne
rect 4410 4164 4764 4262
tri 4764 4164 4862 4262 sw
tri 4862 4164 4960 4262 ne
rect 4960 4164 5314 4262
tri 5314 4164 5412 4262 sw
tri 5412 4164 5510 4262 ne
rect 5510 4164 5864 4262
tri 5864 4164 5962 4262 sw
tri 5962 4164 6060 4262 ne
rect 6060 4164 6414 4262
tri 6414 4164 6512 4262 sw
tri 6512 4164 6610 4262 ne
rect 6610 4164 6964 4262
tri 6964 4164 7062 4262 sw
tri 7062 4164 7160 4262 ne
rect 7160 4164 7514 4262
tri 7514 4164 7612 4262 sw
tri 7612 4164 7710 4262 ne
rect 7710 4164 8064 4262
tri 8064 4164 8162 4262 sw
tri 8162 4164 8260 4262 ne
rect 8260 4164 8614 4262
tri 8614 4164 8712 4262 sw
tri 8712 4164 8810 4262 ne
rect 8810 4164 9164 4262
tri 9164 4164 9262 4262 sw
tri 9262 4164 9360 4262 ne
rect 9360 4164 9714 4262
tri 9714 4164 9812 4262 sw
tri 9812 4164 9910 4262 ne
rect 9910 4164 10264 4262
tri 10264 4164 10362 4262 sw
tri 10362 4164 10460 4262 ne
rect 10460 4164 10814 4262
tri 10814 4164 10912 4262 sw
tri 10912 4164 11010 4262 ne
rect 11010 4164 11364 4262
tri 11364 4164 11462 4262 sw
tri 11462 4164 11560 4262 ne
rect 11560 4164 11914 4262
tri 11914 4164 12012 4262 sw
tri 12012 4164 12110 4262 ne
rect 12110 4164 12464 4262
tri 12464 4164 12562 4262 sw
tri 12562 4164 12660 4262 ne
rect 12660 4164 13014 4262
tri 13014 4164 13112 4262 sw
tri 13112 4164 13210 4262 ne
rect 13210 4164 13564 4262
tri 13564 4164 13662 4262 sw
rect -1025 4160 -88 4164
rect -1025 4040 -310 4160
rect -190 4076 -88 4160
tri -88 4076 0 4164 sw
tri 10 4076 98 4164 ne
rect 98 4160 462 4164
rect 98 4076 240 4160
rect -190 4040 0 4076
rect -1025 4036 0 4040
tri 0 4036 40 4076 sw
tri 98 4036 138 4076 ne
rect 138 4040 240 4076
rect 360 4076 462 4160
tri 462 4076 550 4164 sw
tri 560 4076 648 4164 ne
rect 648 4160 1012 4164
rect 648 4076 790 4160
rect 360 4040 550 4076
rect 138 4036 550 4040
tri -412 3938 -314 4036 ne
rect -314 3938 40 4036
tri 40 3938 138 4036 sw
tri 138 3938 236 4036 ne
rect 236 3988 550 4036
tri 550 3988 638 4076 sw
tri 648 3988 736 4076 ne
rect 736 4040 790 4076
rect 910 4076 1012 4160
tri 1012 4076 1100 4164 sw
tri 1110 4076 1198 4164 ne
rect 1198 4160 1562 4164
rect 1198 4076 1340 4160
rect 910 4040 1100 4076
rect 736 4036 1100 4040
tri 1100 4036 1140 4076 sw
tri 1198 4036 1238 4076 ne
rect 1238 4040 1340 4076
rect 1460 4076 1562 4160
tri 1562 4076 1650 4164 sw
tri 1660 4076 1748 4164 ne
rect 1748 4160 2112 4164
rect 1748 4076 1890 4160
rect 1460 4040 1650 4076
rect 1238 4036 1650 4040
rect 736 3988 1140 4036
rect 236 3938 638 3988
rect -2525 3850 -412 3938
tri -412 3850 -324 3938 sw
tri -314 3850 -226 3938 ne
rect -226 3850 138 3938
tri 138 3850 226 3938 sw
tri 236 3850 324 3938 ne
rect 324 3908 638 3938
tri 638 3908 718 3988 sw
tri 736 3908 816 3988 ne
rect 816 3938 1140 3988
tri 1140 3938 1238 4036 sw
tri 1238 3938 1336 4036 ne
rect 1336 3988 1650 4036
tri 1650 3988 1738 4076 sw
tri 1748 3988 1836 4076 ne
rect 1836 4040 1890 4076
rect 2010 4076 2112 4160
tri 2112 4076 2200 4164 sw
tri 2210 4076 2298 4164 ne
rect 2298 4160 2662 4164
rect 2298 4076 2440 4160
rect 2010 4040 2200 4076
rect 1836 4036 2200 4040
tri 2200 4036 2240 4076 sw
tri 2298 4036 2338 4076 ne
rect 2338 4040 2440 4076
rect 2560 4076 2662 4160
tri 2662 4076 2750 4164 sw
tri 2760 4076 2848 4164 ne
rect 2848 4160 3212 4164
rect 2848 4076 2990 4160
rect 2560 4040 2750 4076
rect 2338 4036 2750 4040
rect 1836 3988 2240 4036
rect 1336 3938 1738 3988
rect 816 3908 1238 3938
rect 324 3850 718 3908
rect -2525 3810 -324 3850
tri -324 3810 -284 3850 sw
tri -226 3810 -186 3850 ne
rect -186 3810 226 3850
tri 226 3810 266 3850 sw
tri 324 3810 364 3850 ne
rect 364 3810 718 3850
tri 718 3810 816 3908 sw
tri 816 3810 914 3908 ne
rect 914 3850 1238 3908
tri 1238 3850 1326 3938 sw
tri 1336 3850 1424 3938 ne
rect 1424 3908 1738 3938
tri 1738 3908 1818 3988 sw
tri 1836 3908 1916 3988 ne
rect 1916 3938 2240 3988
tri 2240 3938 2338 4036 sw
tri 2338 3938 2436 4036 ne
rect 2436 3988 2750 4036
tri 2750 3988 2838 4076 sw
tri 2848 3988 2936 4076 ne
rect 2936 4040 2990 4076
rect 3110 4076 3212 4160
tri 3212 4076 3300 4164 sw
tri 3310 4076 3398 4164 ne
rect 3398 4160 3762 4164
rect 3398 4076 3540 4160
rect 3110 4040 3300 4076
rect 2936 4036 3300 4040
tri 3300 4036 3340 4076 sw
tri 3398 4036 3438 4076 ne
rect 3438 4040 3540 4076
rect 3660 4076 3762 4160
tri 3762 4076 3850 4164 sw
tri 3860 4076 3948 4164 ne
rect 3948 4160 4312 4164
rect 3948 4076 4090 4160
rect 3660 4040 3850 4076
rect 3438 4036 3850 4040
rect 2936 3988 3340 4036
rect 2436 3938 2838 3988
rect 1916 3908 2338 3938
rect 1424 3850 1818 3908
rect 914 3810 1326 3850
tri 1326 3810 1366 3850 sw
tri 1424 3810 1464 3850 ne
rect 1464 3810 1818 3850
tri 1818 3810 1916 3908 sw
tri 1916 3810 2014 3908 ne
rect 2014 3850 2338 3908
tri 2338 3850 2426 3938 sw
tri 2436 3850 2524 3938 ne
rect 2524 3908 2838 3938
tri 2838 3908 2918 3988 sw
tri 2936 3908 3016 3988 ne
rect 3016 3938 3340 3988
tri 3340 3938 3438 4036 sw
tri 3438 3938 3536 4036 ne
rect 3536 3988 3850 4036
tri 3850 3988 3938 4076 sw
tri 3948 3988 4036 4076 ne
rect 4036 4040 4090 4076
rect 4210 4076 4312 4160
tri 4312 4076 4400 4164 sw
tri 4410 4076 4498 4164 ne
rect 4498 4160 4862 4164
rect 4498 4076 4640 4160
rect 4210 4040 4400 4076
rect 4036 4036 4400 4040
tri 4400 4036 4440 4076 sw
tri 4498 4036 4538 4076 ne
rect 4538 4040 4640 4076
rect 4760 4076 4862 4160
tri 4862 4076 4950 4164 sw
tri 4960 4076 5048 4164 ne
rect 5048 4160 5412 4164
rect 5048 4076 5190 4160
rect 4760 4040 4950 4076
rect 4538 4036 4950 4040
rect 4036 3988 4440 4036
rect 3536 3938 3938 3988
rect 3016 3908 3438 3938
rect 2524 3850 2918 3908
rect 2014 3810 2426 3850
tri 2426 3810 2466 3850 sw
tri 2524 3810 2564 3850 ne
rect 2564 3810 2918 3850
tri 2918 3810 3016 3908 sw
tri 3016 3810 3114 3908 ne
rect 3114 3850 3438 3908
tri 3438 3850 3526 3938 sw
tri 3536 3850 3624 3938 ne
rect 3624 3908 3938 3938
tri 3938 3908 4018 3988 sw
tri 4036 3908 4116 3988 ne
rect 4116 3938 4440 3988
tri 4440 3938 4538 4036 sw
tri 4538 3938 4636 4036 ne
rect 4636 3988 4950 4036
tri 4950 3988 5038 4076 sw
tri 5048 3988 5136 4076 ne
rect 5136 4040 5190 4076
rect 5310 4076 5412 4160
tri 5412 4076 5500 4164 sw
tri 5510 4076 5598 4164 ne
rect 5598 4160 5962 4164
rect 5598 4076 5740 4160
rect 5310 4040 5500 4076
rect 5136 4036 5500 4040
tri 5500 4036 5540 4076 sw
tri 5598 4036 5638 4076 ne
rect 5638 4040 5740 4076
rect 5860 4076 5962 4160
tri 5962 4076 6050 4164 sw
tri 6060 4076 6148 4164 ne
rect 6148 4160 6512 4164
rect 6148 4076 6290 4160
rect 5860 4040 6050 4076
rect 5638 4036 6050 4040
rect 5136 3988 5540 4036
rect 4636 3938 5038 3988
rect 4116 3908 4538 3938
rect 3624 3850 4018 3908
rect 3114 3810 3526 3850
tri 3526 3810 3566 3850 sw
tri 3624 3810 3664 3850 ne
rect 3664 3810 4018 3850
tri 4018 3810 4116 3908 sw
tri 4116 3810 4214 3908 ne
rect 4214 3850 4538 3908
tri 4538 3850 4626 3938 sw
tri 4636 3850 4724 3938 ne
rect 4724 3908 5038 3938
tri 5038 3908 5118 3988 sw
tri 5136 3908 5216 3988 ne
rect 5216 3938 5540 3988
tri 5540 3938 5638 4036 sw
tri 5638 3938 5736 4036 ne
rect 5736 3988 6050 4036
tri 6050 3988 6138 4076 sw
tri 6148 3988 6236 4076 ne
rect 6236 4040 6290 4076
rect 6410 4076 6512 4160
tri 6512 4076 6600 4164 sw
tri 6610 4076 6698 4164 ne
rect 6698 4160 7062 4164
rect 6698 4076 6840 4160
rect 6410 4040 6600 4076
rect 6236 4036 6600 4040
tri 6600 4036 6640 4076 sw
tri 6698 4036 6738 4076 ne
rect 6738 4040 6840 4076
rect 6960 4076 7062 4160
tri 7062 4076 7150 4164 sw
tri 7160 4076 7248 4164 ne
rect 7248 4160 7612 4164
rect 7248 4076 7390 4160
rect 6960 4040 7150 4076
rect 6738 4036 7150 4040
rect 6236 3988 6640 4036
rect 5736 3938 6138 3988
rect 5216 3908 5638 3938
rect 4724 3850 5118 3908
rect 4214 3810 4626 3850
tri 4626 3810 4666 3850 sw
tri 4724 3810 4764 3850 ne
rect 4764 3810 5118 3850
tri 5118 3810 5216 3908 sw
tri 5216 3810 5314 3908 ne
rect 5314 3850 5638 3908
tri 5638 3850 5726 3938 sw
tri 5736 3850 5824 3938 ne
rect 5824 3908 6138 3938
tri 6138 3908 6218 3988 sw
tri 6236 3908 6316 3988 ne
rect 6316 3938 6640 3988
tri 6640 3938 6738 4036 sw
tri 6738 3938 6836 4036 ne
rect 6836 3988 7150 4036
tri 7150 3988 7238 4076 sw
tri 7248 3988 7336 4076 ne
rect 7336 4040 7390 4076
rect 7510 4076 7612 4160
tri 7612 4076 7700 4164 sw
tri 7710 4076 7798 4164 ne
rect 7798 4160 8162 4164
rect 7798 4076 7940 4160
rect 7510 4040 7700 4076
rect 7336 4036 7700 4040
tri 7700 4036 7740 4076 sw
tri 7798 4036 7838 4076 ne
rect 7838 4040 7940 4076
rect 8060 4076 8162 4160
tri 8162 4076 8250 4164 sw
tri 8260 4076 8348 4164 ne
rect 8348 4160 8712 4164
rect 8348 4076 8490 4160
rect 8060 4040 8250 4076
rect 7838 4036 8250 4040
rect 7336 3988 7740 4036
rect 6836 3938 7238 3988
rect 6316 3908 6738 3938
rect 5824 3850 6218 3908
rect 5314 3810 5726 3850
tri 5726 3810 5766 3850 sw
tri 5824 3810 5864 3850 ne
rect 5864 3810 6218 3850
tri 6218 3810 6316 3908 sw
tri 6316 3810 6414 3908 ne
rect 6414 3850 6738 3908
tri 6738 3850 6826 3938 sw
tri 6836 3850 6924 3938 ne
rect 6924 3908 7238 3938
tri 7238 3908 7318 3988 sw
tri 7336 3908 7416 3988 ne
rect 7416 3938 7740 3988
tri 7740 3938 7838 4036 sw
tri 7838 3938 7936 4036 ne
rect 7936 3988 8250 4036
tri 8250 3988 8338 4076 sw
tri 8348 3988 8436 4076 ne
rect 8436 4040 8490 4076
rect 8610 4076 8712 4160
tri 8712 4076 8800 4164 sw
tri 8810 4076 8898 4164 ne
rect 8898 4160 9262 4164
rect 8898 4076 9040 4160
rect 8610 4040 8800 4076
rect 8436 4036 8800 4040
tri 8800 4036 8840 4076 sw
tri 8898 4036 8938 4076 ne
rect 8938 4040 9040 4076
rect 9160 4076 9262 4160
tri 9262 4076 9350 4164 sw
tri 9360 4076 9448 4164 ne
rect 9448 4160 9812 4164
rect 9448 4076 9590 4160
rect 9160 4040 9350 4076
rect 8938 4036 9350 4040
rect 8436 3988 8840 4036
rect 7936 3938 8338 3988
rect 7416 3908 7838 3938
rect 6924 3850 7318 3908
rect 6414 3810 6826 3850
tri 6826 3810 6866 3850 sw
tri 6924 3810 6964 3850 ne
rect 6964 3810 7318 3850
tri 7318 3810 7416 3908 sw
tri 7416 3810 7514 3908 ne
rect 7514 3850 7838 3908
tri 7838 3850 7926 3938 sw
tri 7936 3850 8024 3938 ne
rect 8024 3908 8338 3938
tri 8338 3908 8418 3988 sw
tri 8436 3908 8516 3988 ne
rect 8516 3938 8840 3988
tri 8840 3938 8938 4036 sw
tri 8938 3938 9036 4036 ne
rect 9036 3988 9350 4036
tri 9350 3988 9438 4076 sw
tri 9448 3988 9536 4076 ne
rect 9536 4040 9590 4076
rect 9710 4076 9812 4160
tri 9812 4076 9900 4164 sw
tri 9910 4076 9998 4164 ne
rect 9998 4160 10362 4164
rect 9998 4076 10140 4160
rect 9710 4040 9900 4076
rect 9536 4036 9900 4040
tri 9900 4036 9940 4076 sw
tri 9998 4036 10038 4076 ne
rect 10038 4040 10140 4076
rect 10260 4076 10362 4160
tri 10362 4076 10450 4164 sw
tri 10460 4076 10548 4164 ne
rect 10548 4160 10912 4164
rect 10548 4076 10690 4160
rect 10260 4040 10450 4076
rect 10038 4036 10450 4040
rect 9536 3988 9940 4036
rect 9036 3938 9438 3988
rect 8516 3908 8938 3938
rect 8024 3850 8418 3908
rect 7514 3810 7926 3850
tri 7926 3810 7966 3850 sw
tri 8024 3810 8064 3850 ne
rect 8064 3810 8418 3850
tri 8418 3810 8516 3908 sw
tri 8516 3810 8614 3908 ne
rect 8614 3850 8938 3908
tri 8938 3850 9026 3938 sw
tri 9036 3850 9124 3938 ne
rect 9124 3908 9438 3938
tri 9438 3908 9518 3988 sw
tri 9536 3908 9616 3988 ne
rect 9616 3938 9940 3988
tri 9940 3938 10038 4036 sw
tri 10038 3938 10136 4036 ne
rect 10136 3988 10450 4036
tri 10450 3988 10538 4076 sw
tri 10548 3988 10636 4076 ne
rect 10636 4040 10690 4076
rect 10810 4076 10912 4160
tri 10912 4076 11000 4164 sw
tri 11010 4076 11098 4164 ne
rect 11098 4160 11462 4164
rect 11098 4076 11240 4160
rect 10810 4040 11000 4076
rect 10636 4036 11000 4040
tri 11000 4036 11040 4076 sw
tri 11098 4036 11138 4076 ne
rect 11138 4040 11240 4076
rect 11360 4076 11462 4160
tri 11462 4076 11550 4164 sw
tri 11560 4076 11648 4164 ne
rect 11648 4160 12012 4164
rect 11648 4076 11790 4160
rect 11360 4040 11550 4076
rect 11138 4036 11550 4040
rect 10636 3988 11040 4036
rect 10136 3938 10538 3988
rect 9616 3908 10038 3938
rect 9124 3850 9518 3908
rect 8614 3810 9026 3850
tri 9026 3810 9066 3850 sw
tri 9124 3810 9164 3850 ne
rect 9164 3810 9518 3850
tri 9518 3810 9616 3908 sw
tri 9616 3810 9714 3908 ne
rect 9714 3850 10038 3908
tri 10038 3850 10126 3938 sw
tri 10136 3850 10224 3938 ne
rect 10224 3908 10538 3938
tri 10538 3908 10618 3988 sw
tri 10636 3908 10716 3988 ne
rect 10716 3938 11040 3988
tri 11040 3938 11138 4036 sw
tri 11138 3938 11236 4036 ne
rect 11236 3988 11550 4036
tri 11550 3988 11638 4076 sw
tri 11648 3988 11736 4076 ne
rect 11736 4040 11790 4076
rect 11910 4076 12012 4160
tri 12012 4076 12100 4164 sw
tri 12110 4076 12198 4164 ne
rect 12198 4160 12562 4164
rect 12198 4076 12340 4160
rect 11910 4040 12100 4076
rect 11736 4036 12100 4040
tri 12100 4036 12140 4076 sw
tri 12198 4036 12238 4076 ne
rect 12238 4040 12340 4076
rect 12460 4076 12562 4160
tri 12562 4076 12650 4164 sw
tri 12660 4076 12748 4164 ne
rect 12748 4160 13112 4164
rect 12748 4076 12890 4160
rect 12460 4040 12650 4076
rect 12238 4036 12650 4040
rect 11736 3988 12140 4036
rect 11236 3938 11638 3988
rect 10716 3908 11138 3938
rect 10224 3850 10618 3908
rect 9714 3810 10126 3850
tri 10126 3810 10166 3850 sw
tri 10224 3810 10264 3850 ne
rect 10264 3810 10618 3850
tri 10618 3810 10716 3908 sw
tri 10716 3810 10814 3908 ne
rect 10814 3850 11138 3908
tri 11138 3850 11226 3938 sw
tri 11236 3850 11324 3938 ne
rect 11324 3908 11638 3938
tri 11638 3908 11718 3988 sw
tri 11736 3908 11816 3988 ne
rect 11816 3938 12140 3988
tri 12140 3938 12238 4036 sw
tri 12238 3938 12336 4036 ne
rect 12336 3988 12650 4036
tri 12650 3988 12738 4076 sw
tri 12748 3988 12836 4076 ne
rect 12836 4040 12890 4076
rect 13010 4076 13112 4160
tri 13112 4076 13200 4164 sw
tri 13210 4076 13298 4164 ne
rect 13298 4160 14275 4164
rect 13298 4076 13440 4160
rect 13010 4040 13200 4076
rect 12836 4036 13200 4040
tri 13200 4036 13240 4076 sw
tri 13298 4036 13338 4076 ne
rect 13338 4040 13440 4076
rect 13560 4040 14275 4160
rect 13338 4036 14275 4040
rect 12836 3988 13240 4036
rect 12336 3938 12738 3988
rect 11816 3908 12238 3938
rect 11324 3850 11718 3908
rect 10814 3810 11226 3850
tri 11226 3810 11266 3850 sw
tri 11324 3810 11364 3850 ne
rect 11364 3810 11718 3850
tri 11718 3810 11816 3908 sw
tri 11816 3810 11914 3908 ne
rect 11914 3850 12238 3908
tri 12238 3850 12326 3938 sw
tri 12336 3850 12424 3938 ne
rect 12424 3908 12738 3938
tri 12738 3908 12818 3988 sw
tri 12836 3908 12916 3988 ne
rect 12916 3938 13240 3988
tri 13240 3938 13338 4036 sw
tri 13338 3938 13436 4036 ne
rect 13436 3938 14275 4036
rect 12916 3908 13338 3938
rect 12424 3850 12818 3908
rect 11914 3810 12326 3850
tri 12326 3810 12366 3850 sw
tri 12424 3810 12464 3850 ne
rect 12464 3810 12818 3850
tri 12818 3810 12916 3908 sw
tri 12916 3810 13014 3908 ne
rect 13014 3850 13338 3908
tri 13338 3850 13426 3938 sw
tri 13436 3850 13524 3938 ne
rect 13524 3850 14275 3938
rect 13014 3810 13426 3850
tri 13426 3810 13466 3850 sw
tri 13524 3810 13564 3850 ne
rect 13564 3810 14275 3850
rect -2525 3712 -284 3810
tri -284 3712 -186 3810 sw
tri -186 3712 -88 3810 ne
rect -88 3712 266 3810
tri 266 3712 364 3810 sw
tri 364 3712 462 3810 ne
rect 462 3712 816 3810
tri 816 3712 914 3810 sw
tri 914 3712 1012 3810 ne
rect 1012 3712 1366 3810
tri 1366 3712 1464 3810 sw
tri 1464 3712 1562 3810 ne
rect 1562 3712 1916 3810
tri 1916 3712 2014 3810 sw
tri 2014 3712 2112 3810 ne
rect 2112 3712 2466 3810
tri 2466 3712 2564 3810 sw
tri 2564 3712 2662 3810 ne
rect 2662 3712 3016 3810
tri 3016 3712 3114 3810 sw
tri 3114 3712 3212 3810 ne
rect 3212 3712 3566 3810
tri 3566 3712 3664 3810 sw
tri 3664 3712 3762 3810 ne
rect 3762 3712 4116 3810
tri 4116 3712 4214 3810 sw
tri 4214 3712 4312 3810 ne
rect 4312 3712 4666 3810
tri 4666 3712 4764 3810 sw
tri 4764 3712 4862 3810 ne
rect 4862 3712 5216 3810
tri 5216 3712 5314 3810 sw
tri 5314 3712 5412 3810 ne
rect 5412 3712 5766 3810
tri 5766 3712 5864 3810 sw
tri 5864 3712 5962 3810 ne
rect 5962 3712 6316 3810
tri 6316 3712 6414 3810 sw
tri 6414 3712 6512 3810 ne
rect 6512 3712 6866 3810
tri 6866 3712 6964 3810 sw
tri 6964 3712 7062 3810 ne
rect 7062 3712 7416 3810
tri 7416 3712 7514 3810 sw
tri 7514 3712 7612 3810 ne
rect 7612 3712 7966 3810
tri 7966 3712 8064 3810 sw
tri 8064 3712 8162 3810 ne
rect 8162 3712 8516 3810
tri 8516 3712 8614 3810 sw
tri 8614 3712 8712 3810 ne
rect 8712 3712 9066 3810
tri 9066 3712 9164 3810 sw
tri 9164 3712 9262 3810 ne
rect 9262 3712 9616 3810
tri 9616 3712 9714 3810 sw
tri 9714 3712 9812 3810 ne
rect 9812 3712 10166 3810
tri 10166 3712 10264 3810 sw
tri 10264 3712 10362 3810 ne
rect 10362 3712 10716 3810
tri 10716 3712 10814 3810 sw
tri 10814 3712 10912 3810 ne
rect 10912 3712 11266 3810
tri 11266 3712 11364 3810 sw
tri 11364 3712 11462 3810 ne
rect 11462 3712 11816 3810
tri 11816 3712 11914 3810 sw
tri 11914 3712 12012 3810 ne
rect 12012 3712 12366 3810
tri 12366 3712 12464 3810 sw
tri 12464 3712 12562 3810 ne
rect 12562 3712 12916 3810
tri 12916 3712 13014 3810 sw
tri 13014 3712 13112 3810 ne
rect 13112 3712 13466 3810
tri 13466 3712 13564 3810 sw
tri 13564 3712 13662 3810 ne
rect 13662 3712 14275 3810
rect -2525 3614 -186 3712
tri -186 3614 -88 3712 sw
tri -88 3614 10 3712 ne
rect 10 3614 364 3712
tri 364 3614 462 3712 sw
tri 462 3614 560 3712 ne
rect 560 3614 914 3712
tri 914 3614 1012 3712 sw
tri 1012 3614 1110 3712 ne
rect 1110 3614 1464 3712
tri 1464 3614 1562 3712 sw
tri 1562 3614 1660 3712 ne
rect 1660 3614 2014 3712
tri 2014 3614 2112 3712 sw
tri 2112 3614 2210 3712 ne
rect 2210 3614 2564 3712
tri 2564 3614 2662 3712 sw
tri 2662 3614 2760 3712 ne
rect 2760 3614 3114 3712
tri 3114 3614 3212 3712 sw
tri 3212 3614 3310 3712 ne
rect 3310 3614 3664 3712
tri 3664 3614 3762 3712 sw
tri 3762 3614 3860 3712 ne
rect 3860 3614 4214 3712
tri 4214 3614 4312 3712 sw
tri 4312 3614 4410 3712 ne
rect 4410 3614 4764 3712
tri 4764 3614 4862 3712 sw
tri 4862 3614 4960 3712 ne
rect 4960 3614 5314 3712
tri 5314 3614 5412 3712 sw
tri 5412 3614 5510 3712 ne
rect 5510 3614 5864 3712
tri 5864 3614 5962 3712 sw
tri 5962 3614 6060 3712 ne
rect 6060 3614 6414 3712
tri 6414 3614 6512 3712 sw
tri 6512 3614 6610 3712 ne
rect 6610 3614 6964 3712
tri 6964 3614 7062 3712 sw
tri 7062 3614 7160 3712 ne
rect 7160 3614 7514 3712
tri 7514 3614 7612 3712 sw
tri 7612 3614 7710 3712 ne
rect 7710 3614 8064 3712
tri 8064 3614 8162 3712 sw
tri 8162 3614 8260 3712 ne
rect 8260 3614 8614 3712
tri 8614 3614 8712 3712 sw
tri 8712 3614 8810 3712 ne
rect 8810 3614 9164 3712
tri 9164 3614 9262 3712 sw
tri 9262 3614 9360 3712 ne
rect 9360 3614 9714 3712
tri 9714 3614 9812 3712 sw
tri 9812 3614 9910 3712 ne
rect 9910 3614 10264 3712
tri 10264 3614 10362 3712 sw
tri 10362 3614 10460 3712 ne
rect 10460 3614 10814 3712
tri 10814 3614 10912 3712 sw
tri 10912 3614 11010 3712 ne
rect 11010 3614 11364 3712
tri 11364 3614 11462 3712 sw
tri 11462 3614 11560 3712 ne
rect 11560 3614 11914 3712
tri 11914 3614 12012 3712 sw
tri 12012 3614 12110 3712 ne
rect 12110 3614 12464 3712
tri 12464 3614 12562 3712 sw
tri 12562 3614 12660 3712 ne
rect 12660 3614 13014 3712
tri 13014 3614 13112 3712 sw
tri 13112 3614 13210 3712 ne
rect 13210 3614 13564 3712
tri 13564 3614 13662 3712 sw
rect 14775 3614 15775 4262
rect -2525 3610 -88 3614
rect -2525 3490 -310 3610
rect -190 3526 -88 3610
tri -88 3526 0 3614 sw
tri 10 3526 98 3614 ne
rect 98 3610 462 3614
rect 98 3526 240 3610
rect -190 3490 0 3526
rect -2525 3486 0 3490
rect -2525 2838 -1525 3486
tri -412 3388 -314 3486 ne
rect -314 3438 0 3486
tri 0 3438 88 3526 sw
tri 98 3438 186 3526 ne
rect 186 3490 240 3526
rect 360 3526 462 3610
tri 462 3526 550 3614 sw
tri 560 3526 648 3614 ne
rect 648 3610 1012 3614
rect 648 3526 790 3610
rect 360 3490 550 3526
rect 186 3486 550 3490
tri 550 3486 590 3526 sw
tri 648 3486 688 3526 ne
rect 688 3490 790 3526
rect 910 3526 1012 3610
tri 1012 3526 1100 3614 sw
tri 1110 3526 1198 3614 ne
rect 1198 3610 1562 3614
rect 1198 3526 1340 3610
rect 910 3490 1100 3526
rect 688 3486 1100 3490
rect 186 3438 590 3486
rect -314 3388 88 3438
rect -1025 3300 -412 3388
tri -412 3300 -324 3388 sw
tri -314 3300 -226 3388 ne
rect -226 3358 88 3388
tri 88 3358 168 3438 sw
tri 186 3358 266 3438 ne
rect 266 3388 590 3438
tri 590 3388 688 3486 sw
tri 688 3388 786 3486 ne
rect 786 3438 1100 3486
tri 1100 3438 1188 3526 sw
tri 1198 3438 1286 3526 ne
rect 1286 3490 1340 3526
rect 1460 3526 1562 3610
tri 1562 3526 1650 3614 sw
tri 1660 3526 1748 3614 ne
rect 1748 3610 2112 3614
rect 1748 3526 1890 3610
rect 1460 3490 1650 3526
rect 1286 3486 1650 3490
tri 1650 3486 1690 3526 sw
tri 1748 3486 1788 3526 ne
rect 1788 3490 1890 3526
rect 2010 3526 2112 3610
tri 2112 3526 2200 3614 sw
tri 2210 3526 2298 3614 ne
rect 2298 3610 2662 3614
rect 2298 3526 2440 3610
rect 2010 3490 2200 3526
rect 1788 3486 2200 3490
rect 1286 3438 1690 3486
rect 786 3388 1188 3438
rect 266 3358 688 3388
rect -226 3300 168 3358
rect -1025 3260 -324 3300
tri -324 3260 -284 3300 sw
tri -226 3260 -186 3300 ne
rect -186 3260 168 3300
tri 168 3260 266 3358 sw
tri 266 3260 364 3358 ne
rect 364 3300 688 3358
tri 688 3300 776 3388 sw
tri 786 3300 874 3388 ne
rect 874 3358 1188 3388
tri 1188 3358 1268 3438 sw
tri 1286 3358 1366 3438 ne
rect 1366 3388 1690 3438
tri 1690 3388 1788 3486 sw
tri 1788 3388 1886 3486 ne
rect 1886 3438 2200 3486
tri 2200 3438 2288 3526 sw
tri 2298 3438 2386 3526 ne
rect 2386 3490 2440 3526
rect 2560 3526 2662 3610
tri 2662 3526 2750 3614 sw
tri 2760 3526 2848 3614 ne
rect 2848 3610 3212 3614
rect 2848 3526 2990 3610
rect 2560 3490 2750 3526
rect 2386 3486 2750 3490
tri 2750 3486 2790 3526 sw
tri 2848 3486 2888 3526 ne
rect 2888 3490 2990 3526
rect 3110 3526 3212 3610
tri 3212 3526 3300 3614 sw
tri 3310 3526 3398 3614 ne
rect 3398 3610 3762 3614
rect 3398 3526 3540 3610
rect 3110 3490 3300 3526
rect 2888 3486 3300 3490
rect 2386 3438 2790 3486
rect 1886 3388 2288 3438
rect 1366 3358 1788 3388
rect 874 3300 1268 3358
rect 364 3260 776 3300
tri 776 3260 816 3300 sw
tri 874 3260 914 3300 ne
rect 914 3260 1268 3300
tri 1268 3260 1366 3358 sw
tri 1366 3260 1464 3358 ne
rect 1464 3300 1788 3358
tri 1788 3300 1876 3388 sw
tri 1886 3300 1974 3388 ne
rect 1974 3358 2288 3388
tri 2288 3358 2368 3438 sw
tri 2386 3358 2466 3438 ne
rect 2466 3388 2790 3438
tri 2790 3388 2888 3486 sw
tri 2888 3388 2986 3486 ne
rect 2986 3438 3300 3486
tri 3300 3438 3388 3526 sw
tri 3398 3438 3486 3526 ne
rect 3486 3490 3540 3526
rect 3660 3526 3762 3610
tri 3762 3526 3850 3614 sw
tri 3860 3526 3948 3614 ne
rect 3948 3610 4312 3614
rect 3948 3526 4090 3610
rect 3660 3490 3850 3526
rect 3486 3486 3850 3490
tri 3850 3486 3890 3526 sw
tri 3948 3486 3988 3526 ne
rect 3988 3490 4090 3526
rect 4210 3526 4312 3610
tri 4312 3526 4400 3614 sw
tri 4410 3526 4498 3614 ne
rect 4498 3610 4862 3614
rect 4498 3526 4640 3610
rect 4210 3490 4400 3526
rect 3988 3486 4400 3490
rect 3486 3438 3890 3486
rect 2986 3388 3388 3438
rect 2466 3358 2888 3388
rect 1974 3300 2368 3358
rect 1464 3260 1876 3300
tri 1876 3260 1916 3300 sw
tri 1974 3260 2014 3300 ne
rect 2014 3260 2368 3300
tri 2368 3260 2466 3358 sw
tri 2466 3260 2564 3358 ne
rect 2564 3300 2888 3358
tri 2888 3300 2976 3388 sw
tri 2986 3300 3074 3388 ne
rect 3074 3358 3388 3388
tri 3388 3358 3468 3438 sw
tri 3486 3358 3566 3438 ne
rect 3566 3388 3890 3438
tri 3890 3388 3988 3486 sw
tri 3988 3388 4086 3486 ne
rect 4086 3438 4400 3486
tri 4400 3438 4488 3526 sw
tri 4498 3438 4586 3526 ne
rect 4586 3490 4640 3526
rect 4760 3526 4862 3610
tri 4862 3526 4950 3614 sw
tri 4960 3526 5048 3614 ne
rect 5048 3610 5412 3614
rect 5048 3526 5190 3610
rect 4760 3490 4950 3526
rect 4586 3486 4950 3490
tri 4950 3486 4990 3526 sw
tri 5048 3486 5088 3526 ne
rect 5088 3490 5190 3526
rect 5310 3526 5412 3610
tri 5412 3526 5500 3614 sw
tri 5510 3526 5598 3614 ne
rect 5598 3610 5962 3614
rect 5598 3526 5740 3610
rect 5310 3490 5500 3526
rect 5088 3486 5500 3490
rect 4586 3438 4990 3486
rect 4086 3388 4488 3438
rect 3566 3358 3988 3388
rect 3074 3300 3468 3358
rect 2564 3260 2976 3300
tri 2976 3260 3016 3300 sw
tri 3074 3260 3114 3300 ne
rect 3114 3260 3468 3300
tri 3468 3260 3566 3358 sw
tri 3566 3260 3664 3358 ne
rect 3664 3300 3988 3358
tri 3988 3300 4076 3388 sw
tri 4086 3300 4174 3388 ne
rect 4174 3358 4488 3388
tri 4488 3358 4568 3438 sw
tri 4586 3358 4666 3438 ne
rect 4666 3388 4990 3438
tri 4990 3388 5088 3486 sw
tri 5088 3388 5186 3486 ne
rect 5186 3438 5500 3486
tri 5500 3438 5588 3526 sw
tri 5598 3438 5686 3526 ne
rect 5686 3490 5740 3526
rect 5860 3526 5962 3610
tri 5962 3526 6050 3614 sw
tri 6060 3526 6148 3614 ne
rect 6148 3610 6512 3614
rect 6148 3526 6290 3610
rect 5860 3490 6050 3526
rect 5686 3486 6050 3490
tri 6050 3486 6090 3526 sw
tri 6148 3486 6188 3526 ne
rect 6188 3490 6290 3526
rect 6410 3526 6512 3610
tri 6512 3526 6600 3614 sw
tri 6610 3526 6698 3614 ne
rect 6698 3610 7062 3614
rect 6698 3526 6840 3610
rect 6410 3490 6600 3526
rect 6188 3486 6600 3490
rect 5686 3438 6090 3486
rect 5186 3388 5588 3438
rect 4666 3358 5088 3388
rect 4174 3300 4568 3358
rect 3664 3260 4076 3300
tri 4076 3260 4116 3300 sw
tri 4174 3260 4214 3300 ne
rect 4214 3260 4568 3300
tri 4568 3260 4666 3358 sw
tri 4666 3260 4764 3358 ne
rect 4764 3300 5088 3358
tri 5088 3300 5176 3388 sw
tri 5186 3300 5274 3388 ne
rect 5274 3358 5588 3388
tri 5588 3358 5668 3438 sw
tri 5686 3358 5766 3438 ne
rect 5766 3388 6090 3438
tri 6090 3388 6188 3486 sw
tri 6188 3388 6286 3486 ne
rect 6286 3438 6600 3486
tri 6600 3438 6688 3526 sw
tri 6698 3438 6786 3526 ne
rect 6786 3490 6840 3526
rect 6960 3526 7062 3610
tri 7062 3526 7150 3614 sw
tri 7160 3526 7248 3614 ne
rect 7248 3610 7612 3614
rect 7248 3526 7390 3610
rect 6960 3490 7150 3526
rect 6786 3486 7150 3490
tri 7150 3486 7190 3526 sw
tri 7248 3486 7288 3526 ne
rect 7288 3490 7390 3526
rect 7510 3526 7612 3610
tri 7612 3526 7700 3614 sw
tri 7710 3526 7798 3614 ne
rect 7798 3610 8162 3614
rect 7798 3526 7940 3610
rect 7510 3490 7700 3526
rect 7288 3486 7700 3490
rect 6786 3438 7190 3486
rect 6286 3388 6688 3438
rect 5766 3358 6188 3388
rect 5274 3300 5668 3358
rect 4764 3260 5176 3300
tri 5176 3260 5216 3300 sw
tri 5274 3260 5314 3300 ne
rect 5314 3260 5668 3300
tri 5668 3260 5766 3358 sw
tri 5766 3260 5864 3358 ne
rect 5864 3300 6188 3358
tri 6188 3300 6276 3388 sw
tri 6286 3300 6374 3388 ne
rect 6374 3358 6688 3388
tri 6688 3358 6768 3438 sw
tri 6786 3358 6866 3438 ne
rect 6866 3388 7190 3438
tri 7190 3388 7288 3486 sw
tri 7288 3388 7386 3486 ne
rect 7386 3438 7700 3486
tri 7700 3438 7788 3526 sw
tri 7798 3438 7886 3526 ne
rect 7886 3490 7940 3526
rect 8060 3526 8162 3610
tri 8162 3526 8250 3614 sw
tri 8260 3526 8348 3614 ne
rect 8348 3610 8712 3614
rect 8348 3526 8490 3610
rect 8060 3490 8250 3526
rect 7886 3486 8250 3490
tri 8250 3486 8290 3526 sw
tri 8348 3486 8388 3526 ne
rect 8388 3490 8490 3526
rect 8610 3526 8712 3610
tri 8712 3526 8800 3614 sw
tri 8810 3526 8898 3614 ne
rect 8898 3610 9262 3614
rect 8898 3526 9040 3610
rect 8610 3490 8800 3526
rect 8388 3486 8800 3490
rect 7886 3438 8290 3486
rect 7386 3388 7788 3438
rect 6866 3358 7288 3388
rect 6374 3300 6768 3358
rect 5864 3260 6276 3300
tri 6276 3260 6316 3300 sw
tri 6374 3260 6414 3300 ne
rect 6414 3260 6768 3300
tri 6768 3260 6866 3358 sw
tri 6866 3260 6964 3358 ne
rect 6964 3300 7288 3358
tri 7288 3300 7376 3388 sw
tri 7386 3300 7474 3388 ne
rect 7474 3358 7788 3388
tri 7788 3358 7868 3438 sw
tri 7886 3358 7966 3438 ne
rect 7966 3388 8290 3438
tri 8290 3388 8388 3486 sw
tri 8388 3388 8486 3486 ne
rect 8486 3438 8800 3486
tri 8800 3438 8888 3526 sw
tri 8898 3438 8986 3526 ne
rect 8986 3490 9040 3526
rect 9160 3526 9262 3610
tri 9262 3526 9350 3614 sw
tri 9360 3526 9448 3614 ne
rect 9448 3610 9812 3614
rect 9448 3526 9590 3610
rect 9160 3490 9350 3526
rect 8986 3486 9350 3490
tri 9350 3486 9390 3526 sw
tri 9448 3486 9488 3526 ne
rect 9488 3490 9590 3526
rect 9710 3526 9812 3610
tri 9812 3526 9900 3614 sw
tri 9910 3526 9998 3614 ne
rect 9998 3610 10362 3614
rect 9998 3526 10140 3610
rect 9710 3490 9900 3526
rect 9488 3486 9900 3490
rect 8986 3438 9390 3486
rect 8486 3388 8888 3438
rect 7966 3358 8388 3388
rect 7474 3300 7868 3358
rect 6964 3260 7376 3300
tri 7376 3260 7416 3300 sw
tri 7474 3260 7514 3300 ne
rect 7514 3260 7868 3300
tri 7868 3260 7966 3358 sw
tri 7966 3260 8064 3358 ne
rect 8064 3300 8388 3358
tri 8388 3300 8476 3388 sw
tri 8486 3300 8574 3388 ne
rect 8574 3358 8888 3388
tri 8888 3358 8968 3438 sw
tri 8986 3358 9066 3438 ne
rect 9066 3388 9390 3438
tri 9390 3388 9488 3486 sw
tri 9488 3388 9586 3486 ne
rect 9586 3438 9900 3486
tri 9900 3438 9988 3526 sw
tri 9998 3438 10086 3526 ne
rect 10086 3490 10140 3526
rect 10260 3526 10362 3610
tri 10362 3526 10450 3614 sw
tri 10460 3526 10548 3614 ne
rect 10548 3610 10912 3614
rect 10548 3526 10690 3610
rect 10260 3490 10450 3526
rect 10086 3486 10450 3490
tri 10450 3486 10490 3526 sw
tri 10548 3486 10588 3526 ne
rect 10588 3490 10690 3526
rect 10810 3526 10912 3610
tri 10912 3526 11000 3614 sw
tri 11010 3526 11098 3614 ne
rect 11098 3610 11462 3614
rect 11098 3526 11240 3610
rect 10810 3490 11000 3526
rect 10588 3486 11000 3490
rect 10086 3438 10490 3486
rect 9586 3388 9988 3438
rect 9066 3358 9488 3388
rect 8574 3300 8968 3358
rect 8064 3260 8476 3300
tri 8476 3260 8516 3300 sw
tri 8574 3260 8614 3300 ne
rect 8614 3260 8968 3300
tri 8968 3260 9066 3358 sw
tri 9066 3260 9164 3358 ne
rect 9164 3300 9488 3358
tri 9488 3300 9576 3388 sw
tri 9586 3300 9674 3388 ne
rect 9674 3358 9988 3388
tri 9988 3358 10068 3438 sw
tri 10086 3358 10166 3438 ne
rect 10166 3388 10490 3438
tri 10490 3388 10588 3486 sw
tri 10588 3388 10686 3486 ne
rect 10686 3438 11000 3486
tri 11000 3438 11088 3526 sw
tri 11098 3438 11186 3526 ne
rect 11186 3490 11240 3526
rect 11360 3526 11462 3610
tri 11462 3526 11550 3614 sw
tri 11560 3526 11648 3614 ne
rect 11648 3610 12012 3614
rect 11648 3526 11790 3610
rect 11360 3490 11550 3526
rect 11186 3486 11550 3490
tri 11550 3486 11590 3526 sw
tri 11648 3486 11688 3526 ne
rect 11688 3490 11790 3526
rect 11910 3526 12012 3610
tri 12012 3526 12100 3614 sw
tri 12110 3526 12198 3614 ne
rect 12198 3610 12562 3614
rect 12198 3526 12340 3610
rect 11910 3490 12100 3526
rect 11688 3486 12100 3490
rect 11186 3438 11590 3486
rect 10686 3388 11088 3438
rect 10166 3358 10588 3388
rect 9674 3300 10068 3358
rect 9164 3260 9576 3300
tri 9576 3260 9616 3300 sw
tri 9674 3260 9714 3300 ne
rect 9714 3260 10068 3300
tri 10068 3260 10166 3358 sw
tri 10166 3260 10264 3358 ne
rect 10264 3300 10588 3358
tri 10588 3300 10676 3388 sw
tri 10686 3300 10774 3388 ne
rect 10774 3358 11088 3388
tri 11088 3358 11168 3438 sw
tri 11186 3358 11266 3438 ne
rect 11266 3388 11590 3438
tri 11590 3388 11688 3486 sw
tri 11688 3388 11786 3486 ne
rect 11786 3438 12100 3486
tri 12100 3438 12188 3526 sw
tri 12198 3438 12286 3526 ne
rect 12286 3490 12340 3526
rect 12460 3526 12562 3610
tri 12562 3526 12650 3614 sw
tri 12660 3526 12748 3614 ne
rect 12748 3610 13112 3614
rect 12748 3526 12890 3610
rect 12460 3490 12650 3526
rect 12286 3486 12650 3490
tri 12650 3486 12690 3526 sw
tri 12748 3486 12788 3526 ne
rect 12788 3490 12890 3526
rect 13010 3526 13112 3610
tri 13112 3526 13200 3614 sw
tri 13210 3526 13298 3614 ne
rect 13298 3610 15775 3614
rect 13298 3526 13440 3610
rect 13010 3490 13200 3526
rect 12788 3486 13200 3490
rect 12286 3438 12690 3486
rect 11786 3388 12188 3438
rect 11266 3358 11688 3388
rect 10774 3300 11168 3358
rect 10264 3260 10676 3300
tri 10676 3260 10716 3300 sw
tri 10774 3260 10814 3300 ne
rect 10814 3260 11168 3300
tri 11168 3260 11266 3358 sw
tri 11266 3260 11364 3358 ne
rect 11364 3300 11688 3358
tri 11688 3300 11776 3388 sw
tri 11786 3300 11874 3388 ne
rect 11874 3358 12188 3388
tri 12188 3358 12268 3438 sw
tri 12286 3358 12366 3438 ne
rect 12366 3388 12690 3438
tri 12690 3388 12788 3486 sw
tri 12788 3388 12886 3486 ne
rect 12886 3438 13200 3486
tri 13200 3438 13288 3526 sw
tri 13298 3438 13386 3526 ne
rect 13386 3490 13440 3526
rect 13560 3490 15775 3610
rect 13386 3438 15775 3490
rect 12886 3388 13288 3438
rect 12366 3358 12788 3388
rect 11874 3300 12268 3358
rect 11364 3260 11776 3300
tri 11776 3260 11816 3300 sw
tri 11874 3260 11914 3300 ne
rect 11914 3260 12268 3300
tri 12268 3260 12366 3358 sw
tri 12366 3260 12464 3358 ne
rect 12464 3300 12788 3358
tri 12788 3300 12876 3388 sw
tri 12886 3300 12974 3388 ne
rect 12974 3358 13288 3388
tri 13288 3358 13368 3438 sw
tri 13386 3358 13466 3438 ne
rect 13466 3358 14075 3438
rect 12974 3300 13368 3358
rect 12464 3260 12876 3300
tri 12876 3260 12916 3300 sw
tri 12974 3260 13014 3300 ne
rect 13014 3260 13368 3300
tri 13368 3260 13466 3358 sw
tri 13466 3260 13564 3358 ne
rect 13564 3338 14075 3358
rect 14175 3338 15775 3438
rect 13564 3260 15775 3338
rect -1025 3212 -284 3260
rect -1025 3112 -925 3212
rect -825 3162 -284 3212
tri -284 3162 -186 3260 sw
tri -186 3162 -88 3260 ne
rect -88 3162 266 3260
tri 266 3162 364 3260 sw
tri 364 3162 462 3260 ne
rect 462 3162 816 3260
tri 816 3162 914 3260 sw
tri 914 3162 1012 3260 ne
rect 1012 3162 1366 3260
tri 1366 3162 1464 3260 sw
tri 1464 3162 1562 3260 ne
rect 1562 3162 1916 3260
tri 1916 3162 2014 3260 sw
tri 2014 3162 2112 3260 ne
rect 2112 3162 2466 3260
tri 2466 3162 2564 3260 sw
tri 2564 3162 2662 3260 ne
rect 2662 3162 3016 3260
tri 3016 3162 3114 3260 sw
tri 3114 3162 3212 3260 ne
rect 3212 3162 3566 3260
tri 3566 3162 3664 3260 sw
tri 3664 3162 3762 3260 ne
rect 3762 3162 4116 3260
tri 4116 3162 4214 3260 sw
tri 4214 3162 4312 3260 ne
rect 4312 3162 4666 3260
tri 4666 3162 4764 3260 sw
tri 4764 3162 4862 3260 ne
rect 4862 3162 5216 3260
tri 5216 3162 5314 3260 sw
tri 5314 3162 5412 3260 ne
rect 5412 3162 5766 3260
tri 5766 3162 5864 3260 sw
tri 5864 3162 5962 3260 ne
rect 5962 3162 6316 3260
tri 6316 3162 6414 3260 sw
tri 6414 3162 6512 3260 ne
rect 6512 3162 6866 3260
tri 6866 3162 6964 3260 sw
tri 6964 3162 7062 3260 ne
rect 7062 3162 7416 3260
tri 7416 3162 7514 3260 sw
tri 7514 3162 7612 3260 ne
rect 7612 3162 7966 3260
tri 7966 3162 8064 3260 sw
tri 8064 3162 8162 3260 ne
rect 8162 3162 8516 3260
tri 8516 3162 8614 3260 sw
tri 8614 3162 8712 3260 ne
rect 8712 3162 9066 3260
tri 9066 3162 9164 3260 sw
tri 9164 3162 9262 3260 ne
rect 9262 3162 9616 3260
tri 9616 3162 9714 3260 sw
tri 9714 3162 9812 3260 ne
rect 9812 3162 10166 3260
tri 10166 3162 10264 3260 sw
tri 10264 3162 10362 3260 ne
rect 10362 3162 10716 3260
tri 10716 3162 10814 3260 sw
tri 10814 3162 10912 3260 ne
rect 10912 3162 11266 3260
tri 11266 3162 11364 3260 sw
tri 11364 3162 11462 3260 ne
rect 11462 3162 11816 3260
tri 11816 3162 11914 3260 sw
tri 11914 3162 12012 3260 ne
rect 12012 3162 12366 3260
tri 12366 3162 12464 3260 sw
tri 12464 3162 12562 3260 ne
rect 12562 3162 12916 3260
tri 12916 3162 13014 3260 sw
tri 13014 3162 13112 3260 ne
rect 13112 3162 13466 3260
tri 13466 3162 13564 3260 sw
tri 13564 3162 13662 3260 ne
rect 13662 3162 15775 3260
rect -825 3112 -186 3162
rect -1025 3064 -186 3112
tri -186 3064 -88 3162 sw
tri -88 3064 10 3162 ne
rect 10 3064 364 3162
tri 364 3064 462 3162 sw
tri 462 3064 560 3162 ne
rect 560 3064 914 3162
tri 914 3064 1012 3162 sw
tri 1012 3064 1110 3162 ne
rect 1110 3064 1464 3162
tri 1464 3064 1562 3162 sw
tri 1562 3064 1660 3162 ne
rect 1660 3064 2014 3162
tri 2014 3064 2112 3162 sw
tri 2112 3064 2210 3162 ne
rect 2210 3064 2564 3162
tri 2564 3064 2662 3162 sw
tri 2662 3064 2760 3162 ne
rect 2760 3064 3114 3162
tri 3114 3064 3212 3162 sw
tri 3212 3064 3310 3162 ne
rect 3310 3064 3664 3162
tri 3664 3064 3762 3162 sw
tri 3762 3064 3860 3162 ne
rect 3860 3064 4214 3162
tri 4214 3064 4312 3162 sw
tri 4312 3064 4410 3162 ne
rect 4410 3064 4764 3162
tri 4764 3064 4862 3162 sw
tri 4862 3064 4960 3162 ne
rect 4960 3064 5314 3162
tri 5314 3064 5412 3162 sw
tri 5412 3064 5510 3162 ne
rect 5510 3064 5864 3162
tri 5864 3064 5962 3162 sw
tri 5962 3064 6060 3162 ne
rect 6060 3064 6414 3162
tri 6414 3064 6512 3162 sw
tri 6512 3064 6610 3162 ne
rect 6610 3064 6964 3162
tri 6964 3064 7062 3162 sw
tri 7062 3064 7160 3162 ne
rect 7160 3064 7514 3162
tri 7514 3064 7612 3162 sw
tri 7612 3064 7710 3162 ne
rect 7710 3064 8064 3162
tri 8064 3064 8162 3162 sw
tri 8162 3064 8260 3162 ne
rect 8260 3064 8614 3162
tri 8614 3064 8712 3162 sw
tri 8712 3064 8810 3162 ne
rect 8810 3064 9164 3162
tri 9164 3064 9262 3162 sw
tri 9262 3064 9360 3162 ne
rect 9360 3064 9714 3162
tri 9714 3064 9812 3162 sw
tri 9812 3064 9910 3162 ne
rect 9910 3064 10264 3162
tri 10264 3064 10362 3162 sw
tri 10362 3064 10460 3162 ne
rect 10460 3064 10814 3162
tri 10814 3064 10912 3162 sw
tri 10912 3064 11010 3162 ne
rect 11010 3064 11364 3162
tri 11364 3064 11462 3162 sw
tri 11462 3064 11560 3162 ne
rect 11560 3064 11914 3162
tri 11914 3064 12012 3162 sw
tri 12012 3064 12110 3162 ne
rect 12110 3064 12464 3162
tri 12464 3064 12562 3162 sw
tri 12562 3064 12660 3162 ne
rect 12660 3064 13014 3162
tri 13014 3064 13112 3162 sw
tri 13112 3064 13210 3162 ne
rect 13210 3064 13564 3162
tri 13564 3064 13662 3162 sw
rect -1025 3060 -88 3064
rect -1025 2940 -310 3060
rect -190 2976 -88 3060
tri -88 2976 0 3064 sw
tri 10 2976 98 3064 ne
rect 98 3060 462 3064
rect 98 2976 240 3060
rect -190 2940 0 2976
rect -1025 2936 0 2940
tri 0 2936 40 2976 sw
tri 98 2936 138 2976 ne
rect 138 2940 240 2976
rect 360 2976 462 3060
tri 462 2976 550 3064 sw
tri 560 2976 648 3064 ne
rect 648 3060 1012 3064
rect 648 2976 790 3060
rect 360 2940 550 2976
rect 138 2936 550 2940
tri -412 2838 -314 2936 ne
rect -314 2838 40 2936
tri 40 2838 138 2936 sw
tri 138 2838 236 2936 ne
rect 236 2888 550 2936
tri 550 2888 638 2976 sw
tri 648 2888 736 2976 ne
rect 736 2940 790 2976
rect 910 2976 1012 3060
tri 1012 2976 1100 3064 sw
tri 1110 2976 1198 3064 ne
rect 1198 3060 1562 3064
rect 1198 2976 1340 3060
rect 910 2940 1100 2976
rect 736 2936 1100 2940
tri 1100 2936 1140 2976 sw
tri 1198 2936 1238 2976 ne
rect 1238 2940 1340 2976
rect 1460 2976 1562 3060
tri 1562 2976 1650 3064 sw
tri 1660 2976 1748 3064 ne
rect 1748 3060 2112 3064
rect 1748 2976 1890 3060
rect 1460 2940 1650 2976
rect 1238 2936 1650 2940
rect 736 2888 1140 2936
rect 236 2838 638 2888
rect -2525 2750 -412 2838
tri -412 2750 -324 2838 sw
tri -314 2750 -226 2838 ne
rect -226 2750 138 2838
tri 138 2750 226 2838 sw
tri 236 2750 324 2838 ne
rect 324 2808 638 2838
tri 638 2808 718 2888 sw
tri 736 2808 816 2888 ne
rect 816 2838 1140 2888
tri 1140 2838 1238 2936 sw
tri 1238 2838 1336 2936 ne
rect 1336 2888 1650 2936
tri 1650 2888 1738 2976 sw
tri 1748 2888 1836 2976 ne
rect 1836 2940 1890 2976
rect 2010 2976 2112 3060
tri 2112 2976 2200 3064 sw
tri 2210 2976 2298 3064 ne
rect 2298 3060 2662 3064
rect 2298 2976 2440 3060
rect 2010 2940 2200 2976
rect 1836 2936 2200 2940
tri 2200 2936 2240 2976 sw
tri 2298 2936 2338 2976 ne
rect 2338 2940 2440 2976
rect 2560 2976 2662 3060
tri 2662 2976 2750 3064 sw
tri 2760 2976 2848 3064 ne
rect 2848 3060 3212 3064
rect 2848 2976 2990 3060
rect 2560 2940 2750 2976
rect 2338 2936 2750 2940
rect 1836 2888 2240 2936
rect 1336 2838 1738 2888
rect 816 2808 1238 2838
rect 324 2750 718 2808
rect -2525 2710 -324 2750
tri -324 2710 -284 2750 sw
tri -226 2710 -186 2750 ne
rect -186 2710 226 2750
tri 226 2710 266 2750 sw
tri 324 2710 364 2750 ne
rect 364 2710 718 2750
tri 718 2710 816 2808 sw
tri 816 2710 914 2808 ne
rect 914 2750 1238 2808
tri 1238 2750 1326 2838 sw
tri 1336 2750 1424 2838 ne
rect 1424 2808 1738 2838
tri 1738 2808 1818 2888 sw
tri 1836 2808 1916 2888 ne
rect 1916 2838 2240 2888
tri 2240 2838 2338 2936 sw
tri 2338 2838 2436 2936 ne
rect 2436 2888 2750 2936
tri 2750 2888 2838 2976 sw
tri 2848 2888 2936 2976 ne
rect 2936 2940 2990 2976
rect 3110 2976 3212 3060
tri 3212 2976 3300 3064 sw
tri 3310 2976 3398 3064 ne
rect 3398 3060 3762 3064
rect 3398 2976 3540 3060
rect 3110 2940 3300 2976
rect 2936 2936 3300 2940
tri 3300 2936 3340 2976 sw
tri 3398 2936 3438 2976 ne
rect 3438 2940 3540 2976
rect 3660 2976 3762 3060
tri 3762 2976 3850 3064 sw
tri 3860 2976 3948 3064 ne
rect 3948 3060 4312 3064
rect 3948 2976 4090 3060
rect 3660 2940 3850 2976
rect 3438 2936 3850 2940
rect 2936 2888 3340 2936
rect 2436 2838 2838 2888
rect 1916 2808 2338 2838
rect 1424 2750 1818 2808
rect 914 2710 1326 2750
tri 1326 2710 1366 2750 sw
tri 1424 2710 1464 2750 ne
rect 1464 2710 1818 2750
tri 1818 2710 1916 2808 sw
tri 1916 2710 2014 2808 ne
rect 2014 2750 2338 2808
tri 2338 2750 2426 2838 sw
tri 2436 2750 2524 2838 ne
rect 2524 2808 2838 2838
tri 2838 2808 2918 2888 sw
tri 2936 2808 3016 2888 ne
rect 3016 2838 3340 2888
tri 3340 2838 3438 2936 sw
tri 3438 2838 3536 2936 ne
rect 3536 2888 3850 2936
tri 3850 2888 3938 2976 sw
tri 3948 2888 4036 2976 ne
rect 4036 2940 4090 2976
rect 4210 2976 4312 3060
tri 4312 2976 4400 3064 sw
tri 4410 2976 4498 3064 ne
rect 4498 3060 4862 3064
rect 4498 2976 4640 3060
rect 4210 2940 4400 2976
rect 4036 2936 4400 2940
tri 4400 2936 4440 2976 sw
tri 4498 2936 4538 2976 ne
rect 4538 2940 4640 2976
rect 4760 2976 4862 3060
tri 4862 2976 4950 3064 sw
tri 4960 2976 5048 3064 ne
rect 5048 3060 5412 3064
rect 5048 2976 5190 3060
rect 4760 2940 4950 2976
rect 4538 2936 4950 2940
rect 4036 2888 4440 2936
rect 3536 2838 3938 2888
rect 3016 2808 3438 2838
rect 2524 2750 2918 2808
rect 2014 2710 2426 2750
tri 2426 2710 2466 2750 sw
tri 2524 2710 2564 2750 ne
rect 2564 2710 2918 2750
tri 2918 2710 3016 2808 sw
tri 3016 2710 3114 2808 ne
rect 3114 2750 3438 2808
tri 3438 2750 3526 2838 sw
tri 3536 2750 3624 2838 ne
rect 3624 2808 3938 2838
tri 3938 2808 4018 2888 sw
tri 4036 2808 4116 2888 ne
rect 4116 2838 4440 2888
tri 4440 2838 4538 2936 sw
tri 4538 2838 4636 2936 ne
rect 4636 2888 4950 2936
tri 4950 2888 5038 2976 sw
tri 5048 2888 5136 2976 ne
rect 5136 2940 5190 2976
rect 5310 2976 5412 3060
tri 5412 2976 5500 3064 sw
tri 5510 2976 5598 3064 ne
rect 5598 3060 5962 3064
rect 5598 2976 5740 3060
rect 5310 2940 5500 2976
rect 5136 2936 5500 2940
tri 5500 2936 5540 2976 sw
tri 5598 2936 5638 2976 ne
rect 5638 2940 5740 2976
rect 5860 2976 5962 3060
tri 5962 2976 6050 3064 sw
tri 6060 2976 6148 3064 ne
rect 6148 3060 6512 3064
rect 6148 2976 6290 3060
rect 5860 2940 6050 2976
rect 5638 2936 6050 2940
rect 5136 2888 5540 2936
rect 4636 2838 5038 2888
rect 4116 2808 4538 2838
rect 3624 2750 4018 2808
rect 3114 2710 3526 2750
tri 3526 2710 3566 2750 sw
tri 3624 2710 3664 2750 ne
rect 3664 2710 4018 2750
tri 4018 2710 4116 2808 sw
tri 4116 2710 4214 2808 ne
rect 4214 2750 4538 2808
tri 4538 2750 4626 2838 sw
tri 4636 2750 4724 2838 ne
rect 4724 2808 5038 2838
tri 5038 2808 5118 2888 sw
tri 5136 2808 5216 2888 ne
rect 5216 2838 5540 2888
tri 5540 2838 5638 2936 sw
tri 5638 2838 5736 2936 ne
rect 5736 2888 6050 2936
tri 6050 2888 6138 2976 sw
tri 6148 2888 6236 2976 ne
rect 6236 2940 6290 2976
rect 6410 2976 6512 3060
tri 6512 2976 6600 3064 sw
tri 6610 2976 6698 3064 ne
rect 6698 3060 7062 3064
rect 6698 2976 6840 3060
rect 6410 2940 6600 2976
rect 6236 2936 6600 2940
tri 6600 2936 6640 2976 sw
tri 6698 2936 6738 2976 ne
rect 6738 2940 6840 2976
rect 6960 2976 7062 3060
tri 7062 2976 7150 3064 sw
tri 7160 2976 7248 3064 ne
rect 7248 3060 7612 3064
rect 7248 2976 7390 3060
rect 6960 2940 7150 2976
rect 6738 2936 7150 2940
rect 6236 2888 6640 2936
rect 5736 2838 6138 2888
rect 5216 2808 5638 2838
rect 4724 2750 5118 2808
rect 4214 2710 4626 2750
tri 4626 2710 4666 2750 sw
tri 4724 2710 4764 2750 ne
rect 4764 2710 5118 2750
tri 5118 2710 5216 2808 sw
tri 5216 2710 5314 2808 ne
rect 5314 2750 5638 2808
tri 5638 2750 5726 2838 sw
tri 5736 2750 5824 2838 ne
rect 5824 2808 6138 2838
tri 6138 2808 6218 2888 sw
tri 6236 2808 6316 2888 ne
rect 6316 2838 6640 2888
tri 6640 2838 6738 2936 sw
tri 6738 2838 6836 2936 ne
rect 6836 2888 7150 2936
tri 7150 2888 7238 2976 sw
tri 7248 2888 7336 2976 ne
rect 7336 2940 7390 2976
rect 7510 2976 7612 3060
tri 7612 2976 7700 3064 sw
tri 7710 2976 7798 3064 ne
rect 7798 3060 8162 3064
rect 7798 2976 7940 3060
rect 7510 2940 7700 2976
rect 7336 2936 7700 2940
tri 7700 2936 7740 2976 sw
tri 7798 2936 7838 2976 ne
rect 7838 2940 7940 2976
rect 8060 2976 8162 3060
tri 8162 2976 8250 3064 sw
tri 8260 2976 8348 3064 ne
rect 8348 3060 8712 3064
rect 8348 2976 8490 3060
rect 8060 2940 8250 2976
rect 7838 2936 8250 2940
rect 7336 2888 7740 2936
rect 6836 2838 7238 2888
rect 6316 2808 6738 2838
rect 5824 2750 6218 2808
rect 5314 2710 5726 2750
tri 5726 2710 5766 2750 sw
tri 5824 2710 5864 2750 ne
rect 5864 2710 6218 2750
tri 6218 2710 6316 2808 sw
tri 6316 2710 6414 2808 ne
rect 6414 2750 6738 2808
tri 6738 2750 6826 2838 sw
tri 6836 2750 6924 2838 ne
rect 6924 2808 7238 2838
tri 7238 2808 7318 2888 sw
tri 7336 2808 7416 2888 ne
rect 7416 2838 7740 2888
tri 7740 2838 7838 2936 sw
tri 7838 2838 7936 2936 ne
rect 7936 2888 8250 2936
tri 8250 2888 8338 2976 sw
tri 8348 2888 8436 2976 ne
rect 8436 2940 8490 2976
rect 8610 2976 8712 3060
tri 8712 2976 8800 3064 sw
tri 8810 2976 8898 3064 ne
rect 8898 3060 9262 3064
rect 8898 2976 9040 3060
rect 8610 2940 8800 2976
rect 8436 2936 8800 2940
tri 8800 2936 8840 2976 sw
tri 8898 2936 8938 2976 ne
rect 8938 2940 9040 2976
rect 9160 2976 9262 3060
tri 9262 2976 9350 3064 sw
tri 9360 2976 9448 3064 ne
rect 9448 3060 9812 3064
rect 9448 2976 9590 3060
rect 9160 2940 9350 2976
rect 8938 2936 9350 2940
rect 8436 2888 8840 2936
rect 7936 2838 8338 2888
rect 7416 2808 7838 2838
rect 6924 2750 7318 2808
rect 6414 2710 6826 2750
tri 6826 2710 6866 2750 sw
tri 6924 2710 6964 2750 ne
rect 6964 2710 7318 2750
tri 7318 2710 7416 2808 sw
tri 7416 2710 7514 2808 ne
rect 7514 2750 7838 2808
tri 7838 2750 7926 2838 sw
tri 7936 2750 8024 2838 ne
rect 8024 2808 8338 2838
tri 8338 2808 8418 2888 sw
tri 8436 2808 8516 2888 ne
rect 8516 2838 8840 2888
tri 8840 2838 8938 2936 sw
tri 8938 2838 9036 2936 ne
rect 9036 2888 9350 2936
tri 9350 2888 9438 2976 sw
tri 9448 2888 9536 2976 ne
rect 9536 2940 9590 2976
rect 9710 2976 9812 3060
tri 9812 2976 9900 3064 sw
tri 9910 2976 9998 3064 ne
rect 9998 3060 10362 3064
rect 9998 2976 10140 3060
rect 9710 2940 9900 2976
rect 9536 2936 9900 2940
tri 9900 2936 9940 2976 sw
tri 9998 2936 10038 2976 ne
rect 10038 2940 10140 2976
rect 10260 2976 10362 3060
tri 10362 2976 10450 3064 sw
tri 10460 2976 10548 3064 ne
rect 10548 3060 10912 3064
rect 10548 2976 10690 3060
rect 10260 2940 10450 2976
rect 10038 2936 10450 2940
rect 9536 2888 9940 2936
rect 9036 2838 9438 2888
rect 8516 2808 8938 2838
rect 8024 2750 8418 2808
rect 7514 2710 7926 2750
tri 7926 2710 7966 2750 sw
tri 8024 2710 8064 2750 ne
rect 8064 2710 8418 2750
tri 8418 2710 8516 2808 sw
tri 8516 2710 8614 2808 ne
rect 8614 2750 8938 2808
tri 8938 2750 9026 2838 sw
tri 9036 2750 9124 2838 ne
rect 9124 2808 9438 2838
tri 9438 2808 9518 2888 sw
tri 9536 2808 9616 2888 ne
rect 9616 2838 9940 2888
tri 9940 2838 10038 2936 sw
tri 10038 2838 10136 2936 ne
rect 10136 2888 10450 2936
tri 10450 2888 10538 2976 sw
tri 10548 2888 10636 2976 ne
rect 10636 2940 10690 2976
rect 10810 2976 10912 3060
tri 10912 2976 11000 3064 sw
tri 11010 2976 11098 3064 ne
rect 11098 3060 11462 3064
rect 11098 2976 11240 3060
rect 10810 2940 11000 2976
rect 10636 2936 11000 2940
tri 11000 2936 11040 2976 sw
tri 11098 2936 11138 2976 ne
rect 11138 2940 11240 2976
rect 11360 2976 11462 3060
tri 11462 2976 11550 3064 sw
tri 11560 2976 11648 3064 ne
rect 11648 3060 12012 3064
rect 11648 2976 11790 3060
rect 11360 2940 11550 2976
rect 11138 2936 11550 2940
rect 10636 2888 11040 2936
rect 10136 2838 10538 2888
rect 9616 2808 10038 2838
rect 9124 2750 9518 2808
rect 8614 2710 9026 2750
tri 9026 2710 9066 2750 sw
tri 9124 2710 9164 2750 ne
rect 9164 2710 9518 2750
tri 9518 2710 9616 2808 sw
tri 9616 2710 9714 2808 ne
rect 9714 2750 10038 2808
tri 10038 2750 10126 2838 sw
tri 10136 2750 10224 2838 ne
rect 10224 2808 10538 2838
tri 10538 2808 10618 2888 sw
tri 10636 2808 10716 2888 ne
rect 10716 2838 11040 2888
tri 11040 2838 11138 2936 sw
tri 11138 2838 11236 2936 ne
rect 11236 2888 11550 2936
tri 11550 2888 11638 2976 sw
tri 11648 2888 11736 2976 ne
rect 11736 2940 11790 2976
rect 11910 2976 12012 3060
tri 12012 2976 12100 3064 sw
tri 12110 2976 12198 3064 ne
rect 12198 3060 12562 3064
rect 12198 2976 12340 3060
rect 11910 2940 12100 2976
rect 11736 2936 12100 2940
tri 12100 2936 12140 2976 sw
tri 12198 2936 12238 2976 ne
rect 12238 2940 12340 2976
rect 12460 2976 12562 3060
tri 12562 2976 12650 3064 sw
tri 12660 2976 12748 3064 ne
rect 12748 3060 13112 3064
rect 12748 2976 12890 3060
rect 12460 2940 12650 2976
rect 12238 2936 12650 2940
rect 11736 2888 12140 2936
rect 11236 2838 11638 2888
rect 10716 2808 11138 2838
rect 10224 2750 10618 2808
rect 9714 2710 10126 2750
tri 10126 2710 10166 2750 sw
tri 10224 2710 10264 2750 ne
rect 10264 2710 10618 2750
tri 10618 2710 10716 2808 sw
tri 10716 2710 10814 2808 ne
rect 10814 2750 11138 2808
tri 11138 2750 11226 2838 sw
tri 11236 2750 11324 2838 ne
rect 11324 2808 11638 2838
tri 11638 2808 11718 2888 sw
tri 11736 2808 11816 2888 ne
rect 11816 2838 12140 2888
tri 12140 2838 12238 2936 sw
tri 12238 2838 12336 2936 ne
rect 12336 2888 12650 2936
tri 12650 2888 12738 2976 sw
tri 12748 2888 12836 2976 ne
rect 12836 2940 12890 2976
rect 13010 2976 13112 3060
tri 13112 2976 13200 3064 sw
tri 13210 2976 13298 3064 ne
rect 13298 3060 14275 3064
rect 13298 2976 13440 3060
rect 13010 2940 13200 2976
rect 12836 2936 13200 2940
tri 13200 2936 13240 2976 sw
tri 13298 2936 13338 2976 ne
rect 13338 2940 13440 2976
rect 13560 2940 14275 3060
rect 13338 2936 14275 2940
rect 12836 2888 13240 2936
rect 12336 2838 12738 2888
rect 11816 2808 12238 2838
rect 11324 2750 11718 2808
rect 10814 2710 11226 2750
tri 11226 2710 11266 2750 sw
tri 11324 2710 11364 2750 ne
rect 11364 2710 11718 2750
tri 11718 2710 11816 2808 sw
tri 11816 2710 11914 2808 ne
rect 11914 2750 12238 2808
tri 12238 2750 12326 2838 sw
tri 12336 2750 12424 2838 ne
rect 12424 2808 12738 2838
tri 12738 2808 12818 2888 sw
tri 12836 2808 12916 2888 ne
rect 12916 2838 13240 2888
tri 13240 2838 13338 2936 sw
tri 13338 2838 13436 2936 ne
rect 13436 2838 14275 2936
rect 12916 2808 13338 2838
rect 12424 2750 12818 2808
rect 11914 2710 12326 2750
tri 12326 2710 12366 2750 sw
tri 12424 2710 12464 2750 ne
rect 12464 2710 12818 2750
tri 12818 2710 12916 2808 sw
tri 12916 2710 13014 2808 ne
rect 13014 2750 13338 2808
tri 13338 2750 13426 2838 sw
tri 13436 2750 13524 2838 ne
rect 13524 2750 14275 2838
rect 13014 2710 13426 2750
tri 13426 2710 13466 2750 sw
tri 13524 2710 13564 2750 ne
rect 13564 2710 14275 2750
rect -2525 2612 -284 2710
tri -284 2612 -186 2710 sw
tri -186 2612 -88 2710 ne
rect -88 2612 266 2710
tri 266 2612 364 2710 sw
tri 364 2612 462 2710 ne
rect 462 2612 816 2710
tri 816 2612 914 2710 sw
tri 914 2612 1012 2710 ne
rect 1012 2612 1366 2710
tri 1366 2612 1464 2710 sw
tri 1464 2612 1562 2710 ne
rect 1562 2612 1916 2710
tri 1916 2612 2014 2710 sw
tri 2014 2612 2112 2710 ne
rect 2112 2612 2466 2710
tri 2466 2612 2564 2710 sw
tri 2564 2612 2662 2710 ne
rect 2662 2612 3016 2710
tri 3016 2612 3114 2710 sw
tri 3114 2612 3212 2710 ne
rect 3212 2612 3566 2710
tri 3566 2612 3664 2710 sw
tri 3664 2612 3762 2710 ne
rect 3762 2612 4116 2710
tri 4116 2612 4214 2710 sw
tri 4214 2612 4312 2710 ne
rect 4312 2612 4666 2710
tri 4666 2612 4764 2710 sw
tri 4764 2612 4862 2710 ne
rect 4862 2612 5216 2710
tri 5216 2612 5314 2710 sw
tri 5314 2612 5412 2710 ne
rect 5412 2612 5766 2710
tri 5766 2612 5864 2710 sw
tri 5864 2612 5962 2710 ne
rect 5962 2612 6316 2710
tri 6316 2612 6414 2710 sw
tri 6414 2612 6512 2710 ne
rect 6512 2612 6866 2710
tri 6866 2612 6964 2710 sw
tri 6964 2612 7062 2710 ne
rect 7062 2612 7416 2710
tri 7416 2612 7514 2710 sw
tri 7514 2612 7612 2710 ne
rect 7612 2612 7966 2710
tri 7966 2612 8064 2710 sw
tri 8064 2612 8162 2710 ne
rect 8162 2612 8516 2710
tri 8516 2612 8614 2710 sw
tri 8614 2612 8712 2710 ne
rect 8712 2612 9066 2710
tri 9066 2612 9164 2710 sw
tri 9164 2612 9262 2710 ne
rect 9262 2612 9616 2710
tri 9616 2612 9714 2710 sw
tri 9714 2612 9812 2710 ne
rect 9812 2612 10166 2710
tri 10166 2612 10264 2710 sw
tri 10264 2612 10362 2710 ne
rect 10362 2612 10716 2710
tri 10716 2612 10814 2710 sw
tri 10814 2612 10912 2710 ne
rect 10912 2612 11266 2710
tri 11266 2612 11364 2710 sw
tri 11364 2612 11462 2710 ne
rect 11462 2612 11816 2710
tri 11816 2612 11914 2710 sw
tri 11914 2612 12012 2710 ne
rect 12012 2612 12366 2710
tri 12366 2612 12464 2710 sw
tri 12464 2612 12562 2710 ne
rect 12562 2612 12916 2710
tri 12916 2612 13014 2710 sw
tri 13014 2612 13112 2710 ne
rect 13112 2612 13466 2710
tri 13466 2612 13564 2710 sw
tri 13564 2612 13662 2710 ne
rect 13662 2612 14275 2710
rect -2525 2514 -186 2612
tri -186 2514 -88 2612 sw
tri -88 2514 10 2612 ne
rect 10 2514 364 2612
tri 364 2514 462 2612 sw
tri 462 2514 560 2612 ne
rect 560 2514 914 2612
tri 914 2514 1012 2612 sw
tri 1012 2514 1110 2612 ne
rect 1110 2514 1464 2612
tri 1464 2514 1562 2612 sw
tri 1562 2514 1660 2612 ne
rect 1660 2514 2014 2612
tri 2014 2514 2112 2612 sw
tri 2112 2514 2210 2612 ne
rect 2210 2514 2564 2612
tri 2564 2514 2662 2612 sw
tri 2662 2514 2760 2612 ne
rect 2760 2514 3114 2612
tri 3114 2514 3212 2612 sw
tri 3212 2514 3310 2612 ne
rect 3310 2514 3664 2612
tri 3664 2514 3762 2612 sw
tri 3762 2514 3860 2612 ne
rect 3860 2514 4214 2612
tri 4214 2514 4312 2612 sw
tri 4312 2514 4410 2612 ne
rect 4410 2514 4764 2612
tri 4764 2514 4862 2612 sw
tri 4862 2514 4960 2612 ne
rect 4960 2514 5314 2612
tri 5314 2514 5412 2612 sw
tri 5412 2514 5510 2612 ne
rect 5510 2514 5864 2612
tri 5864 2514 5962 2612 sw
tri 5962 2514 6060 2612 ne
rect 6060 2514 6414 2612
tri 6414 2514 6512 2612 sw
tri 6512 2514 6610 2612 ne
rect 6610 2514 6964 2612
tri 6964 2514 7062 2612 sw
tri 7062 2514 7160 2612 ne
rect 7160 2514 7514 2612
tri 7514 2514 7612 2612 sw
tri 7612 2514 7710 2612 ne
rect 7710 2514 8064 2612
tri 8064 2514 8162 2612 sw
tri 8162 2514 8260 2612 ne
rect 8260 2514 8614 2612
tri 8614 2514 8712 2612 sw
tri 8712 2514 8810 2612 ne
rect 8810 2514 9164 2612
tri 9164 2514 9262 2612 sw
tri 9262 2514 9360 2612 ne
rect 9360 2514 9714 2612
tri 9714 2514 9812 2612 sw
tri 9812 2514 9910 2612 ne
rect 9910 2514 10264 2612
tri 10264 2514 10362 2612 sw
tri 10362 2514 10460 2612 ne
rect 10460 2514 10814 2612
tri 10814 2514 10912 2612 sw
tri 10912 2514 11010 2612 ne
rect 11010 2514 11364 2612
tri 11364 2514 11462 2612 sw
tri 11462 2514 11560 2612 ne
rect 11560 2514 11914 2612
tri 11914 2514 12012 2612 sw
tri 12012 2514 12110 2612 ne
rect 12110 2514 12464 2612
tri 12464 2514 12562 2612 sw
tri 12562 2514 12660 2612 ne
rect 12660 2514 13014 2612
tri 13014 2514 13112 2612 sw
tri 13112 2514 13210 2612 ne
rect 13210 2514 13564 2612
tri 13564 2514 13662 2612 sw
rect 14775 2514 15775 3162
rect -2525 2510 -88 2514
rect -2525 2390 -310 2510
rect -190 2426 -88 2510
tri -88 2426 0 2514 sw
tri 10 2426 98 2514 ne
rect 98 2510 462 2514
rect 98 2426 240 2510
rect -190 2390 0 2426
rect -2525 2386 0 2390
rect -2525 1738 -1525 2386
tri -412 2288 -314 2386 ne
rect -314 2338 0 2386
tri 0 2338 88 2426 sw
tri 98 2338 186 2426 ne
rect 186 2390 240 2426
rect 360 2426 462 2510
tri 462 2426 550 2514 sw
tri 560 2426 648 2514 ne
rect 648 2510 1012 2514
rect 648 2426 790 2510
rect 360 2390 550 2426
rect 186 2386 550 2390
tri 550 2386 590 2426 sw
tri 648 2386 688 2426 ne
rect 688 2390 790 2426
rect 910 2426 1012 2510
tri 1012 2426 1100 2514 sw
tri 1110 2426 1198 2514 ne
rect 1198 2510 1562 2514
rect 1198 2426 1340 2510
rect 910 2390 1100 2426
rect 688 2386 1100 2390
rect 186 2338 590 2386
rect -314 2288 88 2338
rect -1025 2200 -412 2288
tri -412 2200 -324 2288 sw
tri -314 2200 -226 2288 ne
rect -226 2258 88 2288
tri 88 2258 168 2338 sw
tri 186 2258 266 2338 ne
rect 266 2288 590 2338
tri 590 2288 688 2386 sw
tri 688 2288 786 2386 ne
rect 786 2338 1100 2386
tri 1100 2338 1188 2426 sw
tri 1198 2338 1286 2426 ne
rect 1286 2390 1340 2426
rect 1460 2426 1562 2510
tri 1562 2426 1650 2514 sw
tri 1660 2426 1748 2514 ne
rect 1748 2510 2112 2514
rect 1748 2426 1890 2510
rect 1460 2390 1650 2426
rect 1286 2386 1650 2390
tri 1650 2386 1690 2426 sw
tri 1748 2386 1788 2426 ne
rect 1788 2390 1890 2426
rect 2010 2426 2112 2510
tri 2112 2426 2200 2514 sw
tri 2210 2426 2298 2514 ne
rect 2298 2510 2662 2514
rect 2298 2426 2440 2510
rect 2010 2390 2200 2426
rect 1788 2386 2200 2390
rect 1286 2338 1690 2386
rect 786 2288 1188 2338
rect 266 2258 688 2288
rect -226 2200 168 2258
rect -1025 2160 -324 2200
tri -324 2160 -284 2200 sw
tri -226 2160 -186 2200 ne
rect -186 2160 168 2200
tri 168 2160 266 2258 sw
tri 266 2160 364 2258 ne
rect 364 2200 688 2258
tri 688 2200 776 2288 sw
tri 786 2200 874 2288 ne
rect 874 2258 1188 2288
tri 1188 2258 1268 2338 sw
tri 1286 2258 1366 2338 ne
rect 1366 2288 1690 2338
tri 1690 2288 1788 2386 sw
tri 1788 2288 1886 2386 ne
rect 1886 2338 2200 2386
tri 2200 2338 2288 2426 sw
tri 2298 2338 2386 2426 ne
rect 2386 2390 2440 2426
rect 2560 2426 2662 2510
tri 2662 2426 2750 2514 sw
tri 2760 2426 2848 2514 ne
rect 2848 2510 3212 2514
rect 2848 2426 2990 2510
rect 2560 2390 2750 2426
rect 2386 2386 2750 2390
tri 2750 2386 2790 2426 sw
tri 2848 2386 2888 2426 ne
rect 2888 2390 2990 2426
rect 3110 2426 3212 2510
tri 3212 2426 3300 2514 sw
tri 3310 2426 3398 2514 ne
rect 3398 2510 3762 2514
rect 3398 2426 3540 2510
rect 3110 2390 3300 2426
rect 2888 2386 3300 2390
rect 2386 2338 2790 2386
rect 1886 2288 2288 2338
rect 1366 2258 1788 2288
rect 874 2200 1268 2258
rect 364 2160 776 2200
tri 776 2160 816 2200 sw
tri 874 2160 914 2200 ne
rect 914 2160 1268 2200
tri 1268 2160 1366 2258 sw
tri 1366 2160 1464 2258 ne
rect 1464 2200 1788 2258
tri 1788 2200 1876 2288 sw
tri 1886 2200 1974 2288 ne
rect 1974 2258 2288 2288
tri 2288 2258 2368 2338 sw
tri 2386 2258 2466 2338 ne
rect 2466 2288 2790 2338
tri 2790 2288 2888 2386 sw
tri 2888 2288 2986 2386 ne
rect 2986 2338 3300 2386
tri 3300 2338 3388 2426 sw
tri 3398 2338 3486 2426 ne
rect 3486 2390 3540 2426
rect 3660 2426 3762 2510
tri 3762 2426 3850 2514 sw
tri 3860 2426 3948 2514 ne
rect 3948 2510 4312 2514
rect 3948 2426 4090 2510
rect 3660 2390 3850 2426
rect 3486 2386 3850 2390
tri 3850 2386 3890 2426 sw
tri 3948 2386 3988 2426 ne
rect 3988 2390 4090 2426
rect 4210 2426 4312 2510
tri 4312 2426 4400 2514 sw
tri 4410 2426 4498 2514 ne
rect 4498 2510 4862 2514
rect 4498 2426 4640 2510
rect 4210 2390 4400 2426
rect 3988 2386 4400 2390
rect 3486 2338 3890 2386
rect 2986 2288 3388 2338
rect 2466 2258 2888 2288
rect 1974 2200 2368 2258
rect 1464 2160 1876 2200
tri 1876 2160 1916 2200 sw
tri 1974 2160 2014 2200 ne
rect 2014 2160 2368 2200
tri 2368 2160 2466 2258 sw
tri 2466 2160 2564 2258 ne
rect 2564 2200 2888 2258
tri 2888 2200 2976 2288 sw
tri 2986 2200 3074 2288 ne
rect 3074 2258 3388 2288
tri 3388 2258 3468 2338 sw
tri 3486 2258 3566 2338 ne
rect 3566 2288 3890 2338
tri 3890 2288 3988 2386 sw
tri 3988 2288 4086 2386 ne
rect 4086 2338 4400 2386
tri 4400 2338 4488 2426 sw
tri 4498 2338 4586 2426 ne
rect 4586 2390 4640 2426
rect 4760 2426 4862 2510
tri 4862 2426 4950 2514 sw
tri 4960 2426 5048 2514 ne
rect 5048 2510 5412 2514
rect 5048 2426 5190 2510
rect 4760 2390 4950 2426
rect 4586 2386 4950 2390
tri 4950 2386 4990 2426 sw
tri 5048 2386 5088 2426 ne
rect 5088 2390 5190 2426
rect 5310 2426 5412 2510
tri 5412 2426 5500 2514 sw
tri 5510 2426 5598 2514 ne
rect 5598 2510 5962 2514
rect 5598 2426 5740 2510
rect 5310 2390 5500 2426
rect 5088 2386 5500 2390
rect 4586 2338 4990 2386
rect 4086 2288 4488 2338
rect 3566 2258 3988 2288
rect 3074 2200 3468 2258
rect 2564 2160 2976 2200
tri 2976 2160 3016 2200 sw
tri 3074 2160 3114 2200 ne
rect 3114 2160 3468 2200
tri 3468 2160 3566 2258 sw
tri 3566 2160 3664 2258 ne
rect 3664 2200 3988 2258
tri 3988 2200 4076 2288 sw
tri 4086 2200 4174 2288 ne
rect 4174 2258 4488 2288
tri 4488 2258 4568 2338 sw
tri 4586 2258 4666 2338 ne
rect 4666 2288 4990 2338
tri 4990 2288 5088 2386 sw
tri 5088 2288 5186 2386 ne
rect 5186 2338 5500 2386
tri 5500 2338 5588 2426 sw
tri 5598 2338 5686 2426 ne
rect 5686 2390 5740 2426
rect 5860 2426 5962 2510
tri 5962 2426 6050 2514 sw
tri 6060 2426 6148 2514 ne
rect 6148 2510 6512 2514
rect 6148 2426 6290 2510
rect 5860 2390 6050 2426
rect 5686 2386 6050 2390
tri 6050 2386 6090 2426 sw
tri 6148 2386 6188 2426 ne
rect 6188 2390 6290 2426
rect 6410 2426 6512 2510
tri 6512 2426 6600 2514 sw
tri 6610 2426 6698 2514 ne
rect 6698 2510 7062 2514
rect 6698 2426 6840 2510
rect 6410 2390 6600 2426
rect 6188 2386 6600 2390
rect 5686 2338 6090 2386
rect 5186 2288 5588 2338
rect 4666 2258 5088 2288
rect 4174 2200 4568 2258
rect 3664 2160 4076 2200
tri 4076 2160 4116 2200 sw
tri 4174 2160 4214 2200 ne
rect 4214 2160 4568 2200
tri 4568 2160 4666 2258 sw
tri 4666 2160 4764 2258 ne
rect 4764 2200 5088 2258
tri 5088 2200 5176 2288 sw
tri 5186 2200 5274 2288 ne
rect 5274 2258 5588 2288
tri 5588 2258 5668 2338 sw
tri 5686 2258 5766 2338 ne
rect 5766 2288 6090 2338
tri 6090 2288 6188 2386 sw
tri 6188 2288 6286 2386 ne
rect 6286 2338 6600 2386
tri 6600 2338 6688 2426 sw
tri 6698 2338 6786 2426 ne
rect 6786 2390 6840 2426
rect 6960 2426 7062 2510
tri 7062 2426 7150 2514 sw
tri 7160 2426 7248 2514 ne
rect 7248 2510 7612 2514
rect 7248 2426 7390 2510
rect 6960 2390 7150 2426
rect 6786 2386 7150 2390
tri 7150 2386 7190 2426 sw
tri 7248 2386 7288 2426 ne
rect 7288 2390 7390 2426
rect 7510 2426 7612 2510
tri 7612 2426 7700 2514 sw
tri 7710 2426 7798 2514 ne
rect 7798 2510 8162 2514
rect 7798 2426 7940 2510
rect 7510 2390 7700 2426
rect 7288 2386 7700 2390
rect 6786 2338 7190 2386
rect 6286 2288 6688 2338
rect 5766 2258 6188 2288
rect 5274 2200 5668 2258
rect 4764 2160 5176 2200
tri 5176 2160 5216 2200 sw
tri 5274 2160 5314 2200 ne
rect 5314 2160 5668 2200
tri 5668 2160 5766 2258 sw
tri 5766 2160 5864 2258 ne
rect 5864 2200 6188 2258
tri 6188 2200 6276 2288 sw
tri 6286 2200 6374 2288 ne
rect 6374 2258 6688 2288
tri 6688 2258 6768 2338 sw
tri 6786 2258 6866 2338 ne
rect 6866 2288 7190 2338
tri 7190 2288 7288 2386 sw
tri 7288 2288 7386 2386 ne
rect 7386 2338 7700 2386
tri 7700 2338 7788 2426 sw
tri 7798 2338 7886 2426 ne
rect 7886 2390 7940 2426
rect 8060 2426 8162 2510
tri 8162 2426 8250 2514 sw
tri 8260 2426 8348 2514 ne
rect 8348 2510 8712 2514
rect 8348 2426 8490 2510
rect 8060 2390 8250 2426
rect 7886 2386 8250 2390
tri 8250 2386 8290 2426 sw
tri 8348 2386 8388 2426 ne
rect 8388 2390 8490 2426
rect 8610 2426 8712 2510
tri 8712 2426 8800 2514 sw
tri 8810 2426 8898 2514 ne
rect 8898 2510 9262 2514
rect 8898 2426 9040 2510
rect 8610 2390 8800 2426
rect 8388 2386 8800 2390
rect 7886 2338 8290 2386
rect 7386 2288 7788 2338
rect 6866 2258 7288 2288
rect 6374 2200 6768 2258
rect 5864 2160 6276 2200
tri 6276 2160 6316 2200 sw
tri 6374 2160 6414 2200 ne
rect 6414 2160 6768 2200
tri 6768 2160 6866 2258 sw
tri 6866 2160 6964 2258 ne
rect 6964 2200 7288 2258
tri 7288 2200 7376 2288 sw
tri 7386 2200 7474 2288 ne
rect 7474 2258 7788 2288
tri 7788 2258 7868 2338 sw
tri 7886 2258 7966 2338 ne
rect 7966 2288 8290 2338
tri 8290 2288 8388 2386 sw
tri 8388 2288 8486 2386 ne
rect 8486 2338 8800 2386
tri 8800 2338 8888 2426 sw
tri 8898 2338 8986 2426 ne
rect 8986 2390 9040 2426
rect 9160 2426 9262 2510
tri 9262 2426 9350 2514 sw
tri 9360 2426 9448 2514 ne
rect 9448 2510 9812 2514
rect 9448 2426 9590 2510
rect 9160 2390 9350 2426
rect 8986 2386 9350 2390
tri 9350 2386 9390 2426 sw
tri 9448 2386 9488 2426 ne
rect 9488 2390 9590 2426
rect 9710 2426 9812 2510
tri 9812 2426 9900 2514 sw
tri 9910 2426 9998 2514 ne
rect 9998 2510 10362 2514
rect 9998 2426 10140 2510
rect 9710 2390 9900 2426
rect 9488 2386 9900 2390
rect 8986 2338 9390 2386
rect 8486 2288 8888 2338
rect 7966 2258 8388 2288
rect 7474 2200 7868 2258
rect 6964 2160 7376 2200
tri 7376 2160 7416 2200 sw
tri 7474 2160 7514 2200 ne
rect 7514 2160 7868 2200
tri 7868 2160 7966 2258 sw
tri 7966 2160 8064 2258 ne
rect 8064 2200 8388 2258
tri 8388 2200 8476 2288 sw
tri 8486 2200 8574 2288 ne
rect 8574 2258 8888 2288
tri 8888 2258 8968 2338 sw
tri 8986 2258 9066 2338 ne
rect 9066 2288 9390 2338
tri 9390 2288 9488 2386 sw
tri 9488 2288 9586 2386 ne
rect 9586 2338 9900 2386
tri 9900 2338 9988 2426 sw
tri 9998 2338 10086 2426 ne
rect 10086 2390 10140 2426
rect 10260 2426 10362 2510
tri 10362 2426 10450 2514 sw
tri 10460 2426 10548 2514 ne
rect 10548 2510 10912 2514
rect 10548 2426 10690 2510
rect 10260 2390 10450 2426
rect 10086 2386 10450 2390
tri 10450 2386 10490 2426 sw
tri 10548 2386 10588 2426 ne
rect 10588 2390 10690 2426
rect 10810 2426 10912 2510
tri 10912 2426 11000 2514 sw
tri 11010 2426 11098 2514 ne
rect 11098 2510 11462 2514
rect 11098 2426 11240 2510
rect 10810 2390 11000 2426
rect 10588 2386 11000 2390
rect 10086 2338 10490 2386
rect 9586 2288 9988 2338
rect 9066 2258 9488 2288
rect 8574 2200 8968 2258
rect 8064 2160 8476 2200
tri 8476 2160 8516 2200 sw
tri 8574 2160 8614 2200 ne
rect 8614 2160 8968 2200
tri 8968 2160 9066 2258 sw
tri 9066 2160 9164 2258 ne
rect 9164 2200 9488 2258
tri 9488 2200 9576 2288 sw
tri 9586 2200 9674 2288 ne
rect 9674 2258 9988 2288
tri 9988 2258 10068 2338 sw
tri 10086 2258 10166 2338 ne
rect 10166 2288 10490 2338
tri 10490 2288 10588 2386 sw
tri 10588 2288 10686 2386 ne
rect 10686 2338 11000 2386
tri 11000 2338 11088 2426 sw
tri 11098 2338 11186 2426 ne
rect 11186 2390 11240 2426
rect 11360 2426 11462 2510
tri 11462 2426 11550 2514 sw
tri 11560 2426 11648 2514 ne
rect 11648 2510 12012 2514
rect 11648 2426 11790 2510
rect 11360 2390 11550 2426
rect 11186 2386 11550 2390
tri 11550 2386 11590 2426 sw
tri 11648 2386 11688 2426 ne
rect 11688 2390 11790 2426
rect 11910 2426 12012 2510
tri 12012 2426 12100 2514 sw
tri 12110 2426 12198 2514 ne
rect 12198 2510 12562 2514
rect 12198 2426 12340 2510
rect 11910 2390 12100 2426
rect 11688 2386 12100 2390
rect 11186 2338 11590 2386
rect 10686 2288 11088 2338
rect 10166 2258 10588 2288
rect 9674 2200 10068 2258
rect 9164 2160 9576 2200
tri 9576 2160 9616 2200 sw
tri 9674 2160 9714 2200 ne
rect 9714 2160 10068 2200
tri 10068 2160 10166 2258 sw
tri 10166 2160 10264 2258 ne
rect 10264 2200 10588 2258
tri 10588 2200 10676 2288 sw
tri 10686 2200 10774 2288 ne
rect 10774 2258 11088 2288
tri 11088 2258 11168 2338 sw
tri 11186 2258 11266 2338 ne
rect 11266 2288 11590 2338
tri 11590 2288 11688 2386 sw
tri 11688 2288 11786 2386 ne
rect 11786 2338 12100 2386
tri 12100 2338 12188 2426 sw
tri 12198 2338 12286 2426 ne
rect 12286 2390 12340 2426
rect 12460 2426 12562 2510
tri 12562 2426 12650 2514 sw
tri 12660 2426 12748 2514 ne
rect 12748 2510 13112 2514
rect 12748 2426 12890 2510
rect 12460 2390 12650 2426
rect 12286 2386 12650 2390
tri 12650 2386 12690 2426 sw
tri 12748 2386 12788 2426 ne
rect 12788 2390 12890 2426
rect 13010 2426 13112 2510
tri 13112 2426 13200 2514 sw
tri 13210 2426 13298 2514 ne
rect 13298 2510 15775 2514
rect 13298 2426 13440 2510
rect 13010 2390 13200 2426
rect 12788 2386 13200 2390
rect 12286 2338 12690 2386
rect 11786 2288 12188 2338
rect 11266 2258 11688 2288
rect 10774 2200 11168 2258
rect 10264 2160 10676 2200
tri 10676 2160 10716 2200 sw
tri 10774 2160 10814 2200 ne
rect 10814 2160 11168 2200
tri 11168 2160 11266 2258 sw
tri 11266 2160 11364 2258 ne
rect 11364 2200 11688 2258
tri 11688 2200 11776 2288 sw
tri 11786 2200 11874 2288 ne
rect 11874 2258 12188 2288
tri 12188 2258 12268 2338 sw
tri 12286 2258 12366 2338 ne
rect 12366 2288 12690 2338
tri 12690 2288 12788 2386 sw
tri 12788 2288 12886 2386 ne
rect 12886 2338 13200 2386
tri 13200 2338 13288 2426 sw
tri 13298 2338 13386 2426 ne
rect 13386 2390 13440 2426
rect 13560 2390 15775 2510
rect 13386 2338 15775 2390
rect 12886 2288 13288 2338
rect 12366 2258 12788 2288
rect 11874 2200 12268 2258
rect 11364 2160 11776 2200
tri 11776 2160 11816 2200 sw
tri 11874 2160 11914 2200 ne
rect 11914 2160 12268 2200
tri 12268 2160 12366 2258 sw
tri 12366 2160 12464 2258 ne
rect 12464 2200 12788 2258
tri 12788 2200 12876 2288 sw
tri 12886 2200 12974 2288 ne
rect 12974 2258 13288 2288
tri 13288 2258 13368 2338 sw
tri 13386 2258 13466 2338 ne
rect 13466 2258 14075 2338
rect 12974 2200 13368 2258
rect 12464 2160 12876 2200
tri 12876 2160 12916 2200 sw
tri 12974 2160 13014 2200 ne
rect 13014 2160 13368 2200
tri 13368 2160 13466 2258 sw
tri 13466 2160 13564 2258 ne
rect 13564 2238 14075 2258
rect 14175 2238 15775 2338
rect 13564 2160 15775 2238
rect -1025 2112 -284 2160
rect -1025 2012 -925 2112
rect -825 2062 -284 2112
tri -284 2062 -186 2160 sw
tri -186 2062 -88 2160 ne
rect -88 2062 266 2160
tri 266 2062 364 2160 sw
tri 364 2062 462 2160 ne
rect 462 2062 816 2160
tri 816 2062 914 2160 sw
tri 914 2062 1012 2160 ne
rect 1012 2062 1366 2160
tri 1366 2062 1464 2160 sw
tri 1464 2062 1562 2160 ne
rect 1562 2062 1916 2160
tri 1916 2062 2014 2160 sw
tri 2014 2062 2112 2160 ne
rect 2112 2062 2466 2160
tri 2466 2062 2564 2160 sw
tri 2564 2062 2662 2160 ne
rect 2662 2062 3016 2160
tri 3016 2062 3114 2160 sw
tri 3114 2062 3212 2160 ne
rect 3212 2062 3566 2160
tri 3566 2062 3664 2160 sw
tri 3664 2062 3762 2160 ne
rect 3762 2062 4116 2160
tri 4116 2062 4214 2160 sw
tri 4214 2062 4312 2160 ne
rect 4312 2062 4666 2160
tri 4666 2062 4764 2160 sw
tri 4764 2062 4862 2160 ne
rect 4862 2062 5216 2160
tri 5216 2062 5314 2160 sw
tri 5314 2062 5412 2160 ne
rect 5412 2062 5766 2160
tri 5766 2062 5864 2160 sw
tri 5864 2062 5962 2160 ne
rect 5962 2062 6316 2160
tri 6316 2062 6414 2160 sw
tri 6414 2062 6512 2160 ne
rect 6512 2062 6866 2160
tri 6866 2062 6964 2160 sw
tri 6964 2062 7062 2160 ne
rect 7062 2062 7416 2160
tri 7416 2062 7514 2160 sw
tri 7514 2062 7612 2160 ne
rect 7612 2062 7966 2160
tri 7966 2062 8064 2160 sw
tri 8064 2062 8162 2160 ne
rect 8162 2062 8516 2160
tri 8516 2062 8614 2160 sw
tri 8614 2062 8712 2160 ne
rect 8712 2062 9066 2160
tri 9066 2062 9164 2160 sw
tri 9164 2062 9262 2160 ne
rect 9262 2062 9616 2160
tri 9616 2062 9714 2160 sw
tri 9714 2062 9812 2160 ne
rect 9812 2062 10166 2160
tri 10166 2062 10264 2160 sw
tri 10264 2062 10362 2160 ne
rect 10362 2062 10716 2160
tri 10716 2062 10814 2160 sw
tri 10814 2062 10912 2160 ne
rect 10912 2062 11266 2160
tri 11266 2062 11364 2160 sw
tri 11364 2062 11462 2160 ne
rect 11462 2062 11816 2160
tri 11816 2062 11914 2160 sw
tri 11914 2062 12012 2160 ne
rect 12012 2062 12366 2160
tri 12366 2062 12464 2160 sw
tri 12464 2062 12562 2160 ne
rect 12562 2062 12916 2160
tri 12916 2062 13014 2160 sw
tri 13014 2062 13112 2160 ne
rect 13112 2062 13466 2160
tri 13466 2062 13564 2160 sw
tri 13564 2062 13662 2160 ne
rect 13662 2062 15775 2160
rect -825 2012 -186 2062
rect -1025 1964 -186 2012
tri -186 1964 -88 2062 sw
tri -88 1964 10 2062 ne
rect 10 1964 364 2062
tri 364 1964 462 2062 sw
tri 462 1964 560 2062 ne
rect 560 1964 914 2062
tri 914 1964 1012 2062 sw
tri 1012 1964 1110 2062 ne
rect 1110 1964 1464 2062
tri 1464 1964 1562 2062 sw
tri 1562 1964 1660 2062 ne
rect 1660 1964 2014 2062
tri 2014 1964 2112 2062 sw
tri 2112 1964 2210 2062 ne
rect 2210 1964 2564 2062
tri 2564 1964 2662 2062 sw
tri 2662 1964 2760 2062 ne
rect 2760 1964 3114 2062
tri 3114 1964 3212 2062 sw
tri 3212 1964 3310 2062 ne
rect 3310 1964 3664 2062
tri 3664 1964 3762 2062 sw
tri 3762 1964 3860 2062 ne
rect 3860 1964 4214 2062
tri 4214 1964 4312 2062 sw
tri 4312 1964 4410 2062 ne
rect 4410 1964 4764 2062
tri 4764 1964 4862 2062 sw
tri 4862 1964 4960 2062 ne
rect 4960 1964 5314 2062
tri 5314 1964 5412 2062 sw
tri 5412 1964 5510 2062 ne
rect 5510 1964 5864 2062
tri 5864 1964 5962 2062 sw
tri 5962 1964 6060 2062 ne
rect 6060 1964 6414 2062
tri 6414 1964 6512 2062 sw
tri 6512 1964 6610 2062 ne
rect 6610 1964 6964 2062
tri 6964 1964 7062 2062 sw
tri 7062 1964 7160 2062 ne
rect 7160 1964 7514 2062
tri 7514 1964 7612 2062 sw
tri 7612 1964 7710 2062 ne
rect 7710 1964 8064 2062
tri 8064 1964 8162 2062 sw
tri 8162 1964 8260 2062 ne
rect 8260 1964 8614 2062
tri 8614 1964 8712 2062 sw
tri 8712 1964 8810 2062 ne
rect 8810 1964 9164 2062
tri 9164 1964 9262 2062 sw
tri 9262 1964 9360 2062 ne
rect 9360 1964 9714 2062
tri 9714 1964 9812 2062 sw
tri 9812 1964 9910 2062 ne
rect 9910 1964 10264 2062
tri 10264 1964 10362 2062 sw
tri 10362 1964 10460 2062 ne
rect 10460 1964 10814 2062
tri 10814 1964 10912 2062 sw
tri 10912 1964 11010 2062 ne
rect 11010 1964 11364 2062
tri 11364 1964 11462 2062 sw
tri 11462 1964 11560 2062 ne
rect 11560 1964 11914 2062
tri 11914 1964 12012 2062 sw
tri 12012 1964 12110 2062 ne
rect 12110 1964 12464 2062
tri 12464 1964 12562 2062 sw
tri 12562 1964 12660 2062 ne
rect 12660 1964 13014 2062
tri 13014 1964 13112 2062 sw
tri 13112 1964 13210 2062 ne
rect 13210 1964 13564 2062
tri 13564 1964 13662 2062 sw
rect -1025 1960 -88 1964
rect -1025 1840 -310 1960
rect -190 1876 -88 1960
tri -88 1876 0 1964 sw
tri 10 1876 98 1964 ne
rect 98 1960 462 1964
rect 98 1876 240 1960
rect -190 1840 0 1876
rect -1025 1836 0 1840
tri 0 1836 40 1876 sw
tri 98 1836 138 1876 ne
rect 138 1840 240 1876
rect 360 1876 462 1960
tri 462 1876 550 1964 sw
tri 560 1876 648 1964 ne
rect 648 1960 1012 1964
rect 648 1876 790 1960
rect 360 1840 550 1876
rect 138 1836 550 1840
tri -412 1738 -314 1836 ne
rect -314 1738 40 1836
tri 40 1738 138 1836 sw
tri 138 1738 236 1836 ne
rect 236 1788 550 1836
tri 550 1788 638 1876 sw
tri 648 1788 736 1876 ne
rect 736 1840 790 1876
rect 910 1876 1012 1960
tri 1012 1876 1100 1964 sw
tri 1110 1876 1198 1964 ne
rect 1198 1960 1562 1964
rect 1198 1876 1340 1960
rect 910 1840 1100 1876
rect 736 1836 1100 1840
tri 1100 1836 1140 1876 sw
tri 1198 1836 1238 1876 ne
rect 1238 1840 1340 1876
rect 1460 1876 1562 1960
tri 1562 1876 1650 1964 sw
tri 1660 1876 1748 1964 ne
rect 1748 1960 2112 1964
rect 1748 1876 1890 1960
rect 1460 1840 1650 1876
rect 1238 1836 1650 1840
rect 736 1788 1140 1836
rect 236 1738 638 1788
rect -2525 1650 -412 1738
tri -412 1650 -324 1738 sw
tri -314 1650 -226 1738 ne
rect -226 1650 138 1738
tri 138 1650 226 1738 sw
tri 236 1650 324 1738 ne
rect 324 1708 638 1738
tri 638 1708 718 1788 sw
tri 736 1708 816 1788 ne
rect 816 1738 1140 1788
tri 1140 1738 1238 1836 sw
tri 1238 1738 1336 1836 ne
rect 1336 1788 1650 1836
tri 1650 1788 1738 1876 sw
tri 1748 1788 1836 1876 ne
rect 1836 1840 1890 1876
rect 2010 1876 2112 1960
tri 2112 1876 2200 1964 sw
tri 2210 1876 2298 1964 ne
rect 2298 1960 2662 1964
rect 2298 1876 2440 1960
rect 2010 1840 2200 1876
rect 1836 1836 2200 1840
tri 2200 1836 2240 1876 sw
tri 2298 1836 2338 1876 ne
rect 2338 1840 2440 1876
rect 2560 1876 2662 1960
tri 2662 1876 2750 1964 sw
tri 2760 1876 2848 1964 ne
rect 2848 1960 3212 1964
rect 2848 1876 2990 1960
rect 2560 1840 2750 1876
rect 2338 1836 2750 1840
rect 1836 1788 2240 1836
rect 1336 1738 1738 1788
rect 816 1708 1238 1738
rect 324 1650 718 1708
rect -2525 1610 -324 1650
tri -324 1610 -284 1650 sw
tri -226 1610 -186 1650 ne
rect -186 1610 226 1650
tri 226 1610 266 1650 sw
tri 324 1610 364 1650 ne
rect 364 1610 718 1650
tri 718 1610 816 1708 sw
tri 816 1610 914 1708 ne
rect 914 1650 1238 1708
tri 1238 1650 1326 1738 sw
tri 1336 1650 1424 1738 ne
rect 1424 1708 1738 1738
tri 1738 1708 1818 1788 sw
tri 1836 1708 1916 1788 ne
rect 1916 1738 2240 1788
tri 2240 1738 2338 1836 sw
tri 2338 1738 2436 1836 ne
rect 2436 1788 2750 1836
tri 2750 1788 2838 1876 sw
tri 2848 1788 2936 1876 ne
rect 2936 1840 2990 1876
rect 3110 1876 3212 1960
tri 3212 1876 3300 1964 sw
tri 3310 1876 3398 1964 ne
rect 3398 1960 3762 1964
rect 3398 1876 3540 1960
rect 3110 1840 3300 1876
rect 2936 1836 3300 1840
tri 3300 1836 3340 1876 sw
tri 3398 1836 3438 1876 ne
rect 3438 1840 3540 1876
rect 3660 1876 3762 1960
tri 3762 1876 3850 1964 sw
tri 3860 1876 3948 1964 ne
rect 3948 1960 4312 1964
rect 3948 1876 4090 1960
rect 3660 1840 3850 1876
rect 3438 1836 3850 1840
rect 2936 1788 3340 1836
rect 2436 1738 2838 1788
rect 1916 1708 2338 1738
rect 1424 1650 1818 1708
rect 914 1610 1326 1650
tri 1326 1610 1366 1650 sw
tri 1424 1610 1464 1650 ne
rect 1464 1610 1818 1650
tri 1818 1610 1916 1708 sw
tri 1916 1610 2014 1708 ne
rect 2014 1650 2338 1708
tri 2338 1650 2426 1738 sw
tri 2436 1650 2524 1738 ne
rect 2524 1708 2838 1738
tri 2838 1708 2918 1788 sw
tri 2936 1708 3016 1788 ne
rect 3016 1738 3340 1788
tri 3340 1738 3438 1836 sw
tri 3438 1738 3536 1836 ne
rect 3536 1788 3850 1836
tri 3850 1788 3938 1876 sw
tri 3948 1788 4036 1876 ne
rect 4036 1840 4090 1876
rect 4210 1876 4312 1960
tri 4312 1876 4400 1964 sw
tri 4410 1876 4498 1964 ne
rect 4498 1960 4862 1964
rect 4498 1876 4640 1960
rect 4210 1840 4400 1876
rect 4036 1836 4400 1840
tri 4400 1836 4440 1876 sw
tri 4498 1836 4538 1876 ne
rect 4538 1840 4640 1876
rect 4760 1876 4862 1960
tri 4862 1876 4950 1964 sw
tri 4960 1876 5048 1964 ne
rect 5048 1960 5412 1964
rect 5048 1876 5190 1960
rect 4760 1840 4950 1876
rect 4538 1836 4950 1840
rect 4036 1788 4440 1836
rect 3536 1738 3938 1788
rect 3016 1708 3438 1738
rect 2524 1650 2918 1708
rect 2014 1610 2426 1650
tri 2426 1610 2466 1650 sw
tri 2524 1610 2564 1650 ne
rect 2564 1610 2918 1650
tri 2918 1610 3016 1708 sw
tri 3016 1610 3114 1708 ne
rect 3114 1650 3438 1708
tri 3438 1650 3526 1738 sw
tri 3536 1650 3624 1738 ne
rect 3624 1708 3938 1738
tri 3938 1708 4018 1788 sw
tri 4036 1708 4116 1788 ne
rect 4116 1738 4440 1788
tri 4440 1738 4538 1836 sw
tri 4538 1738 4636 1836 ne
rect 4636 1788 4950 1836
tri 4950 1788 5038 1876 sw
tri 5048 1788 5136 1876 ne
rect 5136 1840 5190 1876
rect 5310 1876 5412 1960
tri 5412 1876 5500 1964 sw
tri 5510 1876 5598 1964 ne
rect 5598 1960 5962 1964
rect 5598 1876 5740 1960
rect 5310 1840 5500 1876
rect 5136 1836 5500 1840
tri 5500 1836 5540 1876 sw
tri 5598 1836 5638 1876 ne
rect 5638 1840 5740 1876
rect 5860 1876 5962 1960
tri 5962 1876 6050 1964 sw
tri 6060 1876 6148 1964 ne
rect 6148 1960 6512 1964
rect 6148 1876 6290 1960
rect 5860 1840 6050 1876
rect 5638 1836 6050 1840
rect 5136 1788 5540 1836
rect 4636 1738 5038 1788
rect 4116 1708 4538 1738
rect 3624 1650 4018 1708
rect 3114 1610 3526 1650
tri 3526 1610 3566 1650 sw
tri 3624 1610 3664 1650 ne
rect 3664 1610 4018 1650
tri 4018 1610 4116 1708 sw
tri 4116 1610 4214 1708 ne
rect 4214 1650 4538 1708
tri 4538 1650 4626 1738 sw
tri 4636 1650 4724 1738 ne
rect 4724 1708 5038 1738
tri 5038 1708 5118 1788 sw
tri 5136 1708 5216 1788 ne
rect 5216 1738 5540 1788
tri 5540 1738 5638 1836 sw
tri 5638 1738 5736 1836 ne
rect 5736 1788 6050 1836
tri 6050 1788 6138 1876 sw
tri 6148 1788 6236 1876 ne
rect 6236 1840 6290 1876
rect 6410 1876 6512 1960
tri 6512 1876 6600 1964 sw
tri 6610 1876 6698 1964 ne
rect 6698 1960 7062 1964
rect 6698 1876 6840 1960
rect 6410 1840 6600 1876
rect 6236 1836 6600 1840
tri 6600 1836 6640 1876 sw
tri 6698 1836 6738 1876 ne
rect 6738 1840 6840 1876
rect 6960 1876 7062 1960
tri 7062 1876 7150 1964 sw
tri 7160 1876 7248 1964 ne
rect 7248 1960 7612 1964
rect 7248 1876 7390 1960
rect 6960 1840 7150 1876
rect 6738 1836 7150 1840
rect 6236 1788 6640 1836
rect 5736 1738 6138 1788
rect 5216 1708 5638 1738
rect 4724 1650 5118 1708
rect 4214 1610 4626 1650
tri 4626 1610 4666 1650 sw
tri 4724 1610 4764 1650 ne
rect 4764 1610 5118 1650
tri 5118 1610 5216 1708 sw
tri 5216 1610 5314 1708 ne
rect 5314 1650 5638 1708
tri 5638 1650 5726 1738 sw
tri 5736 1650 5824 1738 ne
rect 5824 1708 6138 1738
tri 6138 1708 6218 1788 sw
tri 6236 1708 6316 1788 ne
rect 6316 1738 6640 1788
tri 6640 1738 6738 1836 sw
tri 6738 1738 6836 1836 ne
rect 6836 1788 7150 1836
tri 7150 1788 7238 1876 sw
tri 7248 1788 7336 1876 ne
rect 7336 1840 7390 1876
rect 7510 1876 7612 1960
tri 7612 1876 7700 1964 sw
tri 7710 1876 7798 1964 ne
rect 7798 1960 8162 1964
rect 7798 1876 7940 1960
rect 7510 1840 7700 1876
rect 7336 1836 7700 1840
tri 7700 1836 7740 1876 sw
tri 7798 1836 7838 1876 ne
rect 7838 1840 7940 1876
rect 8060 1876 8162 1960
tri 8162 1876 8250 1964 sw
tri 8260 1876 8348 1964 ne
rect 8348 1960 8712 1964
rect 8348 1876 8490 1960
rect 8060 1840 8250 1876
rect 7838 1836 8250 1840
rect 7336 1788 7740 1836
rect 6836 1738 7238 1788
rect 6316 1708 6738 1738
rect 5824 1650 6218 1708
rect 5314 1610 5726 1650
tri 5726 1610 5766 1650 sw
tri 5824 1610 5864 1650 ne
rect 5864 1610 6218 1650
tri 6218 1610 6316 1708 sw
tri 6316 1610 6414 1708 ne
rect 6414 1650 6738 1708
tri 6738 1650 6826 1738 sw
tri 6836 1650 6924 1738 ne
rect 6924 1708 7238 1738
tri 7238 1708 7318 1788 sw
tri 7336 1708 7416 1788 ne
rect 7416 1738 7740 1788
tri 7740 1738 7838 1836 sw
tri 7838 1738 7936 1836 ne
rect 7936 1788 8250 1836
tri 8250 1788 8338 1876 sw
tri 8348 1788 8436 1876 ne
rect 8436 1840 8490 1876
rect 8610 1876 8712 1960
tri 8712 1876 8800 1964 sw
tri 8810 1876 8898 1964 ne
rect 8898 1960 9262 1964
rect 8898 1876 9040 1960
rect 8610 1840 8800 1876
rect 8436 1836 8800 1840
tri 8800 1836 8840 1876 sw
tri 8898 1836 8938 1876 ne
rect 8938 1840 9040 1876
rect 9160 1876 9262 1960
tri 9262 1876 9350 1964 sw
tri 9360 1876 9448 1964 ne
rect 9448 1960 9812 1964
rect 9448 1876 9590 1960
rect 9160 1840 9350 1876
rect 8938 1836 9350 1840
rect 8436 1788 8840 1836
rect 7936 1738 8338 1788
rect 7416 1708 7838 1738
rect 6924 1650 7318 1708
rect 6414 1610 6826 1650
tri 6826 1610 6866 1650 sw
tri 6924 1610 6964 1650 ne
rect 6964 1610 7318 1650
tri 7318 1610 7416 1708 sw
tri 7416 1610 7514 1708 ne
rect 7514 1650 7838 1708
tri 7838 1650 7926 1738 sw
tri 7936 1650 8024 1738 ne
rect 8024 1708 8338 1738
tri 8338 1708 8418 1788 sw
tri 8436 1708 8516 1788 ne
rect 8516 1738 8840 1788
tri 8840 1738 8938 1836 sw
tri 8938 1738 9036 1836 ne
rect 9036 1788 9350 1836
tri 9350 1788 9438 1876 sw
tri 9448 1788 9536 1876 ne
rect 9536 1840 9590 1876
rect 9710 1876 9812 1960
tri 9812 1876 9900 1964 sw
tri 9910 1876 9998 1964 ne
rect 9998 1960 10362 1964
rect 9998 1876 10140 1960
rect 9710 1840 9900 1876
rect 9536 1836 9900 1840
tri 9900 1836 9940 1876 sw
tri 9998 1836 10038 1876 ne
rect 10038 1840 10140 1876
rect 10260 1876 10362 1960
tri 10362 1876 10450 1964 sw
tri 10460 1876 10548 1964 ne
rect 10548 1960 10912 1964
rect 10548 1876 10690 1960
rect 10260 1840 10450 1876
rect 10038 1836 10450 1840
rect 9536 1788 9940 1836
rect 9036 1738 9438 1788
rect 8516 1708 8938 1738
rect 8024 1650 8418 1708
rect 7514 1610 7926 1650
tri 7926 1610 7966 1650 sw
tri 8024 1610 8064 1650 ne
rect 8064 1610 8418 1650
tri 8418 1610 8516 1708 sw
tri 8516 1610 8614 1708 ne
rect 8614 1650 8938 1708
tri 8938 1650 9026 1738 sw
tri 9036 1650 9124 1738 ne
rect 9124 1708 9438 1738
tri 9438 1708 9518 1788 sw
tri 9536 1708 9616 1788 ne
rect 9616 1738 9940 1788
tri 9940 1738 10038 1836 sw
tri 10038 1738 10136 1836 ne
rect 10136 1788 10450 1836
tri 10450 1788 10538 1876 sw
tri 10548 1788 10636 1876 ne
rect 10636 1840 10690 1876
rect 10810 1876 10912 1960
tri 10912 1876 11000 1964 sw
tri 11010 1876 11098 1964 ne
rect 11098 1960 11462 1964
rect 11098 1876 11240 1960
rect 10810 1840 11000 1876
rect 10636 1836 11000 1840
tri 11000 1836 11040 1876 sw
tri 11098 1836 11138 1876 ne
rect 11138 1840 11240 1876
rect 11360 1876 11462 1960
tri 11462 1876 11550 1964 sw
tri 11560 1876 11648 1964 ne
rect 11648 1960 12012 1964
rect 11648 1876 11790 1960
rect 11360 1840 11550 1876
rect 11138 1836 11550 1840
rect 10636 1788 11040 1836
rect 10136 1738 10538 1788
rect 9616 1708 10038 1738
rect 9124 1650 9518 1708
rect 8614 1610 9026 1650
tri 9026 1610 9066 1650 sw
tri 9124 1610 9164 1650 ne
rect 9164 1610 9518 1650
tri 9518 1610 9616 1708 sw
tri 9616 1610 9714 1708 ne
rect 9714 1650 10038 1708
tri 10038 1650 10126 1738 sw
tri 10136 1650 10224 1738 ne
rect 10224 1708 10538 1738
tri 10538 1708 10618 1788 sw
tri 10636 1708 10716 1788 ne
rect 10716 1738 11040 1788
tri 11040 1738 11138 1836 sw
tri 11138 1738 11236 1836 ne
rect 11236 1788 11550 1836
tri 11550 1788 11638 1876 sw
tri 11648 1788 11736 1876 ne
rect 11736 1840 11790 1876
rect 11910 1876 12012 1960
tri 12012 1876 12100 1964 sw
tri 12110 1876 12198 1964 ne
rect 12198 1960 12562 1964
rect 12198 1876 12340 1960
rect 11910 1840 12100 1876
rect 11736 1836 12100 1840
tri 12100 1836 12140 1876 sw
tri 12198 1836 12238 1876 ne
rect 12238 1840 12340 1876
rect 12460 1876 12562 1960
tri 12562 1876 12650 1964 sw
tri 12660 1876 12748 1964 ne
rect 12748 1960 13112 1964
rect 12748 1876 12890 1960
rect 12460 1840 12650 1876
rect 12238 1836 12650 1840
rect 11736 1788 12140 1836
rect 11236 1738 11638 1788
rect 10716 1708 11138 1738
rect 10224 1650 10618 1708
rect 9714 1610 10126 1650
tri 10126 1610 10166 1650 sw
tri 10224 1610 10264 1650 ne
rect 10264 1610 10618 1650
tri 10618 1610 10716 1708 sw
tri 10716 1610 10814 1708 ne
rect 10814 1650 11138 1708
tri 11138 1650 11226 1738 sw
tri 11236 1650 11324 1738 ne
rect 11324 1708 11638 1738
tri 11638 1708 11718 1788 sw
tri 11736 1708 11816 1788 ne
rect 11816 1738 12140 1788
tri 12140 1738 12238 1836 sw
tri 12238 1738 12336 1836 ne
rect 12336 1788 12650 1836
tri 12650 1788 12738 1876 sw
tri 12748 1788 12836 1876 ne
rect 12836 1840 12890 1876
rect 13010 1876 13112 1960
tri 13112 1876 13200 1964 sw
tri 13210 1876 13298 1964 ne
rect 13298 1960 14275 1964
rect 13298 1876 13440 1960
rect 13010 1840 13200 1876
rect 12836 1836 13200 1840
tri 13200 1836 13240 1876 sw
tri 13298 1836 13338 1876 ne
rect 13338 1840 13440 1876
rect 13560 1840 14275 1960
rect 13338 1836 14275 1840
rect 12836 1788 13240 1836
rect 12336 1738 12738 1788
rect 11816 1708 12238 1738
rect 11324 1650 11718 1708
rect 10814 1610 11226 1650
tri 11226 1610 11266 1650 sw
tri 11324 1610 11364 1650 ne
rect 11364 1610 11718 1650
tri 11718 1610 11816 1708 sw
tri 11816 1610 11914 1708 ne
rect 11914 1650 12238 1708
tri 12238 1650 12326 1738 sw
tri 12336 1650 12424 1738 ne
rect 12424 1708 12738 1738
tri 12738 1708 12818 1788 sw
tri 12836 1708 12916 1788 ne
rect 12916 1738 13240 1788
tri 13240 1738 13338 1836 sw
tri 13338 1738 13436 1836 ne
rect 13436 1738 14275 1836
rect 12916 1708 13338 1738
rect 12424 1650 12818 1708
rect 11914 1610 12326 1650
tri 12326 1610 12366 1650 sw
tri 12424 1610 12464 1650 ne
rect 12464 1610 12818 1650
tri 12818 1610 12916 1708 sw
tri 12916 1610 13014 1708 ne
rect 13014 1650 13338 1708
tri 13338 1650 13426 1738 sw
tri 13436 1650 13524 1738 ne
rect 13524 1650 14275 1738
rect 13014 1610 13426 1650
tri 13426 1610 13466 1650 sw
tri 13524 1610 13564 1650 ne
rect 13564 1610 14275 1650
rect -2525 1512 -284 1610
tri -284 1512 -186 1610 sw
tri -186 1512 -88 1610 ne
rect -88 1512 266 1610
tri 266 1512 364 1610 sw
tri 364 1512 462 1610 ne
rect 462 1512 816 1610
tri 816 1512 914 1610 sw
tri 914 1512 1012 1610 ne
rect 1012 1512 1366 1610
tri 1366 1512 1464 1610 sw
tri 1464 1512 1562 1610 ne
rect 1562 1512 1916 1610
tri 1916 1512 2014 1610 sw
tri 2014 1512 2112 1610 ne
rect 2112 1512 2466 1610
tri 2466 1512 2564 1610 sw
tri 2564 1512 2662 1610 ne
rect 2662 1512 3016 1610
tri 3016 1512 3114 1610 sw
tri 3114 1512 3212 1610 ne
rect 3212 1512 3566 1610
tri 3566 1512 3664 1610 sw
tri 3664 1512 3762 1610 ne
rect 3762 1512 4116 1610
tri 4116 1512 4214 1610 sw
tri 4214 1512 4312 1610 ne
rect 4312 1512 4666 1610
tri 4666 1512 4764 1610 sw
tri 4764 1512 4862 1610 ne
rect 4862 1512 5216 1610
tri 5216 1512 5314 1610 sw
tri 5314 1512 5412 1610 ne
rect 5412 1512 5766 1610
tri 5766 1512 5864 1610 sw
tri 5864 1512 5962 1610 ne
rect 5962 1512 6316 1610
tri 6316 1512 6414 1610 sw
tri 6414 1512 6512 1610 ne
rect 6512 1512 6866 1610
tri 6866 1512 6964 1610 sw
tri 6964 1512 7062 1610 ne
rect 7062 1512 7416 1610
tri 7416 1512 7514 1610 sw
tri 7514 1512 7612 1610 ne
rect 7612 1512 7966 1610
tri 7966 1512 8064 1610 sw
tri 8064 1512 8162 1610 ne
rect 8162 1512 8516 1610
tri 8516 1512 8614 1610 sw
tri 8614 1512 8712 1610 ne
rect 8712 1512 9066 1610
tri 9066 1512 9164 1610 sw
tri 9164 1512 9262 1610 ne
rect 9262 1512 9616 1610
tri 9616 1512 9714 1610 sw
tri 9714 1512 9812 1610 ne
rect 9812 1512 10166 1610
tri 10166 1512 10264 1610 sw
tri 10264 1512 10362 1610 ne
rect 10362 1512 10716 1610
tri 10716 1512 10814 1610 sw
tri 10814 1512 10912 1610 ne
rect 10912 1512 11266 1610
tri 11266 1512 11364 1610 sw
tri 11364 1512 11462 1610 ne
rect 11462 1512 11816 1610
tri 11816 1512 11914 1610 sw
tri 11914 1512 12012 1610 ne
rect 12012 1512 12366 1610
tri 12366 1512 12464 1610 sw
tri 12464 1512 12562 1610 ne
rect 12562 1512 12916 1610
tri 12916 1512 13014 1610 sw
tri 13014 1512 13112 1610 ne
rect 13112 1512 13466 1610
tri 13466 1512 13564 1610 sw
tri 13564 1512 13662 1610 ne
rect 13662 1512 14275 1610
rect -2525 1414 -186 1512
tri -186 1414 -88 1512 sw
tri -88 1414 10 1512 ne
rect 10 1414 364 1512
tri 364 1414 462 1512 sw
tri 462 1414 560 1512 ne
rect 560 1414 914 1512
tri 914 1414 1012 1512 sw
tri 1012 1414 1110 1512 ne
rect 1110 1414 1464 1512
tri 1464 1414 1562 1512 sw
tri 1562 1414 1660 1512 ne
rect 1660 1414 2014 1512
tri 2014 1414 2112 1512 sw
tri 2112 1414 2210 1512 ne
rect 2210 1414 2564 1512
tri 2564 1414 2662 1512 sw
tri 2662 1414 2760 1512 ne
rect 2760 1414 3114 1512
tri 3114 1414 3212 1512 sw
tri 3212 1414 3310 1512 ne
rect 3310 1414 3664 1512
tri 3664 1414 3762 1512 sw
tri 3762 1414 3860 1512 ne
rect 3860 1414 4214 1512
tri 4214 1414 4312 1512 sw
tri 4312 1414 4410 1512 ne
rect 4410 1414 4764 1512
tri 4764 1414 4862 1512 sw
tri 4862 1414 4960 1512 ne
rect 4960 1414 5314 1512
tri 5314 1414 5412 1512 sw
tri 5412 1414 5510 1512 ne
rect 5510 1414 5864 1512
tri 5864 1414 5962 1512 sw
tri 5962 1414 6060 1512 ne
rect 6060 1414 6414 1512
tri 6414 1414 6512 1512 sw
tri 6512 1414 6610 1512 ne
rect 6610 1414 6964 1512
tri 6964 1414 7062 1512 sw
tri 7062 1414 7160 1512 ne
rect 7160 1414 7514 1512
tri 7514 1414 7612 1512 sw
tri 7612 1414 7710 1512 ne
rect 7710 1414 8064 1512
tri 8064 1414 8162 1512 sw
tri 8162 1414 8260 1512 ne
rect 8260 1414 8614 1512
tri 8614 1414 8712 1512 sw
tri 8712 1414 8810 1512 ne
rect 8810 1414 9164 1512
tri 9164 1414 9262 1512 sw
tri 9262 1414 9360 1512 ne
rect 9360 1414 9714 1512
tri 9714 1414 9812 1512 sw
tri 9812 1414 9910 1512 ne
rect 9910 1414 10264 1512
tri 10264 1414 10362 1512 sw
tri 10362 1414 10460 1512 ne
rect 10460 1414 10814 1512
tri 10814 1414 10912 1512 sw
tri 10912 1414 11010 1512 ne
rect 11010 1414 11364 1512
tri 11364 1414 11462 1512 sw
tri 11462 1414 11560 1512 ne
rect 11560 1414 11914 1512
tri 11914 1414 12012 1512 sw
tri 12012 1414 12110 1512 ne
rect 12110 1414 12464 1512
tri 12464 1414 12562 1512 sw
tri 12562 1414 12660 1512 ne
rect 12660 1414 13014 1512
tri 13014 1414 13112 1512 sw
tri 13112 1414 13210 1512 ne
rect 13210 1414 13564 1512
tri 13564 1414 13662 1512 sw
rect 14775 1414 15775 2062
rect -2525 1410 -88 1414
rect -2525 1290 -310 1410
rect -190 1326 -88 1410
tri -88 1326 0 1414 sw
tri 10 1326 98 1414 ne
rect 98 1410 462 1414
rect 98 1326 240 1410
rect -190 1290 0 1326
rect -2525 1286 0 1290
rect -2525 638 -1525 1286
tri -412 1188 -314 1286 ne
rect -314 1238 0 1286
tri 0 1238 88 1326 sw
tri 98 1238 186 1326 ne
rect 186 1290 240 1326
rect 360 1326 462 1410
tri 462 1326 550 1414 sw
tri 560 1326 648 1414 ne
rect 648 1410 1012 1414
rect 648 1326 790 1410
rect 360 1290 550 1326
rect 186 1286 550 1290
tri 550 1286 590 1326 sw
tri 648 1286 688 1326 ne
rect 688 1290 790 1326
rect 910 1326 1012 1410
tri 1012 1326 1100 1414 sw
tri 1110 1326 1198 1414 ne
rect 1198 1410 1562 1414
rect 1198 1326 1340 1410
rect 910 1290 1100 1326
rect 688 1286 1100 1290
rect 186 1238 590 1286
rect -314 1188 88 1238
rect -1025 1100 -412 1188
tri -412 1100 -324 1188 sw
tri -314 1100 -226 1188 ne
rect -226 1158 88 1188
tri 88 1158 168 1238 sw
tri 186 1158 266 1238 ne
rect 266 1188 590 1238
tri 590 1188 688 1286 sw
tri 688 1188 786 1286 ne
rect 786 1238 1100 1286
tri 1100 1238 1188 1326 sw
tri 1198 1238 1286 1326 ne
rect 1286 1290 1340 1326
rect 1460 1326 1562 1410
tri 1562 1326 1650 1414 sw
tri 1660 1326 1748 1414 ne
rect 1748 1410 2112 1414
rect 1748 1326 1890 1410
rect 1460 1290 1650 1326
rect 1286 1286 1650 1290
tri 1650 1286 1690 1326 sw
tri 1748 1286 1788 1326 ne
rect 1788 1290 1890 1326
rect 2010 1326 2112 1410
tri 2112 1326 2200 1414 sw
tri 2210 1326 2298 1414 ne
rect 2298 1410 2662 1414
rect 2298 1326 2440 1410
rect 2010 1290 2200 1326
rect 1788 1286 2200 1290
rect 1286 1238 1690 1286
rect 786 1188 1188 1238
rect 266 1158 688 1188
rect -226 1100 168 1158
rect -1025 1060 -324 1100
tri -324 1060 -284 1100 sw
tri -226 1060 -186 1100 ne
rect -186 1060 168 1100
tri 168 1060 266 1158 sw
tri 266 1060 364 1158 ne
rect 364 1100 688 1158
tri 688 1100 776 1188 sw
tri 786 1100 874 1188 ne
rect 874 1158 1188 1188
tri 1188 1158 1268 1238 sw
tri 1286 1158 1366 1238 ne
rect 1366 1188 1690 1238
tri 1690 1188 1788 1286 sw
tri 1788 1188 1886 1286 ne
rect 1886 1238 2200 1286
tri 2200 1238 2288 1326 sw
tri 2298 1238 2386 1326 ne
rect 2386 1290 2440 1326
rect 2560 1326 2662 1410
tri 2662 1326 2750 1414 sw
tri 2760 1326 2848 1414 ne
rect 2848 1410 3212 1414
rect 2848 1326 2990 1410
rect 2560 1290 2750 1326
rect 2386 1286 2750 1290
tri 2750 1286 2790 1326 sw
tri 2848 1286 2888 1326 ne
rect 2888 1290 2990 1326
rect 3110 1326 3212 1410
tri 3212 1326 3300 1414 sw
tri 3310 1326 3398 1414 ne
rect 3398 1410 3762 1414
rect 3398 1326 3540 1410
rect 3110 1290 3300 1326
rect 2888 1286 3300 1290
rect 2386 1238 2790 1286
rect 1886 1188 2288 1238
rect 1366 1158 1788 1188
rect 874 1100 1268 1158
rect 364 1060 776 1100
tri 776 1060 816 1100 sw
tri 874 1060 914 1100 ne
rect 914 1060 1268 1100
tri 1268 1060 1366 1158 sw
tri 1366 1060 1464 1158 ne
rect 1464 1100 1788 1158
tri 1788 1100 1876 1188 sw
tri 1886 1100 1974 1188 ne
rect 1974 1158 2288 1188
tri 2288 1158 2368 1238 sw
tri 2386 1158 2466 1238 ne
rect 2466 1188 2790 1238
tri 2790 1188 2888 1286 sw
tri 2888 1188 2986 1286 ne
rect 2986 1238 3300 1286
tri 3300 1238 3388 1326 sw
tri 3398 1238 3486 1326 ne
rect 3486 1290 3540 1326
rect 3660 1326 3762 1410
tri 3762 1326 3850 1414 sw
tri 3860 1326 3948 1414 ne
rect 3948 1410 4312 1414
rect 3948 1326 4090 1410
rect 3660 1290 3850 1326
rect 3486 1286 3850 1290
tri 3850 1286 3890 1326 sw
tri 3948 1286 3988 1326 ne
rect 3988 1290 4090 1326
rect 4210 1326 4312 1410
tri 4312 1326 4400 1414 sw
tri 4410 1326 4498 1414 ne
rect 4498 1410 4862 1414
rect 4498 1326 4640 1410
rect 4210 1290 4400 1326
rect 3988 1286 4400 1290
rect 3486 1238 3890 1286
rect 2986 1188 3388 1238
rect 2466 1158 2888 1188
rect 1974 1100 2368 1158
rect 1464 1060 1876 1100
tri 1876 1060 1916 1100 sw
tri 1974 1060 2014 1100 ne
rect 2014 1060 2368 1100
tri 2368 1060 2466 1158 sw
tri 2466 1060 2564 1158 ne
rect 2564 1100 2888 1158
tri 2888 1100 2976 1188 sw
tri 2986 1100 3074 1188 ne
rect 3074 1158 3388 1188
tri 3388 1158 3468 1238 sw
tri 3486 1158 3566 1238 ne
rect 3566 1188 3890 1238
tri 3890 1188 3988 1286 sw
tri 3988 1188 4086 1286 ne
rect 4086 1238 4400 1286
tri 4400 1238 4488 1326 sw
tri 4498 1238 4586 1326 ne
rect 4586 1290 4640 1326
rect 4760 1326 4862 1410
tri 4862 1326 4950 1414 sw
tri 4960 1326 5048 1414 ne
rect 5048 1410 5412 1414
rect 5048 1326 5190 1410
rect 4760 1290 4950 1326
rect 4586 1286 4950 1290
tri 4950 1286 4990 1326 sw
tri 5048 1286 5088 1326 ne
rect 5088 1290 5190 1326
rect 5310 1326 5412 1410
tri 5412 1326 5500 1414 sw
tri 5510 1326 5598 1414 ne
rect 5598 1410 5962 1414
rect 5598 1326 5740 1410
rect 5310 1290 5500 1326
rect 5088 1286 5500 1290
rect 4586 1238 4990 1286
rect 4086 1188 4488 1238
rect 3566 1158 3988 1188
rect 3074 1100 3468 1158
rect 2564 1060 2976 1100
tri 2976 1060 3016 1100 sw
tri 3074 1060 3114 1100 ne
rect 3114 1060 3468 1100
tri 3468 1060 3566 1158 sw
tri 3566 1060 3664 1158 ne
rect 3664 1100 3988 1158
tri 3988 1100 4076 1188 sw
tri 4086 1100 4174 1188 ne
rect 4174 1158 4488 1188
tri 4488 1158 4568 1238 sw
tri 4586 1158 4666 1238 ne
rect 4666 1188 4990 1238
tri 4990 1188 5088 1286 sw
tri 5088 1188 5186 1286 ne
rect 5186 1238 5500 1286
tri 5500 1238 5588 1326 sw
tri 5598 1238 5686 1326 ne
rect 5686 1290 5740 1326
rect 5860 1326 5962 1410
tri 5962 1326 6050 1414 sw
tri 6060 1326 6148 1414 ne
rect 6148 1410 6512 1414
rect 6148 1326 6290 1410
rect 5860 1290 6050 1326
rect 5686 1286 6050 1290
tri 6050 1286 6090 1326 sw
tri 6148 1286 6188 1326 ne
rect 6188 1290 6290 1326
rect 6410 1326 6512 1410
tri 6512 1326 6600 1414 sw
tri 6610 1326 6698 1414 ne
rect 6698 1410 7062 1414
rect 6698 1326 6840 1410
rect 6410 1290 6600 1326
rect 6188 1286 6600 1290
rect 5686 1238 6090 1286
rect 5186 1188 5588 1238
rect 4666 1158 5088 1188
rect 4174 1100 4568 1158
rect 3664 1060 4076 1100
tri 4076 1060 4116 1100 sw
tri 4174 1060 4214 1100 ne
rect 4214 1060 4568 1100
tri 4568 1060 4666 1158 sw
tri 4666 1060 4764 1158 ne
rect 4764 1100 5088 1158
tri 5088 1100 5176 1188 sw
tri 5186 1100 5274 1188 ne
rect 5274 1158 5588 1188
tri 5588 1158 5668 1238 sw
tri 5686 1158 5766 1238 ne
rect 5766 1188 6090 1238
tri 6090 1188 6188 1286 sw
tri 6188 1188 6286 1286 ne
rect 6286 1238 6600 1286
tri 6600 1238 6688 1326 sw
tri 6698 1238 6786 1326 ne
rect 6786 1290 6840 1326
rect 6960 1326 7062 1410
tri 7062 1326 7150 1414 sw
tri 7160 1326 7248 1414 ne
rect 7248 1410 7612 1414
rect 7248 1326 7390 1410
rect 6960 1290 7150 1326
rect 6786 1286 7150 1290
tri 7150 1286 7190 1326 sw
tri 7248 1286 7288 1326 ne
rect 7288 1290 7390 1326
rect 7510 1326 7612 1410
tri 7612 1326 7700 1414 sw
tri 7710 1326 7798 1414 ne
rect 7798 1410 8162 1414
rect 7798 1326 7940 1410
rect 7510 1290 7700 1326
rect 7288 1286 7700 1290
rect 6786 1238 7190 1286
rect 6286 1188 6688 1238
rect 5766 1158 6188 1188
rect 5274 1100 5668 1158
rect 4764 1060 5176 1100
tri 5176 1060 5216 1100 sw
tri 5274 1060 5314 1100 ne
rect 5314 1060 5668 1100
tri 5668 1060 5766 1158 sw
tri 5766 1060 5864 1158 ne
rect 5864 1100 6188 1158
tri 6188 1100 6276 1188 sw
tri 6286 1100 6374 1188 ne
rect 6374 1158 6688 1188
tri 6688 1158 6768 1238 sw
tri 6786 1158 6866 1238 ne
rect 6866 1188 7190 1238
tri 7190 1188 7288 1286 sw
tri 7288 1188 7386 1286 ne
rect 7386 1238 7700 1286
tri 7700 1238 7788 1326 sw
tri 7798 1238 7886 1326 ne
rect 7886 1290 7940 1326
rect 8060 1326 8162 1410
tri 8162 1326 8250 1414 sw
tri 8260 1326 8348 1414 ne
rect 8348 1410 8712 1414
rect 8348 1326 8490 1410
rect 8060 1290 8250 1326
rect 7886 1286 8250 1290
tri 8250 1286 8290 1326 sw
tri 8348 1286 8388 1326 ne
rect 8388 1290 8490 1326
rect 8610 1326 8712 1410
tri 8712 1326 8800 1414 sw
tri 8810 1326 8898 1414 ne
rect 8898 1410 9262 1414
rect 8898 1326 9040 1410
rect 8610 1290 8800 1326
rect 8388 1286 8800 1290
rect 7886 1238 8290 1286
rect 7386 1188 7788 1238
rect 6866 1158 7288 1188
rect 6374 1100 6768 1158
rect 5864 1060 6276 1100
tri 6276 1060 6316 1100 sw
tri 6374 1060 6414 1100 ne
rect 6414 1060 6768 1100
tri 6768 1060 6866 1158 sw
tri 6866 1060 6964 1158 ne
rect 6964 1100 7288 1158
tri 7288 1100 7376 1188 sw
tri 7386 1100 7474 1188 ne
rect 7474 1158 7788 1188
tri 7788 1158 7868 1238 sw
tri 7886 1158 7966 1238 ne
rect 7966 1188 8290 1238
tri 8290 1188 8388 1286 sw
tri 8388 1188 8486 1286 ne
rect 8486 1238 8800 1286
tri 8800 1238 8888 1326 sw
tri 8898 1238 8986 1326 ne
rect 8986 1290 9040 1326
rect 9160 1326 9262 1410
tri 9262 1326 9350 1414 sw
tri 9360 1326 9448 1414 ne
rect 9448 1410 9812 1414
rect 9448 1326 9590 1410
rect 9160 1290 9350 1326
rect 8986 1286 9350 1290
tri 9350 1286 9390 1326 sw
tri 9448 1286 9488 1326 ne
rect 9488 1290 9590 1326
rect 9710 1326 9812 1410
tri 9812 1326 9900 1414 sw
tri 9910 1326 9998 1414 ne
rect 9998 1410 10362 1414
rect 9998 1326 10140 1410
rect 9710 1290 9900 1326
rect 9488 1286 9900 1290
rect 8986 1238 9390 1286
rect 8486 1188 8888 1238
rect 7966 1158 8388 1188
rect 7474 1100 7868 1158
rect 6964 1060 7376 1100
tri 7376 1060 7416 1100 sw
tri 7474 1060 7514 1100 ne
rect 7514 1060 7868 1100
tri 7868 1060 7966 1158 sw
tri 7966 1060 8064 1158 ne
rect 8064 1100 8388 1158
tri 8388 1100 8476 1188 sw
tri 8486 1100 8574 1188 ne
rect 8574 1158 8888 1188
tri 8888 1158 8968 1238 sw
tri 8986 1158 9066 1238 ne
rect 9066 1188 9390 1238
tri 9390 1188 9488 1286 sw
tri 9488 1188 9586 1286 ne
rect 9586 1238 9900 1286
tri 9900 1238 9988 1326 sw
tri 9998 1238 10086 1326 ne
rect 10086 1290 10140 1326
rect 10260 1326 10362 1410
tri 10362 1326 10450 1414 sw
tri 10460 1326 10548 1414 ne
rect 10548 1410 10912 1414
rect 10548 1326 10690 1410
rect 10260 1290 10450 1326
rect 10086 1286 10450 1290
tri 10450 1286 10490 1326 sw
tri 10548 1286 10588 1326 ne
rect 10588 1290 10690 1326
rect 10810 1326 10912 1410
tri 10912 1326 11000 1414 sw
tri 11010 1326 11098 1414 ne
rect 11098 1410 11462 1414
rect 11098 1326 11240 1410
rect 10810 1290 11000 1326
rect 10588 1286 11000 1290
rect 10086 1238 10490 1286
rect 9586 1188 9988 1238
rect 9066 1158 9488 1188
rect 8574 1100 8968 1158
rect 8064 1060 8476 1100
tri 8476 1060 8516 1100 sw
tri 8574 1060 8614 1100 ne
rect 8614 1060 8968 1100
tri 8968 1060 9066 1158 sw
tri 9066 1060 9164 1158 ne
rect 9164 1100 9488 1158
tri 9488 1100 9576 1188 sw
tri 9586 1100 9674 1188 ne
rect 9674 1158 9988 1188
tri 9988 1158 10068 1238 sw
tri 10086 1158 10166 1238 ne
rect 10166 1188 10490 1238
tri 10490 1188 10588 1286 sw
tri 10588 1188 10686 1286 ne
rect 10686 1238 11000 1286
tri 11000 1238 11088 1326 sw
tri 11098 1238 11186 1326 ne
rect 11186 1290 11240 1326
rect 11360 1326 11462 1410
tri 11462 1326 11550 1414 sw
tri 11560 1326 11648 1414 ne
rect 11648 1410 12012 1414
rect 11648 1326 11790 1410
rect 11360 1290 11550 1326
rect 11186 1286 11550 1290
tri 11550 1286 11590 1326 sw
tri 11648 1286 11688 1326 ne
rect 11688 1290 11790 1326
rect 11910 1326 12012 1410
tri 12012 1326 12100 1414 sw
tri 12110 1326 12198 1414 ne
rect 12198 1410 12562 1414
rect 12198 1326 12340 1410
rect 11910 1290 12100 1326
rect 11688 1286 12100 1290
rect 11186 1238 11590 1286
rect 10686 1188 11088 1238
rect 10166 1158 10588 1188
rect 9674 1100 10068 1158
rect 9164 1060 9576 1100
tri 9576 1060 9616 1100 sw
tri 9674 1060 9714 1100 ne
rect 9714 1060 10068 1100
tri 10068 1060 10166 1158 sw
tri 10166 1060 10264 1158 ne
rect 10264 1100 10588 1158
tri 10588 1100 10676 1188 sw
tri 10686 1100 10774 1188 ne
rect 10774 1158 11088 1188
tri 11088 1158 11168 1238 sw
tri 11186 1158 11266 1238 ne
rect 11266 1188 11590 1238
tri 11590 1188 11688 1286 sw
tri 11688 1188 11786 1286 ne
rect 11786 1238 12100 1286
tri 12100 1238 12188 1326 sw
tri 12198 1238 12286 1326 ne
rect 12286 1290 12340 1326
rect 12460 1326 12562 1410
tri 12562 1326 12650 1414 sw
tri 12660 1326 12748 1414 ne
rect 12748 1410 13112 1414
rect 12748 1326 12890 1410
rect 12460 1290 12650 1326
rect 12286 1286 12650 1290
tri 12650 1286 12690 1326 sw
tri 12748 1286 12788 1326 ne
rect 12788 1290 12890 1326
rect 13010 1326 13112 1410
tri 13112 1326 13200 1414 sw
tri 13210 1326 13298 1414 ne
rect 13298 1410 15775 1414
rect 13298 1326 13440 1410
rect 13010 1290 13200 1326
rect 12788 1286 13200 1290
rect 12286 1238 12690 1286
rect 11786 1188 12188 1238
rect 11266 1158 11688 1188
rect 10774 1100 11168 1158
rect 10264 1060 10676 1100
tri 10676 1060 10716 1100 sw
tri 10774 1060 10814 1100 ne
rect 10814 1060 11168 1100
tri 11168 1060 11266 1158 sw
tri 11266 1060 11364 1158 ne
rect 11364 1100 11688 1158
tri 11688 1100 11776 1188 sw
tri 11786 1100 11874 1188 ne
rect 11874 1158 12188 1188
tri 12188 1158 12268 1238 sw
tri 12286 1158 12366 1238 ne
rect 12366 1188 12690 1238
tri 12690 1188 12788 1286 sw
tri 12788 1188 12886 1286 ne
rect 12886 1238 13200 1286
tri 13200 1238 13288 1326 sw
tri 13298 1238 13386 1326 ne
rect 13386 1290 13440 1326
rect 13560 1290 15775 1410
rect 13386 1238 15775 1290
rect 12886 1188 13288 1238
rect 12366 1158 12788 1188
rect 11874 1100 12268 1158
rect 11364 1060 11776 1100
tri 11776 1060 11816 1100 sw
tri 11874 1060 11914 1100 ne
rect 11914 1060 12268 1100
tri 12268 1060 12366 1158 sw
tri 12366 1060 12464 1158 ne
rect 12464 1100 12788 1158
tri 12788 1100 12876 1188 sw
tri 12886 1100 12974 1188 ne
rect 12974 1158 13288 1188
tri 13288 1158 13368 1238 sw
tri 13386 1158 13466 1238 ne
rect 13466 1158 14075 1238
rect 12974 1100 13368 1158
rect 12464 1060 12876 1100
tri 12876 1060 12916 1100 sw
tri 12974 1060 13014 1100 ne
rect 13014 1060 13368 1100
tri 13368 1060 13466 1158 sw
tri 13466 1060 13564 1158 ne
rect 13564 1138 14075 1158
rect 14175 1138 15775 1238
rect 13564 1060 15775 1138
rect -1025 1012 -284 1060
rect -1025 912 -925 1012
rect -825 962 -284 1012
tri -284 962 -186 1060 sw
tri -186 962 -88 1060 ne
rect -88 962 266 1060
tri 266 962 364 1060 sw
tri 364 962 462 1060 ne
rect 462 962 816 1060
tri 816 962 914 1060 sw
tri 914 962 1012 1060 ne
rect 1012 962 1366 1060
tri 1366 962 1464 1060 sw
tri 1464 962 1562 1060 ne
rect 1562 962 1916 1060
tri 1916 962 2014 1060 sw
tri 2014 962 2112 1060 ne
rect 2112 962 2466 1060
tri 2466 962 2564 1060 sw
tri 2564 962 2662 1060 ne
rect 2662 962 3016 1060
tri 3016 962 3114 1060 sw
tri 3114 962 3212 1060 ne
rect 3212 962 3566 1060
tri 3566 962 3664 1060 sw
tri 3664 962 3762 1060 ne
rect 3762 962 4116 1060
tri 4116 962 4214 1060 sw
tri 4214 962 4312 1060 ne
rect 4312 962 4666 1060
tri 4666 962 4764 1060 sw
tri 4764 962 4862 1060 ne
rect 4862 962 5216 1060
tri 5216 962 5314 1060 sw
tri 5314 962 5412 1060 ne
rect 5412 962 5766 1060
tri 5766 962 5864 1060 sw
tri 5864 962 5962 1060 ne
rect 5962 962 6316 1060
tri 6316 962 6414 1060 sw
tri 6414 962 6512 1060 ne
rect 6512 962 6866 1060
tri 6866 962 6964 1060 sw
tri 6964 962 7062 1060 ne
rect 7062 962 7416 1060
tri 7416 962 7514 1060 sw
tri 7514 962 7612 1060 ne
rect 7612 962 7966 1060
tri 7966 962 8064 1060 sw
tri 8064 962 8162 1060 ne
rect 8162 962 8516 1060
tri 8516 962 8614 1060 sw
tri 8614 962 8712 1060 ne
rect 8712 962 9066 1060
tri 9066 962 9164 1060 sw
tri 9164 962 9262 1060 ne
rect 9262 962 9616 1060
tri 9616 962 9714 1060 sw
tri 9714 962 9812 1060 ne
rect 9812 962 10166 1060
tri 10166 962 10264 1060 sw
tri 10264 962 10362 1060 ne
rect 10362 962 10716 1060
tri 10716 962 10814 1060 sw
tri 10814 962 10912 1060 ne
rect 10912 962 11266 1060
tri 11266 962 11364 1060 sw
tri 11364 962 11462 1060 ne
rect 11462 962 11816 1060
tri 11816 962 11914 1060 sw
tri 11914 962 12012 1060 ne
rect 12012 962 12366 1060
tri 12366 962 12464 1060 sw
tri 12464 962 12562 1060 ne
rect 12562 962 12916 1060
tri 12916 962 13014 1060 sw
tri 13014 962 13112 1060 ne
rect 13112 962 13466 1060
tri 13466 962 13564 1060 sw
tri 13564 962 13662 1060 ne
rect 13662 962 15775 1060
rect -825 912 -186 962
rect -1025 864 -186 912
tri -186 864 -88 962 sw
tri -88 864 10 962 ne
rect 10 864 364 962
tri 364 864 462 962 sw
tri 462 864 560 962 ne
rect 560 864 914 962
tri 914 864 1012 962 sw
tri 1012 864 1110 962 ne
rect 1110 864 1464 962
tri 1464 864 1562 962 sw
tri 1562 864 1660 962 ne
rect 1660 864 2014 962
tri 2014 864 2112 962 sw
tri 2112 864 2210 962 ne
rect 2210 864 2564 962
tri 2564 864 2662 962 sw
tri 2662 864 2760 962 ne
rect 2760 864 3114 962
tri 3114 864 3212 962 sw
tri 3212 864 3310 962 ne
rect 3310 864 3664 962
tri 3664 864 3762 962 sw
tri 3762 864 3860 962 ne
rect 3860 864 4214 962
tri 4214 864 4312 962 sw
tri 4312 864 4410 962 ne
rect 4410 864 4764 962
tri 4764 864 4862 962 sw
tri 4862 864 4960 962 ne
rect 4960 864 5314 962
tri 5314 864 5412 962 sw
tri 5412 864 5510 962 ne
rect 5510 864 5864 962
tri 5864 864 5962 962 sw
tri 5962 864 6060 962 ne
rect 6060 864 6414 962
tri 6414 864 6512 962 sw
tri 6512 864 6610 962 ne
rect 6610 864 6964 962
tri 6964 864 7062 962 sw
tri 7062 864 7160 962 ne
rect 7160 864 7514 962
tri 7514 864 7612 962 sw
tri 7612 864 7710 962 ne
rect 7710 864 8064 962
tri 8064 864 8162 962 sw
tri 8162 864 8260 962 ne
rect 8260 864 8614 962
tri 8614 864 8712 962 sw
tri 8712 864 8810 962 ne
rect 8810 864 9164 962
tri 9164 864 9262 962 sw
tri 9262 864 9360 962 ne
rect 9360 864 9714 962
tri 9714 864 9812 962 sw
tri 9812 864 9910 962 ne
rect 9910 864 10264 962
tri 10264 864 10362 962 sw
tri 10362 864 10460 962 ne
rect 10460 864 10814 962
tri 10814 864 10912 962 sw
tri 10912 864 11010 962 ne
rect 11010 864 11364 962
tri 11364 864 11462 962 sw
tri 11462 864 11560 962 ne
rect 11560 864 11914 962
tri 11914 864 12012 962 sw
tri 12012 864 12110 962 ne
rect 12110 864 12464 962
tri 12464 864 12562 962 sw
tri 12562 864 12660 962 ne
rect 12660 864 13014 962
tri 13014 864 13112 962 sw
tri 13112 864 13210 962 ne
rect 13210 864 13564 962
tri 13564 864 13662 962 sw
rect -1025 860 -88 864
rect -1025 740 -310 860
rect -190 776 -88 860
tri -88 776 0 864 sw
tri 10 776 98 864 ne
rect 98 860 462 864
rect 98 776 240 860
rect -190 740 0 776
rect -1025 736 0 740
tri 0 736 40 776 sw
tri 98 736 138 776 ne
rect 138 740 240 776
rect 360 776 462 860
tri 462 776 550 864 sw
tri 560 776 648 864 ne
rect 648 860 1012 864
rect 648 776 790 860
rect 360 740 550 776
rect 138 736 550 740
tri -412 638 -314 736 ne
rect -314 638 40 736
tri 40 638 138 736 sw
tri 138 638 236 736 ne
rect 236 688 550 736
tri 550 688 638 776 sw
tri 648 688 736 776 ne
rect 736 740 790 776
rect 910 776 1012 860
tri 1012 776 1100 864 sw
tri 1110 776 1198 864 ne
rect 1198 860 1562 864
rect 1198 776 1340 860
rect 910 740 1100 776
rect 736 736 1100 740
tri 1100 736 1140 776 sw
tri 1198 736 1238 776 ne
rect 1238 740 1340 776
rect 1460 776 1562 860
tri 1562 776 1650 864 sw
tri 1660 776 1748 864 ne
rect 1748 860 2112 864
rect 1748 776 1890 860
rect 1460 740 1650 776
rect 1238 736 1650 740
rect 736 688 1140 736
rect 236 638 638 688
rect -2525 550 -412 638
tri -412 550 -324 638 sw
tri -314 550 -226 638 ne
rect -226 550 138 638
tri 138 550 226 638 sw
tri 236 550 324 638 ne
rect 324 608 638 638
tri 638 608 718 688 sw
tri 736 608 816 688 ne
rect 816 638 1140 688
tri 1140 638 1238 736 sw
tri 1238 638 1336 736 ne
rect 1336 688 1650 736
tri 1650 688 1738 776 sw
tri 1748 688 1836 776 ne
rect 1836 740 1890 776
rect 2010 776 2112 860
tri 2112 776 2200 864 sw
tri 2210 776 2298 864 ne
rect 2298 860 2662 864
rect 2298 776 2440 860
rect 2010 740 2200 776
rect 1836 736 2200 740
tri 2200 736 2240 776 sw
tri 2298 736 2338 776 ne
rect 2338 740 2440 776
rect 2560 776 2662 860
tri 2662 776 2750 864 sw
tri 2760 776 2848 864 ne
rect 2848 860 3212 864
rect 2848 776 2990 860
rect 2560 740 2750 776
rect 2338 736 2750 740
rect 1836 688 2240 736
rect 1336 638 1738 688
rect 816 608 1238 638
rect 324 550 718 608
rect -2525 510 -324 550
tri -324 510 -284 550 sw
tri -226 510 -186 550 ne
rect -186 510 226 550
tri 226 510 266 550 sw
tri 324 510 364 550 ne
rect 364 510 718 550
tri 718 510 816 608 sw
tri 816 510 914 608 ne
rect 914 550 1238 608
tri 1238 550 1326 638 sw
tri 1336 550 1424 638 ne
rect 1424 608 1738 638
tri 1738 608 1818 688 sw
tri 1836 608 1916 688 ne
rect 1916 638 2240 688
tri 2240 638 2338 736 sw
tri 2338 638 2436 736 ne
rect 2436 688 2750 736
tri 2750 688 2838 776 sw
tri 2848 688 2936 776 ne
rect 2936 740 2990 776
rect 3110 776 3212 860
tri 3212 776 3300 864 sw
tri 3310 776 3398 864 ne
rect 3398 860 3762 864
rect 3398 776 3540 860
rect 3110 740 3300 776
rect 2936 736 3300 740
tri 3300 736 3340 776 sw
tri 3398 736 3438 776 ne
rect 3438 740 3540 776
rect 3660 776 3762 860
tri 3762 776 3850 864 sw
tri 3860 776 3948 864 ne
rect 3948 860 4312 864
rect 3948 776 4090 860
rect 3660 740 3850 776
rect 3438 736 3850 740
rect 2936 688 3340 736
rect 2436 638 2838 688
rect 1916 608 2338 638
rect 1424 550 1818 608
rect 914 510 1326 550
tri 1326 510 1366 550 sw
tri 1424 510 1464 550 ne
rect 1464 510 1818 550
tri 1818 510 1916 608 sw
tri 1916 510 2014 608 ne
rect 2014 550 2338 608
tri 2338 550 2426 638 sw
tri 2436 550 2524 638 ne
rect 2524 608 2838 638
tri 2838 608 2918 688 sw
tri 2936 608 3016 688 ne
rect 3016 638 3340 688
tri 3340 638 3438 736 sw
tri 3438 638 3536 736 ne
rect 3536 688 3850 736
tri 3850 688 3938 776 sw
tri 3948 688 4036 776 ne
rect 4036 740 4090 776
rect 4210 776 4312 860
tri 4312 776 4400 864 sw
tri 4410 776 4498 864 ne
rect 4498 860 4862 864
rect 4498 776 4640 860
rect 4210 740 4400 776
rect 4036 736 4400 740
tri 4400 736 4440 776 sw
tri 4498 736 4538 776 ne
rect 4538 740 4640 776
rect 4760 776 4862 860
tri 4862 776 4950 864 sw
tri 4960 776 5048 864 ne
rect 5048 860 5412 864
rect 5048 776 5190 860
rect 4760 740 4950 776
rect 4538 736 4950 740
rect 4036 688 4440 736
rect 3536 638 3938 688
rect 3016 608 3438 638
rect 2524 550 2918 608
rect 2014 510 2426 550
tri 2426 510 2466 550 sw
tri 2524 510 2564 550 ne
rect 2564 510 2918 550
tri 2918 510 3016 608 sw
tri 3016 510 3114 608 ne
rect 3114 550 3438 608
tri 3438 550 3526 638 sw
tri 3536 550 3624 638 ne
rect 3624 608 3938 638
tri 3938 608 4018 688 sw
tri 4036 608 4116 688 ne
rect 4116 638 4440 688
tri 4440 638 4538 736 sw
tri 4538 638 4636 736 ne
rect 4636 688 4950 736
tri 4950 688 5038 776 sw
tri 5048 688 5136 776 ne
rect 5136 740 5190 776
rect 5310 776 5412 860
tri 5412 776 5500 864 sw
tri 5510 776 5598 864 ne
rect 5598 860 5962 864
rect 5598 776 5740 860
rect 5310 740 5500 776
rect 5136 736 5500 740
tri 5500 736 5540 776 sw
tri 5598 736 5638 776 ne
rect 5638 740 5740 776
rect 5860 776 5962 860
tri 5962 776 6050 864 sw
tri 6060 776 6148 864 ne
rect 6148 860 6512 864
rect 6148 776 6290 860
rect 5860 740 6050 776
rect 5638 736 6050 740
rect 5136 688 5540 736
rect 4636 638 5038 688
rect 4116 608 4538 638
rect 3624 550 4018 608
rect 3114 510 3526 550
tri 3526 510 3566 550 sw
tri 3624 510 3664 550 ne
rect 3664 510 4018 550
tri 4018 510 4116 608 sw
tri 4116 510 4214 608 ne
rect 4214 550 4538 608
tri 4538 550 4626 638 sw
tri 4636 550 4724 638 ne
rect 4724 608 5038 638
tri 5038 608 5118 688 sw
tri 5136 608 5216 688 ne
rect 5216 638 5540 688
tri 5540 638 5638 736 sw
tri 5638 638 5736 736 ne
rect 5736 688 6050 736
tri 6050 688 6138 776 sw
tri 6148 688 6236 776 ne
rect 6236 740 6290 776
rect 6410 776 6512 860
tri 6512 776 6600 864 sw
tri 6610 776 6698 864 ne
rect 6698 860 7062 864
rect 6698 776 6840 860
rect 6410 740 6600 776
rect 6236 736 6600 740
tri 6600 736 6640 776 sw
tri 6698 736 6738 776 ne
rect 6738 740 6840 776
rect 6960 776 7062 860
tri 7062 776 7150 864 sw
tri 7160 776 7248 864 ne
rect 7248 860 7612 864
rect 7248 776 7390 860
rect 6960 740 7150 776
rect 6738 736 7150 740
rect 6236 688 6640 736
rect 5736 638 6138 688
rect 5216 608 5638 638
rect 4724 550 5118 608
rect 4214 510 4626 550
tri 4626 510 4666 550 sw
tri 4724 510 4764 550 ne
rect 4764 510 5118 550
tri 5118 510 5216 608 sw
tri 5216 510 5314 608 ne
rect 5314 550 5638 608
tri 5638 550 5726 638 sw
tri 5736 550 5824 638 ne
rect 5824 608 6138 638
tri 6138 608 6218 688 sw
tri 6236 608 6316 688 ne
rect 6316 638 6640 688
tri 6640 638 6738 736 sw
tri 6738 638 6836 736 ne
rect 6836 688 7150 736
tri 7150 688 7238 776 sw
tri 7248 688 7336 776 ne
rect 7336 740 7390 776
rect 7510 776 7612 860
tri 7612 776 7700 864 sw
tri 7710 776 7798 864 ne
rect 7798 860 8162 864
rect 7798 776 7940 860
rect 7510 740 7700 776
rect 7336 736 7700 740
tri 7700 736 7740 776 sw
tri 7798 736 7838 776 ne
rect 7838 740 7940 776
rect 8060 776 8162 860
tri 8162 776 8250 864 sw
tri 8260 776 8348 864 ne
rect 8348 860 8712 864
rect 8348 776 8490 860
rect 8060 740 8250 776
rect 7838 736 8250 740
rect 7336 688 7740 736
rect 6836 638 7238 688
rect 6316 608 6738 638
rect 5824 550 6218 608
rect 5314 510 5726 550
tri 5726 510 5766 550 sw
tri 5824 510 5864 550 ne
rect 5864 510 6218 550
tri 6218 510 6316 608 sw
tri 6316 510 6414 608 ne
rect 6414 550 6738 608
tri 6738 550 6826 638 sw
tri 6836 550 6924 638 ne
rect 6924 608 7238 638
tri 7238 608 7318 688 sw
tri 7336 608 7416 688 ne
rect 7416 638 7740 688
tri 7740 638 7838 736 sw
tri 7838 638 7936 736 ne
rect 7936 688 8250 736
tri 8250 688 8338 776 sw
tri 8348 688 8436 776 ne
rect 8436 740 8490 776
rect 8610 776 8712 860
tri 8712 776 8800 864 sw
tri 8810 776 8898 864 ne
rect 8898 860 9262 864
rect 8898 776 9040 860
rect 8610 740 8800 776
rect 8436 736 8800 740
tri 8800 736 8840 776 sw
tri 8898 736 8938 776 ne
rect 8938 740 9040 776
rect 9160 776 9262 860
tri 9262 776 9350 864 sw
tri 9360 776 9448 864 ne
rect 9448 860 9812 864
rect 9448 776 9590 860
rect 9160 740 9350 776
rect 8938 736 9350 740
rect 8436 688 8840 736
rect 7936 638 8338 688
rect 7416 608 7838 638
rect 6924 550 7318 608
rect 6414 510 6826 550
tri 6826 510 6866 550 sw
tri 6924 510 6964 550 ne
rect 6964 510 7318 550
tri 7318 510 7416 608 sw
tri 7416 510 7514 608 ne
rect 7514 550 7838 608
tri 7838 550 7926 638 sw
tri 7936 550 8024 638 ne
rect 8024 608 8338 638
tri 8338 608 8418 688 sw
tri 8436 608 8516 688 ne
rect 8516 638 8840 688
tri 8840 638 8938 736 sw
tri 8938 638 9036 736 ne
rect 9036 688 9350 736
tri 9350 688 9438 776 sw
tri 9448 688 9536 776 ne
rect 9536 740 9590 776
rect 9710 776 9812 860
tri 9812 776 9900 864 sw
tri 9910 776 9998 864 ne
rect 9998 860 10362 864
rect 9998 776 10140 860
rect 9710 740 9900 776
rect 9536 736 9900 740
tri 9900 736 9940 776 sw
tri 9998 736 10038 776 ne
rect 10038 740 10140 776
rect 10260 776 10362 860
tri 10362 776 10450 864 sw
tri 10460 776 10548 864 ne
rect 10548 860 10912 864
rect 10548 776 10690 860
rect 10260 740 10450 776
rect 10038 736 10450 740
rect 9536 688 9940 736
rect 9036 638 9438 688
rect 8516 608 8938 638
rect 8024 550 8418 608
rect 7514 510 7926 550
tri 7926 510 7966 550 sw
tri 8024 510 8064 550 ne
rect 8064 510 8418 550
tri 8418 510 8516 608 sw
tri 8516 510 8614 608 ne
rect 8614 550 8938 608
tri 8938 550 9026 638 sw
tri 9036 550 9124 638 ne
rect 9124 608 9438 638
tri 9438 608 9518 688 sw
tri 9536 608 9616 688 ne
rect 9616 638 9940 688
tri 9940 638 10038 736 sw
tri 10038 638 10136 736 ne
rect 10136 688 10450 736
tri 10450 688 10538 776 sw
tri 10548 688 10636 776 ne
rect 10636 740 10690 776
rect 10810 776 10912 860
tri 10912 776 11000 864 sw
tri 11010 776 11098 864 ne
rect 11098 860 11462 864
rect 11098 776 11240 860
rect 10810 740 11000 776
rect 10636 736 11000 740
tri 11000 736 11040 776 sw
tri 11098 736 11138 776 ne
rect 11138 740 11240 776
rect 11360 776 11462 860
tri 11462 776 11550 864 sw
tri 11560 776 11648 864 ne
rect 11648 860 12012 864
rect 11648 776 11790 860
rect 11360 740 11550 776
rect 11138 736 11550 740
rect 10636 688 11040 736
rect 10136 638 10538 688
rect 9616 608 10038 638
rect 9124 550 9518 608
rect 8614 510 9026 550
tri 9026 510 9066 550 sw
tri 9124 510 9164 550 ne
rect 9164 510 9518 550
tri 9518 510 9616 608 sw
tri 9616 510 9714 608 ne
rect 9714 550 10038 608
tri 10038 550 10126 638 sw
tri 10136 550 10224 638 ne
rect 10224 608 10538 638
tri 10538 608 10618 688 sw
tri 10636 608 10716 688 ne
rect 10716 638 11040 688
tri 11040 638 11138 736 sw
tri 11138 638 11236 736 ne
rect 11236 688 11550 736
tri 11550 688 11638 776 sw
tri 11648 688 11736 776 ne
rect 11736 740 11790 776
rect 11910 776 12012 860
tri 12012 776 12100 864 sw
tri 12110 776 12198 864 ne
rect 12198 860 12562 864
rect 12198 776 12340 860
rect 11910 740 12100 776
rect 11736 736 12100 740
tri 12100 736 12140 776 sw
tri 12198 736 12238 776 ne
rect 12238 740 12340 776
rect 12460 776 12562 860
tri 12562 776 12650 864 sw
tri 12660 776 12748 864 ne
rect 12748 860 13112 864
rect 12748 776 12890 860
rect 12460 740 12650 776
rect 12238 736 12650 740
rect 11736 688 12140 736
rect 11236 638 11638 688
rect 10716 608 11138 638
rect 10224 550 10618 608
rect 9714 510 10126 550
tri 10126 510 10166 550 sw
tri 10224 510 10264 550 ne
rect 10264 510 10618 550
tri 10618 510 10716 608 sw
tri 10716 510 10814 608 ne
rect 10814 550 11138 608
tri 11138 550 11226 638 sw
tri 11236 550 11324 638 ne
rect 11324 608 11638 638
tri 11638 608 11718 688 sw
tri 11736 608 11816 688 ne
rect 11816 638 12140 688
tri 12140 638 12238 736 sw
tri 12238 638 12336 736 ne
rect 12336 688 12650 736
tri 12650 688 12738 776 sw
tri 12748 688 12836 776 ne
rect 12836 740 12890 776
rect 13010 776 13112 860
tri 13112 776 13200 864 sw
tri 13210 776 13298 864 ne
rect 13298 860 14275 864
rect 13298 776 13440 860
rect 13010 740 13200 776
rect 12836 736 13200 740
tri 13200 736 13240 776 sw
tri 13298 736 13338 776 ne
rect 13338 740 13440 776
rect 13560 740 14275 860
rect 13338 736 14275 740
rect 12836 688 13240 736
rect 12336 638 12738 688
rect 11816 608 12238 638
rect 11324 550 11718 608
rect 10814 510 11226 550
tri 11226 510 11266 550 sw
tri 11324 510 11364 550 ne
rect 11364 510 11718 550
tri 11718 510 11816 608 sw
tri 11816 510 11914 608 ne
rect 11914 550 12238 608
tri 12238 550 12326 638 sw
tri 12336 550 12424 638 ne
rect 12424 608 12738 638
tri 12738 608 12818 688 sw
tri 12836 608 12916 688 ne
rect 12916 638 13240 688
tri 13240 638 13338 736 sw
tri 13338 638 13436 736 ne
rect 13436 638 14275 736
rect 12916 608 13338 638
rect 12424 550 12818 608
rect 11914 510 12326 550
tri 12326 510 12366 550 sw
tri 12424 510 12464 550 ne
rect 12464 510 12818 550
tri 12818 510 12916 608 sw
tri 12916 510 13014 608 ne
rect 13014 550 13338 608
tri 13338 550 13426 638 sw
tri 13436 550 13524 638 ne
rect 13524 550 14275 638
rect 13014 510 13426 550
tri 13426 510 13466 550 sw
tri 13524 510 13564 550 ne
rect 13564 510 14275 550
rect -2525 412 -284 510
tri -284 412 -186 510 sw
tri -186 412 -88 510 ne
rect -88 412 266 510
tri 266 412 364 510 sw
tri 364 412 462 510 ne
rect 462 412 816 510
tri 816 412 914 510 sw
tri 914 412 1012 510 ne
rect 1012 412 1366 510
tri 1366 412 1464 510 sw
tri 1464 412 1562 510 ne
rect 1562 412 1916 510
tri 1916 412 2014 510 sw
tri 2014 412 2112 510 ne
rect 2112 412 2466 510
tri 2466 412 2564 510 sw
tri 2564 412 2662 510 ne
rect 2662 412 3016 510
tri 3016 412 3114 510 sw
tri 3114 412 3212 510 ne
rect 3212 412 3566 510
tri 3566 412 3664 510 sw
tri 3664 412 3762 510 ne
rect 3762 412 4116 510
tri 4116 412 4214 510 sw
tri 4214 412 4312 510 ne
rect 4312 412 4666 510
tri 4666 412 4764 510 sw
tri 4764 412 4862 510 ne
rect 4862 412 5216 510
tri 5216 412 5314 510 sw
tri 5314 412 5412 510 ne
rect 5412 412 5766 510
tri 5766 412 5864 510 sw
tri 5864 412 5962 510 ne
rect 5962 412 6316 510
tri 6316 412 6414 510 sw
tri 6414 412 6512 510 ne
rect 6512 412 6866 510
tri 6866 412 6964 510 sw
tri 6964 412 7062 510 ne
rect 7062 412 7416 510
tri 7416 412 7514 510 sw
tri 7514 412 7612 510 ne
rect 7612 412 7966 510
tri 7966 412 8064 510 sw
tri 8064 412 8162 510 ne
rect 8162 412 8516 510
tri 8516 412 8614 510 sw
tri 8614 412 8712 510 ne
rect 8712 412 9066 510
tri 9066 412 9164 510 sw
tri 9164 412 9262 510 ne
rect 9262 412 9616 510
tri 9616 412 9714 510 sw
tri 9714 412 9812 510 ne
rect 9812 412 10166 510
tri 10166 412 10264 510 sw
tri 10264 412 10362 510 ne
rect 10362 412 10716 510
tri 10716 412 10814 510 sw
tri 10814 412 10912 510 ne
rect 10912 412 11266 510
tri 11266 412 11364 510 sw
tri 11364 412 11462 510 ne
rect 11462 412 11816 510
tri 11816 412 11914 510 sw
tri 11914 412 12012 510 ne
rect 12012 412 12366 510
tri 12366 412 12464 510 sw
tri 12464 412 12562 510 ne
rect 12562 412 12916 510
tri 12916 412 13014 510 sw
tri 13014 412 13112 510 ne
rect 13112 412 13466 510
tri 13466 412 13564 510 sw
tri 13564 412 13662 510 ne
rect 13662 412 14275 510
rect -2525 314 -186 412
tri -186 314 -88 412 sw
tri -88 314 10 412 ne
rect 10 314 364 412
tri 364 314 462 412 sw
tri 462 314 560 412 ne
rect 560 314 914 412
tri 914 314 1012 412 sw
tri 1012 314 1110 412 ne
rect 1110 314 1464 412
tri 1464 314 1562 412 sw
tri 1562 314 1660 412 ne
rect 1660 314 2014 412
tri 2014 314 2112 412 sw
tri 2112 314 2210 412 ne
rect 2210 314 2564 412
tri 2564 314 2662 412 sw
tri 2662 314 2760 412 ne
rect 2760 314 3114 412
tri 3114 314 3212 412 sw
tri 3212 314 3310 412 ne
rect 3310 314 3664 412
tri 3664 314 3762 412 sw
tri 3762 314 3860 412 ne
rect 3860 314 4214 412
tri 4214 314 4312 412 sw
tri 4312 314 4410 412 ne
rect 4410 314 4764 412
tri 4764 314 4862 412 sw
tri 4862 314 4960 412 ne
rect 4960 314 5314 412
tri 5314 314 5412 412 sw
tri 5412 314 5510 412 ne
rect 5510 314 5864 412
tri 5864 314 5962 412 sw
tri 5962 314 6060 412 ne
rect 6060 314 6414 412
tri 6414 314 6512 412 sw
tri 6512 314 6610 412 ne
rect 6610 314 6964 412
tri 6964 314 7062 412 sw
tri 7062 314 7160 412 ne
rect 7160 314 7514 412
tri 7514 314 7612 412 sw
tri 7612 314 7710 412 ne
rect 7710 314 8064 412
tri 8064 314 8162 412 sw
tri 8162 314 8260 412 ne
rect 8260 314 8614 412
tri 8614 314 8712 412 sw
tri 8712 314 8810 412 ne
rect 8810 314 9164 412
tri 9164 314 9262 412 sw
tri 9262 314 9360 412 ne
rect 9360 314 9714 412
tri 9714 314 9812 412 sw
tri 9812 314 9910 412 ne
rect 9910 314 10264 412
tri 10264 314 10362 412 sw
tri 10362 314 10460 412 ne
rect 10460 314 10814 412
tri 10814 314 10912 412 sw
tri 10912 314 11010 412 ne
rect 11010 314 11364 412
tri 11364 314 11462 412 sw
tri 11462 314 11560 412 ne
rect 11560 314 11914 412
tri 11914 314 12012 412 sw
tri 12012 314 12110 412 ne
rect 12110 314 12464 412
tri 12464 314 12562 412 sw
tri 12562 314 12660 412 ne
rect 12660 314 13014 412
tri 13014 314 13112 412 sw
tri 13112 314 13210 412 ne
rect 13210 314 13564 412
tri 13564 314 13662 412 sw
rect 14775 314 15775 962
rect -2525 310 -88 314
rect -2525 190 -310 310
rect -190 226 -88 310
tri -88 226 0 314 sw
tri 10 226 98 314 ne
rect 98 310 462 314
rect 98 226 240 310
rect -190 190 0 226
rect -2525 186 0 190
rect -2525 -575 -1525 186
tri -412 88 -314 186 ne
rect -314 138 0 186
tri 0 138 88 226 sw
tri 98 138 186 226 ne
rect 186 190 240 226
rect 360 226 462 310
tri 462 226 550 314 sw
tri 560 226 648 314 ne
rect 648 310 1012 314
rect 648 226 790 310
rect 360 190 550 226
rect 186 186 550 190
tri 550 186 590 226 sw
tri 648 186 688 226 ne
rect 688 190 790 226
rect 910 226 1012 310
tri 1012 226 1100 314 sw
tri 1110 226 1198 314 ne
rect 1198 310 1562 314
rect 1198 226 1340 310
rect 910 190 1100 226
rect 688 186 1100 190
rect 186 138 590 186
rect -314 88 88 138
rect -1025 0 -412 88
tri -412 0 -324 88 sw
tri -314 0 -226 88 ne
rect -226 58 88 88
tri 88 58 168 138 sw
tri 186 58 266 138 ne
rect 266 88 590 138
tri 590 88 688 186 sw
tri 688 88 786 186 ne
rect 786 138 1100 186
tri 1100 138 1188 226 sw
tri 1198 138 1286 226 ne
rect 1286 190 1340 226
rect 1460 226 1562 310
tri 1562 226 1650 314 sw
tri 1660 226 1748 314 ne
rect 1748 310 2112 314
rect 1748 226 1890 310
rect 1460 190 1650 226
rect 1286 186 1650 190
tri 1650 186 1690 226 sw
tri 1748 186 1788 226 ne
rect 1788 190 1890 226
rect 2010 226 2112 310
tri 2112 226 2200 314 sw
tri 2210 226 2298 314 ne
rect 2298 310 2662 314
rect 2298 226 2440 310
rect 2010 190 2200 226
rect 1788 186 2200 190
rect 1286 138 1690 186
rect 786 88 1188 138
rect 266 58 688 88
rect -226 0 168 58
tri 168 0 226 58 sw
tri 266 0 324 58 ne
rect 324 0 688 58
tri 688 0 776 88 sw
tri 786 0 874 88 ne
rect 874 58 1188 88
tri 1188 58 1268 138 sw
tri 1286 58 1366 138 ne
rect 1366 88 1690 138
tri 1690 88 1788 186 sw
tri 1788 88 1886 186 ne
rect 1886 138 2200 186
tri 2200 138 2288 226 sw
tri 2298 138 2386 226 ne
rect 2386 190 2440 226
rect 2560 226 2662 310
tri 2662 226 2750 314 sw
tri 2760 226 2848 314 ne
rect 2848 310 3212 314
rect 2848 226 2990 310
rect 2560 190 2750 226
rect 2386 186 2750 190
tri 2750 186 2790 226 sw
tri 2848 186 2888 226 ne
rect 2888 190 2990 226
rect 3110 226 3212 310
tri 3212 226 3300 314 sw
tri 3310 226 3398 314 ne
rect 3398 310 3762 314
rect 3398 226 3540 310
rect 3110 190 3300 226
rect 2888 186 3300 190
rect 2386 138 2790 186
rect 1886 88 2288 138
rect 1366 58 1788 88
rect 874 0 1268 58
tri 1268 0 1326 58 sw
tri 1366 0 1424 58 ne
rect 1424 0 1788 58
tri 1788 0 1876 88 sw
tri 1886 0 1974 88 ne
rect 1974 58 2288 88
tri 2288 58 2368 138 sw
tri 2386 58 2466 138 ne
rect 2466 88 2790 138
tri 2790 88 2888 186 sw
tri 2888 88 2986 186 ne
rect 2986 138 3300 186
tri 3300 138 3388 226 sw
tri 3398 138 3486 226 ne
rect 3486 190 3540 226
rect 3660 226 3762 310
tri 3762 226 3850 314 sw
tri 3860 226 3948 314 ne
rect 3948 310 4312 314
rect 3948 226 4090 310
rect 3660 190 3850 226
rect 3486 186 3850 190
tri 3850 186 3890 226 sw
tri 3948 186 3988 226 ne
rect 3988 190 4090 226
rect 4210 226 4312 310
tri 4312 226 4400 314 sw
tri 4410 226 4498 314 ne
rect 4498 310 4862 314
rect 4498 226 4640 310
rect 4210 190 4400 226
rect 3988 186 4400 190
rect 3486 138 3890 186
rect 2986 88 3388 138
rect 2466 58 2888 88
rect 1974 0 2368 58
tri 2368 0 2426 58 sw
tri 2466 0 2524 58 ne
rect 2524 0 2888 58
tri 2888 0 2976 88 sw
tri 2986 0 3074 88 ne
rect 3074 58 3388 88
tri 3388 58 3468 138 sw
tri 3486 58 3566 138 ne
rect 3566 88 3890 138
tri 3890 88 3988 186 sw
tri 3988 88 4086 186 ne
rect 4086 138 4400 186
tri 4400 138 4488 226 sw
tri 4498 138 4586 226 ne
rect 4586 190 4640 226
rect 4760 226 4862 310
tri 4862 226 4950 314 sw
tri 4960 226 5048 314 ne
rect 5048 310 5412 314
rect 5048 226 5190 310
rect 4760 190 4950 226
rect 4586 186 4950 190
tri 4950 186 4990 226 sw
tri 5048 186 5088 226 ne
rect 5088 190 5190 226
rect 5310 226 5412 310
tri 5412 226 5500 314 sw
tri 5510 226 5598 314 ne
rect 5598 310 5962 314
rect 5598 226 5740 310
rect 5310 190 5500 226
rect 5088 186 5500 190
rect 4586 138 4990 186
rect 4086 88 4488 138
rect 3566 58 3988 88
rect 3074 0 3468 58
tri 3468 0 3526 58 sw
tri 3566 0 3624 58 ne
rect 3624 0 3988 58
tri 3988 0 4076 88 sw
tri 4086 0 4174 88 ne
rect 4174 58 4488 88
tri 4488 58 4568 138 sw
tri 4586 58 4666 138 ne
rect 4666 88 4990 138
tri 4990 88 5088 186 sw
tri 5088 88 5186 186 ne
rect 5186 138 5500 186
tri 5500 138 5588 226 sw
tri 5598 138 5686 226 ne
rect 5686 190 5740 226
rect 5860 226 5962 310
tri 5962 226 6050 314 sw
tri 6060 226 6148 314 ne
rect 6148 310 6512 314
rect 6148 226 6290 310
rect 5860 190 6050 226
rect 5686 186 6050 190
tri 6050 186 6090 226 sw
tri 6148 186 6188 226 ne
rect 6188 190 6290 226
rect 6410 226 6512 310
tri 6512 226 6600 314 sw
tri 6610 226 6698 314 ne
rect 6698 310 7062 314
rect 6698 226 6840 310
rect 6410 190 6600 226
rect 6188 186 6600 190
rect 5686 138 6090 186
rect 5186 88 5588 138
rect 4666 58 5088 88
rect 4174 0 4568 58
tri 4568 0 4626 58 sw
tri 4666 0 4724 58 ne
rect 4724 0 5088 58
tri 5088 0 5176 88 sw
tri 5186 0 5274 88 ne
rect 5274 58 5588 88
tri 5588 58 5668 138 sw
tri 5686 58 5766 138 ne
rect 5766 88 6090 138
tri 6090 88 6188 186 sw
tri 6188 88 6286 186 ne
rect 6286 138 6600 186
tri 6600 138 6688 226 sw
tri 6698 138 6786 226 ne
rect 6786 190 6840 226
rect 6960 226 7062 310
tri 7062 226 7150 314 sw
tri 7160 226 7248 314 ne
rect 7248 310 7612 314
rect 7248 226 7390 310
rect 6960 190 7150 226
rect 6786 186 7150 190
tri 7150 186 7190 226 sw
tri 7248 186 7288 226 ne
rect 7288 190 7390 226
rect 7510 226 7612 310
tri 7612 226 7700 314 sw
tri 7710 226 7798 314 ne
rect 7798 310 8162 314
rect 7798 226 7940 310
rect 7510 190 7700 226
rect 7288 186 7700 190
rect 6786 138 7190 186
rect 6286 88 6688 138
rect 5766 58 6188 88
rect 5274 0 5668 58
tri 5668 0 5726 58 sw
tri 5766 0 5824 58 ne
rect 5824 0 6188 58
tri 6188 0 6276 88 sw
tri 6286 0 6374 88 ne
rect 6374 58 6688 88
tri 6688 58 6768 138 sw
tri 6786 58 6866 138 ne
rect 6866 88 7190 138
tri 7190 88 7288 186 sw
tri 7288 88 7386 186 ne
rect 7386 138 7700 186
tri 7700 138 7788 226 sw
tri 7798 138 7886 226 ne
rect 7886 190 7940 226
rect 8060 226 8162 310
tri 8162 226 8250 314 sw
tri 8260 226 8348 314 ne
rect 8348 310 8712 314
rect 8348 226 8490 310
rect 8060 190 8250 226
rect 7886 186 8250 190
tri 8250 186 8290 226 sw
tri 8348 186 8388 226 ne
rect 8388 190 8490 226
rect 8610 226 8712 310
tri 8712 226 8800 314 sw
tri 8810 226 8898 314 ne
rect 8898 310 9262 314
rect 8898 226 9040 310
rect 8610 190 8800 226
rect 8388 186 8800 190
rect 7886 138 8290 186
rect 7386 88 7788 138
rect 6866 58 7288 88
rect 6374 0 6768 58
tri 6768 0 6826 58 sw
tri 6866 0 6924 58 ne
rect 6924 0 7288 58
tri 7288 0 7376 88 sw
tri 7386 0 7474 88 ne
rect 7474 58 7788 88
tri 7788 58 7868 138 sw
tri 7886 58 7966 138 ne
rect 7966 88 8290 138
tri 8290 88 8388 186 sw
tri 8388 88 8486 186 ne
rect 8486 138 8800 186
tri 8800 138 8888 226 sw
tri 8898 138 8986 226 ne
rect 8986 190 9040 226
rect 9160 226 9262 310
tri 9262 226 9350 314 sw
tri 9360 226 9448 314 ne
rect 9448 310 9812 314
rect 9448 226 9590 310
rect 9160 190 9350 226
rect 8986 186 9350 190
tri 9350 186 9390 226 sw
tri 9448 186 9488 226 ne
rect 9488 190 9590 226
rect 9710 226 9812 310
tri 9812 226 9900 314 sw
tri 9910 226 9998 314 ne
rect 9998 310 10362 314
rect 9998 226 10140 310
rect 9710 190 9900 226
rect 9488 186 9900 190
rect 8986 138 9390 186
rect 8486 88 8888 138
rect 7966 58 8388 88
rect 7474 0 7868 58
tri 7868 0 7926 58 sw
tri 7966 0 8024 58 ne
rect 8024 0 8388 58
tri 8388 0 8476 88 sw
tri 8486 0 8574 88 ne
rect 8574 58 8888 88
tri 8888 58 8968 138 sw
tri 8986 58 9066 138 ne
rect 9066 88 9390 138
tri 9390 88 9488 186 sw
tri 9488 88 9586 186 ne
rect 9586 138 9900 186
tri 9900 138 9988 226 sw
tri 9998 138 10086 226 ne
rect 10086 190 10140 226
rect 10260 226 10362 310
tri 10362 226 10450 314 sw
tri 10460 226 10548 314 ne
rect 10548 310 10912 314
rect 10548 226 10690 310
rect 10260 190 10450 226
rect 10086 186 10450 190
tri 10450 186 10490 226 sw
tri 10548 186 10588 226 ne
rect 10588 190 10690 226
rect 10810 226 10912 310
tri 10912 226 11000 314 sw
tri 11010 226 11098 314 ne
rect 11098 310 11462 314
rect 11098 226 11240 310
rect 10810 190 11000 226
rect 10588 186 11000 190
rect 10086 138 10490 186
rect 9586 88 9988 138
rect 9066 58 9488 88
rect 8574 0 8968 58
tri 8968 0 9026 58 sw
tri 9066 0 9124 58 ne
rect 9124 0 9488 58
tri 9488 0 9576 88 sw
tri 9586 0 9674 88 ne
rect 9674 58 9988 88
tri 9988 58 10068 138 sw
tri 10086 58 10166 138 ne
rect 10166 88 10490 138
tri 10490 88 10588 186 sw
tri 10588 88 10686 186 ne
rect 10686 138 11000 186
tri 11000 138 11088 226 sw
tri 11098 138 11186 226 ne
rect 11186 190 11240 226
rect 11360 226 11462 310
tri 11462 226 11550 314 sw
tri 11560 226 11648 314 ne
rect 11648 310 12012 314
rect 11648 226 11790 310
rect 11360 190 11550 226
rect 11186 186 11550 190
tri 11550 186 11590 226 sw
tri 11648 186 11688 226 ne
rect 11688 190 11790 226
rect 11910 226 12012 310
tri 12012 226 12100 314 sw
tri 12110 226 12198 314 ne
rect 12198 310 12562 314
rect 12198 226 12340 310
rect 11910 190 12100 226
rect 11688 186 12100 190
rect 11186 138 11590 186
rect 10686 88 11088 138
rect 10166 58 10588 88
rect 9674 0 10068 58
tri 10068 0 10126 58 sw
tri 10166 0 10224 58 ne
rect 10224 0 10588 58
tri 10588 0 10676 88 sw
tri 10686 0 10774 88 ne
rect 10774 58 11088 88
tri 11088 58 11168 138 sw
tri 11186 58 11266 138 ne
rect 11266 88 11590 138
tri 11590 88 11688 186 sw
tri 11688 88 11786 186 ne
rect 11786 138 12100 186
tri 12100 138 12188 226 sw
tri 12198 138 12286 226 ne
rect 12286 190 12340 226
rect 12460 226 12562 310
tri 12562 226 12650 314 sw
tri 12660 226 12748 314 ne
rect 12748 310 13112 314
rect 12748 226 12890 310
rect 12460 190 12650 226
rect 12286 186 12650 190
tri 12650 186 12690 226 sw
tri 12748 186 12788 226 ne
rect 12788 190 12890 226
rect 13010 226 13112 310
tri 13112 226 13200 314 sw
tri 13210 226 13298 314 ne
rect 13298 310 15775 314
rect 13298 226 13440 310
rect 13010 190 13200 226
rect 12788 186 13200 190
rect 12286 138 12690 186
rect 11786 88 12188 138
rect 11266 58 11688 88
rect 10774 0 11168 58
tri 11168 0 11226 58 sw
tri 11266 0 11324 58 ne
rect 11324 0 11688 58
tri 11688 0 11776 88 sw
tri 11786 0 11874 88 ne
rect 11874 58 12188 88
tri 12188 58 12268 138 sw
tri 12286 58 12366 138 ne
rect 12366 88 12690 138
tri 12690 88 12788 186 sw
tri 12788 88 12886 186 ne
rect 12886 138 13200 186
tri 13200 138 13288 226 sw
tri 13298 138 13386 226 ne
rect 13386 190 13440 226
rect 13560 190 15775 310
rect 13386 138 15775 190
rect 12886 88 13288 138
rect 12366 58 12788 88
rect 11874 0 12268 58
tri 12268 0 12326 58 sw
tri 12366 0 12424 58 ne
rect 12424 0 12788 58
tri 12788 0 12876 88 sw
tri 12886 0 12974 88 ne
rect 12974 58 13288 88
tri 13288 58 13368 138 sw
tri 13386 58 13466 138 ne
rect 13466 58 14075 138
rect 12974 0 13368 58
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 226 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -98 226 -40
tri 226 -98 324 0 sw
tri 324 -98 422 0 ne
rect 422 -98 776 0
tri 776 -98 874 0 sw
tri 874 -98 972 0 ne
rect 972 -98 1326 0
tri 1326 -98 1424 0 sw
tri 1424 -98 1522 0 ne
rect 1522 -98 1876 0
tri 1876 -98 1974 0 sw
tri 1974 -98 2072 0 ne
rect 2072 -98 2426 0
tri 2426 -98 2524 0 sw
tri 2524 -98 2622 0 ne
rect 2622 -98 2976 0
tri 2976 -98 3074 0 sw
tri 3074 -98 3172 0 ne
rect 3172 -98 3526 0
tri 3526 -98 3624 0 sw
tri 3624 -98 3722 0 ne
rect 3722 -98 4076 0
tri 4076 -98 4174 0 sw
tri 4174 -98 4272 0 ne
rect 4272 -98 4626 0
tri 4626 -98 4724 0 sw
tri 4724 -98 4822 0 ne
rect 4822 -98 5176 0
tri 5176 -98 5274 0 sw
tri 5274 -98 5372 0 ne
rect 5372 -98 5726 0
tri 5726 -98 5824 0 sw
tri 5824 -98 5922 0 ne
rect 5922 -98 6276 0
tri 6276 -98 6374 0 sw
tri 6374 -98 6472 0 ne
rect 6472 -98 6826 0
tri 6826 -98 6924 0 sw
tri 6924 -98 7022 0 ne
rect 7022 -98 7376 0
tri 7376 -98 7474 0 sw
tri 7474 -98 7572 0 ne
rect 7572 -98 7926 0
tri 7926 -98 8024 0 sw
tri 8024 -98 8122 0 ne
rect 8122 -98 8476 0
tri 8476 -98 8574 0 sw
tri 8574 -98 8672 0 ne
rect 8672 -98 9026 0
tri 9026 -98 9124 0 sw
tri 9124 -98 9222 0 ne
rect 9222 -98 9576 0
tri 9576 -98 9674 0 sw
tri 9674 -98 9772 0 ne
rect 9772 -98 10126 0
tri 10126 -98 10224 0 sw
tri 10224 -98 10322 0 ne
rect 10322 -98 10676 0
tri 10676 -98 10774 0 sw
tri 10774 -98 10872 0 ne
rect 10872 -98 11226 0
tri 11226 -98 11324 0 sw
tri 11324 -98 11422 0 ne
rect 11422 -98 11776 0
tri 11776 -98 11874 0 sw
tri 11874 -98 11972 0 ne
rect 11972 -98 12326 0
tri 12326 -98 12424 0 sw
tri 12424 -98 12522 0 ne
rect 12522 -98 12876 0
tri 12876 -98 12974 0 sw
tri 12974 -98 13072 0 ne
rect 13072 -40 13368 0
tri 13368 -40 13466 58 sw
tri 13466 -40 13564 58 ne
rect 13564 38 14075 58
rect 14175 38 15775 138
rect 13564 -40 15775 38
rect 13072 -98 13466 -40
rect -88 -138 324 -98
tri 324 -138 364 -98 sw
tri 422 -138 462 -98 ne
rect 462 -138 874 -98
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -236 10 -138 ne
rect 10 -236 364 -138
tri 364 -236 462 -138 sw
tri 462 -236 560 -138 ne
rect 560 -186 874 -138
tri 874 -186 962 -98 sw
tri 972 -186 1060 -98 ne
rect 1060 -138 1424 -98
tri 1424 -138 1464 -98 sw
tri 1522 -138 1562 -98 ne
rect 1562 -138 1974 -98
rect 1060 -186 1464 -138
rect 560 -236 962 -186
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
tri 10 -324 98 -236 ne
rect 98 -240 462 -236
rect 98 -324 240 -240
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri 0 -364 40 -324 sw
tri 98 -364 138 -324 ne
rect 138 -360 240 -324
rect 360 -324 462 -240
tri 462 -324 550 -236 sw
tri 560 -324 648 -236 ne
rect 648 -240 962 -236
rect 648 -324 790 -240
rect 360 -360 550 -324
rect 138 -364 550 -360
tri 550 -364 590 -324 sw
tri 648 -364 688 -324 ne
rect 688 -360 790 -324
rect 910 -266 962 -240
tri 962 -266 1042 -186 sw
tri 1060 -266 1140 -186 ne
rect 1140 -236 1464 -186
tri 1464 -236 1562 -138 sw
tri 1562 -236 1660 -138 ne
rect 1660 -186 1974 -138
tri 1974 -186 2062 -98 sw
tri 2072 -186 2160 -98 ne
rect 2160 -138 2524 -98
tri 2524 -138 2564 -98 sw
tri 2622 -138 2662 -98 ne
rect 2662 -138 3074 -98
rect 2160 -186 2564 -138
rect 1660 -236 2062 -186
rect 1140 -240 1562 -236
rect 1140 -266 1340 -240
rect 910 -360 1042 -266
rect 688 -364 1042 -360
tri 1042 -364 1140 -266 sw
tri 1140 -364 1238 -266 ne
rect 1238 -360 1340 -266
rect 1460 -324 1562 -240
tri 1562 -324 1650 -236 sw
tri 1660 -324 1748 -236 ne
rect 1748 -240 2062 -236
rect 1748 -324 1890 -240
rect 1460 -360 1650 -324
rect 1238 -364 1650 -360
tri 1650 -364 1690 -324 sw
tri 1748 -364 1788 -324 ne
rect 1788 -360 1890 -324
rect 2010 -266 2062 -240
tri 2062 -266 2142 -186 sw
tri 2160 -266 2240 -186 ne
rect 2240 -236 2564 -186
tri 2564 -236 2662 -138 sw
tri 2662 -236 2760 -138 ne
rect 2760 -186 3074 -138
tri 3074 -186 3162 -98 sw
tri 3172 -186 3260 -98 ne
rect 3260 -138 3624 -98
tri 3624 -138 3664 -98 sw
tri 3722 -138 3762 -98 ne
rect 3762 -138 4174 -98
rect 3260 -186 3664 -138
rect 2760 -236 3162 -186
rect 2240 -240 2662 -236
rect 2240 -266 2440 -240
rect 2010 -360 2142 -266
rect 1788 -364 2142 -360
tri 2142 -364 2240 -266 sw
tri 2240 -324 2298 -266 ne
rect 2298 -324 2440 -266
tri 2298 -364 2338 -324 ne
rect 2338 -360 2440 -324
rect 2560 -324 2662 -240
tri 2662 -324 2750 -236 sw
tri 2760 -324 2848 -236 ne
rect 2848 -240 3162 -236
rect 2848 -324 2990 -240
rect 2560 -360 2750 -324
rect 2338 -364 2750 -360
tri 2750 -364 2790 -324 sw
tri 2848 -364 2888 -324 ne
rect 2888 -360 2990 -324
rect 3110 -266 3162 -240
tri 3162 -266 3242 -186 sw
tri 3260 -266 3340 -186 ne
rect 3340 -236 3664 -186
tri 3664 -236 3762 -138 sw
tri 3762 -236 3860 -138 ne
rect 3860 -186 4174 -138
tri 4174 -186 4262 -98 sw
tri 4272 -186 4360 -98 ne
rect 4360 -138 4724 -98
tri 4724 -138 4764 -98 sw
tri 4822 -138 4862 -98 ne
rect 4862 -138 5274 -98
rect 4360 -186 4764 -138
rect 3860 -236 4262 -186
rect 3340 -240 3762 -236
rect 3340 -266 3540 -240
rect 3110 -360 3242 -266
rect 2888 -364 3242 -360
tri 3242 -364 3340 -266 sw
tri 3340 -324 3398 -266 ne
rect 3398 -324 3540 -266
tri 3398 -364 3438 -324 ne
rect 3438 -360 3540 -324
rect 3660 -324 3762 -240
tri 3762 -324 3850 -236 sw
tri 3860 -324 3948 -236 ne
rect 3948 -240 4262 -236
rect 3948 -324 4090 -240
rect 3660 -360 3850 -324
rect 3438 -364 3850 -360
tri 3850 -364 3890 -324 sw
tri 3948 -364 3988 -324 ne
rect 3988 -360 4090 -324
rect 4210 -266 4262 -240
tri 4262 -266 4342 -186 sw
tri 4360 -266 4440 -186 ne
rect 4440 -236 4764 -186
tri 4764 -236 4862 -138 sw
tri 4862 -236 4960 -138 ne
rect 4960 -186 5274 -138
tri 5274 -186 5362 -98 sw
tri 5372 -186 5460 -98 ne
rect 5460 -138 5824 -98
tri 5824 -138 5864 -98 sw
tri 5922 -138 5962 -98 ne
rect 5962 -138 6374 -98
rect 5460 -186 5864 -138
rect 4960 -236 5362 -186
rect 4440 -240 4862 -236
rect 4440 -266 4640 -240
rect 4210 -360 4342 -266
rect 3988 -364 4342 -360
tri 4342 -364 4440 -266 sw
tri 4440 -364 4538 -266 ne
rect 4538 -360 4640 -266
rect 4760 -324 4862 -240
tri 4862 -324 4950 -236 sw
tri 4960 -324 5048 -236 ne
rect 5048 -240 5362 -236
rect 5048 -324 5190 -240
rect 4760 -360 4950 -324
rect 4538 -364 4950 -360
tri 4950 -364 4990 -324 sw
tri 5048 -364 5088 -324 ne
rect 5088 -360 5190 -324
rect 5310 -266 5362 -240
tri 5362 -266 5442 -186 sw
tri 5460 -266 5540 -186 ne
rect 5540 -236 5864 -186
tri 5864 -236 5962 -138 sw
tri 5962 -236 6060 -138 ne
rect 6060 -186 6374 -138
tri 6374 -186 6462 -98 sw
tri 6472 -186 6560 -98 ne
rect 6560 -138 6924 -98
tri 6924 -138 6964 -98 sw
tri 7022 -138 7062 -98 ne
rect 7062 -138 7474 -98
rect 6560 -186 6964 -138
rect 6060 -236 6462 -186
rect 5540 -240 5962 -236
rect 5540 -266 5740 -240
rect 5310 -360 5442 -266
rect 5088 -364 5442 -360
tri 5442 -364 5540 -266 sw
tri 5540 -324 5598 -266 ne
rect 5598 -324 5740 -266
tri 5598 -364 5638 -324 ne
rect 5638 -360 5740 -324
rect 5860 -324 5962 -240
tri 5962 -324 6050 -236 sw
tri 6060 -324 6148 -236 ne
rect 6148 -240 6462 -236
rect 6148 -324 6290 -240
rect 5860 -360 6050 -324
rect 5638 -364 6050 -360
tri 6050 -364 6090 -324 sw
tri 6148 -364 6188 -324 ne
rect 6188 -360 6290 -324
rect 6410 -266 6462 -240
tri 6462 -266 6542 -186 sw
tri 6560 -266 6640 -186 ne
rect 6640 -236 6964 -186
tri 6964 -236 7062 -138 sw
tri 7062 -236 7160 -138 ne
rect 7160 -186 7474 -138
tri 7474 -186 7562 -98 sw
tri 7572 -186 7660 -98 ne
rect 7660 -138 8024 -98
tri 8024 -138 8064 -98 sw
tri 8122 -138 8162 -98 ne
rect 8162 -138 8574 -98
rect 7660 -186 8064 -138
rect 7160 -236 7562 -186
rect 6640 -240 7062 -236
rect 6640 -266 6840 -240
rect 6410 -360 6542 -266
rect 6188 -364 6542 -360
tri 6542 -364 6640 -266 sw
tri 6640 -324 6698 -266 ne
rect 6698 -324 6840 -266
tri 6698 -364 6738 -324 ne
rect 6738 -360 6840 -324
rect 6960 -324 7062 -240
tri 7062 -324 7150 -236 sw
tri 7160 -324 7248 -236 ne
rect 7248 -240 7562 -236
rect 7248 -324 7390 -240
rect 6960 -360 7150 -324
rect 6738 -364 7150 -360
tri 7150 -364 7190 -324 sw
tri 7248 -364 7288 -324 ne
rect 7288 -360 7390 -324
rect 7510 -266 7562 -240
tri 7562 -266 7642 -186 sw
tri 7660 -266 7740 -186 ne
rect 7740 -236 8064 -186
tri 8064 -236 8162 -138 sw
tri 8162 -236 8260 -138 ne
rect 8260 -186 8574 -138
tri 8574 -186 8662 -98 sw
tri 8672 -186 8760 -98 ne
rect 8760 -138 9124 -98
tri 9124 -138 9164 -98 sw
tri 9222 -138 9262 -98 ne
rect 9262 -138 9674 -98
rect 8760 -186 9164 -138
rect 8260 -236 8662 -186
rect 7740 -240 8162 -236
rect 7740 -266 7940 -240
rect 7510 -360 7642 -266
rect 7288 -364 7642 -360
tri 7642 -364 7740 -266 sw
tri 7740 -364 7838 -266 ne
rect 7838 -360 7940 -266
rect 8060 -324 8162 -240
tri 8162 -324 8250 -236 sw
tri 8260 -324 8348 -236 ne
rect 8348 -240 8662 -236
rect 8348 -324 8490 -240
rect 8060 -360 8250 -324
rect 7838 -364 8250 -360
tri 8250 -364 8290 -324 sw
tri 8348 -364 8388 -324 ne
rect 8388 -360 8490 -324
rect 8610 -266 8662 -240
tri 8662 -266 8742 -186 sw
tri 8760 -266 8840 -186 ne
rect 8840 -236 9164 -186
tri 9164 -236 9262 -138 sw
tri 9262 -236 9360 -138 ne
rect 9360 -186 9674 -138
tri 9674 -186 9762 -98 sw
tri 9772 -186 9860 -98 ne
rect 9860 -138 10224 -98
tri 10224 -138 10264 -98 sw
tri 10322 -138 10362 -98 ne
rect 10362 -138 10774 -98
rect 9860 -186 10264 -138
rect 9360 -236 9762 -186
rect 8840 -240 9262 -236
rect 8840 -266 9040 -240
rect 8610 -360 8742 -266
rect 8388 -364 8742 -360
tri 8742 -364 8840 -266 sw
tri 8840 -324 8898 -266 ne
rect 8898 -324 9040 -266
tri 8898 -364 8938 -324 ne
rect 8938 -360 9040 -324
rect 9160 -324 9262 -240
tri 9262 -324 9350 -236 sw
tri 9360 -324 9448 -236 ne
rect 9448 -240 9762 -236
rect 9448 -324 9590 -240
rect 9160 -360 9350 -324
rect 8938 -364 9350 -360
tri 9350 -364 9390 -324 sw
tri 9448 -364 9488 -324 ne
rect 9488 -360 9590 -324
rect 9710 -266 9762 -240
tri 9762 -266 9842 -186 sw
tri 9860 -266 9940 -186 ne
rect 9940 -236 10264 -186
tri 10264 -236 10362 -138 sw
tri 10362 -236 10460 -138 ne
rect 10460 -186 10774 -138
tri 10774 -186 10862 -98 sw
tri 10872 -186 10960 -98 ne
rect 10960 -138 11324 -98
tri 11324 -138 11364 -98 sw
tri 11422 -138 11462 -98 ne
rect 11462 -138 11874 -98
rect 10960 -186 11364 -138
rect 10460 -236 10862 -186
rect 9940 -240 10362 -236
rect 9940 -266 10140 -240
rect 9710 -360 9842 -266
rect 9488 -364 9842 -360
tri 9842 -364 9940 -266 sw
tri 9940 -324 9998 -266 ne
rect 9998 -324 10140 -266
tri 9998 -364 10038 -324 ne
rect 10038 -360 10140 -324
rect 10260 -324 10362 -240
tri 10362 -324 10450 -236 sw
tri 10460 -324 10548 -236 ne
rect 10548 -240 10862 -236
rect 10548 -324 10690 -240
rect 10260 -360 10450 -324
rect 10038 -364 10450 -360
tri 10450 -364 10490 -324 sw
tri 10548 -364 10588 -324 ne
rect 10588 -360 10690 -324
rect 10810 -266 10862 -240
tri 10862 -266 10942 -186 sw
tri 10960 -266 11040 -186 ne
rect 11040 -236 11364 -186
tri 11364 -236 11462 -138 sw
tri 11462 -236 11560 -138 ne
rect 11560 -186 11874 -138
tri 11874 -186 11962 -98 sw
tri 11972 -186 12060 -98 ne
rect 12060 -138 12424 -98
tri 12424 -138 12464 -98 sw
tri 12522 -138 12562 -98 ne
rect 12562 -138 12974 -98
rect 12060 -186 12464 -138
rect 11560 -236 11962 -186
rect 11040 -240 11462 -236
rect 11040 -266 11240 -240
rect 10810 -360 10942 -266
rect 10588 -364 10942 -360
tri 10942 -364 11040 -266 sw
tri 11040 -364 11138 -266 ne
rect 11138 -360 11240 -266
rect 11360 -324 11462 -240
tri 11462 -324 11550 -236 sw
tri 11560 -324 11648 -236 ne
rect 11648 -240 11962 -236
rect 11648 -324 11790 -240
rect 11360 -360 11550 -324
rect 11138 -364 11550 -360
tri 11550 -364 11590 -324 sw
tri 11648 -364 11688 -324 ne
rect 11688 -360 11790 -324
rect 11910 -266 11962 -240
tri 11962 -266 12042 -186 sw
tri 12060 -266 12140 -186 ne
rect 12140 -236 12464 -186
tri 12464 -236 12562 -138 sw
tri 12562 -236 12660 -138 ne
rect 12660 -186 12974 -138
tri 12974 -186 13062 -98 sw
tri 13072 -186 13160 -98 ne
rect 13160 -138 13466 -98
tri 13466 -138 13564 -40 sw
tri 13564 -138 13662 -40 ne
rect 13662 -138 15775 -40
rect 13160 -186 13564 -138
rect 12660 -236 13062 -186
rect 12140 -240 12562 -236
rect 12140 -266 12340 -240
rect 11910 -360 12042 -266
rect 11688 -364 12042 -360
tri 12042 -364 12140 -266 sw
tri 12140 -324 12198 -266 ne
rect 12198 -324 12340 -266
tri 12198 -364 12238 -324 ne
rect 12238 -360 12340 -324
rect 12460 -324 12562 -240
tri 12562 -324 12650 -236 sw
tri 12660 -324 12748 -236 ne
rect 12748 -240 13062 -236
rect 12748 -324 12890 -240
rect 12460 -360 12650 -324
rect 12238 -364 12650 -360
tri 12650 -364 12690 -324 sw
tri 12748 -364 12788 -324 ne
rect 12788 -360 12890 -324
rect 13010 -266 13062 -240
tri 13062 -266 13142 -186 sw
tri 13160 -266 13240 -186 ne
rect 13240 -236 13564 -186
tri 13564 -236 13662 -138 sw
rect 13240 -240 14275 -236
rect 13240 -266 13440 -240
rect 13010 -360 13142 -266
rect 12788 -364 13142 -360
tri 13142 -364 13240 -266 sw
tri 13240 -324 13298 -266 ne
rect 13298 -324 13440 -266
tri 13298 -364 13338 -324 ne
rect 13338 -360 13440 -324
rect 13560 -360 14275 -240
rect 13338 -364 14275 -360
tri -412 -462 -314 -364 ne
rect -314 -462 40 -364
tri 40 -462 138 -364 sw
tri 138 -462 236 -364 ne
rect 236 -462 590 -364
tri 590 -462 688 -364 sw
tri 688 -462 786 -364 ne
rect 786 -462 1140 -364
tri 1140 -462 1238 -364 sw
tri 1238 -462 1336 -364 ne
rect 1336 -462 1690 -364
tri 1690 -462 1788 -364 sw
tri 1788 -462 1886 -364 ne
rect 1886 -462 2240 -364
tri 2240 -462 2338 -364 sw
tri 2338 -462 2436 -364 ne
rect 2436 -462 2790 -364
tri 2790 -462 2888 -364 sw
tri 2888 -462 2986 -364 ne
rect 2986 -462 3340 -364
tri 3340 -462 3438 -364 sw
tri 3438 -462 3536 -364 ne
rect 3536 -462 3890 -364
tri 3890 -462 3988 -364 sw
tri 3988 -462 4086 -364 ne
rect 4086 -462 4440 -364
tri 4440 -462 4538 -364 sw
tri 4538 -462 4636 -364 ne
rect 4636 -462 4990 -364
tri 4990 -462 5088 -364 sw
tri 5088 -462 5186 -364 ne
rect 5186 -462 5540 -364
tri 5540 -462 5638 -364 sw
tri 5638 -462 5736 -364 ne
rect 5736 -462 6090 -364
tri 6090 -462 6188 -364 sw
tri 6188 -462 6286 -364 ne
rect 6286 -462 6640 -364
tri 6640 -462 6738 -364 sw
tri 6738 -462 6836 -364 ne
rect 6836 -462 7190 -364
tri 7190 -462 7288 -364 sw
tri 7288 -462 7386 -364 ne
rect 7386 -462 7740 -364
tri 7740 -462 7838 -364 sw
tri 7838 -462 7936 -364 ne
rect 7936 -462 8290 -364
tri 8290 -462 8388 -364 sw
tri 8388 -462 8486 -364 ne
rect 8486 -462 8840 -364
tri 8840 -462 8938 -364 sw
tri 8938 -462 9036 -364 ne
rect 9036 -462 9390 -364
tri 9390 -462 9488 -364 sw
tri 9488 -462 9586 -364 ne
rect 9586 -462 9940 -364
tri 9940 -462 10038 -364 sw
tri 10038 -462 10136 -364 ne
rect 10136 -462 10490 -364
tri 10490 -462 10588 -364 sw
tri 10588 -462 10686 -364 ne
rect 10686 -462 11040 -364
tri 11040 -462 11138 -364 sw
tri 11138 -462 11236 -364 ne
rect 11236 -462 11590 -364
tri 11590 -462 11688 -364 sw
tri 11688 -462 11786 -364 ne
rect 11786 -462 12140 -364
tri 12140 -462 12238 -364 sw
tri 12238 -462 12336 -364 ne
rect 12336 -462 12690 -364
tri 12690 -462 12788 -364 sw
tri 12788 -462 12886 -364 ne
rect 12886 -462 13240 -364
tri 13240 -462 13338 -364 sw
tri 13338 -462 13436 -364 ne
rect -314 -875 138 -462
rect -314 -975 -138 -875
rect -38 -975 138 -875
rect -314 -1575 138 -975
rect 236 -1075 688 -462
rect 786 -875 1238 -462
rect 786 -975 962 -875
rect 1062 -975 1238 -875
rect 786 -1575 1238 -975
rect 1336 -1075 1788 -462
rect 1886 -875 2338 -462
rect 1886 -975 2062 -875
rect 2162 -975 2338 -875
rect 1886 -1575 2338 -975
rect 2436 -1075 2888 -462
rect 2986 -875 3438 -462
rect 2986 -975 3162 -875
rect 3262 -975 3438 -875
rect 2986 -1575 3438 -975
rect 3536 -1075 3988 -462
rect 4086 -875 4538 -462
rect 4086 -975 4262 -875
rect 4362 -975 4538 -875
rect 4086 -1575 4538 -975
rect 4636 -1075 5088 -462
rect 5186 -875 5638 -462
rect 5186 -975 5362 -875
rect 5462 -975 5638 -875
rect 5186 -1575 5638 -975
rect 5736 -1075 6188 -462
rect 6286 -875 6738 -462
rect 6286 -975 6462 -875
rect 6562 -975 6738 -875
rect 6286 -1575 6738 -975
rect 6836 -1075 7288 -462
rect 7386 -875 7838 -462
rect 7386 -975 7562 -875
rect 7662 -975 7838 -875
rect 7386 -1575 7838 -975
rect 7936 -1075 8388 -462
rect 8486 -875 8938 -462
rect 8486 -975 8662 -875
rect 8762 -975 8938 -875
rect 8486 -1575 8938 -975
rect 9036 -1075 9488 -462
rect 9586 -875 10038 -462
rect 9586 -975 9762 -875
rect 9862 -975 10038 -875
rect 9586 -1575 10038 -975
rect 10136 -1075 10588 -462
rect 10686 -875 11138 -462
rect 10686 -975 10862 -875
rect 10962 -975 11138 -875
rect 10686 -1575 11138 -975
rect 11236 -1075 11688 -462
rect 11786 -875 12238 -462
rect 11786 -975 11962 -875
rect 12062 -975 12238 -875
rect 11786 -1575 12238 -975
rect 12336 -1075 12788 -462
rect 12886 -875 13338 -462
rect 12886 -975 13062 -875
rect 13162 -975 13338 -875
rect 12886 -1575 13338 -975
rect 13436 -688 14275 -364
rect 13436 -1075 13888 -688
rect 14775 -1575 15775 -138
rect -525 -2575 15775 -1575
<< via3 >>
rect 88 14025 188 14125
rect 1188 14025 1288 14125
rect 2288 14025 2388 14125
rect 3388 14025 3488 14125
rect 4488 14025 4588 14125
rect 5588 14025 5688 14125
rect 6688 14025 6788 14125
rect 7788 14025 7888 14125
rect 8888 14025 8988 14125
rect 9988 14025 10088 14125
rect 11088 14025 11188 14125
rect 12188 14025 12288 14125
rect 13288 14025 13388 14125
rect -310 13390 -190 13510
rect 240 13390 360 13510
rect 790 13390 910 13510
rect 1340 13390 1460 13510
rect 1890 13390 2010 13510
rect 2440 13390 2560 13510
rect 2990 13390 3110 13510
rect 3540 13390 3660 13510
rect 4090 13390 4210 13510
rect 4640 13390 4760 13510
rect 5190 13390 5310 13510
rect 5740 13390 5860 13510
rect 6290 13390 6410 13510
rect 6840 13390 6960 13510
rect 7390 13390 7510 13510
rect 7940 13390 8060 13510
rect 8490 13390 8610 13510
rect 9040 13390 9160 13510
rect 9590 13390 9710 13510
rect 10140 13390 10260 13510
rect 10690 13390 10810 13510
rect 11240 13390 11360 13510
rect 11790 13390 11910 13510
rect 12340 13390 12460 13510
rect 12890 13390 13010 13510
rect 13440 13390 13560 13510
rect 14075 13238 14175 13338
rect -925 13012 -825 13112
rect -310 12840 -190 12960
rect 240 12840 360 12960
rect 790 12840 910 12960
rect 1340 12840 1460 12960
rect 1890 12840 2010 12960
rect 2440 12840 2560 12960
rect 2990 12840 3110 12960
rect 3540 12840 3660 12960
rect 4090 12840 4210 12960
rect 4640 12840 4760 12960
rect 5190 12840 5310 12960
rect 5740 12840 5860 12960
rect 6290 12840 6410 12960
rect 6840 12840 6960 12960
rect 7390 12840 7510 12960
rect 7940 12840 8060 12960
rect 8490 12840 8610 12960
rect 9040 12840 9160 12960
rect 9590 12840 9710 12960
rect 10140 12840 10260 12960
rect 10690 12840 10810 12960
rect 11240 12840 11360 12960
rect 11790 12840 11910 12960
rect 12340 12840 12460 12960
rect 12890 12840 13010 12960
rect 13440 12840 13560 12960
rect -310 12290 -190 12410
rect 240 12290 360 12410
rect 790 12290 910 12410
rect 1340 12290 1460 12410
rect 1890 12290 2010 12410
rect 2440 12290 2560 12410
rect 2990 12290 3110 12410
rect 3540 12290 3660 12410
rect 4090 12290 4210 12410
rect 4640 12290 4760 12410
rect 5190 12290 5310 12410
rect 5740 12290 5860 12410
rect 6290 12290 6410 12410
rect 6840 12290 6960 12410
rect 7390 12290 7510 12410
rect 7940 12290 8060 12410
rect 8490 12290 8610 12410
rect 9040 12290 9160 12410
rect 9590 12290 9710 12410
rect 10140 12290 10260 12410
rect 10690 12290 10810 12410
rect 11240 12290 11360 12410
rect 11790 12290 11910 12410
rect 12340 12290 12460 12410
rect 12890 12290 13010 12410
rect 13440 12290 13560 12410
rect 14075 12138 14175 12238
rect -925 11912 -825 12012
rect -310 11740 -190 11860
rect 240 11740 360 11860
rect 790 11740 910 11860
rect 1340 11740 1460 11860
rect 1890 11740 2010 11860
rect 2440 11740 2560 11860
rect 2990 11740 3110 11860
rect 3540 11740 3660 11860
rect 4090 11740 4210 11860
rect 4640 11740 4760 11860
rect 5190 11740 5310 11860
rect 5740 11740 5860 11860
rect 6290 11740 6410 11860
rect 6840 11740 6960 11860
rect 7390 11740 7510 11860
rect 7940 11740 8060 11860
rect 8490 11740 8610 11860
rect 9040 11740 9160 11860
rect 9590 11740 9710 11860
rect 10140 11740 10260 11860
rect 10690 11740 10810 11860
rect 11240 11740 11360 11860
rect 11790 11740 11910 11860
rect 12340 11740 12460 11860
rect 12890 11740 13010 11860
rect 13440 11740 13560 11860
rect -310 11190 -190 11310
rect 240 11190 360 11310
rect 790 11190 910 11310
rect 1340 11190 1460 11310
rect 1890 11190 2010 11310
rect 2440 11190 2560 11310
rect 2990 11190 3110 11310
rect 3540 11190 3660 11310
rect 4090 11190 4210 11310
rect 4640 11190 4760 11310
rect 5190 11190 5310 11310
rect 5740 11190 5860 11310
rect 6290 11190 6410 11310
rect 6840 11190 6960 11310
rect 7390 11190 7510 11310
rect 7940 11190 8060 11310
rect 8490 11190 8610 11310
rect 9040 11190 9160 11310
rect 9590 11190 9710 11310
rect 10140 11190 10260 11310
rect 10690 11190 10810 11310
rect 11240 11190 11360 11310
rect 11790 11190 11910 11310
rect 12340 11190 12460 11310
rect 12890 11190 13010 11310
rect 13440 11190 13560 11310
rect 14075 11038 14175 11138
rect -925 10812 -825 10912
rect -310 10640 -190 10760
rect 240 10640 360 10760
rect 790 10640 910 10760
rect 1340 10640 1460 10760
rect 1890 10640 2010 10760
rect 2440 10640 2560 10760
rect 2990 10640 3110 10760
rect 3540 10640 3660 10760
rect 4090 10640 4210 10760
rect 4640 10640 4760 10760
rect 5190 10640 5310 10760
rect 5740 10640 5860 10760
rect 6290 10640 6410 10760
rect 6840 10640 6960 10760
rect 7390 10640 7510 10760
rect 7940 10640 8060 10760
rect 8490 10640 8610 10760
rect 9040 10640 9160 10760
rect 9590 10640 9710 10760
rect 10140 10640 10260 10760
rect 10690 10640 10810 10760
rect 11240 10640 11360 10760
rect 11790 10640 11910 10760
rect 12340 10640 12460 10760
rect 12890 10640 13010 10760
rect 13440 10640 13560 10760
rect -310 10090 -190 10210
rect 240 10090 360 10210
rect 790 10090 910 10210
rect 1340 10090 1460 10210
rect 1890 10090 2010 10210
rect 2440 10090 2560 10210
rect 2990 10090 3110 10210
rect 3540 10090 3660 10210
rect 4090 10090 4210 10210
rect 4640 10090 4760 10210
rect 5190 10090 5310 10210
rect 5740 10090 5860 10210
rect 6290 10090 6410 10210
rect 6840 10090 6960 10210
rect 7390 10090 7510 10210
rect 7940 10090 8060 10210
rect 8490 10090 8610 10210
rect 9040 10090 9160 10210
rect 9590 10090 9710 10210
rect 10140 10090 10260 10210
rect 10690 10090 10810 10210
rect 11240 10090 11360 10210
rect 11790 10090 11910 10210
rect 12340 10090 12460 10210
rect 12890 10090 13010 10210
rect 13440 10090 13560 10210
rect 14075 9938 14175 10038
rect -925 9712 -825 9812
rect -310 9540 -190 9660
rect 240 9540 360 9660
rect 790 9540 910 9660
rect 1340 9540 1460 9660
rect 1890 9540 2010 9660
rect 2440 9540 2560 9660
rect 2990 9540 3110 9660
rect 3540 9540 3660 9660
rect 4090 9540 4210 9660
rect 4640 9540 4760 9660
rect 5190 9540 5310 9660
rect 5740 9540 5860 9660
rect 6290 9540 6410 9660
rect 6840 9540 6960 9660
rect 7390 9540 7510 9660
rect 7940 9540 8060 9660
rect 8490 9540 8610 9660
rect 9040 9540 9160 9660
rect 9590 9540 9710 9660
rect 10140 9540 10260 9660
rect 10690 9540 10810 9660
rect 11240 9540 11360 9660
rect 11790 9540 11910 9660
rect 12340 9540 12460 9660
rect 12890 9540 13010 9660
rect 13440 9540 13560 9660
rect -310 8990 -190 9110
rect 240 8990 360 9110
rect 790 8990 910 9110
rect 1340 8990 1460 9110
rect 1890 8990 2010 9110
rect 2440 8990 2560 9110
rect 2990 8990 3110 9110
rect 3540 8990 3660 9110
rect 4090 8990 4210 9110
rect 4640 8990 4760 9110
rect 5190 8990 5310 9110
rect 5740 8990 5860 9110
rect 6290 8990 6410 9110
rect 6840 8990 6960 9110
rect 7390 8990 7510 9110
rect 7940 8990 8060 9110
rect 8490 8990 8610 9110
rect 9040 8990 9160 9110
rect 9590 8990 9710 9110
rect 10140 8990 10260 9110
rect 10690 8990 10810 9110
rect 11240 8990 11360 9110
rect 11790 8990 11910 9110
rect 12340 8990 12460 9110
rect 12890 8990 13010 9110
rect 13440 8990 13560 9110
rect 14075 8838 14175 8938
rect -925 8612 -825 8712
rect -310 8440 -190 8560
rect 240 8440 360 8560
rect 790 8440 910 8560
rect 1340 8440 1460 8560
rect 1890 8440 2010 8560
rect 2440 8440 2560 8560
rect 2990 8440 3110 8560
rect 3540 8440 3660 8560
rect 4090 8440 4210 8560
rect 4640 8440 4760 8560
rect 5190 8440 5310 8560
rect 5740 8440 5860 8560
rect 6290 8440 6410 8560
rect 6840 8440 6960 8560
rect 7390 8440 7510 8560
rect 7940 8440 8060 8560
rect 8490 8440 8610 8560
rect 9040 8440 9160 8560
rect 9590 8440 9710 8560
rect 10140 8440 10260 8560
rect 10690 8440 10810 8560
rect 11240 8440 11360 8560
rect 11790 8440 11910 8560
rect 12340 8440 12460 8560
rect 12890 8440 13010 8560
rect 13440 8440 13560 8560
rect -310 7890 -190 8010
rect 240 7890 360 8010
rect 790 7890 910 8010
rect 1340 7890 1460 8010
rect 1890 7890 2010 8010
rect 2440 7890 2560 8010
rect 2990 7890 3110 8010
rect 3540 7890 3660 8010
rect 4090 7890 4210 8010
rect 4640 7890 4760 8010
rect 5190 7890 5310 8010
rect 5740 7890 5860 8010
rect 6290 7890 6410 8010
rect 6840 7890 6960 8010
rect 7390 7890 7510 8010
rect 7940 7890 8060 8010
rect 8490 7890 8610 8010
rect 9040 7890 9160 8010
rect 9590 7890 9710 8010
rect 10140 7890 10260 8010
rect 10690 7890 10810 8010
rect 11240 7890 11360 8010
rect 11790 7890 11910 8010
rect 12340 7890 12460 8010
rect 12890 7890 13010 8010
rect 13440 7890 13560 8010
rect 14075 7738 14175 7838
rect -925 7512 -825 7612
rect -310 7340 -190 7460
rect 240 7340 360 7460
rect 790 7340 910 7460
rect 1340 7340 1460 7460
rect 1890 7340 2010 7460
rect 2440 7340 2560 7460
rect 2990 7340 3110 7460
rect 3540 7340 3660 7460
rect 4090 7340 4210 7460
rect 4640 7340 4760 7460
rect 5190 7340 5310 7460
rect 5740 7340 5860 7460
rect 6290 7340 6410 7460
rect 6840 7340 6960 7460
rect 7390 7340 7510 7460
rect 7940 7340 8060 7460
rect 8490 7340 8610 7460
rect 9040 7340 9160 7460
rect 9590 7340 9710 7460
rect 10140 7340 10260 7460
rect 10690 7340 10810 7460
rect 11240 7340 11360 7460
rect 11790 7340 11910 7460
rect 12340 7340 12460 7460
rect 12890 7340 13010 7460
rect 13440 7340 13560 7460
rect -310 6790 -190 6910
rect 240 6790 360 6910
rect 790 6790 910 6910
rect 1340 6790 1460 6910
rect 1890 6790 2010 6910
rect 2440 6790 2560 6910
rect 2990 6790 3110 6910
rect 3540 6790 3660 6910
rect 4090 6790 4210 6910
rect 4640 6790 4760 6910
rect 5190 6790 5310 6910
rect 5740 6790 5860 6910
rect 6290 6790 6410 6910
rect 6840 6790 6960 6910
rect 7390 6790 7510 6910
rect 7940 6790 8060 6910
rect 8490 6790 8610 6910
rect 9040 6790 9160 6910
rect 9590 6790 9710 6910
rect 10140 6790 10260 6910
rect 10690 6790 10810 6910
rect 11240 6790 11360 6910
rect 11790 6790 11910 6910
rect 12340 6790 12460 6910
rect 12890 6790 13010 6910
rect 13440 6790 13560 6910
rect 14075 6638 14175 6738
rect -925 6412 -825 6512
rect -310 6240 -190 6360
rect 240 6240 360 6360
rect 790 6240 910 6360
rect 1340 6240 1460 6360
rect 1890 6240 2010 6360
rect 2440 6240 2560 6360
rect 2990 6240 3110 6360
rect 3540 6240 3660 6360
rect 4090 6240 4210 6360
rect 4640 6240 4760 6360
rect 5190 6240 5310 6360
rect 5740 6240 5860 6360
rect 6290 6240 6410 6360
rect 6840 6240 6960 6360
rect 7390 6240 7510 6360
rect 7940 6240 8060 6360
rect 8490 6240 8610 6360
rect 9040 6240 9160 6360
rect 9590 6240 9710 6360
rect 10140 6240 10260 6360
rect 10690 6240 10810 6360
rect 11240 6240 11360 6360
rect 11790 6240 11910 6360
rect 12340 6240 12460 6360
rect 12890 6240 13010 6360
rect 13440 6240 13560 6360
rect -310 5690 -190 5810
rect 240 5690 360 5810
rect 790 5690 910 5810
rect 1340 5690 1460 5810
rect 1890 5690 2010 5810
rect 2440 5690 2560 5810
rect 2990 5690 3110 5810
rect 3540 5690 3660 5810
rect 4090 5690 4210 5810
rect 4640 5690 4760 5810
rect 5190 5690 5310 5810
rect 5740 5690 5860 5810
rect 6290 5690 6410 5810
rect 6840 5690 6960 5810
rect 7390 5690 7510 5810
rect 7940 5690 8060 5810
rect 8490 5690 8610 5810
rect 9040 5690 9160 5810
rect 9590 5690 9710 5810
rect 10140 5690 10260 5810
rect 10690 5690 10810 5810
rect 11240 5690 11360 5810
rect 11790 5690 11910 5810
rect 12340 5690 12460 5810
rect 12890 5690 13010 5810
rect 13440 5690 13560 5810
rect 14075 5538 14175 5638
rect -925 5312 -825 5412
rect -310 5140 -190 5260
rect 240 5140 360 5260
rect 790 5140 910 5260
rect 1340 5140 1460 5260
rect 1890 5140 2010 5260
rect 2440 5140 2560 5260
rect 2990 5140 3110 5260
rect 3540 5140 3660 5260
rect 4090 5140 4210 5260
rect 4640 5140 4760 5260
rect 5190 5140 5310 5260
rect 5740 5140 5860 5260
rect 6290 5140 6410 5260
rect 6840 5140 6960 5260
rect 7390 5140 7510 5260
rect 7940 5140 8060 5260
rect 8490 5140 8610 5260
rect 9040 5140 9160 5260
rect 9590 5140 9710 5260
rect 10140 5140 10260 5260
rect 10690 5140 10810 5260
rect 11240 5140 11360 5260
rect 11790 5140 11910 5260
rect 12340 5140 12460 5260
rect 12890 5140 13010 5260
rect 13440 5140 13560 5260
rect -310 4590 -190 4710
rect 240 4590 360 4710
rect 790 4590 910 4710
rect 1340 4590 1460 4710
rect 1890 4590 2010 4710
rect 2440 4590 2560 4710
rect 2990 4590 3110 4710
rect 3540 4590 3660 4710
rect 4090 4590 4210 4710
rect 4640 4590 4760 4710
rect 5190 4590 5310 4710
rect 5740 4590 5860 4710
rect 6290 4590 6410 4710
rect 6840 4590 6960 4710
rect 7390 4590 7510 4710
rect 7940 4590 8060 4710
rect 8490 4590 8610 4710
rect 9040 4590 9160 4710
rect 9590 4590 9710 4710
rect 10140 4590 10260 4710
rect 10690 4590 10810 4710
rect 11240 4590 11360 4710
rect 11790 4590 11910 4710
rect 12340 4590 12460 4710
rect 12890 4590 13010 4710
rect 13440 4590 13560 4710
rect 14075 4438 14175 4538
rect -925 4212 -825 4312
rect -310 4040 -190 4160
rect 240 4040 360 4160
rect 790 4040 910 4160
rect 1340 4040 1460 4160
rect 1890 4040 2010 4160
rect 2440 4040 2560 4160
rect 2990 4040 3110 4160
rect 3540 4040 3660 4160
rect 4090 4040 4210 4160
rect 4640 4040 4760 4160
rect 5190 4040 5310 4160
rect 5740 4040 5860 4160
rect 6290 4040 6410 4160
rect 6840 4040 6960 4160
rect 7390 4040 7510 4160
rect 7940 4040 8060 4160
rect 8490 4040 8610 4160
rect 9040 4040 9160 4160
rect 9590 4040 9710 4160
rect 10140 4040 10260 4160
rect 10690 4040 10810 4160
rect 11240 4040 11360 4160
rect 11790 4040 11910 4160
rect 12340 4040 12460 4160
rect 12890 4040 13010 4160
rect 13440 4040 13560 4160
rect -310 3490 -190 3610
rect 240 3490 360 3610
rect 790 3490 910 3610
rect 1340 3490 1460 3610
rect 1890 3490 2010 3610
rect 2440 3490 2560 3610
rect 2990 3490 3110 3610
rect 3540 3490 3660 3610
rect 4090 3490 4210 3610
rect 4640 3490 4760 3610
rect 5190 3490 5310 3610
rect 5740 3490 5860 3610
rect 6290 3490 6410 3610
rect 6840 3490 6960 3610
rect 7390 3490 7510 3610
rect 7940 3490 8060 3610
rect 8490 3490 8610 3610
rect 9040 3490 9160 3610
rect 9590 3490 9710 3610
rect 10140 3490 10260 3610
rect 10690 3490 10810 3610
rect 11240 3490 11360 3610
rect 11790 3490 11910 3610
rect 12340 3490 12460 3610
rect 12890 3490 13010 3610
rect 13440 3490 13560 3610
rect 14075 3338 14175 3438
rect -925 3112 -825 3212
rect -310 2940 -190 3060
rect 240 2940 360 3060
rect 790 2940 910 3060
rect 1340 2940 1460 3060
rect 1890 2940 2010 3060
rect 2440 2940 2560 3060
rect 2990 2940 3110 3060
rect 3540 2940 3660 3060
rect 4090 2940 4210 3060
rect 4640 2940 4760 3060
rect 5190 2940 5310 3060
rect 5740 2940 5860 3060
rect 6290 2940 6410 3060
rect 6840 2940 6960 3060
rect 7390 2940 7510 3060
rect 7940 2940 8060 3060
rect 8490 2940 8610 3060
rect 9040 2940 9160 3060
rect 9590 2940 9710 3060
rect 10140 2940 10260 3060
rect 10690 2940 10810 3060
rect 11240 2940 11360 3060
rect 11790 2940 11910 3060
rect 12340 2940 12460 3060
rect 12890 2940 13010 3060
rect 13440 2940 13560 3060
rect -310 2390 -190 2510
rect 240 2390 360 2510
rect 790 2390 910 2510
rect 1340 2390 1460 2510
rect 1890 2390 2010 2510
rect 2440 2390 2560 2510
rect 2990 2390 3110 2510
rect 3540 2390 3660 2510
rect 4090 2390 4210 2510
rect 4640 2390 4760 2510
rect 5190 2390 5310 2510
rect 5740 2390 5860 2510
rect 6290 2390 6410 2510
rect 6840 2390 6960 2510
rect 7390 2390 7510 2510
rect 7940 2390 8060 2510
rect 8490 2390 8610 2510
rect 9040 2390 9160 2510
rect 9590 2390 9710 2510
rect 10140 2390 10260 2510
rect 10690 2390 10810 2510
rect 11240 2390 11360 2510
rect 11790 2390 11910 2510
rect 12340 2390 12460 2510
rect 12890 2390 13010 2510
rect 13440 2390 13560 2510
rect 14075 2238 14175 2338
rect -925 2012 -825 2112
rect -310 1840 -190 1960
rect 240 1840 360 1960
rect 790 1840 910 1960
rect 1340 1840 1460 1960
rect 1890 1840 2010 1960
rect 2440 1840 2560 1960
rect 2990 1840 3110 1960
rect 3540 1840 3660 1960
rect 4090 1840 4210 1960
rect 4640 1840 4760 1960
rect 5190 1840 5310 1960
rect 5740 1840 5860 1960
rect 6290 1840 6410 1960
rect 6840 1840 6960 1960
rect 7390 1840 7510 1960
rect 7940 1840 8060 1960
rect 8490 1840 8610 1960
rect 9040 1840 9160 1960
rect 9590 1840 9710 1960
rect 10140 1840 10260 1960
rect 10690 1840 10810 1960
rect 11240 1840 11360 1960
rect 11790 1840 11910 1960
rect 12340 1840 12460 1960
rect 12890 1840 13010 1960
rect 13440 1840 13560 1960
rect -310 1290 -190 1410
rect 240 1290 360 1410
rect 790 1290 910 1410
rect 1340 1290 1460 1410
rect 1890 1290 2010 1410
rect 2440 1290 2560 1410
rect 2990 1290 3110 1410
rect 3540 1290 3660 1410
rect 4090 1290 4210 1410
rect 4640 1290 4760 1410
rect 5190 1290 5310 1410
rect 5740 1290 5860 1410
rect 6290 1290 6410 1410
rect 6840 1290 6960 1410
rect 7390 1290 7510 1410
rect 7940 1290 8060 1410
rect 8490 1290 8610 1410
rect 9040 1290 9160 1410
rect 9590 1290 9710 1410
rect 10140 1290 10260 1410
rect 10690 1290 10810 1410
rect 11240 1290 11360 1410
rect 11790 1290 11910 1410
rect 12340 1290 12460 1410
rect 12890 1290 13010 1410
rect 13440 1290 13560 1410
rect 14075 1138 14175 1238
rect -925 912 -825 1012
rect -310 740 -190 860
rect 240 740 360 860
rect 790 740 910 860
rect 1340 740 1460 860
rect 1890 740 2010 860
rect 2440 740 2560 860
rect 2990 740 3110 860
rect 3540 740 3660 860
rect 4090 740 4210 860
rect 4640 740 4760 860
rect 5190 740 5310 860
rect 5740 740 5860 860
rect 6290 740 6410 860
rect 6840 740 6960 860
rect 7390 740 7510 860
rect 7940 740 8060 860
rect 8490 740 8610 860
rect 9040 740 9160 860
rect 9590 740 9710 860
rect 10140 740 10260 860
rect 10690 740 10810 860
rect 11240 740 11360 860
rect 11790 740 11910 860
rect 12340 740 12460 860
rect 12890 740 13010 860
rect 13440 740 13560 860
rect -310 190 -190 310
rect 240 190 360 310
rect 790 190 910 310
rect 1340 190 1460 310
rect 1890 190 2010 310
rect 2440 190 2560 310
rect 2990 190 3110 310
rect 3540 190 3660 310
rect 4090 190 4210 310
rect 4640 190 4760 310
rect 5190 190 5310 310
rect 5740 190 5860 310
rect 6290 190 6410 310
rect 6840 190 6960 310
rect 7390 190 7510 310
rect 7940 190 8060 310
rect 8490 190 8610 310
rect 9040 190 9160 310
rect 9590 190 9710 310
rect 10140 190 10260 310
rect 10690 190 10810 310
rect 11240 190 11360 310
rect 11790 190 11910 310
rect 12340 190 12460 310
rect 12890 190 13010 310
rect 13440 190 13560 310
rect -925 -188 -825 -88
rect 14075 38 14175 138
rect -310 -360 -190 -240
rect 240 -360 360 -240
rect 790 -360 910 -240
rect 1340 -360 1460 -240
rect 1890 -360 2010 -240
rect 2440 -360 2560 -240
rect 2990 -360 3110 -240
rect 3540 -360 3660 -240
rect 4090 -360 4210 -240
rect 4640 -360 4760 -240
rect 5190 -360 5310 -240
rect 5740 -360 5860 -240
rect 6290 -360 6410 -240
rect 6840 -360 6960 -240
rect 7390 -360 7510 -240
rect 7940 -360 8060 -240
rect 8490 -360 8610 -240
rect 9040 -360 9160 -240
rect 9590 -360 9710 -240
rect 10140 -360 10260 -240
rect 10690 -360 10810 -240
rect 11240 -360 11360 -240
rect 11790 -360 11910 -240
rect 12340 -360 12460 -240
rect 12890 -360 13010 -240
rect 13440 -360 13560 -240
rect -138 -975 -38 -875
rect 962 -975 1062 -875
rect 2062 -975 2162 -875
rect 3162 -975 3262 -875
rect 4262 -975 4362 -875
rect 5362 -975 5462 -875
rect 6462 -975 6562 -875
rect 7562 -975 7662 -875
rect 8662 -975 8762 -875
rect 9762 -975 9862 -875
rect 10862 -975 10962 -875
rect 11962 -975 12062 -875
rect 13062 -975 13162 -875
<< metal4 >>
rect -2525 14725 13775 15725
rect -2525 13838 -1525 14725
rect -638 13838 -186 14725
rect -2525 13514 -186 13838
rect -88 14125 364 14225
rect -88 14025 88 14125
rect 188 14025 364 14125
rect -88 13612 364 14025
rect 462 13612 914 14725
rect 1012 14125 1464 14225
rect 1012 14025 1188 14125
rect 1288 14025 1464 14125
rect 1012 13612 1464 14025
rect 1562 13612 2014 14725
rect 2112 14125 2564 14225
rect 2112 14025 2288 14125
rect 2388 14025 2564 14125
rect 2112 13612 2564 14025
rect 2662 13612 3114 14725
rect 3212 14125 3664 14225
rect 3212 14025 3388 14125
rect 3488 14025 3664 14125
rect 3212 13612 3664 14025
rect 3762 13612 4214 14725
rect 4312 14125 4764 14225
rect 4312 14025 4488 14125
rect 4588 14025 4764 14125
rect 4312 13612 4764 14025
rect 4862 13612 5314 14725
rect 5412 14125 5864 14225
rect 5412 14025 5588 14125
rect 5688 14025 5864 14125
rect 5412 13612 5864 14025
rect 5962 13612 6414 14725
rect 6512 14125 6964 14225
rect 6512 14025 6688 14125
rect 6788 14025 6964 14125
rect 6512 13612 6964 14025
rect 7062 13612 7514 14725
rect 7612 14125 8064 14225
rect 7612 14025 7788 14125
rect 7888 14025 8064 14125
rect 7612 13612 8064 14025
rect 8162 13612 8614 14725
rect 8712 14125 9164 14225
rect 8712 14025 8888 14125
rect 8988 14025 9164 14125
rect 8712 13612 9164 14025
rect 9262 13612 9714 14725
rect 9812 14125 10264 14225
rect 9812 14025 9988 14125
rect 10088 14025 10264 14125
rect 9812 13612 10264 14025
rect 10362 13612 10814 14725
rect 10912 14125 11364 14225
rect 10912 14025 11088 14125
rect 11188 14025 11364 14125
rect 10912 13612 11364 14025
rect 11462 13612 11914 14725
rect 12012 14125 12464 14225
rect 12012 14025 12188 14125
rect 12288 14025 12464 14125
rect 12012 13612 12464 14025
rect 12562 13612 13014 14725
rect 13112 14125 13564 14225
rect 13112 14025 13288 14125
rect 13388 14025 13564 14125
rect 13112 13612 13564 14025
tri -186 13514 -88 13612 sw
tri -88 13514 10 13612 ne
rect 10 13514 364 13612
tri 364 13514 462 13612 sw
tri 462 13514 560 13612 ne
rect 560 13514 914 13612
tri 914 13514 1012 13612 sw
tri 1012 13514 1110 13612 ne
rect 1110 13514 1464 13612
tri 1464 13514 1562 13612 sw
tri 1562 13514 1660 13612 ne
rect 1660 13514 2014 13612
tri 2014 13514 2112 13612 sw
tri 2112 13514 2210 13612 ne
rect 2210 13514 2564 13612
tri 2564 13514 2662 13612 sw
tri 2662 13514 2760 13612 ne
rect 2760 13514 3114 13612
tri 3114 13514 3212 13612 sw
tri 3212 13514 3310 13612 ne
rect 3310 13514 3664 13612
tri 3664 13514 3762 13612 sw
tri 3762 13514 3860 13612 ne
rect 3860 13514 4214 13612
tri 4214 13514 4312 13612 sw
tri 4312 13514 4410 13612 ne
rect 4410 13514 4764 13612
tri 4764 13514 4862 13612 sw
tri 4862 13514 4960 13612 ne
rect 4960 13514 5314 13612
tri 5314 13514 5412 13612 sw
tri 5412 13514 5510 13612 ne
rect 5510 13514 5864 13612
tri 5864 13514 5962 13612 sw
tri 5962 13514 6060 13612 ne
rect 6060 13514 6414 13612
tri 6414 13514 6512 13612 sw
tri 6512 13514 6610 13612 ne
rect 6610 13514 6964 13612
tri 6964 13514 7062 13612 sw
tri 7062 13514 7160 13612 ne
rect 7160 13514 7514 13612
tri 7514 13514 7612 13612 sw
tri 7612 13514 7710 13612 ne
rect 7710 13514 8064 13612
tri 8064 13514 8162 13612 sw
tri 8162 13514 8260 13612 ne
rect 8260 13514 8614 13612
tri 8614 13514 8712 13612 sw
tri 8712 13514 8810 13612 ne
rect 8810 13514 9164 13612
tri 9164 13514 9262 13612 sw
tri 9262 13514 9360 13612 ne
rect 9360 13514 9714 13612
tri 9714 13514 9812 13612 sw
tri 9812 13514 9910 13612 ne
rect 9910 13514 10264 13612
tri 10264 13514 10362 13612 sw
tri 10362 13514 10460 13612 ne
rect 10460 13514 10814 13612
tri 10814 13514 10912 13612 sw
tri 10912 13514 11010 13612 ne
rect 11010 13514 11364 13612
tri 11364 13514 11462 13612 sw
tri 11462 13514 11560 13612 ne
rect 11560 13514 11914 13612
tri 11914 13514 12012 13612 sw
tri 12012 13514 12110 13612 ne
rect 12110 13514 12464 13612
tri 12464 13514 12562 13612 sw
tri 12562 13514 12660 13612 ne
rect 12660 13514 13014 13612
tri 13014 13514 13112 13612 sw
tri 13112 13514 13210 13612 ne
rect 13210 13514 13564 13612
tri 13564 13514 13662 13612 sw
rect 14775 13514 15775 13725
rect -2525 13510 -88 13514
rect -2525 13390 -310 13510
rect -190 13426 -88 13510
tri -88 13426 0 13514 sw
tri 10 13426 98 13514 ne
rect 98 13510 462 13514
rect 98 13426 240 13510
rect -190 13390 0 13426
rect -2525 13386 0 13390
tri 0 13386 40 13426 sw
tri 98 13386 138 13426 ne
rect 138 13390 240 13426
rect 360 13426 462 13510
tri 462 13426 550 13514 sw
tri 560 13426 648 13514 ne
rect 648 13510 1012 13514
rect 648 13426 790 13510
rect 360 13390 550 13426
rect 138 13386 550 13390
tri 550 13386 590 13426 sw
tri 648 13386 688 13426 ne
rect 688 13390 790 13426
rect 910 13426 1012 13510
tri 1012 13426 1100 13514 sw
tri 1110 13426 1198 13514 ne
rect 1198 13510 1562 13514
rect 1198 13426 1340 13510
rect 910 13390 1100 13426
rect 688 13386 1100 13390
tri 1100 13386 1140 13426 sw
tri 1198 13386 1238 13426 ne
rect 1238 13390 1340 13426
rect 1460 13426 1562 13510
tri 1562 13426 1650 13514 sw
tri 1660 13426 1748 13514 ne
rect 1748 13510 2112 13514
rect 1748 13426 1890 13510
rect 1460 13390 1650 13426
rect 1238 13386 1650 13390
tri 1650 13386 1690 13426 sw
tri 1748 13386 1788 13426 ne
rect 1788 13390 1890 13426
rect 2010 13426 2112 13510
tri 2112 13426 2200 13514 sw
tri 2210 13426 2298 13514 ne
rect 2298 13510 2662 13514
rect 2298 13426 2440 13510
rect 2010 13390 2200 13426
rect 1788 13386 2200 13390
tri 2200 13386 2240 13426 sw
tri 2298 13386 2338 13426 ne
rect 2338 13390 2440 13426
rect 2560 13426 2662 13510
tri 2662 13426 2750 13514 sw
tri 2760 13426 2848 13514 ne
rect 2848 13510 3212 13514
rect 2848 13426 2990 13510
rect 2560 13390 2750 13426
rect 2338 13386 2750 13390
tri 2750 13386 2790 13426 sw
tri 2848 13386 2888 13426 ne
rect 2888 13390 2990 13426
rect 3110 13426 3212 13510
tri 3212 13426 3300 13514 sw
tri 3310 13426 3398 13514 ne
rect 3398 13510 3762 13514
rect 3398 13426 3540 13510
rect 3110 13390 3300 13426
rect 2888 13386 3300 13390
tri 3300 13386 3340 13426 sw
tri 3398 13386 3438 13426 ne
rect 3438 13390 3540 13426
rect 3660 13426 3762 13510
tri 3762 13426 3850 13514 sw
tri 3860 13426 3948 13514 ne
rect 3948 13510 4312 13514
rect 3948 13426 4090 13510
rect 3660 13390 3850 13426
rect 3438 13386 3850 13390
tri 3850 13386 3890 13426 sw
tri 3948 13386 3988 13426 ne
rect 3988 13390 4090 13426
rect 4210 13426 4312 13510
tri 4312 13426 4400 13514 sw
tri 4410 13426 4498 13514 ne
rect 4498 13510 4862 13514
rect 4498 13426 4640 13510
rect 4210 13390 4400 13426
rect 3988 13386 4400 13390
tri 4400 13386 4440 13426 sw
tri 4498 13386 4538 13426 ne
rect 4538 13390 4640 13426
rect 4760 13426 4862 13510
tri 4862 13426 4950 13514 sw
tri 4960 13426 5048 13514 ne
rect 5048 13510 5412 13514
rect 5048 13426 5190 13510
rect 4760 13390 4950 13426
rect 4538 13386 4950 13390
tri 4950 13386 4990 13426 sw
tri 5048 13386 5088 13426 ne
rect 5088 13390 5190 13426
rect 5310 13426 5412 13510
tri 5412 13426 5500 13514 sw
tri 5510 13426 5598 13514 ne
rect 5598 13510 5962 13514
rect 5598 13426 5740 13510
rect 5310 13390 5500 13426
rect 5088 13386 5500 13390
tri 5500 13386 5540 13426 sw
tri 5598 13386 5638 13426 ne
rect 5638 13390 5740 13426
rect 5860 13426 5962 13510
tri 5962 13426 6050 13514 sw
tri 6060 13426 6148 13514 ne
rect 6148 13510 6512 13514
rect 6148 13426 6290 13510
rect 5860 13390 6050 13426
rect 5638 13386 6050 13390
tri 6050 13386 6090 13426 sw
tri 6148 13386 6188 13426 ne
rect 6188 13390 6290 13426
rect 6410 13426 6512 13510
tri 6512 13426 6600 13514 sw
tri 6610 13426 6698 13514 ne
rect 6698 13510 7062 13514
rect 6698 13426 6840 13510
rect 6410 13390 6600 13426
rect 6188 13386 6600 13390
tri 6600 13386 6640 13426 sw
tri 6698 13386 6738 13426 ne
rect 6738 13390 6840 13426
rect 6960 13426 7062 13510
tri 7062 13426 7150 13514 sw
tri 7160 13426 7248 13514 ne
rect 7248 13510 7612 13514
rect 7248 13426 7390 13510
rect 6960 13390 7150 13426
rect 6738 13386 7150 13390
tri 7150 13386 7190 13426 sw
tri 7248 13386 7288 13426 ne
rect 7288 13390 7390 13426
rect 7510 13426 7612 13510
tri 7612 13426 7700 13514 sw
tri 7710 13426 7798 13514 ne
rect 7798 13510 8162 13514
rect 7798 13426 7940 13510
rect 7510 13390 7700 13426
rect 7288 13386 7700 13390
tri 7700 13386 7740 13426 sw
tri 7798 13386 7838 13426 ne
rect 7838 13390 7940 13426
rect 8060 13426 8162 13510
tri 8162 13426 8250 13514 sw
tri 8260 13426 8348 13514 ne
rect 8348 13510 8712 13514
rect 8348 13426 8490 13510
rect 8060 13390 8250 13426
rect 7838 13386 8250 13390
tri 8250 13386 8290 13426 sw
tri 8348 13386 8388 13426 ne
rect 8388 13390 8490 13426
rect 8610 13426 8712 13510
tri 8712 13426 8800 13514 sw
tri 8810 13426 8898 13514 ne
rect 8898 13510 9262 13514
rect 8898 13426 9040 13510
rect 8610 13390 8800 13426
rect 8388 13386 8800 13390
tri 8800 13386 8840 13426 sw
tri 8898 13386 8938 13426 ne
rect 8938 13390 9040 13426
rect 9160 13426 9262 13510
tri 9262 13426 9350 13514 sw
tri 9360 13426 9448 13514 ne
rect 9448 13510 9812 13514
rect 9448 13426 9590 13510
rect 9160 13390 9350 13426
rect 8938 13386 9350 13390
tri 9350 13386 9390 13426 sw
tri 9448 13386 9488 13426 ne
rect 9488 13390 9590 13426
rect 9710 13426 9812 13510
tri 9812 13426 9900 13514 sw
tri 9910 13426 9998 13514 ne
rect 9998 13510 10362 13514
rect 9998 13426 10140 13510
rect 9710 13390 9900 13426
rect 9488 13386 9900 13390
tri 9900 13386 9940 13426 sw
tri 9998 13386 10038 13426 ne
rect 10038 13390 10140 13426
rect 10260 13426 10362 13510
tri 10362 13426 10450 13514 sw
tri 10460 13426 10548 13514 ne
rect 10548 13510 10912 13514
rect 10548 13426 10690 13510
rect 10260 13390 10450 13426
rect 10038 13386 10450 13390
tri 10450 13386 10490 13426 sw
tri 10548 13386 10588 13426 ne
rect 10588 13390 10690 13426
rect 10810 13426 10912 13510
tri 10912 13426 11000 13514 sw
tri 11010 13426 11098 13514 ne
rect 11098 13510 11462 13514
rect 11098 13426 11240 13510
rect 10810 13390 11000 13426
rect 10588 13386 11000 13390
tri 11000 13386 11040 13426 sw
tri 11098 13386 11138 13426 ne
rect 11138 13390 11240 13426
rect 11360 13426 11462 13510
tri 11462 13426 11550 13514 sw
tri 11560 13426 11648 13514 ne
rect 11648 13510 12012 13514
rect 11648 13426 11790 13510
rect 11360 13390 11550 13426
rect 11138 13386 11550 13390
tri 11550 13386 11590 13426 sw
tri 11648 13386 11688 13426 ne
rect 11688 13390 11790 13426
rect 11910 13426 12012 13510
tri 12012 13426 12100 13514 sw
tri 12110 13426 12198 13514 ne
rect 12198 13510 12562 13514
rect 12198 13426 12340 13510
rect 11910 13390 12100 13426
rect 11688 13386 12100 13390
tri 12100 13386 12140 13426 sw
tri 12198 13386 12238 13426 ne
rect 12238 13390 12340 13426
rect 12460 13426 12562 13510
tri 12562 13426 12650 13514 sw
tri 12660 13426 12748 13514 ne
rect 12748 13510 13112 13514
rect 12748 13426 12890 13510
rect 12460 13390 12650 13426
rect 12238 13386 12650 13390
tri 12650 13386 12690 13426 sw
tri 12748 13386 12788 13426 ne
rect 12788 13390 12890 13426
rect 13010 13426 13112 13510
tri 13112 13426 13200 13514 sw
tri 13210 13426 13298 13514 ne
rect 13298 13510 15775 13514
rect 13298 13426 13440 13510
rect 13010 13390 13200 13426
rect 12788 13386 13200 13390
rect -2525 12738 -1525 13386
tri -412 13288 -314 13386 ne
rect -314 13288 40 13386
tri 40 13288 138 13386 sw
tri 138 13288 236 13386 ne
rect 236 13288 590 13386
tri 590 13288 688 13386 sw
tri 688 13288 786 13386 ne
rect 786 13288 1140 13386
tri 1140 13288 1238 13386 sw
tri 1238 13288 1336 13386 ne
rect 1336 13288 1690 13386
tri 1690 13288 1788 13386 sw
tri 1788 13288 1886 13386 ne
rect 1886 13288 2240 13386
tri 2240 13288 2338 13386 sw
tri 2338 13288 2436 13386 ne
rect 2436 13288 2790 13386
tri 2790 13288 2888 13386 sw
tri 2888 13288 2986 13386 ne
rect 2986 13288 3340 13386
tri 3340 13288 3438 13386 sw
tri 3438 13288 3536 13386 ne
rect 3536 13288 3890 13386
tri 3890 13288 3988 13386 sw
tri 3988 13288 4086 13386 ne
rect 4086 13288 4440 13386
tri 4440 13288 4538 13386 sw
tri 4538 13288 4636 13386 ne
rect 4636 13288 4990 13386
tri 4990 13288 5088 13386 sw
tri 5088 13288 5186 13386 ne
rect 5186 13288 5540 13386
tri 5540 13288 5638 13386 sw
tri 5638 13288 5736 13386 ne
rect 5736 13288 6090 13386
tri 6090 13288 6188 13386 sw
tri 6188 13288 6286 13386 ne
rect 6286 13288 6640 13386
tri 6640 13288 6738 13386 sw
tri 6738 13288 6836 13386 ne
rect 6836 13288 7190 13386
tri 7190 13288 7288 13386 sw
tri 7288 13288 7386 13386 ne
rect 7386 13288 7740 13386
tri 7740 13288 7838 13386 sw
tri 7838 13288 7936 13386 ne
rect 7936 13288 8290 13386
tri 8290 13288 8388 13386 sw
tri 8388 13288 8486 13386 ne
rect 8486 13288 8840 13386
tri 8840 13288 8938 13386 sw
tri 8938 13288 9036 13386 ne
rect 9036 13288 9390 13386
tri 9390 13288 9488 13386 sw
tri 9488 13288 9586 13386 ne
rect 9586 13288 9940 13386
tri 9940 13288 10038 13386 sw
tri 10038 13288 10136 13386 ne
rect 10136 13288 10490 13386
tri 10490 13288 10588 13386 sw
tri 10588 13288 10686 13386 ne
rect 10686 13288 11040 13386
tri 11040 13288 11138 13386 sw
tri 11138 13288 11236 13386 ne
rect 11236 13288 11590 13386
tri 11590 13288 11688 13386 sw
tri 11688 13288 11786 13386 ne
rect 11786 13288 12140 13386
tri 12140 13288 12238 13386 sw
tri 12238 13288 12336 13386 ne
rect 12336 13288 12690 13386
tri 12690 13288 12788 13386 sw
tri 12788 13288 12886 13386 ne
rect 12886 13338 13200 13386
tri 13200 13338 13288 13426 sw
tri 13298 13338 13386 13426 ne
rect 13386 13390 13440 13426
rect 13560 13390 15775 13510
rect 13386 13338 15775 13390
rect 12886 13288 13288 13338
rect -1025 13200 -412 13288
tri -412 13200 -324 13288 sw
tri -314 13200 -226 13288 ne
rect -226 13200 138 13288
tri 138 13200 226 13288 sw
tri 236 13200 324 13288 ne
rect 324 13200 688 13288
tri 688 13200 776 13288 sw
tri 786 13200 874 13288 ne
rect 874 13200 1238 13288
tri 1238 13200 1326 13288 sw
tri 1336 13200 1424 13288 ne
rect 1424 13200 1788 13288
tri 1788 13200 1876 13288 sw
tri 1886 13200 1974 13288 ne
rect 1974 13200 2338 13288
tri 2338 13200 2426 13288 sw
tri 2436 13200 2524 13288 ne
rect 2524 13200 2888 13288
tri 2888 13200 2976 13288 sw
tri 2986 13200 3074 13288 ne
rect 3074 13200 3438 13288
tri 3438 13200 3526 13288 sw
tri 3536 13200 3624 13288 ne
rect 3624 13200 3988 13288
tri 3988 13200 4076 13288 sw
tri 4086 13200 4174 13288 ne
rect 4174 13200 4538 13288
tri 4538 13200 4626 13288 sw
tri 4636 13200 4724 13288 ne
rect 4724 13200 5088 13288
tri 5088 13200 5176 13288 sw
tri 5186 13200 5274 13288 ne
rect 5274 13200 5638 13288
tri 5638 13200 5726 13288 sw
tri 5736 13200 5824 13288 ne
rect 5824 13200 6188 13288
tri 6188 13200 6276 13288 sw
tri 6286 13200 6374 13288 ne
rect 6374 13200 6738 13288
tri 6738 13200 6826 13288 sw
tri 6836 13200 6924 13288 ne
rect 6924 13200 7288 13288
tri 7288 13200 7376 13288 sw
tri 7386 13200 7474 13288 ne
rect 7474 13200 7838 13288
tri 7838 13200 7926 13288 sw
tri 7936 13200 8024 13288 ne
rect 8024 13200 8388 13288
tri 8388 13200 8476 13288 sw
tri 8486 13200 8574 13288 ne
rect 8574 13200 8938 13288
tri 8938 13200 9026 13288 sw
tri 9036 13200 9124 13288 ne
rect 9124 13200 9488 13288
tri 9488 13200 9576 13288 sw
tri 9586 13200 9674 13288 ne
rect 9674 13200 10038 13288
tri 10038 13200 10126 13288 sw
tri 10136 13200 10224 13288 ne
rect 10224 13200 10588 13288
tri 10588 13200 10676 13288 sw
tri 10686 13200 10774 13288 ne
rect 10774 13200 11138 13288
tri 11138 13200 11226 13288 sw
tri 11236 13200 11324 13288 ne
rect 11324 13200 11688 13288
tri 11688 13200 11776 13288 sw
tri 11786 13200 11874 13288 ne
rect 11874 13200 12238 13288
tri 12238 13200 12326 13288 sw
tri 12336 13200 12424 13288 ne
rect 12424 13200 12788 13288
tri 12788 13200 12876 13288 sw
tri 12886 13200 12974 13288 ne
rect 12974 13258 13288 13288
tri 13288 13258 13368 13338 sw
tri 13386 13258 13466 13338 ne
rect 13466 13258 14075 13338
rect 12974 13200 13368 13258
rect -1025 13160 -324 13200
tri -324 13160 -284 13200 sw
tri -226 13160 -186 13200 ne
rect -186 13160 226 13200
tri 226 13160 266 13200 sw
tri 324 13160 364 13200 ne
rect 364 13160 776 13200
tri 776 13160 816 13200 sw
tri 874 13160 914 13200 ne
rect 914 13160 1326 13200
tri 1326 13160 1366 13200 sw
tri 1424 13160 1464 13200 ne
rect 1464 13160 1876 13200
tri 1876 13160 1916 13200 sw
tri 1974 13160 2014 13200 ne
rect 2014 13160 2426 13200
tri 2426 13160 2466 13200 sw
tri 2524 13160 2564 13200 ne
rect 2564 13160 2976 13200
tri 2976 13160 3016 13200 sw
tri 3074 13160 3114 13200 ne
rect 3114 13160 3526 13200
tri 3526 13160 3566 13200 sw
tri 3624 13160 3664 13200 ne
rect 3664 13160 4076 13200
tri 4076 13160 4116 13200 sw
tri 4174 13160 4214 13200 ne
rect 4214 13160 4626 13200
tri 4626 13160 4666 13200 sw
tri 4724 13160 4764 13200 ne
rect 4764 13160 5176 13200
tri 5176 13160 5216 13200 sw
tri 5274 13160 5314 13200 ne
rect 5314 13160 5726 13200
tri 5726 13160 5766 13200 sw
tri 5824 13160 5864 13200 ne
rect 5864 13160 6276 13200
tri 6276 13160 6316 13200 sw
tri 6374 13160 6414 13200 ne
rect 6414 13160 6826 13200
tri 6826 13160 6866 13200 sw
tri 6924 13160 6964 13200 ne
rect 6964 13160 7376 13200
tri 7376 13160 7416 13200 sw
tri 7474 13160 7514 13200 ne
rect 7514 13160 7926 13200
tri 7926 13160 7966 13200 sw
tri 8024 13160 8064 13200 ne
rect 8064 13160 8476 13200
tri 8476 13160 8516 13200 sw
tri 8574 13160 8614 13200 ne
rect 8614 13160 9026 13200
tri 9026 13160 9066 13200 sw
tri 9124 13160 9164 13200 ne
rect 9164 13160 9576 13200
tri 9576 13160 9616 13200 sw
tri 9674 13160 9714 13200 ne
rect 9714 13160 10126 13200
tri 10126 13160 10166 13200 sw
tri 10224 13160 10264 13200 ne
rect 10264 13160 10676 13200
tri 10676 13160 10716 13200 sw
tri 10774 13160 10814 13200 ne
rect 10814 13160 11226 13200
tri 11226 13160 11266 13200 sw
tri 11324 13160 11364 13200 ne
rect 11364 13160 11776 13200
tri 11776 13160 11816 13200 sw
tri 11874 13160 11914 13200 ne
rect 11914 13160 12326 13200
tri 12326 13160 12366 13200 sw
tri 12424 13160 12464 13200 ne
rect 12464 13160 12876 13200
tri 12876 13160 12916 13200 sw
tri 12974 13160 13014 13200 ne
rect 13014 13160 13368 13200
tri 13368 13160 13466 13258 sw
tri 13466 13160 13564 13258 ne
rect 13564 13238 14075 13258
rect 14175 13238 15775 13338
rect 13564 13160 15775 13238
rect -1025 13112 -284 13160
rect -1025 13012 -925 13112
rect -825 13062 -284 13112
tri -284 13062 -186 13160 sw
tri -186 13062 -88 13160 ne
rect -88 13062 266 13160
tri 266 13062 364 13160 sw
tri 364 13062 462 13160 ne
rect 462 13062 816 13160
tri 816 13062 914 13160 sw
tri 914 13062 1012 13160 ne
rect 1012 13062 1366 13160
tri 1366 13062 1464 13160 sw
tri 1464 13062 1562 13160 ne
rect 1562 13062 1916 13160
tri 1916 13062 2014 13160 sw
tri 2014 13062 2112 13160 ne
rect 2112 13062 2466 13160
tri 2466 13062 2564 13160 sw
tri 2564 13062 2662 13160 ne
rect 2662 13062 3016 13160
tri 3016 13062 3114 13160 sw
tri 3114 13062 3212 13160 ne
rect 3212 13062 3566 13160
tri 3566 13062 3664 13160 sw
tri 3664 13062 3762 13160 ne
rect 3762 13062 4116 13160
tri 4116 13062 4214 13160 sw
tri 4214 13062 4312 13160 ne
rect 4312 13062 4666 13160
tri 4666 13062 4764 13160 sw
tri 4764 13062 4862 13160 ne
rect 4862 13062 5216 13160
tri 5216 13062 5314 13160 sw
tri 5314 13062 5412 13160 ne
rect 5412 13062 5766 13160
tri 5766 13062 5864 13160 sw
tri 5864 13062 5962 13160 ne
rect 5962 13062 6316 13160
tri 6316 13062 6414 13160 sw
tri 6414 13062 6512 13160 ne
rect 6512 13062 6866 13160
tri 6866 13062 6964 13160 sw
tri 6964 13062 7062 13160 ne
rect 7062 13062 7416 13160
tri 7416 13062 7514 13160 sw
tri 7514 13062 7612 13160 ne
rect 7612 13062 7966 13160
tri 7966 13062 8064 13160 sw
tri 8064 13062 8162 13160 ne
rect 8162 13062 8516 13160
tri 8516 13062 8614 13160 sw
tri 8614 13062 8712 13160 ne
rect 8712 13062 9066 13160
tri 9066 13062 9164 13160 sw
tri 9164 13062 9262 13160 ne
rect 9262 13062 9616 13160
tri 9616 13062 9714 13160 sw
tri 9714 13062 9812 13160 ne
rect 9812 13062 10166 13160
tri 10166 13062 10264 13160 sw
tri 10264 13062 10362 13160 ne
rect 10362 13062 10716 13160
tri 10716 13062 10814 13160 sw
tri 10814 13062 10912 13160 ne
rect 10912 13062 11266 13160
tri 11266 13062 11364 13160 sw
tri 11364 13062 11462 13160 ne
rect 11462 13062 11816 13160
tri 11816 13062 11914 13160 sw
tri 11914 13062 12012 13160 ne
rect 12012 13062 12366 13160
tri 12366 13062 12464 13160 sw
tri 12464 13062 12562 13160 ne
rect 12562 13062 12916 13160
tri 12916 13062 13014 13160 sw
tri 13014 13062 13112 13160 ne
rect 13112 13062 13466 13160
tri 13466 13062 13564 13160 sw
tri 13564 13062 13662 13160 ne
rect 13662 13062 15775 13160
rect -825 13012 -186 13062
rect -1025 12964 -186 13012
tri -186 12964 -88 13062 sw
tri -88 12964 10 13062 ne
rect 10 12964 364 13062
tri 364 12964 462 13062 sw
tri 462 12964 560 13062 ne
rect 560 12964 914 13062
tri 914 12964 1012 13062 sw
tri 1012 12964 1110 13062 ne
rect 1110 12964 1464 13062
tri 1464 12964 1562 13062 sw
tri 1562 12964 1660 13062 ne
rect 1660 12964 2014 13062
tri 2014 12964 2112 13062 sw
tri 2112 12964 2210 13062 ne
rect 2210 12964 2564 13062
tri 2564 12964 2662 13062 sw
tri 2662 12964 2760 13062 ne
rect 2760 12964 3114 13062
tri 3114 12964 3212 13062 sw
tri 3212 12964 3310 13062 ne
rect 3310 12964 3664 13062
tri 3664 12964 3762 13062 sw
tri 3762 12964 3860 13062 ne
rect 3860 12964 4214 13062
tri 4214 12964 4312 13062 sw
tri 4312 12964 4410 13062 ne
rect 4410 12964 4764 13062
tri 4764 12964 4862 13062 sw
tri 4862 12964 4960 13062 ne
rect 4960 12964 5314 13062
tri 5314 12964 5412 13062 sw
tri 5412 12964 5510 13062 ne
rect 5510 12964 5864 13062
tri 5864 12964 5962 13062 sw
tri 5962 12964 6060 13062 ne
rect 6060 12964 6414 13062
tri 6414 12964 6512 13062 sw
tri 6512 12964 6610 13062 ne
rect 6610 12964 6964 13062
tri 6964 12964 7062 13062 sw
tri 7062 12964 7160 13062 ne
rect 7160 12964 7514 13062
tri 7514 12964 7612 13062 sw
tri 7612 12964 7710 13062 ne
rect 7710 12964 8064 13062
tri 8064 12964 8162 13062 sw
tri 8162 12964 8260 13062 ne
rect 8260 12964 8614 13062
tri 8614 12964 8712 13062 sw
tri 8712 12964 8810 13062 ne
rect 8810 12964 9164 13062
tri 9164 12964 9262 13062 sw
tri 9262 12964 9360 13062 ne
rect 9360 12964 9714 13062
tri 9714 12964 9812 13062 sw
tri 9812 12964 9910 13062 ne
rect 9910 12964 10264 13062
tri 10264 12964 10362 13062 sw
tri 10362 12964 10460 13062 ne
rect 10460 12964 10814 13062
tri 10814 12964 10912 13062 sw
tri 10912 12964 11010 13062 ne
rect 11010 12964 11364 13062
tri 11364 12964 11462 13062 sw
tri 11462 12964 11560 13062 ne
rect 11560 12964 11914 13062
tri 11914 12964 12012 13062 sw
tri 12012 12964 12110 13062 ne
rect 12110 12964 12464 13062
tri 12464 12964 12562 13062 sw
tri 12562 12964 12660 13062 ne
rect 12660 12964 13014 13062
tri 13014 12964 13112 13062 sw
tri 13112 12964 13210 13062 ne
rect 13210 12964 13564 13062
tri 13564 12964 13662 13062 sw
rect -1025 12960 -88 12964
rect -1025 12840 -310 12960
rect -190 12876 -88 12960
tri -88 12876 0 12964 sw
tri 10 12876 98 12964 ne
rect 98 12960 462 12964
rect 98 12876 240 12960
rect -190 12840 0 12876
rect -1025 12836 0 12840
tri 0 12836 40 12876 sw
tri 98 12836 138 12876 ne
rect 138 12840 240 12876
rect 360 12876 462 12960
tri 462 12876 550 12964 sw
tri 560 12876 648 12964 ne
rect 648 12960 1012 12964
rect 648 12876 790 12960
rect 360 12840 550 12876
rect 138 12836 550 12840
tri -412 12738 -314 12836 ne
rect -314 12738 40 12836
tri 40 12738 138 12836 sw
tri 138 12738 236 12836 ne
rect 236 12788 550 12836
tri 550 12788 638 12876 sw
tri 648 12788 736 12876 ne
rect 736 12840 790 12876
rect 910 12876 1012 12960
tri 1012 12876 1100 12964 sw
tri 1110 12876 1198 12964 ne
rect 1198 12960 1562 12964
rect 1198 12876 1340 12960
rect 910 12840 1100 12876
rect 736 12836 1100 12840
tri 1100 12836 1140 12876 sw
tri 1198 12836 1238 12876 ne
rect 1238 12840 1340 12876
rect 1460 12876 1562 12960
tri 1562 12876 1650 12964 sw
tri 1660 12876 1748 12964 ne
rect 1748 12960 2112 12964
rect 1748 12876 1890 12960
rect 1460 12840 1650 12876
rect 1238 12836 1650 12840
rect 736 12788 1140 12836
rect 236 12738 638 12788
rect -2525 12650 -412 12738
tri -412 12650 -324 12738 sw
tri -314 12650 -226 12738 ne
rect -226 12650 138 12738
tri 138 12650 226 12738 sw
tri 236 12650 324 12738 ne
rect 324 12708 638 12738
tri 638 12708 718 12788 sw
tri 736 12708 816 12788 ne
rect 816 12738 1140 12788
tri 1140 12738 1238 12836 sw
tri 1238 12738 1336 12836 ne
rect 1336 12788 1650 12836
tri 1650 12788 1738 12876 sw
tri 1748 12788 1836 12876 ne
rect 1836 12840 1890 12876
rect 2010 12876 2112 12960
tri 2112 12876 2200 12964 sw
tri 2210 12876 2298 12964 ne
rect 2298 12960 2662 12964
rect 2298 12876 2440 12960
rect 2010 12840 2200 12876
rect 1836 12836 2200 12840
tri 2200 12836 2240 12876 sw
tri 2298 12836 2338 12876 ne
rect 2338 12840 2440 12876
rect 2560 12876 2662 12960
tri 2662 12876 2750 12964 sw
tri 2760 12876 2848 12964 ne
rect 2848 12960 3212 12964
rect 2848 12876 2990 12960
rect 2560 12840 2750 12876
rect 2338 12836 2750 12840
rect 1836 12788 2240 12836
rect 1336 12738 1738 12788
rect 816 12708 1238 12738
rect 324 12650 718 12708
rect -2525 12610 -324 12650
tri -324 12610 -284 12650 sw
tri -226 12610 -186 12650 ne
rect -186 12610 226 12650
tri 226 12610 266 12650 sw
tri 324 12610 364 12650 ne
rect 364 12610 718 12650
tri 718 12610 816 12708 sw
tri 816 12610 914 12708 ne
rect 914 12650 1238 12708
tri 1238 12650 1326 12738 sw
tri 1336 12650 1424 12738 ne
rect 1424 12708 1738 12738
tri 1738 12708 1818 12788 sw
tri 1836 12708 1916 12788 ne
rect 1916 12738 2240 12788
tri 2240 12738 2338 12836 sw
tri 2338 12738 2436 12836 ne
rect 2436 12788 2750 12836
tri 2750 12788 2838 12876 sw
tri 2848 12788 2936 12876 ne
rect 2936 12840 2990 12876
rect 3110 12876 3212 12960
tri 3212 12876 3300 12964 sw
tri 3310 12876 3398 12964 ne
rect 3398 12960 3762 12964
rect 3398 12876 3540 12960
rect 3110 12840 3300 12876
rect 2936 12836 3300 12840
tri 3300 12836 3340 12876 sw
tri 3398 12836 3438 12876 ne
rect 3438 12840 3540 12876
rect 3660 12876 3762 12960
tri 3762 12876 3850 12964 sw
tri 3860 12876 3948 12964 ne
rect 3948 12960 4312 12964
rect 3948 12876 4090 12960
rect 3660 12840 3850 12876
rect 3438 12836 3850 12840
rect 2936 12788 3340 12836
rect 2436 12738 2838 12788
rect 1916 12708 2338 12738
rect 1424 12650 1818 12708
rect 914 12610 1326 12650
tri 1326 12610 1366 12650 sw
tri 1424 12610 1464 12650 ne
rect 1464 12610 1818 12650
tri 1818 12610 1916 12708 sw
tri 1916 12610 2014 12708 ne
rect 2014 12650 2338 12708
tri 2338 12650 2426 12738 sw
tri 2436 12650 2524 12738 ne
rect 2524 12708 2838 12738
tri 2838 12708 2918 12788 sw
tri 2936 12708 3016 12788 ne
rect 3016 12738 3340 12788
tri 3340 12738 3438 12836 sw
tri 3438 12738 3536 12836 ne
rect 3536 12788 3850 12836
tri 3850 12788 3938 12876 sw
tri 3948 12788 4036 12876 ne
rect 4036 12840 4090 12876
rect 4210 12876 4312 12960
tri 4312 12876 4400 12964 sw
tri 4410 12876 4498 12964 ne
rect 4498 12960 4862 12964
rect 4498 12876 4640 12960
rect 4210 12840 4400 12876
rect 4036 12836 4400 12840
tri 4400 12836 4440 12876 sw
tri 4498 12836 4538 12876 ne
rect 4538 12840 4640 12876
rect 4760 12876 4862 12960
tri 4862 12876 4950 12964 sw
tri 4960 12876 5048 12964 ne
rect 5048 12960 5412 12964
rect 5048 12876 5190 12960
rect 4760 12840 4950 12876
rect 4538 12836 4950 12840
rect 4036 12788 4440 12836
rect 3536 12738 3938 12788
rect 3016 12708 3438 12738
rect 2524 12650 2918 12708
rect 2014 12610 2426 12650
tri 2426 12610 2466 12650 sw
tri 2524 12610 2564 12650 ne
rect 2564 12610 2918 12650
tri 2918 12610 3016 12708 sw
tri 3016 12610 3114 12708 ne
rect 3114 12650 3438 12708
tri 3438 12650 3526 12738 sw
tri 3536 12650 3624 12738 ne
rect 3624 12708 3938 12738
tri 3938 12708 4018 12788 sw
tri 4036 12708 4116 12788 ne
rect 4116 12738 4440 12788
tri 4440 12738 4538 12836 sw
tri 4538 12738 4636 12836 ne
rect 4636 12788 4950 12836
tri 4950 12788 5038 12876 sw
tri 5048 12788 5136 12876 ne
rect 5136 12840 5190 12876
rect 5310 12876 5412 12960
tri 5412 12876 5500 12964 sw
tri 5510 12876 5598 12964 ne
rect 5598 12960 5962 12964
rect 5598 12876 5740 12960
rect 5310 12840 5500 12876
rect 5136 12836 5500 12840
tri 5500 12836 5540 12876 sw
tri 5598 12836 5638 12876 ne
rect 5638 12840 5740 12876
rect 5860 12876 5962 12960
tri 5962 12876 6050 12964 sw
tri 6060 12876 6148 12964 ne
rect 6148 12960 6512 12964
rect 6148 12876 6290 12960
rect 5860 12840 6050 12876
rect 5638 12836 6050 12840
rect 5136 12788 5540 12836
rect 4636 12738 5038 12788
rect 4116 12708 4538 12738
rect 3624 12650 4018 12708
rect 3114 12610 3526 12650
tri 3526 12610 3566 12650 sw
tri 3624 12610 3664 12650 ne
rect 3664 12610 4018 12650
tri 4018 12610 4116 12708 sw
tri 4116 12610 4214 12708 ne
rect 4214 12650 4538 12708
tri 4538 12650 4626 12738 sw
tri 4636 12650 4724 12738 ne
rect 4724 12708 5038 12738
tri 5038 12708 5118 12788 sw
tri 5136 12708 5216 12788 ne
rect 5216 12738 5540 12788
tri 5540 12738 5638 12836 sw
tri 5638 12738 5736 12836 ne
rect 5736 12788 6050 12836
tri 6050 12788 6138 12876 sw
tri 6148 12788 6236 12876 ne
rect 6236 12840 6290 12876
rect 6410 12876 6512 12960
tri 6512 12876 6600 12964 sw
tri 6610 12876 6698 12964 ne
rect 6698 12960 7062 12964
rect 6698 12876 6840 12960
rect 6410 12840 6600 12876
rect 6236 12836 6600 12840
tri 6600 12836 6640 12876 sw
tri 6698 12836 6738 12876 ne
rect 6738 12840 6840 12876
rect 6960 12876 7062 12960
tri 7062 12876 7150 12964 sw
tri 7160 12876 7248 12964 ne
rect 7248 12960 7612 12964
rect 7248 12876 7390 12960
rect 6960 12840 7150 12876
rect 6738 12836 7150 12840
rect 6236 12788 6640 12836
rect 5736 12738 6138 12788
rect 5216 12708 5638 12738
rect 4724 12650 5118 12708
rect 4214 12610 4626 12650
tri 4626 12610 4666 12650 sw
tri 4724 12610 4764 12650 ne
rect 4764 12610 5118 12650
tri 5118 12610 5216 12708 sw
tri 5216 12610 5314 12708 ne
rect 5314 12650 5638 12708
tri 5638 12650 5726 12738 sw
tri 5736 12650 5824 12738 ne
rect 5824 12708 6138 12738
tri 6138 12708 6218 12788 sw
tri 6236 12708 6316 12788 ne
rect 6316 12738 6640 12788
tri 6640 12738 6738 12836 sw
tri 6738 12738 6836 12836 ne
rect 6836 12788 7150 12836
tri 7150 12788 7238 12876 sw
tri 7248 12788 7336 12876 ne
rect 7336 12840 7390 12876
rect 7510 12876 7612 12960
tri 7612 12876 7700 12964 sw
tri 7710 12876 7798 12964 ne
rect 7798 12960 8162 12964
rect 7798 12876 7940 12960
rect 7510 12840 7700 12876
rect 7336 12836 7700 12840
tri 7700 12836 7740 12876 sw
tri 7798 12836 7838 12876 ne
rect 7838 12840 7940 12876
rect 8060 12876 8162 12960
tri 8162 12876 8250 12964 sw
tri 8260 12876 8348 12964 ne
rect 8348 12960 8712 12964
rect 8348 12876 8490 12960
rect 8060 12840 8250 12876
rect 7838 12836 8250 12840
rect 7336 12788 7740 12836
rect 6836 12738 7238 12788
rect 6316 12708 6738 12738
rect 5824 12650 6218 12708
rect 5314 12610 5726 12650
tri 5726 12610 5766 12650 sw
tri 5824 12610 5864 12650 ne
rect 5864 12610 6218 12650
tri 6218 12610 6316 12708 sw
tri 6316 12610 6414 12708 ne
rect 6414 12650 6738 12708
tri 6738 12650 6826 12738 sw
tri 6836 12650 6924 12738 ne
rect 6924 12708 7238 12738
tri 7238 12708 7318 12788 sw
tri 7336 12708 7416 12788 ne
rect 7416 12738 7740 12788
tri 7740 12738 7838 12836 sw
tri 7838 12738 7936 12836 ne
rect 7936 12788 8250 12836
tri 8250 12788 8338 12876 sw
tri 8348 12788 8436 12876 ne
rect 8436 12840 8490 12876
rect 8610 12876 8712 12960
tri 8712 12876 8800 12964 sw
tri 8810 12876 8898 12964 ne
rect 8898 12960 9262 12964
rect 8898 12876 9040 12960
rect 8610 12840 8800 12876
rect 8436 12836 8800 12840
tri 8800 12836 8840 12876 sw
tri 8898 12836 8938 12876 ne
rect 8938 12840 9040 12876
rect 9160 12876 9262 12960
tri 9262 12876 9350 12964 sw
tri 9360 12876 9448 12964 ne
rect 9448 12960 9812 12964
rect 9448 12876 9590 12960
rect 9160 12840 9350 12876
rect 8938 12836 9350 12840
rect 8436 12788 8840 12836
rect 7936 12738 8338 12788
rect 7416 12708 7838 12738
rect 6924 12650 7318 12708
rect 6414 12610 6826 12650
tri 6826 12610 6866 12650 sw
tri 6924 12610 6964 12650 ne
rect 6964 12610 7318 12650
tri 7318 12610 7416 12708 sw
tri 7416 12610 7514 12708 ne
rect 7514 12650 7838 12708
tri 7838 12650 7926 12738 sw
tri 7936 12650 8024 12738 ne
rect 8024 12708 8338 12738
tri 8338 12708 8418 12788 sw
tri 8436 12708 8516 12788 ne
rect 8516 12738 8840 12788
tri 8840 12738 8938 12836 sw
tri 8938 12738 9036 12836 ne
rect 9036 12788 9350 12836
tri 9350 12788 9438 12876 sw
tri 9448 12788 9536 12876 ne
rect 9536 12840 9590 12876
rect 9710 12876 9812 12960
tri 9812 12876 9900 12964 sw
tri 9910 12876 9998 12964 ne
rect 9998 12960 10362 12964
rect 9998 12876 10140 12960
rect 9710 12840 9900 12876
rect 9536 12836 9900 12840
tri 9900 12836 9940 12876 sw
tri 9998 12836 10038 12876 ne
rect 10038 12840 10140 12876
rect 10260 12876 10362 12960
tri 10362 12876 10450 12964 sw
tri 10460 12876 10548 12964 ne
rect 10548 12960 10912 12964
rect 10548 12876 10690 12960
rect 10260 12840 10450 12876
rect 10038 12836 10450 12840
rect 9536 12788 9940 12836
rect 9036 12738 9438 12788
rect 8516 12708 8938 12738
rect 8024 12650 8418 12708
rect 7514 12610 7926 12650
tri 7926 12610 7966 12650 sw
tri 8024 12610 8064 12650 ne
rect 8064 12610 8418 12650
tri 8418 12610 8516 12708 sw
tri 8516 12610 8614 12708 ne
rect 8614 12650 8938 12708
tri 8938 12650 9026 12738 sw
tri 9036 12650 9124 12738 ne
rect 9124 12708 9438 12738
tri 9438 12708 9518 12788 sw
tri 9536 12708 9616 12788 ne
rect 9616 12738 9940 12788
tri 9940 12738 10038 12836 sw
tri 10038 12738 10136 12836 ne
rect 10136 12788 10450 12836
tri 10450 12788 10538 12876 sw
tri 10548 12788 10636 12876 ne
rect 10636 12840 10690 12876
rect 10810 12876 10912 12960
tri 10912 12876 11000 12964 sw
tri 11010 12876 11098 12964 ne
rect 11098 12960 11462 12964
rect 11098 12876 11240 12960
rect 10810 12840 11000 12876
rect 10636 12836 11000 12840
tri 11000 12836 11040 12876 sw
tri 11098 12836 11138 12876 ne
rect 11138 12840 11240 12876
rect 11360 12876 11462 12960
tri 11462 12876 11550 12964 sw
tri 11560 12876 11648 12964 ne
rect 11648 12960 12012 12964
rect 11648 12876 11790 12960
rect 11360 12840 11550 12876
rect 11138 12836 11550 12840
rect 10636 12788 11040 12836
rect 10136 12738 10538 12788
rect 9616 12708 10038 12738
rect 9124 12650 9518 12708
rect 8614 12610 9026 12650
tri 9026 12610 9066 12650 sw
tri 9124 12610 9164 12650 ne
rect 9164 12610 9518 12650
tri 9518 12610 9616 12708 sw
tri 9616 12610 9714 12708 ne
rect 9714 12650 10038 12708
tri 10038 12650 10126 12738 sw
tri 10136 12650 10224 12738 ne
rect 10224 12708 10538 12738
tri 10538 12708 10618 12788 sw
tri 10636 12708 10716 12788 ne
rect 10716 12738 11040 12788
tri 11040 12738 11138 12836 sw
tri 11138 12738 11236 12836 ne
rect 11236 12788 11550 12836
tri 11550 12788 11638 12876 sw
tri 11648 12788 11736 12876 ne
rect 11736 12840 11790 12876
rect 11910 12876 12012 12960
tri 12012 12876 12100 12964 sw
tri 12110 12876 12198 12964 ne
rect 12198 12960 12562 12964
rect 12198 12876 12340 12960
rect 11910 12840 12100 12876
rect 11736 12836 12100 12840
tri 12100 12836 12140 12876 sw
tri 12198 12836 12238 12876 ne
rect 12238 12840 12340 12876
rect 12460 12876 12562 12960
tri 12562 12876 12650 12964 sw
tri 12660 12876 12748 12964 ne
rect 12748 12960 13112 12964
rect 12748 12876 12890 12960
rect 12460 12840 12650 12876
rect 12238 12836 12650 12840
rect 11736 12788 12140 12836
rect 11236 12738 11638 12788
rect 10716 12708 11138 12738
rect 10224 12650 10618 12708
rect 9714 12610 10126 12650
tri 10126 12610 10166 12650 sw
tri 10224 12610 10264 12650 ne
rect 10264 12610 10618 12650
tri 10618 12610 10716 12708 sw
tri 10716 12610 10814 12708 ne
rect 10814 12650 11138 12708
tri 11138 12650 11226 12738 sw
tri 11236 12650 11324 12738 ne
rect 11324 12708 11638 12738
tri 11638 12708 11718 12788 sw
tri 11736 12708 11816 12788 ne
rect 11816 12738 12140 12788
tri 12140 12738 12238 12836 sw
tri 12238 12738 12336 12836 ne
rect 12336 12788 12650 12836
tri 12650 12788 12738 12876 sw
tri 12748 12788 12836 12876 ne
rect 12836 12840 12890 12876
rect 13010 12876 13112 12960
tri 13112 12876 13200 12964 sw
tri 13210 12876 13298 12964 ne
rect 13298 12960 14275 12964
rect 13298 12876 13440 12960
rect 13010 12840 13200 12876
rect 12836 12836 13200 12840
tri 13200 12836 13240 12876 sw
tri 13298 12836 13338 12876 ne
rect 13338 12840 13440 12876
rect 13560 12840 14275 12960
rect 13338 12836 14275 12840
rect 12836 12788 13240 12836
rect 12336 12738 12738 12788
rect 11816 12708 12238 12738
rect 11324 12650 11718 12708
rect 10814 12610 11226 12650
tri 11226 12610 11266 12650 sw
tri 11324 12610 11364 12650 ne
rect 11364 12610 11718 12650
tri 11718 12610 11816 12708 sw
tri 11816 12610 11914 12708 ne
rect 11914 12650 12238 12708
tri 12238 12650 12326 12738 sw
tri 12336 12650 12424 12738 ne
rect 12424 12708 12738 12738
tri 12738 12708 12818 12788 sw
tri 12836 12708 12916 12788 ne
rect 12916 12738 13240 12788
tri 13240 12738 13338 12836 sw
tri 13338 12738 13436 12836 ne
rect 13436 12738 14275 12836
rect 12916 12708 13338 12738
rect 12424 12650 12818 12708
rect 11914 12610 12326 12650
tri 12326 12610 12366 12650 sw
tri 12424 12610 12464 12650 ne
rect 12464 12610 12818 12650
tri 12818 12610 12916 12708 sw
tri 12916 12610 13014 12708 ne
rect 13014 12650 13338 12708
tri 13338 12650 13426 12738 sw
tri 13436 12650 13524 12738 ne
rect 13524 12650 14275 12738
rect 13014 12610 13426 12650
tri 13426 12610 13466 12650 sw
tri 13524 12610 13564 12650 ne
rect 13564 12610 14275 12650
rect -2525 12512 -284 12610
tri -284 12512 -186 12610 sw
tri -186 12512 -88 12610 ne
rect -88 12512 266 12610
tri 266 12512 364 12610 sw
tri 364 12512 462 12610 ne
rect 462 12512 816 12610
tri 816 12512 914 12610 sw
tri 914 12512 1012 12610 ne
rect 1012 12512 1366 12610
tri 1366 12512 1464 12610 sw
tri 1464 12512 1562 12610 ne
rect 1562 12512 1916 12610
tri 1916 12512 2014 12610 sw
tri 2014 12512 2112 12610 ne
rect 2112 12512 2466 12610
tri 2466 12512 2564 12610 sw
tri 2564 12512 2662 12610 ne
rect 2662 12512 3016 12610
tri 3016 12512 3114 12610 sw
tri 3114 12512 3212 12610 ne
rect 3212 12512 3566 12610
tri 3566 12512 3664 12610 sw
tri 3664 12512 3762 12610 ne
rect 3762 12512 4116 12610
tri 4116 12512 4214 12610 sw
tri 4214 12512 4312 12610 ne
rect 4312 12512 4666 12610
tri 4666 12512 4764 12610 sw
tri 4764 12512 4862 12610 ne
rect 4862 12512 5216 12610
tri 5216 12512 5314 12610 sw
tri 5314 12512 5412 12610 ne
rect 5412 12512 5766 12610
tri 5766 12512 5864 12610 sw
tri 5864 12512 5962 12610 ne
rect 5962 12512 6316 12610
tri 6316 12512 6414 12610 sw
tri 6414 12512 6512 12610 ne
rect 6512 12512 6866 12610
tri 6866 12512 6964 12610 sw
tri 6964 12512 7062 12610 ne
rect 7062 12512 7416 12610
tri 7416 12512 7514 12610 sw
tri 7514 12512 7612 12610 ne
rect 7612 12512 7966 12610
tri 7966 12512 8064 12610 sw
tri 8064 12512 8162 12610 ne
rect 8162 12512 8516 12610
tri 8516 12512 8614 12610 sw
tri 8614 12512 8712 12610 ne
rect 8712 12512 9066 12610
tri 9066 12512 9164 12610 sw
tri 9164 12512 9262 12610 ne
rect 9262 12512 9616 12610
tri 9616 12512 9714 12610 sw
tri 9714 12512 9812 12610 ne
rect 9812 12512 10166 12610
tri 10166 12512 10264 12610 sw
tri 10264 12512 10362 12610 ne
rect 10362 12512 10716 12610
tri 10716 12512 10814 12610 sw
tri 10814 12512 10912 12610 ne
rect 10912 12512 11266 12610
tri 11266 12512 11364 12610 sw
tri 11364 12512 11462 12610 ne
rect 11462 12512 11816 12610
tri 11816 12512 11914 12610 sw
tri 11914 12512 12012 12610 ne
rect 12012 12512 12366 12610
tri 12366 12512 12464 12610 sw
tri 12464 12512 12562 12610 ne
rect 12562 12512 12916 12610
tri 12916 12512 13014 12610 sw
tri 13014 12512 13112 12610 ne
rect 13112 12512 13466 12610
tri 13466 12512 13564 12610 sw
tri 13564 12512 13662 12610 ne
rect 13662 12512 14275 12610
rect -2525 12414 -186 12512
tri -186 12414 -88 12512 sw
tri -88 12414 10 12512 ne
rect 10 12414 364 12512
tri 364 12414 462 12512 sw
tri 462 12414 560 12512 ne
rect 560 12414 914 12512
tri 914 12414 1012 12512 sw
tri 1012 12414 1110 12512 ne
rect 1110 12414 1464 12512
tri 1464 12414 1562 12512 sw
tri 1562 12414 1660 12512 ne
rect 1660 12414 2014 12512
tri 2014 12414 2112 12512 sw
tri 2112 12414 2210 12512 ne
rect 2210 12414 2564 12512
tri 2564 12414 2662 12512 sw
tri 2662 12414 2760 12512 ne
rect 2760 12414 3114 12512
tri 3114 12414 3212 12512 sw
tri 3212 12414 3310 12512 ne
rect 3310 12414 3664 12512
tri 3664 12414 3762 12512 sw
tri 3762 12414 3860 12512 ne
rect 3860 12414 4214 12512
tri 4214 12414 4312 12512 sw
tri 4312 12414 4410 12512 ne
rect 4410 12414 4764 12512
tri 4764 12414 4862 12512 sw
tri 4862 12414 4960 12512 ne
rect 4960 12414 5314 12512
tri 5314 12414 5412 12512 sw
tri 5412 12414 5510 12512 ne
rect 5510 12414 5864 12512
tri 5864 12414 5962 12512 sw
tri 5962 12414 6060 12512 ne
rect 6060 12414 6414 12512
tri 6414 12414 6512 12512 sw
tri 6512 12414 6610 12512 ne
rect 6610 12414 6964 12512
tri 6964 12414 7062 12512 sw
tri 7062 12414 7160 12512 ne
rect 7160 12414 7514 12512
tri 7514 12414 7612 12512 sw
tri 7612 12414 7710 12512 ne
rect 7710 12414 8064 12512
tri 8064 12414 8162 12512 sw
tri 8162 12414 8260 12512 ne
rect 8260 12414 8614 12512
tri 8614 12414 8712 12512 sw
tri 8712 12414 8810 12512 ne
rect 8810 12414 9164 12512
tri 9164 12414 9262 12512 sw
tri 9262 12414 9360 12512 ne
rect 9360 12414 9714 12512
tri 9714 12414 9812 12512 sw
tri 9812 12414 9910 12512 ne
rect 9910 12414 10264 12512
tri 10264 12414 10362 12512 sw
tri 10362 12414 10460 12512 ne
rect 10460 12414 10814 12512
tri 10814 12414 10912 12512 sw
tri 10912 12414 11010 12512 ne
rect 11010 12414 11364 12512
tri 11364 12414 11462 12512 sw
tri 11462 12414 11560 12512 ne
rect 11560 12414 11914 12512
tri 11914 12414 12012 12512 sw
tri 12012 12414 12110 12512 ne
rect 12110 12414 12464 12512
tri 12464 12414 12562 12512 sw
tri 12562 12414 12660 12512 ne
rect 12660 12414 13014 12512
tri 13014 12414 13112 12512 sw
tri 13112 12414 13210 12512 ne
rect 13210 12414 13564 12512
tri 13564 12414 13662 12512 sw
rect 14775 12414 15775 13062
rect -2525 12410 -88 12414
rect -2525 12290 -310 12410
rect -190 12326 -88 12410
tri -88 12326 0 12414 sw
tri 10 12326 98 12414 ne
rect 98 12410 462 12414
rect 98 12326 240 12410
rect -190 12290 0 12326
rect -2525 12286 0 12290
rect -2525 11638 -1525 12286
tri -412 12188 -314 12286 ne
rect -314 12238 0 12286
tri 0 12238 88 12326 sw
tri 98 12238 186 12326 ne
rect 186 12290 240 12326
rect 360 12326 462 12410
tri 462 12326 550 12414 sw
tri 560 12326 648 12414 ne
rect 648 12410 1012 12414
rect 648 12326 790 12410
rect 360 12290 550 12326
rect 186 12286 550 12290
tri 550 12286 590 12326 sw
tri 648 12286 688 12326 ne
rect 688 12290 790 12326
rect 910 12326 1012 12410
tri 1012 12326 1100 12414 sw
tri 1110 12326 1198 12414 ne
rect 1198 12410 1562 12414
rect 1198 12326 1340 12410
rect 910 12290 1100 12326
rect 688 12286 1100 12290
rect 186 12238 590 12286
rect -314 12188 88 12238
rect -1025 12100 -412 12188
tri -412 12100 -324 12188 sw
tri -314 12100 -226 12188 ne
rect -226 12158 88 12188
tri 88 12158 168 12238 sw
tri 186 12158 266 12238 ne
rect 266 12188 590 12238
tri 590 12188 688 12286 sw
tri 688 12188 786 12286 ne
rect 786 12238 1100 12286
tri 1100 12238 1188 12326 sw
tri 1198 12238 1286 12326 ne
rect 1286 12290 1340 12326
rect 1460 12326 1562 12410
tri 1562 12326 1650 12414 sw
tri 1660 12326 1748 12414 ne
rect 1748 12410 2112 12414
rect 1748 12326 1890 12410
rect 1460 12290 1650 12326
rect 1286 12286 1650 12290
tri 1650 12286 1690 12326 sw
tri 1748 12286 1788 12326 ne
rect 1788 12290 1890 12326
rect 2010 12326 2112 12410
tri 2112 12326 2200 12414 sw
tri 2210 12326 2298 12414 ne
rect 2298 12410 2662 12414
rect 2298 12326 2440 12410
rect 2010 12290 2200 12326
rect 1788 12286 2200 12290
rect 1286 12238 1690 12286
rect 786 12188 1188 12238
rect 266 12158 688 12188
rect -226 12100 168 12158
rect -1025 12060 -324 12100
tri -324 12060 -284 12100 sw
tri -226 12060 -186 12100 ne
rect -186 12060 168 12100
tri 168 12060 266 12158 sw
tri 266 12060 364 12158 ne
rect 364 12100 688 12158
tri 688 12100 776 12188 sw
tri 786 12100 874 12188 ne
rect 874 12158 1188 12188
tri 1188 12158 1268 12238 sw
tri 1286 12158 1366 12238 ne
rect 1366 12188 1690 12238
tri 1690 12188 1788 12286 sw
tri 1788 12188 1886 12286 ne
rect 1886 12238 2200 12286
tri 2200 12238 2288 12326 sw
tri 2298 12238 2386 12326 ne
rect 2386 12290 2440 12326
rect 2560 12326 2662 12410
tri 2662 12326 2750 12414 sw
tri 2760 12326 2848 12414 ne
rect 2848 12410 3212 12414
rect 2848 12326 2990 12410
rect 2560 12290 2750 12326
rect 2386 12286 2750 12290
tri 2750 12286 2790 12326 sw
tri 2848 12286 2888 12326 ne
rect 2888 12290 2990 12326
rect 3110 12326 3212 12410
tri 3212 12326 3300 12414 sw
tri 3310 12326 3398 12414 ne
rect 3398 12410 3762 12414
rect 3398 12326 3540 12410
rect 3110 12290 3300 12326
rect 2888 12286 3300 12290
rect 2386 12238 2790 12286
rect 1886 12188 2288 12238
rect 1366 12158 1788 12188
rect 874 12100 1268 12158
rect 364 12060 776 12100
tri 776 12060 816 12100 sw
tri 874 12060 914 12100 ne
rect 914 12060 1268 12100
tri 1268 12060 1366 12158 sw
tri 1366 12060 1464 12158 ne
rect 1464 12100 1788 12158
tri 1788 12100 1876 12188 sw
tri 1886 12100 1974 12188 ne
rect 1974 12158 2288 12188
tri 2288 12158 2368 12238 sw
tri 2386 12158 2466 12238 ne
rect 2466 12188 2790 12238
tri 2790 12188 2888 12286 sw
tri 2888 12188 2986 12286 ne
rect 2986 12238 3300 12286
tri 3300 12238 3388 12326 sw
tri 3398 12238 3486 12326 ne
rect 3486 12290 3540 12326
rect 3660 12326 3762 12410
tri 3762 12326 3850 12414 sw
tri 3860 12326 3948 12414 ne
rect 3948 12410 4312 12414
rect 3948 12326 4090 12410
rect 3660 12290 3850 12326
rect 3486 12286 3850 12290
tri 3850 12286 3890 12326 sw
tri 3948 12286 3988 12326 ne
rect 3988 12290 4090 12326
rect 4210 12326 4312 12410
tri 4312 12326 4400 12414 sw
tri 4410 12326 4498 12414 ne
rect 4498 12410 4862 12414
rect 4498 12326 4640 12410
rect 4210 12290 4400 12326
rect 3988 12286 4400 12290
rect 3486 12238 3890 12286
rect 2986 12188 3388 12238
rect 2466 12158 2888 12188
rect 1974 12100 2368 12158
rect 1464 12060 1876 12100
tri 1876 12060 1916 12100 sw
tri 1974 12060 2014 12100 ne
rect 2014 12060 2368 12100
tri 2368 12060 2466 12158 sw
tri 2466 12060 2564 12158 ne
rect 2564 12100 2888 12158
tri 2888 12100 2976 12188 sw
tri 2986 12100 3074 12188 ne
rect 3074 12158 3388 12188
tri 3388 12158 3468 12238 sw
tri 3486 12158 3566 12238 ne
rect 3566 12188 3890 12238
tri 3890 12188 3988 12286 sw
tri 3988 12188 4086 12286 ne
rect 4086 12238 4400 12286
tri 4400 12238 4488 12326 sw
tri 4498 12238 4586 12326 ne
rect 4586 12290 4640 12326
rect 4760 12326 4862 12410
tri 4862 12326 4950 12414 sw
tri 4960 12326 5048 12414 ne
rect 5048 12410 5412 12414
rect 5048 12326 5190 12410
rect 4760 12290 4950 12326
rect 4586 12286 4950 12290
tri 4950 12286 4990 12326 sw
tri 5048 12286 5088 12326 ne
rect 5088 12290 5190 12326
rect 5310 12326 5412 12410
tri 5412 12326 5500 12414 sw
tri 5510 12326 5598 12414 ne
rect 5598 12410 5962 12414
rect 5598 12326 5740 12410
rect 5310 12290 5500 12326
rect 5088 12286 5500 12290
rect 4586 12238 4990 12286
rect 4086 12188 4488 12238
rect 3566 12158 3988 12188
rect 3074 12100 3468 12158
rect 2564 12060 2976 12100
tri 2976 12060 3016 12100 sw
tri 3074 12060 3114 12100 ne
rect 3114 12060 3468 12100
tri 3468 12060 3566 12158 sw
tri 3566 12060 3664 12158 ne
rect 3664 12100 3988 12158
tri 3988 12100 4076 12188 sw
tri 4086 12100 4174 12188 ne
rect 4174 12158 4488 12188
tri 4488 12158 4568 12238 sw
tri 4586 12158 4666 12238 ne
rect 4666 12188 4990 12238
tri 4990 12188 5088 12286 sw
tri 5088 12188 5186 12286 ne
rect 5186 12238 5500 12286
tri 5500 12238 5588 12326 sw
tri 5598 12238 5686 12326 ne
rect 5686 12290 5740 12326
rect 5860 12326 5962 12410
tri 5962 12326 6050 12414 sw
tri 6060 12326 6148 12414 ne
rect 6148 12410 6512 12414
rect 6148 12326 6290 12410
rect 5860 12290 6050 12326
rect 5686 12286 6050 12290
tri 6050 12286 6090 12326 sw
tri 6148 12286 6188 12326 ne
rect 6188 12290 6290 12326
rect 6410 12326 6512 12410
tri 6512 12326 6600 12414 sw
tri 6610 12326 6698 12414 ne
rect 6698 12410 7062 12414
rect 6698 12326 6840 12410
rect 6410 12290 6600 12326
rect 6188 12286 6600 12290
rect 5686 12238 6090 12286
rect 5186 12188 5588 12238
rect 4666 12158 5088 12188
rect 4174 12100 4568 12158
rect 3664 12060 4076 12100
tri 4076 12060 4116 12100 sw
tri 4174 12060 4214 12100 ne
rect 4214 12060 4568 12100
tri 4568 12060 4666 12158 sw
tri 4666 12060 4764 12158 ne
rect 4764 12100 5088 12158
tri 5088 12100 5176 12188 sw
tri 5186 12100 5274 12188 ne
rect 5274 12158 5588 12188
tri 5588 12158 5668 12238 sw
tri 5686 12158 5766 12238 ne
rect 5766 12188 6090 12238
tri 6090 12188 6188 12286 sw
tri 6188 12188 6286 12286 ne
rect 6286 12238 6600 12286
tri 6600 12238 6688 12326 sw
tri 6698 12238 6786 12326 ne
rect 6786 12290 6840 12326
rect 6960 12326 7062 12410
tri 7062 12326 7150 12414 sw
tri 7160 12326 7248 12414 ne
rect 7248 12410 7612 12414
rect 7248 12326 7390 12410
rect 6960 12290 7150 12326
rect 6786 12286 7150 12290
tri 7150 12286 7190 12326 sw
tri 7248 12286 7288 12326 ne
rect 7288 12290 7390 12326
rect 7510 12326 7612 12410
tri 7612 12326 7700 12414 sw
tri 7710 12326 7798 12414 ne
rect 7798 12410 8162 12414
rect 7798 12326 7940 12410
rect 7510 12290 7700 12326
rect 7288 12286 7700 12290
rect 6786 12238 7190 12286
rect 6286 12188 6688 12238
rect 5766 12158 6188 12188
rect 5274 12100 5668 12158
rect 4764 12060 5176 12100
tri 5176 12060 5216 12100 sw
tri 5274 12060 5314 12100 ne
rect 5314 12060 5668 12100
tri 5668 12060 5766 12158 sw
tri 5766 12060 5864 12158 ne
rect 5864 12100 6188 12158
tri 6188 12100 6276 12188 sw
tri 6286 12100 6374 12188 ne
rect 6374 12158 6688 12188
tri 6688 12158 6768 12238 sw
tri 6786 12158 6866 12238 ne
rect 6866 12188 7190 12238
tri 7190 12188 7288 12286 sw
tri 7288 12188 7386 12286 ne
rect 7386 12238 7700 12286
tri 7700 12238 7788 12326 sw
tri 7798 12238 7886 12326 ne
rect 7886 12290 7940 12326
rect 8060 12326 8162 12410
tri 8162 12326 8250 12414 sw
tri 8260 12326 8348 12414 ne
rect 8348 12410 8712 12414
rect 8348 12326 8490 12410
rect 8060 12290 8250 12326
rect 7886 12286 8250 12290
tri 8250 12286 8290 12326 sw
tri 8348 12286 8388 12326 ne
rect 8388 12290 8490 12326
rect 8610 12326 8712 12410
tri 8712 12326 8800 12414 sw
tri 8810 12326 8898 12414 ne
rect 8898 12410 9262 12414
rect 8898 12326 9040 12410
rect 8610 12290 8800 12326
rect 8388 12286 8800 12290
rect 7886 12238 8290 12286
rect 7386 12188 7788 12238
rect 6866 12158 7288 12188
rect 6374 12100 6768 12158
rect 5864 12060 6276 12100
tri 6276 12060 6316 12100 sw
tri 6374 12060 6414 12100 ne
rect 6414 12060 6768 12100
tri 6768 12060 6866 12158 sw
tri 6866 12060 6964 12158 ne
rect 6964 12100 7288 12158
tri 7288 12100 7376 12188 sw
tri 7386 12100 7474 12188 ne
rect 7474 12158 7788 12188
tri 7788 12158 7868 12238 sw
tri 7886 12158 7966 12238 ne
rect 7966 12188 8290 12238
tri 8290 12188 8388 12286 sw
tri 8388 12188 8486 12286 ne
rect 8486 12238 8800 12286
tri 8800 12238 8888 12326 sw
tri 8898 12238 8986 12326 ne
rect 8986 12290 9040 12326
rect 9160 12326 9262 12410
tri 9262 12326 9350 12414 sw
tri 9360 12326 9448 12414 ne
rect 9448 12410 9812 12414
rect 9448 12326 9590 12410
rect 9160 12290 9350 12326
rect 8986 12286 9350 12290
tri 9350 12286 9390 12326 sw
tri 9448 12286 9488 12326 ne
rect 9488 12290 9590 12326
rect 9710 12326 9812 12410
tri 9812 12326 9900 12414 sw
tri 9910 12326 9998 12414 ne
rect 9998 12410 10362 12414
rect 9998 12326 10140 12410
rect 9710 12290 9900 12326
rect 9488 12286 9900 12290
rect 8986 12238 9390 12286
rect 8486 12188 8888 12238
rect 7966 12158 8388 12188
rect 7474 12100 7868 12158
rect 6964 12060 7376 12100
tri 7376 12060 7416 12100 sw
tri 7474 12060 7514 12100 ne
rect 7514 12060 7868 12100
tri 7868 12060 7966 12158 sw
tri 7966 12060 8064 12158 ne
rect 8064 12100 8388 12158
tri 8388 12100 8476 12188 sw
tri 8486 12100 8574 12188 ne
rect 8574 12158 8888 12188
tri 8888 12158 8968 12238 sw
tri 8986 12158 9066 12238 ne
rect 9066 12188 9390 12238
tri 9390 12188 9488 12286 sw
tri 9488 12188 9586 12286 ne
rect 9586 12238 9900 12286
tri 9900 12238 9988 12326 sw
tri 9998 12238 10086 12326 ne
rect 10086 12290 10140 12326
rect 10260 12326 10362 12410
tri 10362 12326 10450 12414 sw
tri 10460 12326 10548 12414 ne
rect 10548 12410 10912 12414
rect 10548 12326 10690 12410
rect 10260 12290 10450 12326
rect 10086 12286 10450 12290
tri 10450 12286 10490 12326 sw
tri 10548 12286 10588 12326 ne
rect 10588 12290 10690 12326
rect 10810 12326 10912 12410
tri 10912 12326 11000 12414 sw
tri 11010 12326 11098 12414 ne
rect 11098 12410 11462 12414
rect 11098 12326 11240 12410
rect 10810 12290 11000 12326
rect 10588 12286 11000 12290
rect 10086 12238 10490 12286
rect 9586 12188 9988 12238
rect 9066 12158 9488 12188
rect 8574 12100 8968 12158
rect 8064 12060 8476 12100
tri 8476 12060 8516 12100 sw
tri 8574 12060 8614 12100 ne
rect 8614 12060 8968 12100
tri 8968 12060 9066 12158 sw
tri 9066 12060 9164 12158 ne
rect 9164 12100 9488 12158
tri 9488 12100 9576 12188 sw
tri 9586 12100 9674 12188 ne
rect 9674 12158 9988 12188
tri 9988 12158 10068 12238 sw
tri 10086 12158 10166 12238 ne
rect 10166 12188 10490 12238
tri 10490 12188 10588 12286 sw
tri 10588 12188 10686 12286 ne
rect 10686 12238 11000 12286
tri 11000 12238 11088 12326 sw
tri 11098 12238 11186 12326 ne
rect 11186 12290 11240 12326
rect 11360 12326 11462 12410
tri 11462 12326 11550 12414 sw
tri 11560 12326 11648 12414 ne
rect 11648 12410 12012 12414
rect 11648 12326 11790 12410
rect 11360 12290 11550 12326
rect 11186 12286 11550 12290
tri 11550 12286 11590 12326 sw
tri 11648 12286 11688 12326 ne
rect 11688 12290 11790 12326
rect 11910 12326 12012 12410
tri 12012 12326 12100 12414 sw
tri 12110 12326 12198 12414 ne
rect 12198 12410 12562 12414
rect 12198 12326 12340 12410
rect 11910 12290 12100 12326
rect 11688 12286 12100 12290
rect 11186 12238 11590 12286
rect 10686 12188 11088 12238
rect 10166 12158 10588 12188
rect 9674 12100 10068 12158
rect 9164 12060 9576 12100
tri 9576 12060 9616 12100 sw
tri 9674 12060 9714 12100 ne
rect 9714 12060 10068 12100
tri 10068 12060 10166 12158 sw
tri 10166 12060 10264 12158 ne
rect 10264 12100 10588 12158
tri 10588 12100 10676 12188 sw
tri 10686 12100 10774 12188 ne
rect 10774 12158 11088 12188
tri 11088 12158 11168 12238 sw
tri 11186 12158 11266 12238 ne
rect 11266 12188 11590 12238
tri 11590 12188 11688 12286 sw
tri 11688 12188 11786 12286 ne
rect 11786 12238 12100 12286
tri 12100 12238 12188 12326 sw
tri 12198 12238 12286 12326 ne
rect 12286 12290 12340 12326
rect 12460 12326 12562 12410
tri 12562 12326 12650 12414 sw
tri 12660 12326 12748 12414 ne
rect 12748 12410 13112 12414
rect 12748 12326 12890 12410
rect 12460 12290 12650 12326
rect 12286 12286 12650 12290
tri 12650 12286 12690 12326 sw
tri 12748 12286 12788 12326 ne
rect 12788 12290 12890 12326
rect 13010 12326 13112 12410
tri 13112 12326 13200 12414 sw
tri 13210 12326 13298 12414 ne
rect 13298 12410 15775 12414
rect 13298 12326 13440 12410
rect 13010 12290 13200 12326
rect 12788 12286 13200 12290
rect 12286 12238 12690 12286
rect 11786 12188 12188 12238
rect 11266 12158 11688 12188
rect 10774 12100 11168 12158
rect 10264 12060 10676 12100
tri 10676 12060 10716 12100 sw
tri 10774 12060 10814 12100 ne
rect 10814 12060 11168 12100
tri 11168 12060 11266 12158 sw
tri 11266 12060 11364 12158 ne
rect 11364 12100 11688 12158
tri 11688 12100 11776 12188 sw
tri 11786 12100 11874 12188 ne
rect 11874 12158 12188 12188
tri 12188 12158 12268 12238 sw
tri 12286 12158 12366 12238 ne
rect 12366 12188 12690 12238
tri 12690 12188 12788 12286 sw
tri 12788 12188 12886 12286 ne
rect 12886 12238 13200 12286
tri 13200 12238 13288 12326 sw
tri 13298 12238 13386 12326 ne
rect 13386 12290 13440 12326
rect 13560 12290 15775 12410
rect 13386 12238 15775 12290
rect 12886 12188 13288 12238
rect 12366 12158 12788 12188
rect 11874 12100 12268 12158
rect 11364 12060 11776 12100
tri 11776 12060 11816 12100 sw
tri 11874 12060 11914 12100 ne
rect 11914 12060 12268 12100
tri 12268 12060 12366 12158 sw
tri 12366 12060 12464 12158 ne
rect 12464 12100 12788 12158
tri 12788 12100 12876 12188 sw
tri 12886 12100 12974 12188 ne
rect 12974 12158 13288 12188
tri 13288 12158 13368 12238 sw
tri 13386 12158 13466 12238 ne
rect 13466 12158 14075 12238
rect 12974 12100 13368 12158
rect 12464 12060 12876 12100
tri 12876 12060 12916 12100 sw
tri 12974 12060 13014 12100 ne
rect 13014 12060 13368 12100
tri 13368 12060 13466 12158 sw
tri 13466 12060 13564 12158 ne
rect 13564 12138 14075 12158
rect 14175 12138 15775 12238
rect 13564 12060 15775 12138
rect -1025 12012 -284 12060
rect -1025 11912 -925 12012
rect -825 11962 -284 12012
tri -284 11962 -186 12060 sw
tri -186 11962 -88 12060 ne
rect -88 11962 266 12060
tri 266 11962 364 12060 sw
tri 364 11962 462 12060 ne
rect 462 11962 816 12060
tri 816 11962 914 12060 sw
tri 914 11962 1012 12060 ne
rect 1012 11962 1366 12060
tri 1366 11962 1464 12060 sw
tri 1464 11962 1562 12060 ne
rect 1562 11962 1916 12060
tri 1916 11962 2014 12060 sw
tri 2014 11962 2112 12060 ne
rect 2112 11962 2466 12060
tri 2466 11962 2564 12060 sw
tri 2564 11962 2662 12060 ne
rect 2662 11962 3016 12060
tri 3016 11962 3114 12060 sw
tri 3114 11962 3212 12060 ne
rect 3212 11962 3566 12060
tri 3566 11962 3664 12060 sw
tri 3664 11962 3762 12060 ne
rect 3762 11962 4116 12060
tri 4116 11962 4214 12060 sw
tri 4214 11962 4312 12060 ne
rect 4312 11962 4666 12060
tri 4666 11962 4764 12060 sw
tri 4764 11962 4862 12060 ne
rect 4862 11962 5216 12060
tri 5216 11962 5314 12060 sw
tri 5314 11962 5412 12060 ne
rect 5412 11962 5766 12060
tri 5766 11962 5864 12060 sw
tri 5864 11962 5962 12060 ne
rect 5962 11962 6316 12060
tri 6316 11962 6414 12060 sw
tri 6414 11962 6512 12060 ne
rect 6512 11962 6866 12060
tri 6866 11962 6964 12060 sw
tri 6964 11962 7062 12060 ne
rect 7062 11962 7416 12060
tri 7416 11962 7514 12060 sw
tri 7514 11962 7612 12060 ne
rect 7612 11962 7966 12060
tri 7966 11962 8064 12060 sw
tri 8064 11962 8162 12060 ne
rect 8162 11962 8516 12060
tri 8516 11962 8614 12060 sw
tri 8614 11962 8712 12060 ne
rect 8712 11962 9066 12060
tri 9066 11962 9164 12060 sw
tri 9164 11962 9262 12060 ne
rect 9262 11962 9616 12060
tri 9616 11962 9714 12060 sw
tri 9714 11962 9812 12060 ne
rect 9812 11962 10166 12060
tri 10166 11962 10264 12060 sw
tri 10264 11962 10362 12060 ne
rect 10362 11962 10716 12060
tri 10716 11962 10814 12060 sw
tri 10814 11962 10912 12060 ne
rect 10912 11962 11266 12060
tri 11266 11962 11364 12060 sw
tri 11364 11962 11462 12060 ne
rect 11462 11962 11816 12060
tri 11816 11962 11914 12060 sw
tri 11914 11962 12012 12060 ne
rect 12012 11962 12366 12060
tri 12366 11962 12464 12060 sw
tri 12464 11962 12562 12060 ne
rect 12562 11962 12916 12060
tri 12916 11962 13014 12060 sw
tri 13014 11962 13112 12060 ne
rect 13112 11962 13466 12060
tri 13466 11962 13564 12060 sw
tri 13564 11962 13662 12060 ne
rect 13662 11962 15775 12060
rect -825 11912 -186 11962
rect -1025 11864 -186 11912
tri -186 11864 -88 11962 sw
tri -88 11864 10 11962 ne
rect 10 11864 364 11962
tri 364 11864 462 11962 sw
tri 462 11864 560 11962 ne
rect 560 11864 914 11962
tri 914 11864 1012 11962 sw
tri 1012 11864 1110 11962 ne
rect 1110 11864 1464 11962
tri 1464 11864 1562 11962 sw
tri 1562 11864 1660 11962 ne
rect 1660 11864 2014 11962
tri 2014 11864 2112 11962 sw
tri 2112 11864 2210 11962 ne
rect 2210 11864 2564 11962
tri 2564 11864 2662 11962 sw
tri 2662 11864 2760 11962 ne
rect 2760 11864 3114 11962
tri 3114 11864 3212 11962 sw
tri 3212 11864 3310 11962 ne
rect 3310 11864 3664 11962
tri 3664 11864 3762 11962 sw
tri 3762 11864 3860 11962 ne
rect 3860 11864 4214 11962
tri 4214 11864 4312 11962 sw
tri 4312 11864 4410 11962 ne
rect 4410 11864 4764 11962
tri 4764 11864 4862 11962 sw
tri 4862 11864 4960 11962 ne
rect 4960 11864 5314 11962
tri 5314 11864 5412 11962 sw
tri 5412 11864 5510 11962 ne
rect 5510 11864 5864 11962
tri 5864 11864 5962 11962 sw
tri 5962 11864 6060 11962 ne
rect 6060 11864 6414 11962
tri 6414 11864 6512 11962 sw
tri 6512 11864 6610 11962 ne
rect 6610 11864 6964 11962
tri 6964 11864 7062 11962 sw
tri 7062 11864 7160 11962 ne
rect 7160 11864 7514 11962
tri 7514 11864 7612 11962 sw
tri 7612 11864 7710 11962 ne
rect 7710 11864 8064 11962
tri 8064 11864 8162 11962 sw
tri 8162 11864 8260 11962 ne
rect 8260 11864 8614 11962
tri 8614 11864 8712 11962 sw
tri 8712 11864 8810 11962 ne
rect 8810 11864 9164 11962
tri 9164 11864 9262 11962 sw
tri 9262 11864 9360 11962 ne
rect 9360 11864 9714 11962
tri 9714 11864 9812 11962 sw
tri 9812 11864 9910 11962 ne
rect 9910 11864 10264 11962
tri 10264 11864 10362 11962 sw
tri 10362 11864 10460 11962 ne
rect 10460 11864 10814 11962
tri 10814 11864 10912 11962 sw
tri 10912 11864 11010 11962 ne
rect 11010 11864 11364 11962
tri 11364 11864 11462 11962 sw
tri 11462 11864 11560 11962 ne
rect 11560 11864 11914 11962
tri 11914 11864 12012 11962 sw
tri 12012 11864 12110 11962 ne
rect 12110 11864 12464 11962
tri 12464 11864 12562 11962 sw
tri 12562 11864 12660 11962 ne
rect 12660 11864 13014 11962
tri 13014 11864 13112 11962 sw
tri 13112 11864 13210 11962 ne
rect 13210 11864 13564 11962
tri 13564 11864 13662 11962 sw
rect -1025 11860 -88 11864
rect -1025 11740 -310 11860
rect -190 11776 -88 11860
tri -88 11776 0 11864 sw
tri 10 11776 98 11864 ne
rect 98 11860 462 11864
rect 98 11776 240 11860
rect -190 11740 0 11776
rect -1025 11736 0 11740
tri 0 11736 40 11776 sw
tri 98 11736 138 11776 ne
rect 138 11740 240 11776
rect 360 11776 462 11860
tri 462 11776 550 11864 sw
tri 560 11776 648 11864 ne
rect 648 11860 1012 11864
rect 648 11776 790 11860
rect 360 11740 550 11776
rect 138 11736 550 11740
tri -412 11638 -314 11736 ne
rect -314 11638 40 11736
tri 40 11638 138 11736 sw
tri 138 11638 236 11736 ne
rect 236 11688 550 11736
tri 550 11688 638 11776 sw
tri 648 11688 736 11776 ne
rect 736 11740 790 11776
rect 910 11776 1012 11860
tri 1012 11776 1100 11864 sw
tri 1110 11776 1198 11864 ne
rect 1198 11860 1562 11864
rect 1198 11776 1340 11860
rect 910 11740 1100 11776
rect 736 11736 1100 11740
tri 1100 11736 1140 11776 sw
tri 1198 11736 1238 11776 ne
rect 1238 11740 1340 11776
rect 1460 11776 1562 11860
tri 1562 11776 1650 11864 sw
tri 1660 11776 1748 11864 ne
rect 1748 11860 2112 11864
rect 1748 11776 1890 11860
rect 1460 11740 1650 11776
rect 1238 11736 1650 11740
rect 736 11688 1140 11736
rect 236 11638 638 11688
rect -2525 11550 -412 11638
tri -412 11550 -324 11638 sw
tri -314 11550 -226 11638 ne
rect -226 11550 138 11638
tri 138 11550 226 11638 sw
tri 236 11550 324 11638 ne
rect 324 11608 638 11638
tri 638 11608 718 11688 sw
tri 736 11608 816 11688 ne
rect 816 11638 1140 11688
tri 1140 11638 1238 11736 sw
tri 1238 11638 1336 11736 ne
rect 1336 11688 1650 11736
tri 1650 11688 1738 11776 sw
tri 1748 11688 1836 11776 ne
rect 1836 11740 1890 11776
rect 2010 11776 2112 11860
tri 2112 11776 2200 11864 sw
tri 2210 11776 2298 11864 ne
rect 2298 11860 2662 11864
rect 2298 11776 2440 11860
rect 2010 11740 2200 11776
rect 1836 11736 2200 11740
tri 2200 11736 2240 11776 sw
tri 2298 11736 2338 11776 ne
rect 2338 11740 2440 11776
rect 2560 11776 2662 11860
tri 2662 11776 2750 11864 sw
tri 2760 11776 2848 11864 ne
rect 2848 11860 3212 11864
rect 2848 11776 2990 11860
rect 2560 11740 2750 11776
rect 2338 11736 2750 11740
rect 1836 11688 2240 11736
rect 1336 11638 1738 11688
rect 816 11608 1238 11638
rect 324 11550 718 11608
rect -2525 11510 -324 11550
tri -324 11510 -284 11550 sw
tri -226 11510 -186 11550 ne
rect -186 11510 226 11550
tri 226 11510 266 11550 sw
tri 324 11510 364 11550 ne
rect 364 11510 718 11550
tri 718 11510 816 11608 sw
tri 816 11510 914 11608 ne
rect 914 11550 1238 11608
tri 1238 11550 1326 11638 sw
tri 1336 11550 1424 11638 ne
rect 1424 11608 1738 11638
tri 1738 11608 1818 11688 sw
tri 1836 11608 1916 11688 ne
rect 1916 11638 2240 11688
tri 2240 11638 2338 11736 sw
tri 2338 11638 2436 11736 ne
rect 2436 11688 2750 11736
tri 2750 11688 2838 11776 sw
tri 2848 11688 2936 11776 ne
rect 2936 11740 2990 11776
rect 3110 11776 3212 11860
tri 3212 11776 3300 11864 sw
tri 3310 11776 3398 11864 ne
rect 3398 11860 3762 11864
rect 3398 11776 3540 11860
rect 3110 11740 3300 11776
rect 2936 11736 3300 11740
tri 3300 11736 3340 11776 sw
tri 3398 11736 3438 11776 ne
rect 3438 11740 3540 11776
rect 3660 11776 3762 11860
tri 3762 11776 3850 11864 sw
tri 3860 11776 3948 11864 ne
rect 3948 11860 4312 11864
rect 3948 11776 4090 11860
rect 3660 11740 3850 11776
rect 3438 11736 3850 11740
rect 2936 11688 3340 11736
rect 2436 11638 2838 11688
rect 1916 11608 2338 11638
rect 1424 11550 1818 11608
rect 914 11510 1326 11550
tri 1326 11510 1366 11550 sw
tri 1424 11510 1464 11550 ne
rect 1464 11510 1818 11550
tri 1818 11510 1916 11608 sw
tri 1916 11510 2014 11608 ne
rect 2014 11550 2338 11608
tri 2338 11550 2426 11638 sw
tri 2436 11550 2524 11638 ne
rect 2524 11608 2838 11638
tri 2838 11608 2918 11688 sw
tri 2936 11608 3016 11688 ne
rect 3016 11638 3340 11688
tri 3340 11638 3438 11736 sw
tri 3438 11638 3536 11736 ne
rect 3536 11688 3850 11736
tri 3850 11688 3938 11776 sw
tri 3948 11688 4036 11776 ne
rect 4036 11740 4090 11776
rect 4210 11776 4312 11860
tri 4312 11776 4400 11864 sw
tri 4410 11776 4498 11864 ne
rect 4498 11860 4862 11864
rect 4498 11776 4640 11860
rect 4210 11740 4400 11776
rect 4036 11736 4400 11740
tri 4400 11736 4440 11776 sw
tri 4498 11736 4538 11776 ne
rect 4538 11740 4640 11776
rect 4760 11776 4862 11860
tri 4862 11776 4950 11864 sw
tri 4960 11776 5048 11864 ne
rect 5048 11860 5412 11864
rect 5048 11776 5190 11860
rect 4760 11740 4950 11776
rect 4538 11736 4950 11740
rect 4036 11688 4440 11736
rect 3536 11638 3938 11688
rect 3016 11608 3438 11638
rect 2524 11550 2918 11608
rect 2014 11510 2426 11550
tri 2426 11510 2466 11550 sw
tri 2524 11510 2564 11550 ne
rect 2564 11510 2918 11550
tri 2918 11510 3016 11608 sw
tri 3016 11510 3114 11608 ne
rect 3114 11550 3438 11608
tri 3438 11550 3526 11638 sw
tri 3536 11550 3624 11638 ne
rect 3624 11608 3938 11638
tri 3938 11608 4018 11688 sw
tri 4036 11608 4116 11688 ne
rect 4116 11638 4440 11688
tri 4440 11638 4538 11736 sw
tri 4538 11638 4636 11736 ne
rect 4636 11688 4950 11736
tri 4950 11688 5038 11776 sw
tri 5048 11688 5136 11776 ne
rect 5136 11740 5190 11776
rect 5310 11776 5412 11860
tri 5412 11776 5500 11864 sw
tri 5510 11776 5598 11864 ne
rect 5598 11860 5962 11864
rect 5598 11776 5740 11860
rect 5310 11740 5500 11776
rect 5136 11736 5500 11740
tri 5500 11736 5540 11776 sw
tri 5598 11736 5638 11776 ne
rect 5638 11740 5740 11776
rect 5860 11776 5962 11860
tri 5962 11776 6050 11864 sw
tri 6060 11776 6148 11864 ne
rect 6148 11860 6512 11864
rect 6148 11776 6290 11860
rect 5860 11740 6050 11776
rect 5638 11736 6050 11740
rect 5136 11688 5540 11736
rect 4636 11638 5038 11688
rect 4116 11608 4538 11638
rect 3624 11550 4018 11608
rect 3114 11510 3526 11550
tri 3526 11510 3566 11550 sw
tri 3624 11510 3664 11550 ne
rect 3664 11510 4018 11550
tri 4018 11510 4116 11608 sw
tri 4116 11510 4214 11608 ne
rect 4214 11550 4538 11608
tri 4538 11550 4626 11638 sw
tri 4636 11550 4724 11638 ne
rect 4724 11608 5038 11638
tri 5038 11608 5118 11688 sw
tri 5136 11608 5216 11688 ne
rect 5216 11638 5540 11688
tri 5540 11638 5638 11736 sw
tri 5638 11638 5736 11736 ne
rect 5736 11688 6050 11736
tri 6050 11688 6138 11776 sw
tri 6148 11688 6236 11776 ne
rect 6236 11740 6290 11776
rect 6410 11776 6512 11860
tri 6512 11776 6600 11864 sw
tri 6610 11776 6698 11864 ne
rect 6698 11860 7062 11864
rect 6698 11776 6840 11860
rect 6410 11740 6600 11776
rect 6236 11736 6600 11740
tri 6600 11736 6640 11776 sw
tri 6698 11736 6738 11776 ne
rect 6738 11740 6840 11776
rect 6960 11776 7062 11860
tri 7062 11776 7150 11864 sw
tri 7160 11776 7248 11864 ne
rect 7248 11860 7612 11864
rect 7248 11776 7390 11860
rect 6960 11740 7150 11776
rect 6738 11736 7150 11740
rect 6236 11688 6640 11736
rect 5736 11638 6138 11688
rect 5216 11608 5638 11638
rect 4724 11550 5118 11608
rect 4214 11510 4626 11550
tri 4626 11510 4666 11550 sw
tri 4724 11510 4764 11550 ne
rect 4764 11510 5118 11550
tri 5118 11510 5216 11608 sw
tri 5216 11510 5314 11608 ne
rect 5314 11550 5638 11608
tri 5638 11550 5726 11638 sw
tri 5736 11550 5824 11638 ne
rect 5824 11608 6138 11638
tri 6138 11608 6218 11688 sw
tri 6236 11608 6316 11688 ne
rect 6316 11638 6640 11688
tri 6640 11638 6738 11736 sw
tri 6738 11638 6836 11736 ne
rect 6836 11688 7150 11736
tri 7150 11688 7238 11776 sw
tri 7248 11688 7336 11776 ne
rect 7336 11740 7390 11776
rect 7510 11776 7612 11860
tri 7612 11776 7700 11864 sw
tri 7710 11776 7798 11864 ne
rect 7798 11860 8162 11864
rect 7798 11776 7940 11860
rect 7510 11740 7700 11776
rect 7336 11736 7700 11740
tri 7700 11736 7740 11776 sw
tri 7798 11736 7838 11776 ne
rect 7838 11740 7940 11776
rect 8060 11776 8162 11860
tri 8162 11776 8250 11864 sw
tri 8260 11776 8348 11864 ne
rect 8348 11860 8712 11864
rect 8348 11776 8490 11860
rect 8060 11740 8250 11776
rect 7838 11736 8250 11740
rect 7336 11688 7740 11736
rect 6836 11638 7238 11688
rect 6316 11608 6738 11638
rect 5824 11550 6218 11608
rect 5314 11510 5726 11550
tri 5726 11510 5766 11550 sw
tri 5824 11510 5864 11550 ne
rect 5864 11510 6218 11550
tri 6218 11510 6316 11608 sw
tri 6316 11510 6414 11608 ne
rect 6414 11550 6738 11608
tri 6738 11550 6826 11638 sw
tri 6836 11550 6924 11638 ne
rect 6924 11608 7238 11638
tri 7238 11608 7318 11688 sw
tri 7336 11608 7416 11688 ne
rect 7416 11638 7740 11688
tri 7740 11638 7838 11736 sw
tri 7838 11638 7936 11736 ne
rect 7936 11688 8250 11736
tri 8250 11688 8338 11776 sw
tri 8348 11688 8436 11776 ne
rect 8436 11740 8490 11776
rect 8610 11776 8712 11860
tri 8712 11776 8800 11864 sw
tri 8810 11776 8898 11864 ne
rect 8898 11860 9262 11864
rect 8898 11776 9040 11860
rect 8610 11740 8800 11776
rect 8436 11736 8800 11740
tri 8800 11736 8840 11776 sw
tri 8898 11736 8938 11776 ne
rect 8938 11740 9040 11776
rect 9160 11776 9262 11860
tri 9262 11776 9350 11864 sw
tri 9360 11776 9448 11864 ne
rect 9448 11860 9812 11864
rect 9448 11776 9590 11860
rect 9160 11740 9350 11776
rect 8938 11736 9350 11740
rect 8436 11688 8840 11736
rect 7936 11638 8338 11688
rect 7416 11608 7838 11638
rect 6924 11550 7318 11608
rect 6414 11510 6826 11550
tri 6826 11510 6866 11550 sw
tri 6924 11510 6964 11550 ne
rect 6964 11510 7318 11550
tri 7318 11510 7416 11608 sw
tri 7416 11510 7514 11608 ne
rect 7514 11550 7838 11608
tri 7838 11550 7926 11638 sw
tri 7936 11550 8024 11638 ne
rect 8024 11608 8338 11638
tri 8338 11608 8418 11688 sw
tri 8436 11608 8516 11688 ne
rect 8516 11638 8840 11688
tri 8840 11638 8938 11736 sw
tri 8938 11638 9036 11736 ne
rect 9036 11688 9350 11736
tri 9350 11688 9438 11776 sw
tri 9448 11688 9536 11776 ne
rect 9536 11740 9590 11776
rect 9710 11776 9812 11860
tri 9812 11776 9900 11864 sw
tri 9910 11776 9998 11864 ne
rect 9998 11860 10362 11864
rect 9998 11776 10140 11860
rect 9710 11740 9900 11776
rect 9536 11736 9900 11740
tri 9900 11736 9940 11776 sw
tri 9998 11736 10038 11776 ne
rect 10038 11740 10140 11776
rect 10260 11776 10362 11860
tri 10362 11776 10450 11864 sw
tri 10460 11776 10548 11864 ne
rect 10548 11860 10912 11864
rect 10548 11776 10690 11860
rect 10260 11740 10450 11776
rect 10038 11736 10450 11740
rect 9536 11688 9940 11736
rect 9036 11638 9438 11688
rect 8516 11608 8938 11638
rect 8024 11550 8418 11608
rect 7514 11510 7926 11550
tri 7926 11510 7966 11550 sw
tri 8024 11510 8064 11550 ne
rect 8064 11510 8418 11550
tri 8418 11510 8516 11608 sw
tri 8516 11510 8614 11608 ne
rect 8614 11550 8938 11608
tri 8938 11550 9026 11638 sw
tri 9036 11550 9124 11638 ne
rect 9124 11608 9438 11638
tri 9438 11608 9518 11688 sw
tri 9536 11608 9616 11688 ne
rect 9616 11638 9940 11688
tri 9940 11638 10038 11736 sw
tri 10038 11638 10136 11736 ne
rect 10136 11688 10450 11736
tri 10450 11688 10538 11776 sw
tri 10548 11688 10636 11776 ne
rect 10636 11740 10690 11776
rect 10810 11776 10912 11860
tri 10912 11776 11000 11864 sw
tri 11010 11776 11098 11864 ne
rect 11098 11860 11462 11864
rect 11098 11776 11240 11860
rect 10810 11740 11000 11776
rect 10636 11736 11000 11740
tri 11000 11736 11040 11776 sw
tri 11098 11736 11138 11776 ne
rect 11138 11740 11240 11776
rect 11360 11776 11462 11860
tri 11462 11776 11550 11864 sw
tri 11560 11776 11648 11864 ne
rect 11648 11860 12012 11864
rect 11648 11776 11790 11860
rect 11360 11740 11550 11776
rect 11138 11736 11550 11740
rect 10636 11688 11040 11736
rect 10136 11638 10538 11688
rect 9616 11608 10038 11638
rect 9124 11550 9518 11608
rect 8614 11510 9026 11550
tri 9026 11510 9066 11550 sw
tri 9124 11510 9164 11550 ne
rect 9164 11510 9518 11550
tri 9518 11510 9616 11608 sw
tri 9616 11510 9714 11608 ne
rect 9714 11550 10038 11608
tri 10038 11550 10126 11638 sw
tri 10136 11550 10224 11638 ne
rect 10224 11608 10538 11638
tri 10538 11608 10618 11688 sw
tri 10636 11608 10716 11688 ne
rect 10716 11638 11040 11688
tri 11040 11638 11138 11736 sw
tri 11138 11638 11236 11736 ne
rect 11236 11688 11550 11736
tri 11550 11688 11638 11776 sw
tri 11648 11688 11736 11776 ne
rect 11736 11740 11790 11776
rect 11910 11776 12012 11860
tri 12012 11776 12100 11864 sw
tri 12110 11776 12198 11864 ne
rect 12198 11860 12562 11864
rect 12198 11776 12340 11860
rect 11910 11740 12100 11776
rect 11736 11736 12100 11740
tri 12100 11736 12140 11776 sw
tri 12198 11736 12238 11776 ne
rect 12238 11740 12340 11776
rect 12460 11776 12562 11860
tri 12562 11776 12650 11864 sw
tri 12660 11776 12748 11864 ne
rect 12748 11860 13112 11864
rect 12748 11776 12890 11860
rect 12460 11740 12650 11776
rect 12238 11736 12650 11740
rect 11736 11688 12140 11736
rect 11236 11638 11638 11688
rect 10716 11608 11138 11638
rect 10224 11550 10618 11608
rect 9714 11510 10126 11550
tri 10126 11510 10166 11550 sw
tri 10224 11510 10264 11550 ne
rect 10264 11510 10618 11550
tri 10618 11510 10716 11608 sw
tri 10716 11510 10814 11608 ne
rect 10814 11550 11138 11608
tri 11138 11550 11226 11638 sw
tri 11236 11550 11324 11638 ne
rect 11324 11608 11638 11638
tri 11638 11608 11718 11688 sw
tri 11736 11608 11816 11688 ne
rect 11816 11638 12140 11688
tri 12140 11638 12238 11736 sw
tri 12238 11638 12336 11736 ne
rect 12336 11688 12650 11736
tri 12650 11688 12738 11776 sw
tri 12748 11688 12836 11776 ne
rect 12836 11740 12890 11776
rect 13010 11776 13112 11860
tri 13112 11776 13200 11864 sw
tri 13210 11776 13298 11864 ne
rect 13298 11860 14275 11864
rect 13298 11776 13440 11860
rect 13010 11740 13200 11776
rect 12836 11736 13200 11740
tri 13200 11736 13240 11776 sw
tri 13298 11736 13338 11776 ne
rect 13338 11740 13440 11776
rect 13560 11740 14275 11860
rect 13338 11736 14275 11740
rect 12836 11688 13240 11736
rect 12336 11638 12738 11688
rect 11816 11608 12238 11638
rect 11324 11550 11718 11608
rect 10814 11510 11226 11550
tri 11226 11510 11266 11550 sw
tri 11324 11510 11364 11550 ne
rect 11364 11510 11718 11550
tri 11718 11510 11816 11608 sw
tri 11816 11510 11914 11608 ne
rect 11914 11550 12238 11608
tri 12238 11550 12326 11638 sw
tri 12336 11550 12424 11638 ne
rect 12424 11608 12738 11638
tri 12738 11608 12818 11688 sw
tri 12836 11608 12916 11688 ne
rect 12916 11638 13240 11688
tri 13240 11638 13338 11736 sw
tri 13338 11638 13436 11736 ne
rect 13436 11638 14275 11736
rect 12916 11608 13338 11638
rect 12424 11550 12818 11608
rect 11914 11510 12326 11550
tri 12326 11510 12366 11550 sw
tri 12424 11510 12464 11550 ne
rect 12464 11510 12818 11550
tri 12818 11510 12916 11608 sw
tri 12916 11510 13014 11608 ne
rect 13014 11550 13338 11608
tri 13338 11550 13426 11638 sw
tri 13436 11550 13524 11638 ne
rect 13524 11550 14275 11638
rect 13014 11510 13426 11550
tri 13426 11510 13466 11550 sw
tri 13524 11510 13564 11550 ne
rect 13564 11510 14275 11550
rect -2525 11412 -284 11510
tri -284 11412 -186 11510 sw
tri -186 11412 -88 11510 ne
rect -88 11412 266 11510
tri 266 11412 364 11510 sw
tri 364 11412 462 11510 ne
rect 462 11412 816 11510
tri 816 11412 914 11510 sw
tri 914 11412 1012 11510 ne
rect 1012 11412 1366 11510
tri 1366 11412 1464 11510 sw
tri 1464 11412 1562 11510 ne
rect 1562 11412 1916 11510
tri 1916 11412 2014 11510 sw
tri 2014 11412 2112 11510 ne
rect 2112 11412 2466 11510
tri 2466 11412 2564 11510 sw
tri 2564 11412 2662 11510 ne
rect 2662 11412 3016 11510
tri 3016 11412 3114 11510 sw
tri 3114 11412 3212 11510 ne
rect 3212 11412 3566 11510
tri 3566 11412 3664 11510 sw
tri 3664 11412 3762 11510 ne
rect 3762 11412 4116 11510
tri 4116 11412 4214 11510 sw
tri 4214 11412 4312 11510 ne
rect 4312 11412 4666 11510
tri 4666 11412 4764 11510 sw
tri 4764 11412 4862 11510 ne
rect 4862 11412 5216 11510
tri 5216 11412 5314 11510 sw
tri 5314 11412 5412 11510 ne
rect 5412 11412 5766 11510
tri 5766 11412 5864 11510 sw
tri 5864 11412 5962 11510 ne
rect 5962 11412 6316 11510
tri 6316 11412 6414 11510 sw
tri 6414 11412 6512 11510 ne
rect 6512 11412 6866 11510
tri 6866 11412 6964 11510 sw
tri 6964 11412 7062 11510 ne
rect 7062 11412 7416 11510
tri 7416 11412 7514 11510 sw
tri 7514 11412 7612 11510 ne
rect 7612 11412 7966 11510
tri 7966 11412 8064 11510 sw
tri 8064 11412 8162 11510 ne
rect 8162 11412 8516 11510
tri 8516 11412 8614 11510 sw
tri 8614 11412 8712 11510 ne
rect 8712 11412 9066 11510
tri 9066 11412 9164 11510 sw
tri 9164 11412 9262 11510 ne
rect 9262 11412 9616 11510
tri 9616 11412 9714 11510 sw
tri 9714 11412 9812 11510 ne
rect 9812 11412 10166 11510
tri 10166 11412 10264 11510 sw
tri 10264 11412 10362 11510 ne
rect 10362 11412 10716 11510
tri 10716 11412 10814 11510 sw
tri 10814 11412 10912 11510 ne
rect 10912 11412 11266 11510
tri 11266 11412 11364 11510 sw
tri 11364 11412 11462 11510 ne
rect 11462 11412 11816 11510
tri 11816 11412 11914 11510 sw
tri 11914 11412 12012 11510 ne
rect 12012 11412 12366 11510
tri 12366 11412 12464 11510 sw
tri 12464 11412 12562 11510 ne
rect 12562 11412 12916 11510
tri 12916 11412 13014 11510 sw
tri 13014 11412 13112 11510 ne
rect 13112 11412 13466 11510
tri 13466 11412 13564 11510 sw
tri 13564 11412 13662 11510 ne
rect 13662 11412 14275 11510
rect -2525 11314 -186 11412
tri -186 11314 -88 11412 sw
tri -88 11314 10 11412 ne
rect 10 11314 364 11412
tri 364 11314 462 11412 sw
tri 462 11314 560 11412 ne
rect 560 11314 914 11412
tri 914 11314 1012 11412 sw
tri 1012 11314 1110 11412 ne
rect 1110 11314 1464 11412
tri 1464 11314 1562 11412 sw
tri 1562 11314 1660 11412 ne
rect 1660 11314 2014 11412
tri 2014 11314 2112 11412 sw
tri 2112 11314 2210 11412 ne
rect 2210 11314 2564 11412
tri 2564 11314 2662 11412 sw
tri 2662 11314 2760 11412 ne
rect 2760 11314 3114 11412
tri 3114 11314 3212 11412 sw
tri 3212 11314 3310 11412 ne
rect 3310 11314 3664 11412
tri 3664 11314 3762 11412 sw
tri 3762 11314 3860 11412 ne
rect 3860 11314 4214 11412
tri 4214 11314 4312 11412 sw
tri 4312 11314 4410 11412 ne
rect 4410 11314 4764 11412
tri 4764 11314 4862 11412 sw
tri 4862 11314 4960 11412 ne
rect 4960 11314 5314 11412
tri 5314 11314 5412 11412 sw
tri 5412 11314 5510 11412 ne
rect 5510 11314 5864 11412
tri 5864 11314 5962 11412 sw
tri 5962 11314 6060 11412 ne
rect 6060 11314 6414 11412
tri 6414 11314 6512 11412 sw
tri 6512 11314 6610 11412 ne
rect 6610 11314 6964 11412
tri 6964 11314 7062 11412 sw
tri 7062 11314 7160 11412 ne
rect 7160 11314 7514 11412
tri 7514 11314 7612 11412 sw
tri 7612 11314 7710 11412 ne
rect 7710 11314 8064 11412
tri 8064 11314 8162 11412 sw
tri 8162 11314 8260 11412 ne
rect 8260 11314 8614 11412
tri 8614 11314 8712 11412 sw
tri 8712 11314 8810 11412 ne
rect 8810 11314 9164 11412
tri 9164 11314 9262 11412 sw
tri 9262 11314 9360 11412 ne
rect 9360 11314 9714 11412
tri 9714 11314 9812 11412 sw
tri 9812 11314 9910 11412 ne
rect 9910 11314 10264 11412
tri 10264 11314 10362 11412 sw
tri 10362 11314 10460 11412 ne
rect 10460 11314 10814 11412
tri 10814 11314 10912 11412 sw
tri 10912 11314 11010 11412 ne
rect 11010 11314 11364 11412
tri 11364 11314 11462 11412 sw
tri 11462 11314 11560 11412 ne
rect 11560 11314 11914 11412
tri 11914 11314 12012 11412 sw
tri 12012 11314 12110 11412 ne
rect 12110 11314 12464 11412
tri 12464 11314 12562 11412 sw
tri 12562 11314 12660 11412 ne
rect 12660 11314 13014 11412
tri 13014 11314 13112 11412 sw
tri 13112 11314 13210 11412 ne
rect 13210 11314 13564 11412
tri 13564 11314 13662 11412 sw
rect 14775 11314 15775 11962
rect -2525 11310 -88 11314
rect -2525 11190 -310 11310
rect -190 11226 -88 11310
tri -88 11226 0 11314 sw
tri 10 11226 98 11314 ne
rect 98 11310 462 11314
rect 98 11226 240 11310
rect -190 11190 0 11226
rect -2525 11186 0 11190
rect -2525 10538 -1525 11186
tri -412 11088 -314 11186 ne
rect -314 11138 0 11186
tri 0 11138 88 11226 sw
tri 98 11138 186 11226 ne
rect 186 11190 240 11226
rect 360 11226 462 11310
tri 462 11226 550 11314 sw
tri 560 11226 648 11314 ne
rect 648 11310 1012 11314
rect 648 11226 790 11310
rect 360 11190 550 11226
rect 186 11186 550 11190
tri 550 11186 590 11226 sw
tri 648 11186 688 11226 ne
rect 688 11190 790 11226
rect 910 11226 1012 11310
tri 1012 11226 1100 11314 sw
tri 1110 11226 1198 11314 ne
rect 1198 11310 1562 11314
rect 1198 11226 1340 11310
rect 910 11190 1100 11226
rect 688 11186 1100 11190
rect 186 11138 590 11186
rect -314 11088 88 11138
rect -1025 11000 -412 11088
tri -412 11000 -324 11088 sw
tri -314 11000 -226 11088 ne
rect -226 11058 88 11088
tri 88 11058 168 11138 sw
tri 186 11058 266 11138 ne
rect 266 11088 590 11138
tri 590 11088 688 11186 sw
tri 688 11088 786 11186 ne
rect 786 11138 1100 11186
tri 1100 11138 1188 11226 sw
tri 1198 11138 1286 11226 ne
rect 1286 11190 1340 11226
rect 1460 11226 1562 11310
tri 1562 11226 1650 11314 sw
tri 1660 11226 1748 11314 ne
rect 1748 11310 2112 11314
rect 1748 11226 1890 11310
rect 1460 11190 1650 11226
rect 1286 11186 1650 11190
tri 1650 11186 1690 11226 sw
tri 1748 11186 1788 11226 ne
rect 1788 11190 1890 11226
rect 2010 11226 2112 11310
tri 2112 11226 2200 11314 sw
tri 2210 11226 2298 11314 ne
rect 2298 11310 2662 11314
rect 2298 11226 2440 11310
rect 2010 11190 2200 11226
rect 1788 11186 2200 11190
rect 1286 11138 1690 11186
rect 786 11088 1188 11138
rect 266 11058 688 11088
rect -226 11000 168 11058
rect -1025 10960 -324 11000
tri -324 10960 -284 11000 sw
tri -226 10960 -186 11000 ne
rect -186 10960 168 11000
tri 168 10960 266 11058 sw
tri 266 10960 364 11058 ne
rect 364 11000 688 11058
tri 688 11000 776 11088 sw
tri 786 11000 874 11088 ne
rect 874 11058 1188 11088
tri 1188 11058 1268 11138 sw
tri 1286 11058 1366 11138 ne
rect 1366 11088 1690 11138
tri 1690 11088 1788 11186 sw
tri 1788 11088 1886 11186 ne
rect 1886 11138 2200 11186
tri 2200 11138 2288 11226 sw
tri 2298 11138 2386 11226 ne
rect 2386 11190 2440 11226
rect 2560 11226 2662 11310
tri 2662 11226 2750 11314 sw
tri 2760 11226 2848 11314 ne
rect 2848 11310 3212 11314
rect 2848 11226 2990 11310
rect 2560 11190 2750 11226
rect 2386 11186 2750 11190
tri 2750 11186 2790 11226 sw
tri 2848 11186 2888 11226 ne
rect 2888 11190 2990 11226
rect 3110 11226 3212 11310
tri 3212 11226 3300 11314 sw
tri 3310 11226 3398 11314 ne
rect 3398 11310 3762 11314
rect 3398 11226 3540 11310
rect 3110 11190 3300 11226
rect 2888 11186 3300 11190
rect 2386 11138 2790 11186
rect 1886 11088 2288 11138
rect 1366 11058 1788 11088
rect 874 11000 1268 11058
rect 364 10960 776 11000
tri 776 10960 816 11000 sw
tri 874 10960 914 11000 ne
rect 914 10960 1268 11000
tri 1268 10960 1366 11058 sw
tri 1366 10960 1464 11058 ne
rect 1464 11000 1788 11058
tri 1788 11000 1876 11088 sw
tri 1886 11000 1974 11088 ne
rect 1974 11058 2288 11088
tri 2288 11058 2368 11138 sw
tri 2386 11058 2466 11138 ne
rect 2466 11088 2790 11138
tri 2790 11088 2888 11186 sw
tri 2888 11088 2986 11186 ne
rect 2986 11138 3300 11186
tri 3300 11138 3388 11226 sw
tri 3398 11138 3486 11226 ne
rect 3486 11190 3540 11226
rect 3660 11226 3762 11310
tri 3762 11226 3850 11314 sw
tri 3860 11226 3948 11314 ne
rect 3948 11310 4312 11314
rect 3948 11226 4090 11310
rect 3660 11190 3850 11226
rect 3486 11186 3850 11190
tri 3850 11186 3890 11226 sw
tri 3948 11186 3988 11226 ne
rect 3988 11190 4090 11226
rect 4210 11226 4312 11310
tri 4312 11226 4400 11314 sw
tri 4410 11226 4498 11314 ne
rect 4498 11310 4862 11314
rect 4498 11226 4640 11310
rect 4210 11190 4400 11226
rect 3988 11186 4400 11190
rect 3486 11138 3890 11186
rect 2986 11088 3388 11138
rect 2466 11058 2888 11088
rect 1974 11000 2368 11058
rect 1464 10960 1876 11000
tri 1876 10960 1916 11000 sw
tri 1974 10960 2014 11000 ne
rect 2014 10960 2368 11000
tri 2368 10960 2466 11058 sw
tri 2466 10960 2564 11058 ne
rect 2564 11000 2888 11058
tri 2888 11000 2976 11088 sw
tri 2986 11000 3074 11088 ne
rect 3074 11058 3388 11088
tri 3388 11058 3468 11138 sw
tri 3486 11058 3566 11138 ne
rect 3566 11088 3890 11138
tri 3890 11088 3988 11186 sw
tri 3988 11088 4086 11186 ne
rect 4086 11138 4400 11186
tri 4400 11138 4488 11226 sw
tri 4498 11138 4586 11226 ne
rect 4586 11190 4640 11226
rect 4760 11226 4862 11310
tri 4862 11226 4950 11314 sw
tri 4960 11226 5048 11314 ne
rect 5048 11310 5412 11314
rect 5048 11226 5190 11310
rect 4760 11190 4950 11226
rect 4586 11186 4950 11190
tri 4950 11186 4990 11226 sw
tri 5048 11186 5088 11226 ne
rect 5088 11190 5190 11226
rect 5310 11226 5412 11310
tri 5412 11226 5500 11314 sw
tri 5510 11226 5598 11314 ne
rect 5598 11310 5962 11314
rect 5598 11226 5740 11310
rect 5310 11190 5500 11226
rect 5088 11186 5500 11190
rect 4586 11138 4990 11186
rect 4086 11088 4488 11138
rect 3566 11058 3988 11088
rect 3074 11000 3468 11058
rect 2564 10960 2976 11000
tri 2976 10960 3016 11000 sw
tri 3074 10960 3114 11000 ne
rect 3114 10960 3468 11000
tri 3468 10960 3566 11058 sw
tri 3566 10960 3664 11058 ne
rect 3664 11000 3988 11058
tri 3988 11000 4076 11088 sw
tri 4086 11000 4174 11088 ne
rect 4174 11058 4488 11088
tri 4488 11058 4568 11138 sw
tri 4586 11058 4666 11138 ne
rect 4666 11088 4990 11138
tri 4990 11088 5088 11186 sw
tri 5088 11088 5186 11186 ne
rect 5186 11138 5500 11186
tri 5500 11138 5588 11226 sw
tri 5598 11138 5686 11226 ne
rect 5686 11190 5740 11226
rect 5860 11226 5962 11310
tri 5962 11226 6050 11314 sw
tri 6060 11226 6148 11314 ne
rect 6148 11310 6512 11314
rect 6148 11226 6290 11310
rect 5860 11190 6050 11226
rect 5686 11186 6050 11190
tri 6050 11186 6090 11226 sw
tri 6148 11186 6188 11226 ne
rect 6188 11190 6290 11226
rect 6410 11226 6512 11310
tri 6512 11226 6600 11314 sw
tri 6610 11226 6698 11314 ne
rect 6698 11310 7062 11314
rect 6698 11226 6840 11310
rect 6410 11190 6600 11226
rect 6188 11186 6600 11190
rect 5686 11138 6090 11186
rect 5186 11088 5588 11138
rect 4666 11058 5088 11088
rect 4174 11000 4568 11058
rect 3664 10960 4076 11000
tri 4076 10960 4116 11000 sw
tri 4174 10960 4214 11000 ne
rect 4214 10960 4568 11000
tri 4568 10960 4666 11058 sw
tri 4666 10960 4764 11058 ne
rect 4764 11000 5088 11058
tri 5088 11000 5176 11088 sw
tri 5186 11000 5274 11088 ne
rect 5274 11058 5588 11088
tri 5588 11058 5668 11138 sw
tri 5686 11058 5766 11138 ne
rect 5766 11088 6090 11138
tri 6090 11088 6188 11186 sw
tri 6188 11088 6286 11186 ne
rect 6286 11138 6600 11186
tri 6600 11138 6688 11226 sw
tri 6698 11138 6786 11226 ne
rect 6786 11190 6840 11226
rect 6960 11226 7062 11310
tri 7062 11226 7150 11314 sw
tri 7160 11226 7248 11314 ne
rect 7248 11310 7612 11314
rect 7248 11226 7390 11310
rect 6960 11190 7150 11226
rect 6786 11186 7150 11190
tri 7150 11186 7190 11226 sw
tri 7248 11186 7288 11226 ne
rect 7288 11190 7390 11226
rect 7510 11226 7612 11310
tri 7612 11226 7700 11314 sw
tri 7710 11226 7798 11314 ne
rect 7798 11310 8162 11314
rect 7798 11226 7940 11310
rect 7510 11190 7700 11226
rect 7288 11186 7700 11190
rect 6786 11138 7190 11186
rect 6286 11088 6688 11138
rect 5766 11058 6188 11088
rect 5274 11000 5668 11058
rect 4764 10960 5176 11000
tri 5176 10960 5216 11000 sw
tri 5274 10960 5314 11000 ne
rect 5314 10960 5668 11000
tri 5668 10960 5766 11058 sw
tri 5766 10960 5864 11058 ne
rect 5864 11000 6188 11058
tri 6188 11000 6276 11088 sw
tri 6286 11000 6374 11088 ne
rect 6374 11058 6688 11088
tri 6688 11058 6768 11138 sw
tri 6786 11058 6866 11138 ne
rect 6866 11088 7190 11138
tri 7190 11088 7288 11186 sw
tri 7288 11088 7386 11186 ne
rect 7386 11138 7700 11186
tri 7700 11138 7788 11226 sw
tri 7798 11138 7886 11226 ne
rect 7886 11190 7940 11226
rect 8060 11226 8162 11310
tri 8162 11226 8250 11314 sw
tri 8260 11226 8348 11314 ne
rect 8348 11310 8712 11314
rect 8348 11226 8490 11310
rect 8060 11190 8250 11226
rect 7886 11186 8250 11190
tri 8250 11186 8290 11226 sw
tri 8348 11186 8388 11226 ne
rect 8388 11190 8490 11226
rect 8610 11226 8712 11310
tri 8712 11226 8800 11314 sw
tri 8810 11226 8898 11314 ne
rect 8898 11310 9262 11314
rect 8898 11226 9040 11310
rect 8610 11190 8800 11226
rect 8388 11186 8800 11190
rect 7886 11138 8290 11186
rect 7386 11088 7788 11138
rect 6866 11058 7288 11088
rect 6374 11000 6768 11058
rect 5864 10960 6276 11000
tri 6276 10960 6316 11000 sw
tri 6374 10960 6414 11000 ne
rect 6414 10960 6768 11000
tri 6768 10960 6866 11058 sw
tri 6866 10960 6964 11058 ne
rect 6964 11000 7288 11058
tri 7288 11000 7376 11088 sw
tri 7386 11000 7474 11088 ne
rect 7474 11058 7788 11088
tri 7788 11058 7868 11138 sw
tri 7886 11058 7966 11138 ne
rect 7966 11088 8290 11138
tri 8290 11088 8388 11186 sw
tri 8388 11088 8486 11186 ne
rect 8486 11138 8800 11186
tri 8800 11138 8888 11226 sw
tri 8898 11138 8986 11226 ne
rect 8986 11190 9040 11226
rect 9160 11226 9262 11310
tri 9262 11226 9350 11314 sw
tri 9360 11226 9448 11314 ne
rect 9448 11310 9812 11314
rect 9448 11226 9590 11310
rect 9160 11190 9350 11226
rect 8986 11186 9350 11190
tri 9350 11186 9390 11226 sw
tri 9448 11186 9488 11226 ne
rect 9488 11190 9590 11226
rect 9710 11226 9812 11310
tri 9812 11226 9900 11314 sw
tri 9910 11226 9998 11314 ne
rect 9998 11310 10362 11314
rect 9998 11226 10140 11310
rect 9710 11190 9900 11226
rect 9488 11186 9900 11190
rect 8986 11138 9390 11186
rect 8486 11088 8888 11138
rect 7966 11058 8388 11088
rect 7474 11000 7868 11058
rect 6964 10960 7376 11000
tri 7376 10960 7416 11000 sw
tri 7474 10960 7514 11000 ne
rect 7514 10960 7868 11000
tri 7868 10960 7966 11058 sw
tri 7966 10960 8064 11058 ne
rect 8064 11000 8388 11058
tri 8388 11000 8476 11088 sw
tri 8486 11000 8574 11088 ne
rect 8574 11058 8888 11088
tri 8888 11058 8968 11138 sw
tri 8986 11058 9066 11138 ne
rect 9066 11088 9390 11138
tri 9390 11088 9488 11186 sw
tri 9488 11088 9586 11186 ne
rect 9586 11138 9900 11186
tri 9900 11138 9988 11226 sw
tri 9998 11138 10086 11226 ne
rect 10086 11190 10140 11226
rect 10260 11226 10362 11310
tri 10362 11226 10450 11314 sw
tri 10460 11226 10548 11314 ne
rect 10548 11310 10912 11314
rect 10548 11226 10690 11310
rect 10260 11190 10450 11226
rect 10086 11186 10450 11190
tri 10450 11186 10490 11226 sw
tri 10548 11186 10588 11226 ne
rect 10588 11190 10690 11226
rect 10810 11226 10912 11310
tri 10912 11226 11000 11314 sw
tri 11010 11226 11098 11314 ne
rect 11098 11310 11462 11314
rect 11098 11226 11240 11310
rect 10810 11190 11000 11226
rect 10588 11186 11000 11190
rect 10086 11138 10490 11186
rect 9586 11088 9988 11138
rect 9066 11058 9488 11088
rect 8574 11000 8968 11058
rect 8064 10960 8476 11000
tri 8476 10960 8516 11000 sw
tri 8574 10960 8614 11000 ne
rect 8614 10960 8968 11000
tri 8968 10960 9066 11058 sw
tri 9066 10960 9164 11058 ne
rect 9164 11000 9488 11058
tri 9488 11000 9576 11088 sw
tri 9586 11000 9674 11088 ne
rect 9674 11058 9988 11088
tri 9988 11058 10068 11138 sw
tri 10086 11058 10166 11138 ne
rect 10166 11088 10490 11138
tri 10490 11088 10588 11186 sw
tri 10588 11088 10686 11186 ne
rect 10686 11138 11000 11186
tri 11000 11138 11088 11226 sw
tri 11098 11138 11186 11226 ne
rect 11186 11190 11240 11226
rect 11360 11226 11462 11310
tri 11462 11226 11550 11314 sw
tri 11560 11226 11648 11314 ne
rect 11648 11310 12012 11314
rect 11648 11226 11790 11310
rect 11360 11190 11550 11226
rect 11186 11186 11550 11190
tri 11550 11186 11590 11226 sw
tri 11648 11186 11688 11226 ne
rect 11688 11190 11790 11226
rect 11910 11226 12012 11310
tri 12012 11226 12100 11314 sw
tri 12110 11226 12198 11314 ne
rect 12198 11310 12562 11314
rect 12198 11226 12340 11310
rect 11910 11190 12100 11226
rect 11688 11186 12100 11190
rect 11186 11138 11590 11186
rect 10686 11088 11088 11138
rect 10166 11058 10588 11088
rect 9674 11000 10068 11058
rect 9164 10960 9576 11000
tri 9576 10960 9616 11000 sw
tri 9674 10960 9714 11000 ne
rect 9714 10960 10068 11000
tri 10068 10960 10166 11058 sw
tri 10166 10960 10264 11058 ne
rect 10264 11000 10588 11058
tri 10588 11000 10676 11088 sw
tri 10686 11000 10774 11088 ne
rect 10774 11058 11088 11088
tri 11088 11058 11168 11138 sw
tri 11186 11058 11266 11138 ne
rect 11266 11088 11590 11138
tri 11590 11088 11688 11186 sw
tri 11688 11088 11786 11186 ne
rect 11786 11138 12100 11186
tri 12100 11138 12188 11226 sw
tri 12198 11138 12286 11226 ne
rect 12286 11190 12340 11226
rect 12460 11226 12562 11310
tri 12562 11226 12650 11314 sw
tri 12660 11226 12748 11314 ne
rect 12748 11310 13112 11314
rect 12748 11226 12890 11310
rect 12460 11190 12650 11226
rect 12286 11186 12650 11190
tri 12650 11186 12690 11226 sw
tri 12748 11186 12788 11226 ne
rect 12788 11190 12890 11226
rect 13010 11226 13112 11310
tri 13112 11226 13200 11314 sw
tri 13210 11226 13298 11314 ne
rect 13298 11310 15775 11314
rect 13298 11226 13440 11310
rect 13010 11190 13200 11226
rect 12788 11186 13200 11190
rect 12286 11138 12690 11186
rect 11786 11088 12188 11138
rect 11266 11058 11688 11088
rect 10774 11000 11168 11058
rect 10264 10960 10676 11000
tri 10676 10960 10716 11000 sw
tri 10774 10960 10814 11000 ne
rect 10814 10960 11168 11000
tri 11168 10960 11266 11058 sw
tri 11266 10960 11364 11058 ne
rect 11364 11000 11688 11058
tri 11688 11000 11776 11088 sw
tri 11786 11000 11874 11088 ne
rect 11874 11058 12188 11088
tri 12188 11058 12268 11138 sw
tri 12286 11058 12366 11138 ne
rect 12366 11088 12690 11138
tri 12690 11088 12788 11186 sw
tri 12788 11088 12886 11186 ne
rect 12886 11138 13200 11186
tri 13200 11138 13288 11226 sw
tri 13298 11138 13386 11226 ne
rect 13386 11190 13440 11226
rect 13560 11190 15775 11310
rect 13386 11138 15775 11190
rect 12886 11088 13288 11138
rect 12366 11058 12788 11088
rect 11874 11000 12268 11058
rect 11364 10960 11776 11000
tri 11776 10960 11816 11000 sw
tri 11874 10960 11914 11000 ne
rect 11914 10960 12268 11000
tri 12268 10960 12366 11058 sw
tri 12366 10960 12464 11058 ne
rect 12464 11000 12788 11058
tri 12788 11000 12876 11088 sw
tri 12886 11000 12974 11088 ne
rect 12974 11058 13288 11088
tri 13288 11058 13368 11138 sw
tri 13386 11058 13466 11138 ne
rect 13466 11058 14075 11138
rect 12974 11000 13368 11058
rect 12464 10960 12876 11000
tri 12876 10960 12916 11000 sw
tri 12974 10960 13014 11000 ne
rect 13014 10960 13368 11000
tri 13368 10960 13466 11058 sw
tri 13466 10960 13564 11058 ne
rect 13564 11038 14075 11058
rect 14175 11038 15775 11138
rect 13564 10960 15775 11038
rect -1025 10912 -284 10960
rect -1025 10812 -925 10912
rect -825 10862 -284 10912
tri -284 10862 -186 10960 sw
tri -186 10862 -88 10960 ne
rect -88 10862 266 10960
tri 266 10862 364 10960 sw
tri 364 10862 462 10960 ne
rect 462 10862 816 10960
tri 816 10862 914 10960 sw
tri 914 10862 1012 10960 ne
rect 1012 10862 1366 10960
tri 1366 10862 1464 10960 sw
tri 1464 10862 1562 10960 ne
rect 1562 10862 1916 10960
tri 1916 10862 2014 10960 sw
tri 2014 10862 2112 10960 ne
rect 2112 10862 2466 10960
tri 2466 10862 2564 10960 sw
tri 2564 10862 2662 10960 ne
rect 2662 10862 3016 10960
tri 3016 10862 3114 10960 sw
tri 3114 10862 3212 10960 ne
rect 3212 10862 3566 10960
tri 3566 10862 3664 10960 sw
tri 3664 10862 3762 10960 ne
rect 3762 10862 4116 10960
tri 4116 10862 4214 10960 sw
tri 4214 10862 4312 10960 ne
rect 4312 10862 4666 10960
tri 4666 10862 4764 10960 sw
tri 4764 10862 4862 10960 ne
rect 4862 10862 5216 10960
tri 5216 10862 5314 10960 sw
tri 5314 10862 5412 10960 ne
rect 5412 10862 5766 10960
tri 5766 10862 5864 10960 sw
tri 5864 10862 5962 10960 ne
rect 5962 10862 6316 10960
tri 6316 10862 6414 10960 sw
tri 6414 10862 6512 10960 ne
rect 6512 10862 6866 10960
tri 6866 10862 6964 10960 sw
tri 6964 10862 7062 10960 ne
rect 7062 10862 7416 10960
tri 7416 10862 7514 10960 sw
tri 7514 10862 7612 10960 ne
rect 7612 10862 7966 10960
tri 7966 10862 8064 10960 sw
tri 8064 10862 8162 10960 ne
rect 8162 10862 8516 10960
tri 8516 10862 8614 10960 sw
tri 8614 10862 8712 10960 ne
rect 8712 10862 9066 10960
tri 9066 10862 9164 10960 sw
tri 9164 10862 9262 10960 ne
rect 9262 10862 9616 10960
tri 9616 10862 9714 10960 sw
tri 9714 10862 9812 10960 ne
rect 9812 10862 10166 10960
tri 10166 10862 10264 10960 sw
tri 10264 10862 10362 10960 ne
rect 10362 10862 10716 10960
tri 10716 10862 10814 10960 sw
tri 10814 10862 10912 10960 ne
rect 10912 10862 11266 10960
tri 11266 10862 11364 10960 sw
tri 11364 10862 11462 10960 ne
rect 11462 10862 11816 10960
tri 11816 10862 11914 10960 sw
tri 11914 10862 12012 10960 ne
rect 12012 10862 12366 10960
tri 12366 10862 12464 10960 sw
tri 12464 10862 12562 10960 ne
rect 12562 10862 12916 10960
tri 12916 10862 13014 10960 sw
tri 13014 10862 13112 10960 ne
rect 13112 10862 13466 10960
tri 13466 10862 13564 10960 sw
tri 13564 10862 13662 10960 ne
rect 13662 10862 15775 10960
rect -825 10812 -186 10862
rect -1025 10764 -186 10812
tri -186 10764 -88 10862 sw
tri -88 10764 10 10862 ne
rect 10 10764 364 10862
tri 364 10764 462 10862 sw
tri 462 10764 560 10862 ne
rect 560 10764 914 10862
tri 914 10764 1012 10862 sw
tri 1012 10764 1110 10862 ne
rect 1110 10764 1464 10862
tri 1464 10764 1562 10862 sw
tri 1562 10764 1660 10862 ne
rect 1660 10764 2014 10862
tri 2014 10764 2112 10862 sw
tri 2112 10764 2210 10862 ne
rect 2210 10764 2564 10862
tri 2564 10764 2662 10862 sw
tri 2662 10764 2760 10862 ne
rect 2760 10764 3114 10862
tri 3114 10764 3212 10862 sw
tri 3212 10764 3310 10862 ne
rect 3310 10764 3664 10862
tri 3664 10764 3762 10862 sw
tri 3762 10764 3860 10862 ne
rect 3860 10764 4214 10862
tri 4214 10764 4312 10862 sw
tri 4312 10764 4410 10862 ne
rect 4410 10764 4764 10862
tri 4764 10764 4862 10862 sw
tri 4862 10764 4960 10862 ne
rect 4960 10764 5314 10862
tri 5314 10764 5412 10862 sw
tri 5412 10764 5510 10862 ne
rect 5510 10764 5864 10862
tri 5864 10764 5962 10862 sw
tri 5962 10764 6060 10862 ne
rect 6060 10764 6414 10862
tri 6414 10764 6512 10862 sw
tri 6512 10764 6610 10862 ne
rect 6610 10764 6964 10862
tri 6964 10764 7062 10862 sw
tri 7062 10764 7160 10862 ne
rect 7160 10764 7514 10862
tri 7514 10764 7612 10862 sw
tri 7612 10764 7710 10862 ne
rect 7710 10764 8064 10862
tri 8064 10764 8162 10862 sw
tri 8162 10764 8260 10862 ne
rect 8260 10764 8614 10862
tri 8614 10764 8712 10862 sw
tri 8712 10764 8810 10862 ne
rect 8810 10764 9164 10862
tri 9164 10764 9262 10862 sw
tri 9262 10764 9360 10862 ne
rect 9360 10764 9714 10862
tri 9714 10764 9812 10862 sw
tri 9812 10764 9910 10862 ne
rect 9910 10764 10264 10862
tri 10264 10764 10362 10862 sw
tri 10362 10764 10460 10862 ne
rect 10460 10764 10814 10862
tri 10814 10764 10912 10862 sw
tri 10912 10764 11010 10862 ne
rect 11010 10764 11364 10862
tri 11364 10764 11462 10862 sw
tri 11462 10764 11560 10862 ne
rect 11560 10764 11914 10862
tri 11914 10764 12012 10862 sw
tri 12012 10764 12110 10862 ne
rect 12110 10764 12464 10862
tri 12464 10764 12562 10862 sw
tri 12562 10764 12660 10862 ne
rect 12660 10764 13014 10862
tri 13014 10764 13112 10862 sw
tri 13112 10764 13210 10862 ne
rect 13210 10764 13564 10862
tri 13564 10764 13662 10862 sw
rect -1025 10760 -88 10764
rect -1025 10640 -310 10760
rect -190 10676 -88 10760
tri -88 10676 0 10764 sw
tri 10 10676 98 10764 ne
rect 98 10760 462 10764
rect 98 10676 240 10760
rect -190 10640 0 10676
rect -1025 10636 0 10640
tri 0 10636 40 10676 sw
tri 98 10636 138 10676 ne
rect 138 10640 240 10676
rect 360 10676 462 10760
tri 462 10676 550 10764 sw
tri 560 10676 648 10764 ne
rect 648 10760 1012 10764
rect 648 10676 790 10760
rect 360 10640 550 10676
rect 138 10636 550 10640
tri -412 10538 -314 10636 ne
rect -314 10538 40 10636
tri 40 10538 138 10636 sw
tri 138 10538 236 10636 ne
rect 236 10588 550 10636
tri 550 10588 638 10676 sw
tri 648 10588 736 10676 ne
rect 736 10640 790 10676
rect 910 10676 1012 10760
tri 1012 10676 1100 10764 sw
tri 1110 10676 1198 10764 ne
rect 1198 10760 1562 10764
rect 1198 10676 1340 10760
rect 910 10640 1100 10676
rect 736 10636 1100 10640
tri 1100 10636 1140 10676 sw
tri 1198 10636 1238 10676 ne
rect 1238 10640 1340 10676
rect 1460 10676 1562 10760
tri 1562 10676 1650 10764 sw
tri 1660 10676 1748 10764 ne
rect 1748 10760 2112 10764
rect 1748 10676 1890 10760
rect 1460 10640 1650 10676
rect 1238 10636 1650 10640
rect 736 10588 1140 10636
rect 236 10538 638 10588
rect -2525 10450 -412 10538
tri -412 10450 -324 10538 sw
tri -314 10450 -226 10538 ne
rect -226 10450 138 10538
tri 138 10450 226 10538 sw
tri 236 10450 324 10538 ne
rect 324 10508 638 10538
tri 638 10508 718 10588 sw
tri 736 10508 816 10588 ne
rect 816 10538 1140 10588
tri 1140 10538 1238 10636 sw
tri 1238 10538 1336 10636 ne
rect 1336 10588 1650 10636
tri 1650 10588 1738 10676 sw
tri 1748 10588 1836 10676 ne
rect 1836 10640 1890 10676
rect 2010 10676 2112 10760
tri 2112 10676 2200 10764 sw
tri 2210 10676 2298 10764 ne
rect 2298 10760 2662 10764
rect 2298 10676 2440 10760
rect 2010 10640 2200 10676
rect 1836 10636 2200 10640
tri 2200 10636 2240 10676 sw
tri 2298 10636 2338 10676 ne
rect 2338 10640 2440 10676
rect 2560 10676 2662 10760
tri 2662 10676 2750 10764 sw
tri 2760 10676 2848 10764 ne
rect 2848 10760 3212 10764
rect 2848 10676 2990 10760
rect 2560 10640 2750 10676
rect 2338 10636 2750 10640
rect 1836 10588 2240 10636
rect 1336 10538 1738 10588
rect 816 10508 1238 10538
rect 324 10450 718 10508
rect -2525 10410 -324 10450
tri -324 10410 -284 10450 sw
tri -226 10410 -186 10450 ne
rect -186 10410 226 10450
tri 226 10410 266 10450 sw
tri 324 10410 364 10450 ne
rect 364 10410 718 10450
tri 718 10410 816 10508 sw
tri 816 10410 914 10508 ne
rect 914 10450 1238 10508
tri 1238 10450 1326 10538 sw
tri 1336 10450 1424 10538 ne
rect 1424 10508 1738 10538
tri 1738 10508 1818 10588 sw
tri 1836 10508 1916 10588 ne
rect 1916 10538 2240 10588
tri 2240 10538 2338 10636 sw
tri 2338 10538 2436 10636 ne
rect 2436 10588 2750 10636
tri 2750 10588 2838 10676 sw
tri 2848 10588 2936 10676 ne
rect 2936 10640 2990 10676
rect 3110 10676 3212 10760
tri 3212 10676 3300 10764 sw
tri 3310 10676 3398 10764 ne
rect 3398 10760 3762 10764
rect 3398 10676 3540 10760
rect 3110 10640 3300 10676
rect 2936 10636 3300 10640
tri 3300 10636 3340 10676 sw
tri 3398 10636 3438 10676 ne
rect 3438 10640 3540 10676
rect 3660 10676 3762 10760
tri 3762 10676 3850 10764 sw
tri 3860 10676 3948 10764 ne
rect 3948 10760 4312 10764
rect 3948 10676 4090 10760
rect 3660 10640 3850 10676
rect 3438 10636 3850 10640
rect 2936 10588 3340 10636
rect 2436 10538 2838 10588
rect 1916 10508 2338 10538
rect 1424 10450 1818 10508
rect 914 10410 1326 10450
tri 1326 10410 1366 10450 sw
tri 1424 10410 1464 10450 ne
rect 1464 10410 1818 10450
tri 1818 10410 1916 10508 sw
tri 1916 10410 2014 10508 ne
rect 2014 10450 2338 10508
tri 2338 10450 2426 10538 sw
tri 2436 10450 2524 10538 ne
rect 2524 10508 2838 10538
tri 2838 10508 2918 10588 sw
tri 2936 10508 3016 10588 ne
rect 3016 10538 3340 10588
tri 3340 10538 3438 10636 sw
tri 3438 10538 3536 10636 ne
rect 3536 10588 3850 10636
tri 3850 10588 3938 10676 sw
tri 3948 10588 4036 10676 ne
rect 4036 10640 4090 10676
rect 4210 10676 4312 10760
tri 4312 10676 4400 10764 sw
tri 4410 10676 4498 10764 ne
rect 4498 10760 4862 10764
rect 4498 10676 4640 10760
rect 4210 10640 4400 10676
rect 4036 10636 4400 10640
tri 4400 10636 4440 10676 sw
tri 4498 10636 4538 10676 ne
rect 4538 10640 4640 10676
rect 4760 10676 4862 10760
tri 4862 10676 4950 10764 sw
tri 4960 10676 5048 10764 ne
rect 5048 10760 5412 10764
rect 5048 10676 5190 10760
rect 4760 10640 4950 10676
rect 4538 10636 4950 10640
rect 4036 10588 4440 10636
rect 3536 10538 3938 10588
rect 3016 10508 3438 10538
rect 2524 10450 2918 10508
rect 2014 10410 2426 10450
tri 2426 10410 2466 10450 sw
tri 2524 10410 2564 10450 ne
rect 2564 10410 2918 10450
tri 2918 10410 3016 10508 sw
tri 3016 10410 3114 10508 ne
rect 3114 10450 3438 10508
tri 3438 10450 3526 10538 sw
tri 3536 10450 3624 10538 ne
rect 3624 10508 3938 10538
tri 3938 10508 4018 10588 sw
tri 4036 10508 4116 10588 ne
rect 4116 10538 4440 10588
tri 4440 10538 4538 10636 sw
tri 4538 10538 4636 10636 ne
rect 4636 10588 4950 10636
tri 4950 10588 5038 10676 sw
tri 5048 10588 5136 10676 ne
rect 5136 10640 5190 10676
rect 5310 10676 5412 10760
tri 5412 10676 5500 10764 sw
tri 5510 10676 5598 10764 ne
rect 5598 10760 5962 10764
rect 5598 10676 5740 10760
rect 5310 10640 5500 10676
rect 5136 10636 5500 10640
tri 5500 10636 5540 10676 sw
tri 5598 10636 5638 10676 ne
rect 5638 10640 5740 10676
rect 5860 10676 5962 10760
tri 5962 10676 6050 10764 sw
tri 6060 10676 6148 10764 ne
rect 6148 10760 6512 10764
rect 6148 10676 6290 10760
rect 5860 10640 6050 10676
rect 5638 10636 6050 10640
rect 5136 10588 5540 10636
rect 4636 10538 5038 10588
rect 4116 10508 4538 10538
rect 3624 10450 4018 10508
rect 3114 10410 3526 10450
tri 3526 10410 3566 10450 sw
tri 3624 10410 3664 10450 ne
rect 3664 10410 4018 10450
tri 4018 10410 4116 10508 sw
tri 4116 10410 4214 10508 ne
rect 4214 10450 4538 10508
tri 4538 10450 4626 10538 sw
tri 4636 10450 4724 10538 ne
rect 4724 10508 5038 10538
tri 5038 10508 5118 10588 sw
tri 5136 10508 5216 10588 ne
rect 5216 10538 5540 10588
tri 5540 10538 5638 10636 sw
tri 5638 10538 5736 10636 ne
rect 5736 10588 6050 10636
tri 6050 10588 6138 10676 sw
tri 6148 10588 6236 10676 ne
rect 6236 10640 6290 10676
rect 6410 10676 6512 10760
tri 6512 10676 6600 10764 sw
tri 6610 10676 6698 10764 ne
rect 6698 10760 7062 10764
rect 6698 10676 6840 10760
rect 6410 10640 6600 10676
rect 6236 10636 6600 10640
tri 6600 10636 6640 10676 sw
tri 6698 10636 6738 10676 ne
rect 6738 10640 6840 10676
rect 6960 10676 7062 10760
tri 7062 10676 7150 10764 sw
tri 7160 10676 7248 10764 ne
rect 7248 10760 7612 10764
rect 7248 10676 7390 10760
rect 6960 10640 7150 10676
rect 6738 10636 7150 10640
rect 6236 10588 6640 10636
rect 5736 10538 6138 10588
rect 5216 10508 5638 10538
rect 4724 10450 5118 10508
rect 4214 10410 4626 10450
tri 4626 10410 4666 10450 sw
tri 4724 10410 4764 10450 ne
rect 4764 10410 5118 10450
tri 5118 10410 5216 10508 sw
tri 5216 10410 5314 10508 ne
rect 5314 10450 5638 10508
tri 5638 10450 5726 10538 sw
tri 5736 10450 5824 10538 ne
rect 5824 10508 6138 10538
tri 6138 10508 6218 10588 sw
tri 6236 10508 6316 10588 ne
rect 6316 10538 6640 10588
tri 6640 10538 6738 10636 sw
tri 6738 10538 6836 10636 ne
rect 6836 10588 7150 10636
tri 7150 10588 7238 10676 sw
tri 7248 10588 7336 10676 ne
rect 7336 10640 7390 10676
rect 7510 10676 7612 10760
tri 7612 10676 7700 10764 sw
tri 7710 10676 7798 10764 ne
rect 7798 10760 8162 10764
rect 7798 10676 7940 10760
rect 7510 10640 7700 10676
rect 7336 10636 7700 10640
tri 7700 10636 7740 10676 sw
tri 7798 10636 7838 10676 ne
rect 7838 10640 7940 10676
rect 8060 10676 8162 10760
tri 8162 10676 8250 10764 sw
tri 8260 10676 8348 10764 ne
rect 8348 10760 8712 10764
rect 8348 10676 8490 10760
rect 8060 10640 8250 10676
rect 7838 10636 8250 10640
rect 7336 10588 7740 10636
rect 6836 10538 7238 10588
rect 6316 10508 6738 10538
rect 5824 10450 6218 10508
rect 5314 10410 5726 10450
tri 5726 10410 5766 10450 sw
tri 5824 10410 5864 10450 ne
rect 5864 10410 6218 10450
tri 6218 10410 6316 10508 sw
tri 6316 10410 6414 10508 ne
rect 6414 10450 6738 10508
tri 6738 10450 6826 10538 sw
tri 6836 10450 6924 10538 ne
rect 6924 10508 7238 10538
tri 7238 10508 7318 10588 sw
tri 7336 10508 7416 10588 ne
rect 7416 10538 7740 10588
tri 7740 10538 7838 10636 sw
tri 7838 10538 7936 10636 ne
rect 7936 10588 8250 10636
tri 8250 10588 8338 10676 sw
tri 8348 10588 8436 10676 ne
rect 8436 10640 8490 10676
rect 8610 10676 8712 10760
tri 8712 10676 8800 10764 sw
tri 8810 10676 8898 10764 ne
rect 8898 10760 9262 10764
rect 8898 10676 9040 10760
rect 8610 10640 8800 10676
rect 8436 10636 8800 10640
tri 8800 10636 8840 10676 sw
tri 8898 10636 8938 10676 ne
rect 8938 10640 9040 10676
rect 9160 10676 9262 10760
tri 9262 10676 9350 10764 sw
tri 9360 10676 9448 10764 ne
rect 9448 10760 9812 10764
rect 9448 10676 9590 10760
rect 9160 10640 9350 10676
rect 8938 10636 9350 10640
rect 8436 10588 8840 10636
rect 7936 10538 8338 10588
rect 7416 10508 7838 10538
rect 6924 10450 7318 10508
rect 6414 10410 6826 10450
tri 6826 10410 6866 10450 sw
tri 6924 10410 6964 10450 ne
rect 6964 10410 7318 10450
tri 7318 10410 7416 10508 sw
tri 7416 10410 7514 10508 ne
rect 7514 10450 7838 10508
tri 7838 10450 7926 10538 sw
tri 7936 10450 8024 10538 ne
rect 8024 10508 8338 10538
tri 8338 10508 8418 10588 sw
tri 8436 10508 8516 10588 ne
rect 8516 10538 8840 10588
tri 8840 10538 8938 10636 sw
tri 8938 10538 9036 10636 ne
rect 9036 10588 9350 10636
tri 9350 10588 9438 10676 sw
tri 9448 10588 9536 10676 ne
rect 9536 10640 9590 10676
rect 9710 10676 9812 10760
tri 9812 10676 9900 10764 sw
tri 9910 10676 9998 10764 ne
rect 9998 10760 10362 10764
rect 9998 10676 10140 10760
rect 9710 10640 9900 10676
rect 9536 10636 9900 10640
tri 9900 10636 9940 10676 sw
tri 9998 10636 10038 10676 ne
rect 10038 10640 10140 10676
rect 10260 10676 10362 10760
tri 10362 10676 10450 10764 sw
tri 10460 10676 10548 10764 ne
rect 10548 10760 10912 10764
rect 10548 10676 10690 10760
rect 10260 10640 10450 10676
rect 10038 10636 10450 10640
rect 9536 10588 9940 10636
rect 9036 10538 9438 10588
rect 8516 10508 8938 10538
rect 8024 10450 8418 10508
rect 7514 10410 7926 10450
tri 7926 10410 7966 10450 sw
tri 8024 10410 8064 10450 ne
rect 8064 10410 8418 10450
tri 8418 10410 8516 10508 sw
tri 8516 10410 8614 10508 ne
rect 8614 10450 8938 10508
tri 8938 10450 9026 10538 sw
tri 9036 10450 9124 10538 ne
rect 9124 10508 9438 10538
tri 9438 10508 9518 10588 sw
tri 9536 10508 9616 10588 ne
rect 9616 10538 9940 10588
tri 9940 10538 10038 10636 sw
tri 10038 10538 10136 10636 ne
rect 10136 10588 10450 10636
tri 10450 10588 10538 10676 sw
tri 10548 10588 10636 10676 ne
rect 10636 10640 10690 10676
rect 10810 10676 10912 10760
tri 10912 10676 11000 10764 sw
tri 11010 10676 11098 10764 ne
rect 11098 10760 11462 10764
rect 11098 10676 11240 10760
rect 10810 10640 11000 10676
rect 10636 10636 11000 10640
tri 11000 10636 11040 10676 sw
tri 11098 10636 11138 10676 ne
rect 11138 10640 11240 10676
rect 11360 10676 11462 10760
tri 11462 10676 11550 10764 sw
tri 11560 10676 11648 10764 ne
rect 11648 10760 12012 10764
rect 11648 10676 11790 10760
rect 11360 10640 11550 10676
rect 11138 10636 11550 10640
rect 10636 10588 11040 10636
rect 10136 10538 10538 10588
rect 9616 10508 10038 10538
rect 9124 10450 9518 10508
rect 8614 10410 9026 10450
tri 9026 10410 9066 10450 sw
tri 9124 10410 9164 10450 ne
rect 9164 10410 9518 10450
tri 9518 10410 9616 10508 sw
tri 9616 10410 9714 10508 ne
rect 9714 10450 10038 10508
tri 10038 10450 10126 10538 sw
tri 10136 10450 10224 10538 ne
rect 10224 10508 10538 10538
tri 10538 10508 10618 10588 sw
tri 10636 10508 10716 10588 ne
rect 10716 10538 11040 10588
tri 11040 10538 11138 10636 sw
tri 11138 10538 11236 10636 ne
rect 11236 10588 11550 10636
tri 11550 10588 11638 10676 sw
tri 11648 10588 11736 10676 ne
rect 11736 10640 11790 10676
rect 11910 10676 12012 10760
tri 12012 10676 12100 10764 sw
tri 12110 10676 12198 10764 ne
rect 12198 10760 12562 10764
rect 12198 10676 12340 10760
rect 11910 10640 12100 10676
rect 11736 10636 12100 10640
tri 12100 10636 12140 10676 sw
tri 12198 10636 12238 10676 ne
rect 12238 10640 12340 10676
rect 12460 10676 12562 10760
tri 12562 10676 12650 10764 sw
tri 12660 10676 12748 10764 ne
rect 12748 10760 13112 10764
rect 12748 10676 12890 10760
rect 12460 10640 12650 10676
rect 12238 10636 12650 10640
rect 11736 10588 12140 10636
rect 11236 10538 11638 10588
rect 10716 10508 11138 10538
rect 10224 10450 10618 10508
rect 9714 10410 10126 10450
tri 10126 10410 10166 10450 sw
tri 10224 10410 10264 10450 ne
rect 10264 10410 10618 10450
tri 10618 10410 10716 10508 sw
tri 10716 10410 10814 10508 ne
rect 10814 10450 11138 10508
tri 11138 10450 11226 10538 sw
tri 11236 10450 11324 10538 ne
rect 11324 10508 11638 10538
tri 11638 10508 11718 10588 sw
tri 11736 10508 11816 10588 ne
rect 11816 10538 12140 10588
tri 12140 10538 12238 10636 sw
tri 12238 10538 12336 10636 ne
rect 12336 10588 12650 10636
tri 12650 10588 12738 10676 sw
tri 12748 10588 12836 10676 ne
rect 12836 10640 12890 10676
rect 13010 10676 13112 10760
tri 13112 10676 13200 10764 sw
tri 13210 10676 13298 10764 ne
rect 13298 10760 14275 10764
rect 13298 10676 13440 10760
rect 13010 10640 13200 10676
rect 12836 10636 13200 10640
tri 13200 10636 13240 10676 sw
tri 13298 10636 13338 10676 ne
rect 13338 10640 13440 10676
rect 13560 10640 14275 10760
rect 13338 10636 14275 10640
rect 12836 10588 13240 10636
rect 12336 10538 12738 10588
rect 11816 10508 12238 10538
rect 11324 10450 11718 10508
rect 10814 10410 11226 10450
tri 11226 10410 11266 10450 sw
tri 11324 10410 11364 10450 ne
rect 11364 10410 11718 10450
tri 11718 10410 11816 10508 sw
tri 11816 10410 11914 10508 ne
rect 11914 10450 12238 10508
tri 12238 10450 12326 10538 sw
tri 12336 10450 12424 10538 ne
rect 12424 10508 12738 10538
tri 12738 10508 12818 10588 sw
tri 12836 10508 12916 10588 ne
rect 12916 10538 13240 10588
tri 13240 10538 13338 10636 sw
tri 13338 10538 13436 10636 ne
rect 13436 10538 14275 10636
rect 12916 10508 13338 10538
rect 12424 10450 12818 10508
rect 11914 10410 12326 10450
tri 12326 10410 12366 10450 sw
tri 12424 10410 12464 10450 ne
rect 12464 10410 12818 10450
tri 12818 10410 12916 10508 sw
tri 12916 10410 13014 10508 ne
rect 13014 10450 13338 10508
tri 13338 10450 13426 10538 sw
tri 13436 10450 13524 10538 ne
rect 13524 10450 14275 10538
rect 13014 10410 13426 10450
tri 13426 10410 13466 10450 sw
tri 13524 10410 13564 10450 ne
rect 13564 10410 14275 10450
rect -2525 10312 -284 10410
tri -284 10312 -186 10410 sw
tri -186 10312 -88 10410 ne
rect -88 10312 266 10410
tri 266 10312 364 10410 sw
tri 364 10312 462 10410 ne
rect 462 10312 816 10410
tri 816 10312 914 10410 sw
tri 914 10312 1012 10410 ne
rect 1012 10312 1366 10410
tri 1366 10312 1464 10410 sw
tri 1464 10312 1562 10410 ne
rect 1562 10312 1916 10410
tri 1916 10312 2014 10410 sw
tri 2014 10312 2112 10410 ne
rect 2112 10312 2466 10410
tri 2466 10312 2564 10410 sw
tri 2564 10312 2662 10410 ne
rect 2662 10312 3016 10410
tri 3016 10312 3114 10410 sw
tri 3114 10312 3212 10410 ne
rect 3212 10312 3566 10410
tri 3566 10312 3664 10410 sw
tri 3664 10312 3762 10410 ne
rect 3762 10312 4116 10410
tri 4116 10312 4214 10410 sw
tri 4214 10312 4312 10410 ne
rect 4312 10312 4666 10410
tri 4666 10312 4764 10410 sw
tri 4764 10312 4862 10410 ne
rect 4862 10312 5216 10410
tri 5216 10312 5314 10410 sw
tri 5314 10312 5412 10410 ne
rect 5412 10312 5766 10410
tri 5766 10312 5864 10410 sw
tri 5864 10312 5962 10410 ne
rect 5962 10312 6316 10410
tri 6316 10312 6414 10410 sw
tri 6414 10312 6512 10410 ne
rect 6512 10312 6866 10410
tri 6866 10312 6964 10410 sw
tri 6964 10312 7062 10410 ne
rect 7062 10312 7416 10410
tri 7416 10312 7514 10410 sw
tri 7514 10312 7612 10410 ne
rect 7612 10312 7966 10410
tri 7966 10312 8064 10410 sw
tri 8064 10312 8162 10410 ne
rect 8162 10312 8516 10410
tri 8516 10312 8614 10410 sw
tri 8614 10312 8712 10410 ne
rect 8712 10312 9066 10410
tri 9066 10312 9164 10410 sw
tri 9164 10312 9262 10410 ne
rect 9262 10312 9616 10410
tri 9616 10312 9714 10410 sw
tri 9714 10312 9812 10410 ne
rect 9812 10312 10166 10410
tri 10166 10312 10264 10410 sw
tri 10264 10312 10362 10410 ne
rect 10362 10312 10716 10410
tri 10716 10312 10814 10410 sw
tri 10814 10312 10912 10410 ne
rect 10912 10312 11266 10410
tri 11266 10312 11364 10410 sw
tri 11364 10312 11462 10410 ne
rect 11462 10312 11816 10410
tri 11816 10312 11914 10410 sw
tri 11914 10312 12012 10410 ne
rect 12012 10312 12366 10410
tri 12366 10312 12464 10410 sw
tri 12464 10312 12562 10410 ne
rect 12562 10312 12916 10410
tri 12916 10312 13014 10410 sw
tri 13014 10312 13112 10410 ne
rect 13112 10312 13466 10410
tri 13466 10312 13564 10410 sw
tri 13564 10312 13662 10410 ne
rect 13662 10312 14275 10410
rect -2525 10214 -186 10312
tri -186 10214 -88 10312 sw
tri -88 10214 10 10312 ne
rect 10 10214 364 10312
tri 364 10214 462 10312 sw
tri 462 10214 560 10312 ne
rect 560 10214 914 10312
tri 914 10214 1012 10312 sw
tri 1012 10214 1110 10312 ne
rect 1110 10214 1464 10312
tri 1464 10214 1562 10312 sw
tri 1562 10214 1660 10312 ne
rect 1660 10214 2014 10312
tri 2014 10214 2112 10312 sw
tri 2112 10214 2210 10312 ne
rect 2210 10214 2564 10312
tri 2564 10214 2662 10312 sw
tri 2662 10214 2760 10312 ne
rect 2760 10214 3114 10312
tri 3114 10214 3212 10312 sw
tri 3212 10214 3310 10312 ne
rect 3310 10214 3664 10312
tri 3664 10214 3762 10312 sw
tri 3762 10214 3860 10312 ne
rect 3860 10214 4214 10312
tri 4214 10214 4312 10312 sw
tri 4312 10214 4410 10312 ne
rect 4410 10214 4764 10312
tri 4764 10214 4862 10312 sw
tri 4862 10214 4960 10312 ne
rect 4960 10214 5314 10312
tri 5314 10214 5412 10312 sw
tri 5412 10214 5510 10312 ne
rect 5510 10214 5864 10312
tri 5864 10214 5962 10312 sw
tri 5962 10214 6060 10312 ne
rect 6060 10214 6414 10312
tri 6414 10214 6512 10312 sw
tri 6512 10214 6610 10312 ne
rect 6610 10214 6964 10312
tri 6964 10214 7062 10312 sw
tri 7062 10214 7160 10312 ne
rect 7160 10214 7514 10312
tri 7514 10214 7612 10312 sw
tri 7612 10214 7710 10312 ne
rect 7710 10214 8064 10312
tri 8064 10214 8162 10312 sw
tri 8162 10214 8260 10312 ne
rect 8260 10214 8614 10312
tri 8614 10214 8712 10312 sw
tri 8712 10214 8810 10312 ne
rect 8810 10214 9164 10312
tri 9164 10214 9262 10312 sw
tri 9262 10214 9360 10312 ne
rect 9360 10214 9714 10312
tri 9714 10214 9812 10312 sw
tri 9812 10214 9910 10312 ne
rect 9910 10214 10264 10312
tri 10264 10214 10362 10312 sw
tri 10362 10214 10460 10312 ne
rect 10460 10214 10814 10312
tri 10814 10214 10912 10312 sw
tri 10912 10214 11010 10312 ne
rect 11010 10214 11364 10312
tri 11364 10214 11462 10312 sw
tri 11462 10214 11560 10312 ne
rect 11560 10214 11914 10312
tri 11914 10214 12012 10312 sw
tri 12012 10214 12110 10312 ne
rect 12110 10214 12464 10312
tri 12464 10214 12562 10312 sw
tri 12562 10214 12660 10312 ne
rect 12660 10214 13014 10312
tri 13014 10214 13112 10312 sw
tri 13112 10214 13210 10312 ne
rect 13210 10214 13564 10312
tri 13564 10214 13662 10312 sw
rect 14775 10214 15775 10862
rect -2525 10210 -88 10214
rect -2525 10090 -310 10210
rect -190 10126 -88 10210
tri -88 10126 0 10214 sw
tri 10 10126 98 10214 ne
rect 98 10210 462 10214
rect 98 10126 240 10210
rect -190 10090 0 10126
rect -2525 10086 0 10090
rect -2525 9438 -1525 10086
tri -412 9988 -314 10086 ne
rect -314 10038 0 10086
tri 0 10038 88 10126 sw
tri 98 10038 186 10126 ne
rect 186 10090 240 10126
rect 360 10126 462 10210
tri 462 10126 550 10214 sw
tri 560 10126 648 10214 ne
rect 648 10210 1012 10214
rect 648 10126 790 10210
rect 360 10090 550 10126
rect 186 10086 550 10090
tri 550 10086 590 10126 sw
tri 648 10086 688 10126 ne
rect 688 10090 790 10126
rect 910 10126 1012 10210
tri 1012 10126 1100 10214 sw
tri 1110 10126 1198 10214 ne
rect 1198 10210 1562 10214
rect 1198 10126 1340 10210
rect 910 10090 1100 10126
rect 688 10086 1100 10090
rect 186 10038 590 10086
rect -314 9988 88 10038
rect -1025 9900 -412 9988
tri -412 9900 -324 9988 sw
tri -314 9900 -226 9988 ne
rect -226 9958 88 9988
tri 88 9958 168 10038 sw
tri 186 9958 266 10038 ne
rect 266 9988 590 10038
tri 590 9988 688 10086 sw
tri 688 9988 786 10086 ne
rect 786 10038 1100 10086
tri 1100 10038 1188 10126 sw
tri 1198 10038 1286 10126 ne
rect 1286 10090 1340 10126
rect 1460 10126 1562 10210
tri 1562 10126 1650 10214 sw
tri 1660 10126 1748 10214 ne
rect 1748 10210 2112 10214
rect 1748 10126 1890 10210
rect 1460 10090 1650 10126
rect 1286 10086 1650 10090
tri 1650 10086 1690 10126 sw
tri 1748 10086 1788 10126 ne
rect 1788 10090 1890 10126
rect 2010 10126 2112 10210
tri 2112 10126 2200 10214 sw
tri 2210 10126 2298 10214 ne
rect 2298 10210 2662 10214
rect 2298 10126 2440 10210
rect 2010 10090 2200 10126
rect 1788 10086 2200 10090
rect 1286 10038 1690 10086
rect 786 9988 1188 10038
rect 266 9958 688 9988
rect -226 9900 168 9958
rect -1025 9860 -324 9900
tri -324 9860 -284 9900 sw
tri -226 9860 -186 9900 ne
rect -186 9860 168 9900
tri 168 9860 266 9958 sw
tri 266 9860 364 9958 ne
rect 364 9900 688 9958
tri 688 9900 776 9988 sw
tri 786 9900 874 9988 ne
rect 874 9958 1188 9988
tri 1188 9958 1268 10038 sw
tri 1286 9958 1366 10038 ne
rect 1366 9988 1690 10038
tri 1690 9988 1788 10086 sw
tri 1788 9988 1886 10086 ne
rect 1886 10038 2200 10086
tri 2200 10038 2288 10126 sw
tri 2298 10038 2386 10126 ne
rect 2386 10090 2440 10126
rect 2560 10126 2662 10210
tri 2662 10126 2750 10214 sw
tri 2760 10126 2848 10214 ne
rect 2848 10210 3212 10214
rect 2848 10126 2990 10210
rect 2560 10090 2750 10126
rect 2386 10086 2750 10090
tri 2750 10086 2790 10126 sw
tri 2848 10086 2888 10126 ne
rect 2888 10090 2990 10126
rect 3110 10126 3212 10210
tri 3212 10126 3300 10214 sw
tri 3310 10126 3398 10214 ne
rect 3398 10210 3762 10214
rect 3398 10126 3540 10210
rect 3110 10090 3300 10126
rect 2888 10086 3300 10090
rect 2386 10038 2790 10086
rect 1886 9988 2288 10038
rect 1366 9958 1788 9988
rect 874 9900 1268 9958
rect 364 9860 776 9900
tri 776 9860 816 9900 sw
tri 874 9860 914 9900 ne
rect 914 9860 1268 9900
tri 1268 9860 1366 9958 sw
tri 1366 9860 1464 9958 ne
rect 1464 9900 1788 9958
tri 1788 9900 1876 9988 sw
tri 1886 9900 1974 9988 ne
rect 1974 9958 2288 9988
tri 2288 9958 2368 10038 sw
tri 2386 9958 2466 10038 ne
rect 2466 9988 2790 10038
tri 2790 9988 2888 10086 sw
tri 2888 9988 2986 10086 ne
rect 2986 10038 3300 10086
tri 3300 10038 3388 10126 sw
tri 3398 10038 3486 10126 ne
rect 3486 10090 3540 10126
rect 3660 10126 3762 10210
tri 3762 10126 3850 10214 sw
tri 3860 10126 3948 10214 ne
rect 3948 10210 4312 10214
rect 3948 10126 4090 10210
rect 3660 10090 3850 10126
rect 3486 10086 3850 10090
tri 3850 10086 3890 10126 sw
tri 3948 10086 3988 10126 ne
rect 3988 10090 4090 10126
rect 4210 10126 4312 10210
tri 4312 10126 4400 10214 sw
tri 4410 10126 4498 10214 ne
rect 4498 10210 4862 10214
rect 4498 10126 4640 10210
rect 4210 10090 4400 10126
rect 3988 10086 4400 10090
rect 3486 10038 3890 10086
rect 2986 9988 3388 10038
rect 2466 9958 2888 9988
rect 1974 9900 2368 9958
rect 1464 9860 1876 9900
tri 1876 9860 1916 9900 sw
tri 1974 9860 2014 9900 ne
rect 2014 9860 2368 9900
tri 2368 9860 2466 9958 sw
tri 2466 9860 2564 9958 ne
rect 2564 9900 2888 9958
tri 2888 9900 2976 9988 sw
tri 2986 9900 3074 9988 ne
rect 3074 9958 3388 9988
tri 3388 9958 3468 10038 sw
tri 3486 9958 3566 10038 ne
rect 3566 9988 3890 10038
tri 3890 9988 3988 10086 sw
tri 3988 9988 4086 10086 ne
rect 4086 10038 4400 10086
tri 4400 10038 4488 10126 sw
tri 4498 10038 4586 10126 ne
rect 4586 10090 4640 10126
rect 4760 10126 4862 10210
tri 4862 10126 4950 10214 sw
tri 4960 10126 5048 10214 ne
rect 5048 10210 5412 10214
rect 5048 10126 5190 10210
rect 4760 10090 4950 10126
rect 4586 10086 4950 10090
tri 4950 10086 4990 10126 sw
tri 5048 10086 5088 10126 ne
rect 5088 10090 5190 10126
rect 5310 10126 5412 10210
tri 5412 10126 5500 10214 sw
tri 5510 10126 5598 10214 ne
rect 5598 10210 5962 10214
rect 5598 10126 5740 10210
rect 5310 10090 5500 10126
rect 5088 10086 5500 10090
rect 4586 10038 4990 10086
rect 4086 9988 4488 10038
rect 3566 9958 3988 9988
rect 3074 9900 3468 9958
rect 2564 9860 2976 9900
tri 2976 9860 3016 9900 sw
tri 3074 9860 3114 9900 ne
rect 3114 9860 3468 9900
tri 3468 9860 3566 9958 sw
tri 3566 9860 3664 9958 ne
rect 3664 9900 3988 9958
tri 3988 9900 4076 9988 sw
tri 4086 9900 4174 9988 ne
rect 4174 9958 4488 9988
tri 4488 9958 4568 10038 sw
tri 4586 9958 4666 10038 ne
rect 4666 9988 4990 10038
tri 4990 9988 5088 10086 sw
tri 5088 9988 5186 10086 ne
rect 5186 10038 5500 10086
tri 5500 10038 5588 10126 sw
tri 5598 10038 5686 10126 ne
rect 5686 10090 5740 10126
rect 5860 10126 5962 10210
tri 5962 10126 6050 10214 sw
tri 6060 10126 6148 10214 ne
rect 6148 10210 6512 10214
rect 6148 10126 6290 10210
rect 5860 10090 6050 10126
rect 5686 10086 6050 10090
tri 6050 10086 6090 10126 sw
tri 6148 10086 6188 10126 ne
rect 6188 10090 6290 10126
rect 6410 10126 6512 10210
tri 6512 10126 6600 10214 sw
tri 6610 10126 6698 10214 ne
rect 6698 10210 7062 10214
rect 6698 10126 6840 10210
rect 6410 10090 6600 10126
rect 6188 10086 6600 10090
rect 5686 10038 6090 10086
rect 5186 9988 5588 10038
rect 4666 9958 5088 9988
rect 4174 9900 4568 9958
rect 3664 9860 4076 9900
tri 4076 9860 4116 9900 sw
tri 4174 9860 4214 9900 ne
rect 4214 9860 4568 9900
tri 4568 9860 4666 9958 sw
tri 4666 9860 4764 9958 ne
rect 4764 9900 5088 9958
tri 5088 9900 5176 9988 sw
tri 5186 9900 5274 9988 ne
rect 5274 9958 5588 9988
tri 5588 9958 5668 10038 sw
tri 5686 9958 5766 10038 ne
rect 5766 9988 6090 10038
tri 6090 9988 6188 10086 sw
tri 6188 9988 6286 10086 ne
rect 6286 10038 6600 10086
tri 6600 10038 6688 10126 sw
tri 6698 10038 6786 10126 ne
rect 6786 10090 6840 10126
rect 6960 10126 7062 10210
tri 7062 10126 7150 10214 sw
tri 7160 10126 7248 10214 ne
rect 7248 10210 7612 10214
rect 7248 10126 7390 10210
rect 6960 10090 7150 10126
rect 6786 10086 7150 10090
tri 7150 10086 7190 10126 sw
tri 7248 10086 7288 10126 ne
rect 7288 10090 7390 10126
rect 7510 10126 7612 10210
tri 7612 10126 7700 10214 sw
tri 7710 10126 7798 10214 ne
rect 7798 10210 8162 10214
rect 7798 10126 7940 10210
rect 7510 10090 7700 10126
rect 7288 10086 7700 10090
rect 6786 10038 7190 10086
rect 6286 9988 6688 10038
rect 5766 9958 6188 9988
rect 5274 9900 5668 9958
rect 4764 9860 5176 9900
tri 5176 9860 5216 9900 sw
tri 5274 9860 5314 9900 ne
rect 5314 9860 5668 9900
tri 5668 9860 5766 9958 sw
tri 5766 9860 5864 9958 ne
rect 5864 9900 6188 9958
tri 6188 9900 6276 9988 sw
tri 6286 9900 6374 9988 ne
rect 6374 9958 6688 9988
tri 6688 9958 6768 10038 sw
tri 6786 9958 6866 10038 ne
rect 6866 9988 7190 10038
tri 7190 9988 7288 10086 sw
tri 7288 9988 7386 10086 ne
rect 7386 10038 7700 10086
tri 7700 10038 7788 10126 sw
tri 7798 10038 7886 10126 ne
rect 7886 10090 7940 10126
rect 8060 10126 8162 10210
tri 8162 10126 8250 10214 sw
tri 8260 10126 8348 10214 ne
rect 8348 10210 8712 10214
rect 8348 10126 8490 10210
rect 8060 10090 8250 10126
rect 7886 10086 8250 10090
tri 8250 10086 8290 10126 sw
tri 8348 10086 8388 10126 ne
rect 8388 10090 8490 10126
rect 8610 10126 8712 10210
tri 8712 10126 8800 10214 sw
tri 8810 10126 8898 10214 ne
rect 8898 10210 9262 10214
rect 8898 10126 9040 10210
rect 8610 10090 8800 10126
rect 8388 10086 8800 10090
rect 7886 10038 8290 10086
rect 7386 9988 7788 10038
rect 6866 9958 7288 9988
rect 6374 9900 6768 9958
rect 5864 9860 6276 9900
tri 6276 9860 6316 9900 sw
tri 6374 9860 6414 9900 ne
rect 6414 9860 6768 9900
tri 6768 9860 6866 9958 sw
tri 6866 9860 6964 9958 ne
rect 6964 9900 7288 9958
tri 7288 9900 7376 9988 sw
tri 7386 9900 7474 9988 ne
rect 7474 9958 7788 9988
tri 7788 9958 7868 10038 sw
tri 7886 9958 7966 10038 ne
rect 7966 9988 8290 10038
tri 8290 9988 8388 10086 sw
tri 8388 9988 8486 10086 ne
rect 8486 10038 8800 10086
tri 8800 10038 8888 10126 sw
tri 8898 10038 8986 10126 ne
rect 8986 10090 9040 10126
rect 9160 10126 9262 10210
tri 9262 10126 9350 10214 sw
tri 9360 10126 9448 10214 ne
rect 9448 10210 9812 10214
rect 9448 10126 9590 10210
rect 9160 10090 9350 10126
rect 8986 10086 9350 10090
tri 9350 10086 9390 10126 sw
tri 9448 10086 9488 10126 ne
rect 9488 10090 9590 10126
rect 9710 10126 9812 10210
tri 9812 10126 9900 10214 sw
tri 9910 10126 9998 10214 ne
rect 9998 10210 10362 10214
rect 9998 10126 10140 10210
rect 9710 10090 9900 10126
rect 9488 10086 9900 10090
rect 8986 10038 9390 10086
rect 8486 9988 8888 10038
rect 7966 9958 8388 9988
rect 7474 9900 7868 9958
rect 6964 9860 7376 9900
tri 7376 9860 7416 9900 sw
tri 7474 9860 7514 9900 ne
rect 7514 9860 7868 9900
tri 7868 9860 7966 9958 sw
tri 7966 9860 8064 9958 ne
rect 8064 9900 8388 9958
tri 8388 9900 8476 9988 sw
tri 8486 9900 8574 9988 ne
rect 8574 9958 8888 9988
tri 8888 9958 8968 10038 sw
tri 8986 9958 9066 10038 ne
rect 9066 9988 9390 10038
tri 9390 9988 9488 10086 sw
tri 9488 9988 9586 10086 ne
rect 9586 10038 9900 10086
tri 9900 10038 9988 10126 sw
tri 9998 10038 10086 10126 ne
rect 10086 10090 10140 10126
rect 10260 10126 10362 10210
tri 10362 10126 10450 10214 sw
tri 10460 10126 10548 10214 ne
rect 10548 10210 10912 10214
rect 10548 10126 10690 10210
rect 10260 10090 10450 10126
rect 10086 10086 10450 10090
tri 10450 10086 10490 10126 sw
tri 10548 10086 10588 10126 ne
rect 10588 10090 10690 10126
rect 10810 10126 10912 10210
tri 10912 10126 11000 10214 sw
tri 11010 10126 11098 10214 ne
rect 11098 10210 11462 10214
rect 11098 10126 11240 10210
rect 10810 10090 11000 10126
rect 10588 10086 11000 10090
rect 10086 10038 10490 10086
rect 9586 9988 9988 10038
rect 9066 9958 9488 9988
rect 8574 9900 8968 9958
rect 8064 9860 8476 9900
tri 8476 9860 8516 9900 sw
tri 8574 9860 8614 9900 ne
rect 8614 9860 8968 9900
tri 8968 9860 9066 9958 sw
tri 9066 9860 9164 9958 ne
rect 9164 9900 9488 9958
tri 9488 9900 9576 9988 sw
tri 9586 9900 9674 9988 ne
rect 9674 9958 9988 9988
tri 9988 9958 10068 10038 sw
tri 10086 9958 10166 10038 ne
rect 10166 9988 10490 10038
tri 10490 9988 10588 10086 sw
tri 10588 9988 10686 10086 ne
rect 10686 10038 11000 10086
tri 11000 10038 11088 10126 sw
tri 11098 10038 11186 10126 ne
rect 11186 10090 11240 10126
rect 11360 10126 11462 10210
tri 11462 10126 11550 10214 sw
tri 11560 10126 11648 10214 ne
rect 11648 10210 12012 10214
rect 11648 10126 11790 10210
rect 11360 10090 11550 10126
rect 11186 10086 11550 10090
tri 11550 10086 11590 10126 sw
tri 11648 10086 11688 10126 ne
rect 11688 10090 11790 10126
rect 11910 10126 12012 10210
tri 12012 10126 12100 10214 sw
tri 12110 10126 12198 10214 ne
rect 12198 10210 12562 10214
rect 12198 10126 12340 10210
rect 11910 10090 12100 10126
rect 11688 10086 12100 10090
rect 11186 10038 11590 10086
rect 10686 9988 11088 10038
rect 10166 9958 10588 9988
rect 9674 9900 10068 9958
rect 9164 9860 9576 9900
tri 9576 9860 9616 9900 sw
tri 9674 9860 9714 9900 ne
rect 9714 9860 10068 9900
tri 10068 9860 10166 9958 sw
tri 10166 9860 10264 9958 ne
rect 10264 9900 10588 9958
tri 10588 9900 10676 9988 sw
tri 10686 9900 10774 9988 ne
rect 10774 9958 11088 9988
tri 11088 9958 11168 10038 sw
tri 11186 9958 11266 10038 ne
rect 11266 9988 11590 10038
tri 11590 9988 11688 10086 sw
tri 11688 9988 11786 10086 ne
rect 11786 10038 12100 10086
tri 12100 10038 12188 10126 sw
tri 12198 10038 12286 10126 ne
rect 12286 10090 12340 10126
rect 12460 10126 12562 10210
tri 12562 10126 12650 10214 sw
tri 12660 10126 12748 10214 ne
rect 12748 10210 13112 10214
rect 12748 10126 12890 10210
rect 12460 10090 12650 10126
rect 12286 10086 12650 10090
tri 12650 10086 12690 10126 sw
tri 12748 10086 12788 10126 ne
rect 12788 10090 12890 10126
rect 13010 10126 13112 10210
tri 13112 10126 13200 10214 sw
tri 13210 10126 13298 10214 ne
rect 13298 10210 15775 10214
rect 13298 10126 13440 10210
rect 13010 10090 13200 10126
rect 12788 10086 13200 10090
rect 12286 10038 12690 10086
rect 11786 9988 12188 10038
rect 11266 9958 11688 9988
rect 10774 9900 11168 9958
rect 10264 9860 10676 9900
tri 10676 9860 10716 9900 sw
tri 10774 9860 10814 9900 ne
rect 10814 9860 11168 9900
tri 11168 9860 11266 9958 sw
tri 11266 9860 11364 9958 ne
rect 11364 9900 11688 9958
tri 11688 9900 11776 9988 sw
tri 11786 9900 11874 9988 ne
rect 11874 9958 12188 9988
tri 12188 9958 12268 10038 sw
tri 12286 9958 12366 10038 ne
rect 12366 9988 12690 10038
tri 12690 9988 12788 10086 sw
tri 12788 9988 12886 10086 ne
rect 12886 10038 13200 10086
tri 13200 10038 13288 10126 sw
tri 13298 10038 13386 10126 ne
rect 13386 10090 13440 10126
rect 13560 10090 15775 10210
rect 13386 10038 15775 10090
rect 12886 9988 13288 10038
rect 12366 9958 12788 9988
rect 11874 9900 12268 9958
rect 11364 9860 11776 9900
tri 11776 9860 11816 9900 sw
tri 11874 9860 11914 9900 ne
rect 11914 9860 12268 9900
tri 12268 9860 12366 9958 sw
tri 12366 9860 12464 9958 ne
rect 12464 9900 12788 9958
tri 12788 9900 12876 9988 sw
tri 12886 9900 12974 9988 ne
rect 12974 9958 13288 9988
tri 13288 9958 13368 10038 sw
tri 13386 9958 13466 10038 ne
rect 13466 9958 14075 10038
rect 12974 9900 13368 9958
rect 12464 9860 12876 9900
tri 12876 9860 12916 9900 sw
tri 12974 9860 13014 9900 ne
rect 13014 9860 13368 9900
tri 13368 9860 13466 9958 sw
tri 13466 9860 13564 9958 ne
rect 13564 9938 14075 9958
rect 14175 9938 15775 10038
rect 13564 9860 15775 9938
rect -1025 9812 -284 9860
rect -1025 9712 -925 9812
rect -825 9762 -284 9812
tri -284 9762 -186 9860 sw
tri -186 9762 -88 9860 ne
rect -88 9762 266 9860
tri 266 9762 364 9860 sw
tri 364 9762 462 9860 ne
rect 462 9762 816 9860
tri 816 9762 914 9860 sw
tri 914 9762 1012 9860 ne
rect 1012 9762 1366 9860
tri 1366 9762 1464 9860 sw
tri 1464 9762 1562 9860 ne
rect 1562 9762 1916 9860
tri 1916 9762 2014 9860 sw
tri 2014 9762 2112 9860 ne
rect 2112 9762 2466 9860
tri 2466 9762 2564 9860 sw
tri 2564 9762 2662 9860 ne
rect 2662 9762 3016 9860
tri 3016 9762 3114 9860 sw
tri 3114 9762 3212 9860 ne
rect 3212 9762 3566 9860
tri 3566 9762 3664 9860 sw
tri 3664 9762 3762 9860 ne
rect 3762 9762 4116 9860
tri 4116 9762 4214 9860 sw
tri 4214 9762 4312 9860 ne
rect 4312 9762 4666 9860
tri 4666 9762 4764 9860 sw
tri 4764 9762 4862 9860 ne
rect 4862 9762 5216 9860
tri 5216 9762 5314 9860 sw
tri 5314 9762 5412 9860 ne
rect 5412 9762 5766 9860
tri 5766 9762 5864 9860 sw
tri 5864 9762 5962 9860 ne
rect 5962 9762 6316 9860
tri 6316 9762 6414 9860 sw
tri 6414 9762 6512 9860 ne
rect 6512 9762 6866 9860
tri 6866 9762 6964 9860 sw
tri 6964 9762 7062 9860 ne
rect 7062 9762 7416 9860
tri 7416 9762 7514 9860 sw
tri 7514 9762 7612 9860 ne
rect 7612 9762 7966 9860
tri 7966 9762 8064 9860 sw
tri 8064 9762 8162 9860 ne
rect 8162 9762 8516 9860
tri 8516 9762 8614 9860 sw
tri 8614 9762 8712 9860 ne
rect 8712 9762 9066 9860
tri 9066 9762 9164 9860 sw
tri 9164 9762 9262 9860 ne
rect 9262 9762 9616 9860
tri 9616 9762 9714 9860 sw
tri 9714 9762 9812 9860 ne
rect 9812 9762 10166 9860
tri 10166 9762 10264 9860 sw
tri 10264 9762 10362 9860 ne
rect 10362 9762 10716 9860
tri 10716 9762 10814 9860 sw
tri 10814 9762 10912 9860 ne
rect 10912 9762 11266 9860
tri 11266 9762 11364 9860 sw
tri 11364 9762 11462 9860 ne
rect 11462 9762 11816 9860
tri 11816 9762 11914 9860 sw
tri 11914 9762 12012 9860 ne
rect 12012 9762 12366 9860
tri 12366 9762 12464 9860 sw
tri 12464 9762 12562 9860 ne
rect 12562 9762 12916 9860
tri 12916 9762 13014 9860 sw
tri 13014 9762 13112 9860 ne
rect 13112 9762 13466 9860
tri 13466 9762 13564 9860 sw
tri 13564 9762 13662 9860 ne
rect 13662 9762 15775 9860
rect -825 9712 -186 9762
rect -1025 9664 -186 9712
tri -186 9664 -88 9762 sw
tri -88 9664 10 9762 ne
rect 10 9664 364 9762
tri 364 9664 462 9762 sw
tri 462 9664 560 9762 ne
rect 560 9664 914 9762
tri 914 9664 1012 9762 sw
tri 1012 9664 1110 9762 ne
rect 1110 9664 1464 9762
tri 1464 9664 1562 9762 sw
tri 1562 9664 1660 9762 ne
rect 1660 9664 2014 9762
tri 2014 9664 2112 9762 sw
tri 2112 9664 2210 9762 ne
rect 2210 9664 2564 9762
tri 2564 9664 2662 9762 sw
tri 2662 9664 2760 9762 ne
rect 2760 9664 3114 9762
tri 3114 9664 3212 9762 sw
tri 3212 9664 3310 9762 ne
rect 3310 9664 3664 9762
tri 3664 9664 3762 9762 sw
tri 3762 9664 3860 9762 ne
rect 3860 9664 4214 9762
tri 4214 9664 4312 9762 sw
tri 4312 9664 4410 9762 ne
rect 4410 9664 4764 9762
tri 4764 9664 4862 9762 sw
tri 4862 9664 4960 9762 ne
rect 4960 9664 5314 9762
tri 5314 9664 5412 9762 sw
tri 5412 9664 5510 9762 ne
rect 5510 9664 5864 9762
tri 5864 9664 5962 9762 sw
tri 5962 9664 6060 9762 ne
rect 6060 9664 6414 9762
tri 6414 9664 6512 9762 sw
tri 6512 9664 6610 9762 ne
rect 6610 9664 6964 9762
tri 6964 9664 7062 9762 sw
tri 7062 9664 7160 9762 ne
rect 7160 9664 7514 9762
tri 7514 9664 7612 9762 sw
tri 7612 9664 7710 9762 ne
rect 7710 9664 8064 9762
tri 8064 9664 8162 9762 sw
tri 8162 9664 8260 9762 ne
rect 8260 9664 8614 9762
tri 8614 9664 8712 9762 sw
tri 8712 9664 8810 9762 ne
rect 8810 9664 9164 9762
tri 9164 9664 9262 9762 sw
tri 9262 9664 9360 9762 ne
rect 9360 9664 9714 9762
tri 9714 9664 9812 9762 sw
tri 9812 9664 9910 9762 ne
rect 9910 9664 10264 9762
tri 10264 9664 10362 9762 sw
tri 10362 9664 10460 9762 ne
rect 10460 9664 10814 9762
tri 10814 9664 10912 9762 sw
tri 10912 9664 11010 9762 ne
rect 11010 9664 11364 9762
tri 11364 9664 11462 9762 sw
tri 11462 9664 11560 9762 ne
rect 11560 9664 11914 9762
tri 11914 9664 12012 9762 sw
tri 12012 9664 12110 9762 ne
rect 12110 9664 12464 9762
tri 12464 9664 12562 9762 sw
tri 12562 9664 12660 9762 ne
rect 12660 9664 13014 9762
tri 13014 9664 13112 9762 sw
tri 13112 9664 13210 9762 ne
rect 13210 9664 13564 9762
tri 13564 9664 13662 9762 sw
rect -1025 9660 -88 9664
rect -1025 9540 -310 9660
rect -190 9576 -88 9660
tri -88 9576 0 9664 sw
tri 10 9576 98 9664 ne
rect 98 9660 462 9664
rect 98 9576 240 9660
rect -190 9540 0 9576
rect -1025 9536 0 9540
tri 0 9536 40 9576 sw
tri 98 9536 138 9576 ne
rect 138 9540 240 9576
rect 360 9576 462 9660
tri 462 9576 550 9664 sw
tri 560 9576 648 9664 ne
rect 648 9660 1012 9664
rect 648 9576 790 9660
rect 360 9540 550 9576
rect 138 9536 550 9540
tri -412 9438 -314 9536 ne
rect -314 9438 40 9536
tri 40 9438 138 9536 sw
tri 138 9438 236 9536 ne
rect 236 9488 550 9536
tri 550 9488 638 9576 sw
tri 648 9488 736 9576 ne
rect 736 9540 790 9576
rect 910 9576 1012 9660
tri 1012 9576 1100 9664 sw
tri 1110 9576 1198 9664 ne
rect 1198 9660 1562 9664
rect 1198 9576 1340 9660
rect 910 9540 1100 9576
rect 736 9536 1100 9540
tri 1100 9536 1140 9576 sw
tri 1198 9536 1238 9576 ne
rect 1238 9540 1340 9576
rect 1460 9576 1562 9660
tri 1562 9576 1650 9664 sw
tri 1660 9576 1748 9664 ne
rect 1748 9660 2112 9664
rect 1748 9576 1890 9660
rect 1460 9540 1650 9576
rect 1238 9536 1650 9540
rect 736 9488 1140 9536
rect 236 9438 638 9488
rect -2525 9350 -412 9438
tri -412 9350 -324 9438 sw
tri -314 9350 -226 9438 ne
rect -226 9350 138 9438
tri 138 9350 226 9438 sw
tri 236 9350 324 9438 ne
rect 324 9408 638 9438
tri 638 9408 718 9488 sw
tri 736 9408 816 9488 ne
rect 816 9438 1140 9488
tri 1140 9438 1238 9536 sw
tri 1238 9438 1336 9536 ne
rect 1336 9488 1650 9536
tri 1650 9488 1738 9576 sw
tri 1748 9488 1836 9576 ne
rect 1836 9540 1890 9576
rect 2010 9576 2112 9660
tri 2112 9576 2200 9664 sw
tri 2210 9576 2298 9664 ne
rect 2298 9660 2662 9664
rect 2298 9576 2440 9660
rect 2010 9540 2200 9576
rect 1836 9536 2200 9540
tri 2200 9536 2240 9576 sw
tri 2298 9536 2338 9576 ne
rect 2338 9540 2440 9576
rect 2560 9576 2662 9660
tri 2662 9576 2750 9664 sw
tri 2760 9576 2848 9664 ne
rect 2848 9660 3212 9664
rect 2848 9576 2990 9660
rect 2560 9540 2750 9576
rect 2338 9536 2750 9540
rect 1836 9488 2240 9536
rect 1336 9438 1738 9488
rect 816 9408 1238 9438
rect 324 9350 718 9408
rect -2525 9310 -324 9350
tri -324 9310 -284 9350 sw
tri -226 9310 -186 9350 ne
rect -186 9310 226 9350
tri 226 9310 266 9350 sw
tri 324 9310 364 9350 ne
rect 364 9310 718 9350
tri 718 9310 816 9408 sw
tri 816 9310 914 9408 ne
rect 914 9350 1238 9408
tri 1238 9350 1326 9438 sw
tri 1336 9350 1424 9438 ne
rect 1424 9408 1738 9438
tri 1738 9408 1818 9488 sw
tri 1836 9408 1916 9488 ne
rect 1916 9438 2240 9488
tri 2240 9438 2338 9536 sw
tri 2338 9438 2436 9536 ne
rect 2436 9488 2750 9536
tri 2750 9488 2838 9576 sw
tri 2848 9488 2936 9576 ne
rect 2936 9540 2990 9576
rect 3110 9576 3212 9660
tri 3212 9576 3300 9664 sw
tri 3310 9576 3398 9664 ne
rect 3398 9660 3762 9664
rect 3398 9576 3540 9660
rect 3110 9540 3300 9576
rect 2936 9536 3300 9540
tri 3300 9536 3340 9576 sw
tri 3398 9536 3438 9576 ne
rect 3438 9540 3540 9576
rect 3660 9576 3762 9660
tri 3762 9576 3850 9664 sw
tri 3860 9576 3948 9664 ne
rect 3948 9660 4312 9664
rect 3948 9576 4090 9660
rect 3660 9540 3850 9576
rect 3438 9536 3850 9540
rect 2936 9488 3340 9536
rect 2436 9438 2838 9488
rect 1916 9408 2338 9438
rect 1424 9350 1818 9408
rect 914 9310 1326 9350
tri 1326 9310 1366 9350 sw
tri 1424 9310 1464 9350 ne
rect 1464 9310 1818 9350
tri 1818 9310 1916 9408 sw
tri 1916 9310 2014 9408 ne
rect 2014 9350 2338 9408
tri 2338 9350 2426 9438 sw
tri 2436 9350 2524 9438 ne
rect 2524 9408 2838 9438
tri 2838 9408 2918 9488 sw
tri 2936 9408 3016 9488 ne
rect 3016 9438 3340 9488
tri 3340 9438 3438 9536 sw
tri 3438 9438 3536 9536 ne
rect 3536 9488 3850 9536
tri 3850 9488 3938 9576 sw
tri 3948 9488 4036 9576 ne
rect 4036 9540 4090 9576
rect 4210 9576 4312 9660
tri 4312 9576 4400 9664 sw
tri 4410 9576 4498 9664 ne
rect 4498 9660 4862 9664
rect 4498 9576 4640 9660
rect 4210 9540 4400 9576
rect 4036 9536 4400 9540
tri 4400 9536 4440 9576 sw
tri 4498 9536 4538 9576 ne
rect 4538 9540 4640 9576
rect 4760 9576 4862 9660
tri 4862 9576 4950 9664 sw
tri 4960 9576 5048 9664 ne
rect 5048 9660 5412 9664
rect 5048 9576 5190 9660
rect 4760 9540 4950 9576
rect 4538 9536 4950 9540
rect 4036 9488 4440 9536
rect 3536 9438 3938 9488
rect 3016 9408 3438 9438
rect 2524 9350 2918 9408
rect 2014 9310 2426 9350
tri 2426 9310 2466 9350 sw
tri 2524 9310 2564 9350 ne
rect 2564 9310 2918 9350
tri 2918 9310 3016 9408 sw
tri 3016 9310 3114 9408 ne
rect 3114 9350 3438 9408
tri 3438 9350 3526 9438 sw
tri 3536 9350 3624 9438 ne
rect 3624 9408 3938 9438
tri 3938 9408 4018 9488 sw
tri 4036 9408 4116 9488 ne
rect 4116 9438 4440 9488
tri 4440 9438 4538 9536 sw
tri 4538 9438 4636 9536 ne
rect 4636 9488 4950 9536
tri 4950 9488 5038 9576 sw
tri 5048 9488 5136 9576 ne
rect 5136 9540 5190 9576
rect 5310 9576 5412 9660
tri 5412 9576 5500 9664 sw
tri 5510 9576 5598 9664 ne
rect 5598 9660 5962 9664
rect 5598 9576 5740 9660
rect 5310 9540 5500 9576
rect 5136 9536 5500 9540
tri 5500 9536 5540 9576 sw
tri 5598 9536 5638 9576 ne
rect 5638 9540 5740 9576
rect 5860 9576 5962 9660
tri 5962 9576 6050 9664 sw
tri 6060 9576 6148 9664 ne
rect 6148 9660 6512 9664
rect 6148 9576 6290 9660
rect 5860 9540 6050 9576
rect 5638 9536 6050 9540
rect 5136 9488 5540 9536
rect 4636 9438 5038 9488
rect 4116 9408 4538 9438
rect 3624 9350 4018 9408
rect 3114 9310 3526 9350
tri 3526 9310 3566 9350 sw
tri 3624 9310 3664 9350 ne
rect 3664 9310 4018 9350
tri 4018 9310 4116 9408 sw
tri 4116 9310 4214 9408 ne
rect 4214 9350 4538 9408
tri 4538 9350 4626 9438 sw
tri 4636 9350 4724 9438 ne
rect 4724 9408 5038 9438
tri 5038 9408 5118 9488 sw
tri 5136 9408 5216 9488 ne
rect 5216 9438 5540 9488
tri 5540 9438 5638 9536 sw
tri 5638 9438 5736 9536 ne
rect 5736 9488 6050 9536
tri 6050 9488 6138 9576 sw
tri 6148 9488 6236 9576 ne
rect 6236 9540 6290 9576
rect 6410 9576 6512 9660
tri 6512 9576 6600 9664 sw
tri 6610 9576 6698 9664 ne
rect 6698 9660 7062 9664
rect 6698 9576 6840 9660
rect 6410 9540 6600 9576
rect 6236 9536 6600 9540
tri 6600 9536 6640 9576 sw
tri 6698 9536 6738 9576 ne
rect 6738 9540 6840 9576
rect 6960 9576 7062 9660
tri 7062 9576 7150 9664 sw
tri 7160 9576 7248 9664 ne
rect 7248 9660 7612 9664
rect 7248 9576 7390 9660
rect 6960 9540 7150 9576
rect 6738 9536 7150 9540
rect 6236 9488 6640 9536
rect 5736 9438 6138 9488
rect 5216 9408 5638 9438
rect 4724 9350 5118 9408
rect 4214 9310 4626 9350
tri 4626 9310 4666 9350 sw
tri 4724 9310 4764 9350 ne
rect 4764 9310 5118 9350
tri 5118 9310 5216 9408 sw
tri 5216 9310 5314 9408 ne
rect 5314 9350 5638 9408
tri 5638 9350 5726 9438 sw
tri 5736 9350 5824 9438 ne
rect 5824 9408 6138 9438
tri 6138 9408 6218 9488 sw
tri 6236 9408 6316 9488 ne
rect 6316 9438 6640 9488
tri 6640 9438 6738 9536 sw
tri 6738 9438 6836 9536 ne
rect 6836 9488 7150 9536
tri 7150 9488 7238 9576 sw
tri 7248 9488 7336 9576 ne
rect 7336 9540 7390 9576
rect 7510 9576 7612 9660
tri 7612 9576 7700 9664 sw
tri 7710 9576 7798 9664 ne
rect 7798 9660 8162 9664
rect 7798 9576 7940 9660
rect 7510 9540 7700 9576
rect 7336 9536 7700 9540
tri 7700 9536 7740 9576 sw
tri 7798 9536 7838 9576 ne
rect 7838 9540 7940 9576
rect 8060 9576 8162 9660
tri 8162 9576 8250 9664 sw
tri 8260 9576 8348 9664 ne
rect 8348 9660 8712 9664
rect 8348 9576 8490 9660
rect 8060 9540 8250 9576
rect 7838 9536 8250 9540
rect 7336 9488 7740 9536
rect 6836 9438 7238 9488
rect 6316 9408 6738 9438
rect 5824 9350 6218 9408
rect 5314 9310 5726 9350
tri 5726 9310 5766 9350 sw
tri 5824 9310 5864 9350 ne
rect 5864 9310 6218 9350
tri 6218 9310 6316 9408 sw
tri 6316 9310 6414 9408 ne
rect 6414 9350 6738 9408
tri 6738 9350 6826 9438 sw
tri 6836 9350 6924 9438 ne
rect 6924 9408 7238 9438
tri 7238 9408 7318 9488 sw
tri 7336 9408 7416 9488 ne
rect 7416 9438 7740 9488
tri 7740 9438 7838 9536 sw
tri 7838 9438 7936 9536 ne
rect 7936 9488 8250 9536
tri 8250 9488 8338 9576 sw
tri 8348 9488 8436 9576 ne
rect 8436 9540 8490 9576
rect 8610 9576 8712 9660
tri 8712 9576 8800 9664 sw
tri 8810 9576 8898 9664 ne
rect 8898 9660 9262 9664
rect 8898 9576 9040 9660
rect 8610 9540 8800 9576
rect 8436 9536 8800 9540
tri 8800 9536 8840 9576 sw
tri 8898 9536 8938 9576 ne
rect 8938 9540 9040 9576
rect 9160 9576 9262 9660
tri 9262 9576 9350 9664 sw
tri 9360 9576 9448 9664 ne
rect 9448 9660 9812 9664
rect 9448 9576 9590 9660
rect 9160 9540 9350 9576
rect 8938 9536 9350 9540
rect 8436 9488 8840 9536
rect 7936 9438 8338 9488
rect 7416 9408 7838 9438
rect 6924 9350 7318 9408
rect 6414 9310 6826 9350
tri 6826 9310 6866 9350 sw
tri 6924 9310 6964 9350 ne
rect 6964 9310 7318 9350
tri 7318 9310 7416 9408 sw
tri 7416 9310 7514 9408 ne
rect 7514 9350 7838 9408
tri 7838 9350 7926 9438 sw
tri 7936 9350 8024 9438 ne
rect 8024 9408 8338 9438
tri 8338 9408 8418 9488 sw
tri 8436 9408 8516 9488 ne
rect 8516 9438 8840 9488
tri 8840 9438 8938 9536 sw
tri 8938 9438 9036 9536 ne
rect 9036 9488 9350 9536
tri 9350 9488 9438 9576 sw
tri 9448 9488 9536 9576 ne
rect 9536 9540 9590 9576
rect 9710 9576 9812 9660
tri 9812 9576 9900 9664 sw
tri 9910 9576 9998 9664 ne
rect 9998 9660 10362 9664
rect 9998 9576 10140 9660
rect 9710 9540 9900 9576
rect 9536 9536 9900 9540
tri 9900 9536 9940 9576 sw
tri 9998 9536 10038 9576 ne
rect 10038 9540 10140 9576
rect 10260 9576 10362 9660
tri 10362 9576 10450 9664 sw
tri 10460 9576 10548 9664 ne
rect 10548 9660 10912 9664
rect 10548 9576 10690 9660
rect 10260 9540 10450 9576
rect 10038 9536 10450 9540
rect 9536 9488 9940 9536
rect 9036 9438 9438 9488
rect 8516 9408 8938 9438
rect 8024 9350 8418 9408
rect 7514 9310 7926 9350
tri 7926 9310 7966 9350 sw
tri 8024 9310 8064 9350 ne
rect 8064 9310 8418 9350
tri 8418 9310 8516 9408 sw
tri 8516 9310 8614 9408 ne
rect 8614 9350 8938 9408
tri 8938 9350 9026 9438 sw
tri 9036 9350 9124 9438 ne
rect 9124 9408 9438 9438
tri 9438 9408 9518 9488 sw
tri 9536 9408 9616 9488 ne
rect 9616 9438 9940 9488
tri 9940 9438 10038 9536 sw
tri 10038 9438 10136 9536 ne
rect 10136 9488 10450 9536
tri 10450 9488 10538 9576 sw
tri 10548 9488 10636 9576 ne
rect 10636 9540 10690 9576
rect 10810 9576 10912 9660
tri 10912 9576 11000 9664 sw
tri 11010 9576 11098 9664 ne
rect 11098 9660 11462 9664
rect 11098 9576 11240 9660
rect 10810 9540 11000 9576
rect 10636 9536 11000 9540
tri 11000 9536 11040 9576 sw
tri 11098 9536 11138 9576 ne
rect 11138 9540 11240 9576
rect 11360 9576 11462 9660
tri 11462 9576 11550 9664 sw
tri 11560 9576 11648 9664 ne
rect 11648 9660 12012 9664
rect 11648 9576 11790 9660
rect 11360 9540 11550 9576
rect 11138 9536 11550 9540
rect 10636 9488 11040 9536
rect 10136 9438 10538 9488
rect 9616 9408 10038 9438
rect 9124 9350 9518 9408
rect 8614 9310 9026 9350
tri 9026 9310 9066 9350 sw
tri 9124 9310 9164 9350 ne
rect 9164 9310 9518 9350
tri 9518 9310 9616 9408 sw
tri 9616 9310 9714 9408 ne
rect 9714 9350 10038 9408
tri 10038 9350 10126 9438 sw
tri 10136 9350 10224 9438 ne
rect 10224 9408 10538 9438
tri 10538 9408 10618 9488 sw
tri 10636 9408 10716 9488 ne
rect 10716 9438 11040 9488
tri 11040 9438 11138 9536 sw
tri 11138 9438 11236 9536 ne
rect 11236 9488 11550 9536
tri 11550 9488 11638 9576 sw
tri 11648 9488 11736 9576 ne
rect 11736 9540 11790 9576
rect 11910 9576 12012 9660
tri 12012 9576 12100 9664 sw
tri 12110 9576 12198 9664 ne
rect 12198 9660 12562 9664
rect 12198 9576 12340 9660
rect 11910 9540 12100 9576
rect 11736 9536 12100 9540
tri 12100 9536 12140 9576 sw
tri 12198 9536 12238 9576 ne
rect 12238 9540 12340 9576
rect 12460 9576 12562 9660
tri 12562 9576 12650 9664 sw
tri 12660 9576 12748 9664 ne
rect 12748 9660 13112 9664
rect 12748 9576 12890 9660
rect 12460 9540 12650 9576
rect 12238 9536 12650 9540
rect 11736 9488 12140 9536
rect 11236 9438 11638 9488
rect 10716 9408 11138 9438
rect 10224 9350 10618 9408
rect 9714 9310 10126 9350
tri 10126 9310 10166 9350 sw
tri 10224 9310 10264 9350 ne
rect 10264 9310 10618 9350
tri 10618 9310 10716 9408 sw
tri 10716 9310 10814 9408 ne
rect 10814 9350 11138 9408
tri 11138 9350 11226 9438 sw
tri 11236 9350 11324 9438 ne
rect 11324 9408 11638 9438
tri 11638 9408 11718 9488 sw
tri 11736 9408 11816 9488 ne
rect 11816 9438 12140 9488
tri 12140 9438 12238 9536 sw
tri 12238 9438 12336 9536 ne
rect 12336 9488 12650 9536
tri 12650 9488 12738 9576 sw
tri 12748 9488 12836 9576 ne
rect 12836 9540 12890 9576
rect 13010 9576 13112 9660
tri 13112 9576 13200 9664 sw
tri 13210 9576 13298 9664 ne
rect 13298 9660 14275 9664
rect 13298 9576 13440 9660
rect 13010 9540 13200 9576
rect 12836 9536 13200 9540
tri 13200 9536 13240 9576 sw
tri 13298 9536 13338 9576 ne
rect 13338 9540 13440 9576
rect 13560 9540 14275 9660
rect 13338 9536 14275 9540
rect 12836 9488 13240 9536
rect 12336 9438 12738 9488
rect 11816 9408 12238 9438
rect 11324 9350 11718 9408
rect 10814 9310 11226 9350
tri 11226 9310 11266 9350 sw
tri 11324 9310 11364 9350 ne
rect 11364 9310 11718 9350
tri 11718 9310 11816 9408 sw
tri 11816 9310 11914 9408 ne
rect 11914 9350 12238 9408
tri 12238 9350 12326 9438 sw
tri 12336 9350 12424 9438 ne
rect 12424 9408 12738 9438
tri 12738 9408 12818 9488 sw
tri 12836 9408 12916 9488 ne
rect 12916 9438 13240 9488
tri 13240 9438 13338 9536 sw
tri 13338 9438 13436 9536 ne
rect 13436 9438 14275 9536
rect 12916 9408 13338 9438
rect 12424 9350 12818 9408
rect 11914 9310 12326 9350
tri 12326 9310 12366 9350 sw
tri 12424 9310 12464 9350 ne
rect 12464 9310 12818 9350
tri 12818 9310 12916 9408 sw
tri 12916 9310 13014 9408 ne
rect 13014 9350 13338 9408
tri 13338 9350 13426 9438 sw
tri 13436 9350 13524 9438 ne
rect 13524 9350 14275 9438
rect 13014 9310 13426 9350
tri 13426 9310 13466 9350 sw
tri 13524 9310 13564 9350 ne
rect 13564 9310 14275 9350
rect -2525 9212 -284 9310
tri -284 9212 -186 9310 sw
tri -186 9212 -88 9310 ne
rect -88 9212 266 9310
tri 266 9212 364 9310 sw
tri 364 9212 462 9310 ne
rect 462 9212 816 9310
tri 816 9212 914 9310 sw
tri 914 9212 1012 9310 ne
rect 1012 9212 1366 9310
tri 1366 9212 1464 9310 sw
tri 1464 9212 1562 9310 ne
rect 1562 9212 1916 9310
tri 1916 9212 2014 9310 sw
tri 2014 9212 2112 9310 ne
rect 2112 9212 2466 9310
tri 2466 9212 2564 9310 sw
tri 2564 9212 2662 9310 ne
rect 2662 9212 3016 9310
tri 3016 9212 3114 9310 sw
tri 3114 9212 3212 9310 ne
rect 3212 9212 3566 9310
tri 3566 9212 3664 9310 sw
tri 3664 9212 3762 9310 ne
rect 3762 9212 4116 9310
tri 4116 9212 4214 9310 sw
tri 4214 9212 4312 9310 ne
rect 4312 9212 4666 9310
tri 4666 9212 4764 9310 sw
tri 4764 9212 4862 9310 ne
rect 4862 9212 5216 9310
tri 5216 9212 5314 9310 sw
tri 5314 9212 5412 9310 ne
rect 5412 9212 5766 9310
tri 5766 9212 5864 9310 sw
tri 5864 9212 5962 9310 ne
rect 5962 9212 6316 9310
tri 6316 9212 6414 9310 sw
tri 6414 9212 6512 9310 ne
rect 6512 9212 6866 9310
tri 6866 9212 6964 9310 sw
tri 6964 9212 7062 9310 ne
rect 7062 9212 7416 9310
tri 7416 9212 7514 9310 sw
tri 7514 9212 7612 9310 ne
rect 7612 9212 7966 9310
tri 7966 9212 8064 9310 sw
tri 8064 9212 8162 9310 ne
rect 8162 9212 8516 9310
tri 8516 9212 8614 9310 sw
tri 8614 9212 8712 9310 ne
rect 8712 9212 9066 9310
tri 9066 9212 9164 9310 sw
tri 9164 9212 9262 9310 ne
rect 9262 9212 9616 9310
tri 9616 9212 9714 9310 sw
tri 9714 9212 9812 9310 ne
rect 9812 9212 10166 9310
tri 10166 9212 10264 9310 sw
tri 10264 9212 10362 9310 ne
rect 10362 9212 10716 9310
tri 10716 9212 10814 9310 sw
tri 10814 9212 10912 9310 ne
rect 10912 9212 11266 9310
tri 11266 9212 11364 9310 sw
tri 11364 9212 11462 9310 ne
rect 11462 9212 11816 9310
tri 11816 9212 11914 9310 sw
tri 11914 9212 12012 9310 ne
rect 12012 9212 12366 9310
tri 12366 9212 12464 9310 sw
tri 12464 9212 12562 9310 ne
rect 12562 9212 12916 9310
tri 12916 9212 13014 9310 sw
tri 13014 9212 13112 9310 ne
rect 13112 9212 13466 9310
tri 13466 9212 13564 9310 sw
tri 13564 9212 13662 9310 ne
rect 13662 9212 14275 9310
rect -2525 9114 -186 9212
tri -186 9114 -88 9212 sw
tri -88 9114 10 9212 ne
rect 10 9114 364 9212
tri 364 9114 462 9212 sw
tri 462 9114 560 9212 ne
rect 560 9114 914 9212
tri 914 9114 1012 9212 sw
tri 1012 9114 1110 9212 ne
rect 1110 9114 1464 9212
tri 1464 9114 1562 9212 sw
tri 1562 9114 1660 9212 ne
rect 1660 9114 2014 9212
tri 2014 9114 2112 9212 sw
tri 2112 9114 2210 9212 ne
rect 2210 9114 2564 9212
tri 2564 9114 2662 9212 sw
tri 2662 9114 2760 9212 ne
rect 2760 9114 3114 9212
tri 3114 9114 3212 9212 sw
tri 3212 9114 3310 9212 ne
rect 3310 9114 3664 9212
tri 3664 9114 3762 9212 sw
tri 3762 9114 3860 9212 ne
rect 3860 9114 4214 9212
tri 4214 9114 4312 9212 sw
tri 4312 9114 4410 9212 ne
rect 4410 9114 4764 9212
tri 4764 9114 4862 9212 sw
tri 4862 9114 4960 9212 ne
rect 4960 9114 5314 9212
tri 5314 9114 5412 9212 sw
tri 5412 9114 5510 9212 ne
rect 5510 9114 5864 9212
tri 5864 9114 5962 9212 sw
tri 5962 9114 6060 9212 ne
rect 6060 9114 6414 9212
tri 6414 9114 6512 9212 sw
tri 6512 9114 6610 9212 ne
rect 6610 9114 6964 9212
tri 6964 9114 7062 9212 sw
tri 7062 9114 7160 9212 ne
rect 7160 9114 7514 9212
tri 7514 9114 7612 9212 sw
tri 7612 9114 7710 9212 ne
rect 7710 9114 8064 9212
tri 8064 9114 8162 9212 sw
tri 8162 9114 8260 9212 ne
rect 8260 9114 8614 9212
tri 8614 9114 8712 9212 sw
tri 8712 9114 8810 9212 ne
rect 8810 9114 9164 9212
tri 9164 9114 9262 9212 sw
tri 9262 9114 9360 9212 ne
rect 9360 9114 9714 9212
tri 9714 9114 9812 9212 sw
tri 9812 9114 9910 9212 ne
rect 9910 9114 10264 9212
tri 10264 9114 10362 9212 sw
tri 10362 9114 10460 9212 ne
rect 10460 9114 10814 9212
tri 10814 9114 10912 9212 sw
tri 10912 9114 11010 9212 ne
rect 11010 9114 11364 9212
tri 11364 9114 11462 9212 sw
tri 11462 9114 11560 9212 ne
rect 11560 9114 11914 9212
tri 11914 9114 12012 9212 sw
tri 12012 9114 12110 9212 ne
rect 12110 9114 12464 9212
tri 12464 9114 12562 9212 sw
tri 12562 9114 12660 9212 ne
rect 12660 9114 13014 9212
tri 13014 9114 13112 9212 sw
tri 13112 9114 13210 9212 ne
rect 13210 9114 13564 9212
tri 13564 9114 13662 9212 sw
rect 14775 9114 15775 9762
rect -2525 9110 -88 9114
rect -2525 8990 -310 9110
rect -190 9026 -88 9110
tri -88 9026 0 9114 sw
tri 10 9026 98 9114 ne
rect 98 9110 462 9114
rect 98 9026 240 9110
rect -190 8990 0 9026
rect -2525 8986 0 8990
rect -2525 8338 -1525 8986
tri -412 8888 -314 8986 ne
rect -314 8938 0 8986
tri 0 8938 88 9026 sw
tri 98 8938 186 9026 ne
rect 186 8990 240 9026
rect 360 9026 462 9110
tri 462 9026 550 9114 sw
tri 560 9026 648 9114 ne
rect 648 9110 1012 9114
rect 648 9026 790 9110
rect 360 8990 550 9026
rect 186 8986 550 8990
tri 550 8986 590 9026 sw
tri 648 8986 688 9026 ne
rect 688 8990 790 9026
rect 910 9026 1012 9110
tri 1012 9026 1100 9114 sw
tri 1110 9026 1198 9114 ne
rect 1198 9110 1562 9114
rect 1198 9026 1340 9110
rect 910 8990 1100 9026
rect 688 8986 1100 8990
rect 186 8938 590 8986
rect -314 8888 88 8938
rect -1025 8800 -412 8888
tri -412 8800 -324 8888 sw
tri -314 8800 -226 8888 ne
rect -226 8858 88 8888
tri 88 8858 168 8938 sw
tri 186 8858 266 8938 ne
rect 266 8888 590 8938
tri 590 8888 688 8986 sw
tri 688 8888 786 8986 ne
rect 786 8938 1100 8986
tri 1100 8938 1188 9026 sw
tri 1198 8938 1286 9026 ne
rect 1286 8990 1340 9026
rect 1460 9026 1562 9110
tri 1562 9026 1650 9114 sw
tri 1660 9026 1748 9114 ne
rect 1748 9110 2112 9114
rect 1748 9026 1890 9110
rect 1460 8990 1650 9026
rect 1286 8986 1650 8990
tri 1650 8986 1690 9026 sw
tri 1748 8986 1788 9026 ne
rect 1788 8990 1890 9026
rect 2010 9026 2112 9110
tri 2112 9026 2200 9114 sw
tri 2210 9026 2298 9114 ne
rect 2298 9110 2662 9114
rect 2298 9026 2440 9110
rect 2010 8990 2200 9026
rect 1788 8986 2200 8990
rect 1286 8938 1690 8986
rect 786 8888 1188 8938
rect 266 8858 688 8888
rect -226 8800 168 8858
rect -1025 8760 -324 8800
tri -324 8760 -284 8800 sw
tri -226 8760 -186 8800 ne
rect -186 8760 168 8800
tri 168 8760 266 8858 sw
tri 266 8760 364 8858 ne
rect 364 8800 688 8858
tri 688 8800 776 8888 sw
tri 786 8800 874 8888 ne
rect 874 8858 1188 8888
tri 1188 8858 1268 8938 sw
tri 1286 8858 1366 8938 ne
rect 1366 8888 1690 8938
tri 1690 8888 1788 8986 sw
tri 1788 8888 1886 8986 ne
rect 1886 8938 2200 8986
tri 2200 8938 2288 9026 sw
tri 2298 8938 2386 9026 ne
rect 2386 8990 2440 9026
rect 2560 9026 2662 9110
tri 2662 9026 2750 9114 sw
tri 2760 9026 2848 9114 ne
rect 2848 9110 3212 9114
rect 2848 9026 2990 9110
rect 2560 8990 2750 9026
rect 2386 8986 2750 8990
tri 2750 8986 2790 9026 sw
tri 2848 8986 2888 9026 ne
rect 2888 8990 2990 9026
rect 3110 9026 3212 9110
tri 3212 9026 3300 9114 sw
tri 3310 9026 3398 9114 ne
rect 3398 9110 3762 9114
rect 3398 9026 3540 9110
rect 3110 8990 3300 9026
rect 2888 8986 3300 8990
rect 2386 8938 2790 8986
rect 1886 8888 2288 8938
rect 1366 8858 1788 8888
rect 874 8800 1268 8858
rect 364 8760 776 8800
tri 776 8760 816 8800 sw
tri 874 8760 914 8800 ne
rect 914 8760 1268 8800
tri 1268 8760 1366 8858 sw
tri 1366 8760 1464 8858 ne
rect 1464 8800 1788 8858
tri 1788 8800 1876 8888 sw
tri 1886 8800 1974 8888 ne
rect 1974 8858 2288 8888
tri 2288 8858 2368 8938 sw
tri 2386 8858 2466 8938 ne
rect 2466 8888 2790 8938
tri 2790 8888 2888 8986 sw
tri 2888 8888 2986 8986 ne
rect 2986 8938 3300 8986
tri 3300 8938 3388 9026 sw
tri 3398 8938 3486 9026 ne
rect 3486 8990 3540 9026
rect 3660 9026 3762 9110
tri 3762 9026 3850 9114 sw
tri 3860 9026 3948 9114 ne
rect 3948 9110 4312 9114
rect 3948 9026 4090 9110
rect 3660 8990 3850 9026
rect 3486 8986 3850 8990
tri 3850 8986 3890 9026 sw
tri 3948 8986 3988 9026 ne
rect 3988 8990 4090 9026
rect 4210 9026 4312 9110
tri 4312 9026 4400 9114 sw
tri 4410 9026 4498 9114 ne
rect 4498 9110 4862 9114
rect 4498 9026 4640 9110
rect 4210 8990 4400 9026
rect 3988 8986 4400 8990
rect 3486 8938 3890 8986
rect 2986 8888 3388 8938
rect 2466 8858 2888 8888
rect 1974 8800 2368 8858
rect 1464 8760 1876 8800
tri 1876 8760 1916 8800 sw
tri 1974 8760 2014 8800 ne
rect 2014 8760 2368 8800
tri 2368 8760 2466 8858 sw
tri 2466 8760 2564 8858 ne
rect 2564 8800 2888 8858
tri 2888 8800 2976 8888 sw
tri 2986 8800 3074 8888 ne
rect 3074 8858 3388 8888
tri 3388 8858 3468 8938 sw
tri 3486 8858 3566 8938 ne
rect 3566 8888 3890 8938
tri 3890 8888 3988 8986 sw
tri 3988 8888 4086 8986 ne
rect 4086 8938 4400 8986
tri 4400 8938 4488 9026 sw
tri 4498 8938 4586 9026 ne
rect 4586 8990 4640 9026
rect 4760 9026 4862 9110
tri 4862 9026 4950 9114 sw
tri 4960 9026 5048 9114 ne
rect 5048 9110 5412 9114
rect 5048 9026 5190 9110
rect 4760 8990 4950 9026
rect 4586 8986 4950 8990
tri 4950 8986 4990 9026 sw
tri 5048 8986 5088 9026 ne
rect 5088 8990 5190 9026
rect 5310 9026 5412 9110
tri 5412 9026 5500 9114 sw
tri 5510 9026 5598 9114 ne
rect 5598 9110 5962 9114
rect 5598 9026 5740 9110
rect 5310 8990 5500 9026
rect 5088 8986 5500 8990
rect 4586 8938 4990 8986
rect 4086 8888 4488 8938
rect 3566 8858 3988 8888
rect 3074 8800 3468 8858
rect 2564 8760 2976 8800
tri 2976 8760 3016 8800 sw
tri 3074 8760 3114 8800 ne
rect 3114 8760 3468 8800
tri 3468 8760 3566 8858 sw
tri 3566 8760 3664 8858 ne
rect 3664 8800 3988 8858
tri 3988 8800 4076 8888 sw
tri 4086 8800 4174 8888 ne
rect 4174 8858 4488 8888
tri 4488 8858 4568 8938 sw
tri 4586 8858 4666 8938 ne
rect 4666 8888 4990 8938
tri 4990 8888 5088 8986 sw
tri 5088 8888 5186 8986 ne
rect 5186 8938 5500 8986
tri 5500 8938 5588 9026 sw
tri 5598 8938 5686 9026 ne
rect 5686 8990 5740 9026
rect 5860 9026 5962 9110
tri 5962 9026 6050 9114 sw
tri 6060 9026 6148 9114 ne
rect 6148 9110 6512 9114
rect 6148 9026 6290 9110
rect 5860 8990 6050 9026
rect 5686 8986 6050 8990
tri 6050 8986 6090 9026 sw
tri 6148 8986 6188 9026 ne
rect 6188 8990 6290 9026
rect 6410 9026 6512 9110
tri 6512 9026 6600 9114 sw
tri 6610 9026 6698 9114 ne
rect 6698 9110 7062 9114
rect 6698 9026 6840 9110
rect 6410 8990 6600 9026
rect 6188 8986 6600 8990
rect 5686 8938 6090 8986
rect 5186 8888 5588 8938
rect 4666 8858 5088 8888
rect 4174 8800 4568 8858
rect 3664 8760 4076 8800
tri 4076 8760 4116 8800 sw
tri 4174 8760 4214 8800 ne
rect 4214 8760 4568 8800
tri 4568 8760 4666 8858 sw
tri 4666 8760 4764 8858 ne
rect 4764 8800 5088 8858
tri 5088 8800 5176 8888 sw
tri 5186 8800 5274 8888 ne
rect 5274 8858 5588 8888
tri 5588 8858 5668 8938 sw
tri 5686 8858 5766 8938 ne
rect 5766 8888 6090 8938
tri 6090 8888 6188 8986 sw
tri 6188 8888 6286 8986 ne
rect 6286 8938 6600 8986
tri 6600 8938 6688 9026 sw
tri 6698 8938 6786 9026 ne
rect 6786 8990 6840 9026
rect 6960 9026 7062 9110
tri 7062 9026 7150 9114 sw
tri 7160 9026 7248 9114 ne
rect 7248 9110 7612 9114
rect 7248 9026 7390 9110
rect 6960 8990 7150 9026
rect 6786 8986 7150 8990
tri 7150 8986 7190 9026 sw
tri 7248 8986 7288 9026 ne
rect 7288 8990 7390 9026
rect 7510 9026 7612 9110
tri 7612 9026 7700 9114 sw
tri 7710 9026 7798 9114 ne
rect 7798 9110 8162 9114
rect 7798 9026 7940 9110
rect 7510 8990 7700 9026
rect 7288 8986 7700 8990
rect 6786 8938 7190 8986
rect 6286 8888 6688 8938
rect 5766 8858 6188 8888
rect 5274 8800 5668 8858
rect 4764 8760 5176 8800
tri 5176 8760 5216 8800 sw
tri 5274 8760 5314 8800 ne
rect 5314 8760 5668 8800
tri 5668 8760 5766 8858 sw
tri 5766 8760 5864 8858 ne
rect 5864 8800 6188 8858
tri 6188 8800 6276 8888 sw
tri 6286 8800 6374 8888 ne
rect 6374 8858 6688 8888
tri 6688 8858 6768 8938 sw
tri 6786 8858 6866 8938 ne
rect 6866 8888 7190 8938
tri 7190 8888 7288 8986 sw
tri 7288 8888 7386 8986 ne
rect 7386 8938 7700 8986
tri 7700 8938 7788 9026 sw
tri 7798 8938 7886 9026 ne
rect 7886 8990 7940 9026
rect 8060 9026 8162 9110
tri 8162 9026 8250 9114 sw
tri 8260 9026 8348 9114 ne
rect 8348 9110 8712 9114
rect 8348 9026 8490 9110
rect 8060 8990 8250 9026
rect 7886 8986 8250 8990
tri 8250 8986 8290 9026 sw
tri 8348 8986 8388 9026 ne
rect 8388 8990 8490 9026
rect 8610 9026 8712 9110
tri 8712 9026 8800 9114 sw
tri 8810 9026 8898 9114 ne
rect 8898 9110 9262 9114
rect 8898 9026 9040 9110
rect 8610 8990 8800 9026
rect 8388 8986 8800 8990
rect 7886 8938 8290 8986
rect 7386 8888 7788 8938
rect 6866 8858 7288 8888
rect 6374 8800 6768 8858
rect 5864 8760 6276 8800
tri 6276 8760 6316 8800 sw
tri 6374 8760 6414 8800 ne
rect 6414 8760 6768 8800
tri 6768 8760 6866 8858 sw
tri 6866 8760 6964 8858 ne
rect 6964 8800 7288 8858
tri 7288 8800 7376 8888 sw
tri 7386 8800 7474 8888 ne
rect 7474 8858 7788 8888
tri 7788 8858 7868 8938 sw
tri 7886 8858 7966 8938 ne
rect 7966 8888 8290 8938
tri 8290 8888 8388 8986 sw
tri 8388 8888 8486 8986 ne
rect 8486 8938 8800 8986
tri 8800 8938 8888 9026 sw
tri 8898 8938 8986 9026 ne
rect 8986 8990 9040 9026
rect 9160 9026 9262 9110
tri 9262 9026 9350 9114 sw
tri 9360 9026 9448 9114 ne
rect 9448 9110 9812 9114
rect 9448 9026 9590 9110
rect 9160 8990 9350 9026
rect 8986 8986 9350 8990
tri 9350 8986 9390 9026 sw
tri 9448 8986 9488 9026 ne
rect 9488 8990 9590 9026
rect 9710 9026 9812 9110
tri 9812 9026 9900 9114 sw
tri 9910 9026 9998 9114 ne
rect 9998 9110 10362 9114
rect 9998 9026 10140 9110
rect 9710 8990 9900 9026
rect 9488 8986 9900 8990
rect 8986 8938 9390 8986
rect 8486 8888 8888 8938
rect 7966 8858 8388 8888
rect 7474 8800 7868 8858
rect 6964 8760 7376 8800
tri 7376 8760 7416 8800 sw
tri 7474 8760 7514 8800 ne
rect 7514 8760 7868 8800
tri 7868 8760 7966 8858 sw
tri 7966 8760 8064 8858 ne
rect 8064 8800 8388 8858
tri 8388 8800 8476 8888 sw
tri 8486 8800 8574 8888 ne
rect 8574 8858 8888 8888
tri 8888 8858 8968 8938 sw
tri 8986 8858 9066 8938 ne
rect 9066 8888 9390 8938
tri 9390 8888 9488 8986 sw
tri 9488 8888 9586 8986 ne
rect 9586 8938 9900 8986
tri 9900 8938 9988 9026 sw
tri 9998 8938 10086 9026 ne
rect 10086 8990 10140 9026
rect 10260 9026 10362 9110
tri 10362 9026 10450 9114 sw
tri 10460 9026 10548 9114 ne
rect 10548 9110 10912 9114
rect 10548 9026 10690 9110
rect 10260 8990 10450 9026
rect 10086 8986 10450 8990
tri 10450 8986 10490 9026 sw
tri 10548 8986 10588 9026 ne
rect 10588 8990 10690 9026
rect 10810 9026 10912 9110
tri 10912 9026 11000 9114 sw
tri 11010 9026 11098 9114 ne
rect 11098 9110 11462 9114
rect 11098 9026 11240 9110
rect 10810 8990 11000 9026
rect 10588 8986 11000 8990
rect 10086 8938 10490 8986
rect 9586 8888 9988 8938
rect 9066 8858 9488 8888
rect 8574 8800 8968 8858
rect 8064 8760 8476 8800
tri 8476 8760 8516 8800 sw
tri 8574 8760 8614 8800 ne
rect 8614 8760 8968 8800
tri 8968 8760 9066 8858 sw
tri 9066 8760 9164 8858 ne
rect 9164 8800 9488 8858
tri 9488 8800 9576 8888 sw
tri 9586 8800 9674 8888 ne
rect 9674 8858 9988 8888
tri 9988 8858 10068 8938 sw
tri 10086 8858 10166 8938 ne
rect 10166 8888 10490 8938
tri 10490 8888 10588 8986 sw
tri 10588 8888 10686 8986 ne
rect 10686 8938 11000 8986
tri 11000 8938 11088 9026 sw
tri 11098 8938 11186 9026 ne
rect 11186 8990 11240 9026
rect 11360 9026 11462 9110
tri 11462 9026 11550 9114 sw
tri 11560 9026 11648 9114 ne
rect 11648 9110 12012 9114
rect 11648 9026 11790 9110
rect 11360 8990 11550 9026
rect 11186 8986 11550 8990
tri 11550 8986 11590 9026 sw
tri 11648 8986 11688 9026 ne
rect 11688 8990 11790 9026
rect 11910 9026 12012 9110
tri 12012 9026 12100 9114 sw
tri 12110 9026 12198 9114 ne
rect 12198 9110 12562 9114
rect 12198 9026 12340 9110
rect 11910 8990 12100 9026
rect 11688 8986 12100 8990
rect 11186 8938 11590 8986
rect 10686 8888 11088 8938
rect 10166 8858 10588 8888
rect 9674 8800 10068 8858
rect 9164 8760 9576 8800
tri 9576 8760 9616 8800 sw
tri 9674 8760 9714 8800 ne
rect 9714 8760 10068 8800
tri 10068 8760 10166 8858 sw
tri 10166 8760 10264 8858 ne
rect 10264 8800 10588 8858
tri 10588 8800 10676 8888 sw
tri 10686 8800 10774 8888 ne
rect 10774 8858 11088 8888
tri 11088 8858 11168 8938 sw
tri 11186 8858 11266 8938 ne
rect 11266 8888 11590 8938
tri 11590 8888 11688 8986 sw
tri 11688 8888 11786 8986 ne
rect 11786 8938 12100 8986
tri 12100 8938 12188 9026 sw
tri 12198 8938 12286 9026 ne
rect 12286 8990 12340 9026
rect 12460 9026 12562 9110
tri 12562 9026 12650 9114 sw
tri 12660 9026 12748 9114 ne
rect 12748 9110 13112 9114
rect 12748 9026 12890 9110
rect 12460 8990 12650 9026
rect 12286 8986 12650 8990
tri 12650 8986 12690 9026 sw
tri 12748 8986 12788 9026 ne
rect 12788 8990 12890 9026
rect 13010 9026 13112 9110
tri 13112 9026 13200 9114 sw
tri 13210 9026 13298 9114 ne
rect 13298 9110 15775 9114
rect 13298 9026 13440 9110
rect 13010 8990 13200 9026
rect 12788 8986 13200 8990
rect 12286 8938 12690 8986
rect 11786 8888 12188 8938
rect 11266 8858 11688 8888
rect 10774 8800 11168 8858
rect 10264 8760 10676 8800
tri 10676 8760 10716 8800 sw
tri 10774 8760 10814 8800 ne
rect 10814 8760 11168 8800
tri 11168 8760 11266 8858 sw
tri 11266 8760 11364 8858 ne
rect 11364 8800 11688 8858
tri 11688 8800 11776 8888 sw
tri 11786 8800 11874 8888 ne
rect 11874 8858 12188 8888
tri 12188 8858 12268 8938 sw
tri 12286 8858 12366 8938 ne
rect 12366 8888 12690 8938
tri 12690 8888 12788 8986 sw
tri 12788 8888 12886 8986 ne
rect 12886 8938 13200 8986
tri 13200 8938 13288 9026 sw
tri 13298 8938 13386 9026 ne
rect 13386 8990 13440 9026
rect 13560 8990 15775 9110
rect 13386 8938 15775 8990
rect 12886 8888 13288 8938
rect 12366 8858 12788 8888
rect 11874 8800 12268 8858
rect 11364 8760 11776 8800
tri 11776 8760 11816 8800 sw
tri 11874 8760 11914 8800 ne
rect 11914 8760 12268 8800
tri 12268 8760 12366 8858 sw
tri 12366 8760 12464 8858 ne
rect 12464 8800 12788 8858
tri 12788 8800 12876 8888 sw
tri 12886 8800 12974 8888 ne
rect 12974 8858 13288 8888
tri 13288 8858 13368 8938 sw
tri 13386 8858 13466 8938 ne
rect 13466 8858 14075 8938
rect 12974 8800 13368 8858
rect 12464 8760 12876 8800
tri 12876 8760 12916 8800 sw
tri 12974 8760 13014 8800 ne
rect 13014 8760 13368 8800
tri 13368 8760 13466 8858 sw
tri 13466 8760 13564 8858 ne
rect 13564 8838 14075 8858
rect 14175 8838 15775 8938
rect 13564 8760 15775 8838
rect -1025 8712 -284 8760
rect -1025 8612 -925 8712
rect -825 8662 -284 8712
tri -284 8662 -186 8760 sw
tri -186 8662 -88 8760 ne
rect -88 8662 266 8760
tri 266 8662 364 8760 sw
tri 364 8662 462 8760 ne
rect 462 8662 816 8760
tri 816 8662 914 8760 sw
tri 914 8662 1012 8760 ne
rect 1012 8662 1366 8760
tri 1366 8662 1464 8760 sw
tri 1464 8662 1562 8760 ne
rect 1562 8662 1916 8760
tri 1916 8662 2014 8760 sw
tri 2014 8662 2112 8760 ne
rect 2112 8662 2466 8760
tri 2466 8662 2564 8760 sw
tri 2564 8662 2662 8760 ne
rect 2662 8662 3016 8760
tri 3016 8662 3114 8760 sw
tri 3114 8662 3212 8760 ne
rect 3212 8662 3566 8760
tri 3566 8662 3664 8760 sw
tri 3664 8662 3762 8760 ne
rect 3762 8662 4116 8760
tri 4116 8662 4214 8760 sw
tri 4214 8662 4312 8760 ne
rect 4312 8662 4666 8760
tri 4666 8662 4764 8760 sw
tri 4764 8662 4862 8760 ne
rect 4862 8662 5216 8760
tri 5216 8662 5314 8760 sw
tri 5314 8662 5412 8760 ne
rect 5412 8662 5766 8760
tri 5766 8662 5864 8760 sw
tri 5864 8662 5962 8760 ne
rect 5962 8662 6316 8760
tri 6316 8662 6414 8760 sw
tri 6414 8662 6512 8760 ne
rect 6512 8662 6866 8760
tri 6866 8662 6964 8760 sw
tri 6964 8662 7062 8760 ne
rect 7062 8662 7416 8760
tri 7416 8662 7514 8760 sw
tri 7514 8662 7612 8760 ne
rect 7612 8662 7966 8760
tri 7966 8662 8064 8760 sw
tri 8064 8662 8162 8760 ne
rect 8162 8662 8516 8760
tri 8516 8662 8614 8760 sw
tri 8614 8662 8712 8760 ne
rect 8712 8662 9066 8760
tri 9066 8662 9164 8760 sw
tri 9164 8662 9262 8760 ne
rect 9262 8662 9616 8760
tri 9616 8662 9714 8760 sw
tri 9714 8662 9812 8760 ne
rect 9812 8662 10166 8760
tri 10166 8662 10264 8760 sw
tri 10264 8662 10362 8760 ne
rect 10362 8662 10716 8760
tri 10716 8662 10814 8760 sw
tri 10814 8662 10912 8760 ne
rect 10912 8662 11266 8760
tri 11266 8662 11364 8760 sw
tri 11364 8662 11462 8760 ne
rect 11462 8662 11816 8760
tri 11816 8662 11914 8760 sw
tri 11914 8662 12012 8760 ne
rect 12012 8662 12366 8760
tri 12366 8662 12464 8760 sw
tri 12464 8662 12562 8760 ne
rect 12562 8662 12916 8760
tri 12916 8662 13014 8760 sw
tri 13014 8662 13112 8760 ne
rect 13112 8662 13466 8760
tri 13466 8662 13564 8760 sw
tri 13564 8662 13662 8760 ne
rect 13662 8662 15775 8760
rect -825 8612 -186 8662
rect -1025 8564 -186 8612
tri -186 8564 -88 8662 sw
tri -88 8564 10 8662 ne
rect 10 8564 364 8662
tri 364 8564 462 8662 sw
tri 462 8564 560 8662 ne
rect 560 8564 914 8662
tri 914 8564 1012 8662 sw
tri 1012 8564 1110 8662 ne
rect 1110 8564 1464 8662
tri 1464 8564 1562 8662 sw
tri 1562 8564 1660 8662 ne
rect 1660 8564 2014 8662
tri 2014 8564 2112 8662 sw
tri 2112 8564 2210 8662 ne
rect 2210 8564 2564 8662
tri 2564 8564 2662 8662 sw
tri 2662 8564 2760 8662 ne
rect 2760 8564 3114 8662
tri 3114 8564 3212 8662 sw
tri 3212 8564 3310 8662 ne
rect 3310 8564 3664 8662
tri 3664 8564 3762 8662 sw
tri 3762 8564 3860 8662 ne
rect 3860 8564 4214 8662
tri 4214 8564 4312 8662 sw
tri 4312 8564 4410 8662 ne
rect 4410 8564 4764 8662
tri 4764 8564 4862 8662 sw
tri 4862 8564 4960 8662 ne
rect 4960 8564 5314 8662
tri 5314 8564 5412 8662 sw
tri 5412 8564 5510 8662 ne
rect 5510 8564 5864 8662
tri 5864 8564 5962 8662 sw
tri 5962 8564 6060 8662 ne
rect 6060 8564 6414 8662
tri 6414 8564 6512 8662 sw
tri 6512 8564 6610 8662 ne
rect 6610 8564 6964 8662
tri 6964 8564 7062 8662 sw
tri 7062 8564 7160 8662 ne
rect 7160 8564 7514 8662
tri 7514 8564 7612 8662 sw
tri 7612 8564 7710 8662 ne
rect 7710 8564 8064 8662
tri 8064 8564 8162 8662 sw
tri 8162 8564 8260 8662 ne
rect 8260 8564 8614 8662
tri 8614 8564 8712 8662 sw
tri 8712 8564 8810 8662 ne
rect 8810 8564 9164 8662
tri 9164 8564 9262 8662 sw
tri 9262 8564 9360 8662 ne
rect 9360 8564 9714 8662
tri 9714 8564 9812 8662 sw
tri 9812 8564 9910 8662 ne
rect 9910 8564 10264 8662
tri 10264 8564 10362 8662 sw
tri 10362 8564 10460 8662 ne
rect 10460 8564 10814 8662
tri 10814 8564 10912 8662 sw
tri 10912 8564 11010 8662 ne
rect 11010 8564 11364 8662
tri 11364 8564 11462 8662 sw
tri 11462 8564 11560 8662 ne
rect 11560 8564 11914 8662
tri 11914 8564 12012 8662 sw
tri 12012 8564 12110 8662 ne
rect 12110 8564 12464 8662
tri 12464 8564 12562 8662 sw
tri 12562 8564 12660 8662 ne
rect 12660 8564 13014 8662
tri 13014 8564 13112 8662 sw
tri 13112 8564 13210 8662 ne
rect 13210 8564 13564 8662
tri 13564 8564 13662 8662 sw
rect -1025 8560 -88 8564
rect -1025 8440 -310 8560
rect -190 8476 -88 8560
tri -88 8476 0 8564 sw
tri 10 8476 98 8564 ne
rect 98 8560 462 8564
rect 98 8476 240 8560
rect -190 8440 0 8476
rect -1025 8436 0 8440
tri 0 8436 40 8476 sw
tri 98 8436 138 8476 ne
rect 138 8440 240 8476
rect 360 8476 462 8560
tri 462 8476 550 8564 sw
tri 560 8476 648 8564 ne
rect 648 8560 1012 8564
rect 648 8476 790 8560
rect 360 8440 550 8476
rect 138 8436 550 8440
tri -412 8338 -314 8436 ne
rect -314 8338 40 8436
tri 40 8338 138 8436 sw
tri 138 8338 236 8436 ne
rect 236 8388 550 8436
tri 550 8388 638 8476 sw
tri 648 8388 736 8476 ne
rect 736 8440 790 8476
rect 910 8476 1012 8560
tri 1012 8476 1100 8564 sw
tri 1110 8476 1198 8564 ne
rect 1198 8560 1562 8564
rect 1198 8476 1340 8560
rect 910 8440 1100 8476
rect 736 8436 1100 8440
tri 1100 8436 1140 8476 sw
tri 1198 8436 1238 8476 ne
rect 1238 8440 1340 8476
rect 1460 8476 1562 8560
tri 1562 8476 1650 8564 sw
tri 1660 8476 1748 8564 ne
rect 1748 8560 2112 8564
rect 1748 8476 1890 8560
rect 1460 8440 1650 8476
rect 1238 8436 1650 8440
rect 736 8388 1140 8436
rect 236 8338 638 8388
rect -2525 8250 -412 8338
tri -412 8250 -324 8338 sw
tri -314 8250 -226 8338 ne
rect -226 8250 138 8338
tri 138 8250 226 8338 sw
tri 236 8250 324 8338 ne
rect 324 8308 638 8338
tri 638 8308 718 8388 sw
tri 736 8308 816 8388 ne
rect 816 8338 1140 8388
tri 1140 8338 1238 8436 sw
tri 1238 8338 1336 8436 ne
rect 1336 8388 1650 8436
tri 1650 8388 1738 8476 sw
tri 1748 8388 1836 8476 ne
rect 1836 8440 1890 8476
rect 2010 8476 2112 8560
tri 2112 8476 2200 8564 sw
tri 2210 8476 2298 8564 ne
rect 2298 8560 2662 8564
rect 2298 8476 2440 8560
rect 2010 8440 2200 8476
rect 1836 8436 2200 8440
tri 2200 8436 2240 8476 sw
tri 2298 8436 2338 8476 ne
rect 2338 8440 2440 8476
rect 2560 8476 2662 8560
tri 2662 8476 2750 8564 sw
tri 2760 8476 2848 8564 ne
rect 2848 8560 3212 8564
rect 2848 8476 2990 8560
rect 2560 8440 2750 8476
rect 2338 8436 2750 8440
rect 1836 8388 2240 8436
rect 1336 8338 1738 8388
rect 816 8308 1238 8338
rect 324 8250 718 8308
rect -2525 8210 -324 8250
tri -324 8210 -284 8250 sw
tri -226 8210 -186 8250 ne
rect -186 8210 226 8250
tri 226 8210 266 8250 sw
tri 324 8210 364 8250 ne
rect 364 8210 718 8250
tri 718 8210 816 8308 sw
tri 816 8210 914 8308 ne
rect 914 8250 1238 8308
tri 1238 8250 1326 8338 sw
tri 1336 8250 1424 8338 ne
rect 1424 8308 1738 8338
tri 1738 8308 1818 8388 sw
tri 1836 8308 1916 8388 ne
rect 1916 8338 2240 8388
tri 2240 8338 2338 8436 sw
tri 2338 8338 2436 8436 ne
rect 2436 8388 2750 8436
tri 2750 8388 2838 8476 sw
tri 2848 8388 2936 8476 ne
rect 2936 8440 2990 8476
rect 3110 8476 3212 8560
tri 3212 8476 3300 8564 sw
tri 3310 8476 3398 8564 ne
rect 3398 8560 3762 8564
rect 3398 8476 3540 8560
rect 3110 8440 3300 8476
rect 2936 8436 3300 8440
tri 3300 8436 3340 8476 sw
tri 3398 8436 3438 8476 ne
rect 3438 8440 3540 8476
rect 3660 8476 3762 8560
tri 3762 8476 3850 8564 sw
tri 3860 8476 3948 8564 ne
rect 3948 8560 4312 8564
rect 3948 8476 4090 8560
rect 3660 8440 3850 8476
rect 3438 8436 3850 8440
rect 2936 8388 3340 8436
rect 2436 8338 2838 8388
rect 1916 8308 2338 8338
rect 1424 8250 1818 8308
rect 914 8210 1326 8250
tri 1326 8210 1366 8250 sw
tri 1424 8210 1464 8250 ne
rect 1464 8210 1818 8250
tri 1818 8210 1916 8308 sw
tri 1916 8210 2014 8308 ne
rect 2014 8250 2338 8308
tri 2338 8250 2426 8338 sw
tri 2436 8250 2524 8338 ne
rect 2524 8308 2838 8338
tri 2838 8308 2918 8388 sw
tri 2936 8308 3016 8388 ne
rect 3016 8338 3340 8388
tri 3340 8338 3438 8436 sw
tri 3438 8338 3536 8436 ne
rect 3536 8388 3850 8436
tri 3850 8388 3938 8476 sw
tri 3948 8388 4036 8476 ne
rect 4036 8440 4090 8476
rect 4210 8476 4312 8560
tri 4312 8476 4400 8564 sw
tri 4410 8476 4498 8564 ne
rect 4498 8560 4862 8564
rect 4498 8476 4640 8560
rect 4210 8440 4400 8476
rect 4036 8436 4400 8440
tri 4400 8436 4440 8476 sw
tri 4498 8436 4538 8476 ne
rect 4538 8440 4640 8476
rect 4760 8476 4862 8560
tri 4862 8476 4950 8564 sw
tri 4960 8476 5048 8564 ne
rect 5048 8560 5412 8564
rect 5048 8476 5190 8560
rect 4760 8440 4950 8476
rect 4538 8436 4950 8440
rect 4036 8388 4440 8436
rect 3536 8338 3938 8388
rect 3016 8308 3438 8338
rect 2524 8250 2918 8308
rect 2014 8210 2426 8250
tri 2426 8210 2466 8250 sw
tri 2524 8210 2564 8250 ne
rect 2564 8210 2918 8250
tri 2918 8210 3016 8308 sw
tri 3016 8210 3114 8308 ne
rect 3114 8250 3438 8308
tri 3438 8250 3526 8338 sw
tri 3536 8250 3624 8338 ne
rect 3624 8308 3938 8338
tri 3938 8308 4018 8388 sw
tri 4036 8308 4116 8388 ne
rect 4116 8338 4440 8388
tri 4440 8338 4538 8436 sw
tri 4538 8338 4636 8436 ne
rect 4636 8388 4950 8436
tri 4950 8388 5038 8476 sw
tri 5048 8388 5136 8476 ne
rect 5136 8440 5190 8476
rect 5310 8476 5412 8560
tri 5412 8476 5500 8564 sw
tri 5510 8476 5598 8564 ne
rect 5598 8560 5962 8564
rect 5598 8476 5740 8560
rect 5310 8440 5500 8476
rect 5136 8436 5500 8440
tri 5500 8436 5540 8476 sw
tri 5598 8436 5638 8476 ne
rect 5638 8440 5740 8476
rect 5860 8476 5962 8560
tri 5962 8476 6050 8564 sw
tri 6060 8476 6148 8564 ne
rect 6148 8560 6512 8564
rect 6148 8476 6290 8560
rect 5860 8440 6050 8476
rect 5638 8436 6050 8440
rect 5136 8388 5540 8436
rect 4636 8338 5038 8388
rect 4116 8308 4538 8338
rect 3624 8250 4018 8308
rect 3114 8210 3526 8250
tri 3526 8210 3566 8250 sw
tri 3624 8210 3664 8250 ne
rect 3664 8210 4018 8250
tri 4018 8210 4116 8308 sw
tri 4116 8210 4214 8308 ne
rect 4214 8250 4538 8308
tri 4538 8250 4626 8338 sw
tri 4636 8250 4724 8338 ne
rect 4724 8308 5038 8338
tri 5038 8308 5118 8388 sw
tri 5136 8308 5216 8388 ne
rect 5216 8338 5540 8388
tri 5540 8338 5638 8436 sw
tri 5638 8338 5736 8436 ne
rect 5736 8388 6050 8436
tri 6050 8388 6138 8476 sw
tri 6148 8388 6236 8476 ne
rect 6236 8440 6290 8476
rect 6410 8476 6512 8560
tri 6512 8476 6600 8564 sw
tri 6610 8476 6698 8564 ne
rect 6698 8560 7062 8564
rect 6698 8476 6840 8560
rect 6410 8440 6600 8476
rect 6236 8436 6600 8440
tri 6600 8436 6640 8476 sw
tri 6698 8436 6738 8476 ne
rect 6738 8440 6840 8476
rect 6960 8476 7062 8560
tri 7062 8476 7150 8564 sw
tri 7160 8476 7248 8564 ne
rect 7248 8560 7612 8564
rect 7248 8476 7390 8560
rect 6960 8440 7150 8476
rect 6738 8436 7150 8440
rect 6236 8388 6640 8436
rect 5736 8338 6138 8388
rect 5216 8308 5638 8338
rect 4724 8250 5118 8308
rect 4214 8210 4626 8250
tri 4626 8210 4666 8250 sw
tri 4724 8210 4764 8250 ne
rect 4764 8210 5118 8250
tri 5118 8210 5216 8308 sw
tri 5216 8210 5314 8308 ne
rect 5314 8250 5638 8308
tri 5638 8250 5726 8338 sw
tri 5736 8250 5824 8338 ne
rect 5824 8308 6138 8338
tri 6138 8308 6218 8388 sw
tri 6236 8308 6316 8388 ne
rect 6316 8338 6640 8388
tri 6640 8338 6738 8436 sw
tri 6738 8338 6836 8436 ne
rect 6836 8388 7150 8436
tri 7150 8388 7238 8476 sw
tri 7248 8388 7336 8476 ne
rect 7336 8440 7390 8476
rect 7510 8476 7612 8560
tri 7612 8476 7700 8564 sw
tri 7710 8476 7798 8564 ne
rect 7798 8560 8162 8564
rect 7798 8476 7940 8560
rect 7510 8440 7700 8476
rect 7336 8436 7700 8440
tri 7700 8436 7740 8476 sw
tri 7798 8436 7838 8476 ne
rect 7838 8440 7940 8476
rect 8060 8476 8162 8560
tri 8162 8476 8250 8564 sw
tri 8260 8476 8348 8564 ne
rect 8348 8560 8712 8564
rect 8348 8476 8490 8560
rect 8060 8440 8250 8476
rect 7838 8436 8250 8440
rect 7336 8388 7740 8436
rect 6836 8338 7238 8388
rect 6316 8308 6738 8338
rect 5824 8250 6218 8308
rect 5314 8210 5726 8250
tri 5726 8210 5766 8250 sw
tri 5824 8210 5864 8250 ne
rect 5864 8210 6218 8250
tri 6218 8210 6316 8308 sw
tri 6316 8210 6414 8308 ne
rect 6414 8250 6738 8308
tri 6738 8250 6826 8338 sw
tri 6836 8250 6924 8338 ne
rect 6924 8308 7238 8338
tri 7238 8308 7318 8388 sw
tri 7336 8308 7416 8388 ne
rect 7416 8338 7740 8388
tri 7740 8338 7838 8436 sw
tri 7838 8338 7936 8436 ne
rect 7936 8388 8250 8436
tri 8250 8388 8338 8476 sw
tri 8348 8388 8436 8476 ne
rect 8436 8440 8490 8476
rect 8610 8476 8712 8560
tri 8712 8476 8800 8564 sw
tri 8810 8476 8898 8564 ne
rect 8898 8560 9262 8564
rect 8898 8476 9040 8560
rect 8610 8440 8800 8476
rect 8436 8436 8800 8440
tri 8800 8436 8840 8476 sw
tri 8898 8436 8938 8476 ne
rect 8938 8440 9040 8476
rect 9160 8476 9262 8560
tri 9262 8476 9350 8564 sw
tri 9360 8476 9448 8564 ne
rect 9448 8560 9812 8564
rect 9448 8476 9590 8560
rect 9160 8440 9350 8476
rect 8938 8436 9350 8440
rect 8436 8388 8840 8436
rect 7936 8338 8338 8388
rect 7416 8308 7838 8338
rect 6924 8250 7318 8308
rect 6414 8210 6826 8250
tri 6826 8210 6866 8250 sw
tri 6924 8210 6964 8250 ne
rect 6964 8210 7318 8250
tri 7318 8210 7416 8308 sw
tri 7416 8210 7514 8308 ne
rect 7514 8250 7838 8308
tri 7838 8250 7926 8338 sw
tri 7936 8250 8024 8338 ne
rect 8024 8308 8338 8338
tri 8338 8308 8418 8388 sw
tri 8436 8308 8516 8388 ne
rect 8516 8338 8840 8388
tri 8840 8338 8938 8436 sw
tri 8938 8338 9036 8436 ne
rect 9036 8388 9350 8436
tri 9350 8388 9438 8476 sw
tri 9448 8388 9536 8476 ne
rect 9536 8440 9590 8476
rect 9710 8476 9812 8560
tri 9812 8476 9900 8564 sw
tri 9910 8476 9998 8564 ne
rect 9998 8560 10362 8564
rect 9998 8476 10140 8560
rect 9710 8440 9900 8476
rect 9536 8436 9900 8440
tri 9900 8436 9940 8476 sw
tri 9998 8436 10038 8476 ne
rect 10038 8440 10140 8476
rect 10260 8476 10362 8560
tri 10362 8476 10450 8564 sw
tri 10460 8476 10548 8564 ne
rect 10548 8560 10912 8564
rect 10548 8476 10690 8560
rect 10260 8440 10450 8476
rect 10038 8436 10450 8440
rect 9536 8388 9940 8436
rect 9036 8338 9438 8388
rect 8516 8308 8938 8338
rect 8024 8250 8418 8308
rect 7514 8210 7926 8250
tri 7926 8210 7966 8250 sw
tri 8024 8210 8064 8250 ne
rect 8064 8210 8418 8250
tri 8418 8210 8516 8308 sw
tri 8516 8210 8614 8308 ne
rect 8614 8250 8938 8308
tri 8938 8250 9026 8338 sw
tri 9036 8250 9124 8338 ne
rect 9124 8308 9438 8338
tri 9438 8308 9518 8388 sw
tri 9536 8308 9616 8388 ne
rect 9616 8338 9940 8388
tri 9940 8338 10038 8436 sw
tri 10038 8338 10136 8436 ne
rect 10136 8388 10450 8436
tri 10450 8388 10538 8476 sw
tri 10548 8388 10636 8476 ne
rect 10636 8440 10690 8476
rect 10810 8476 10912 8560
tri 10912 8476 11000 8564 sw
tri 11010 8476 11098 8564 ne
rect 11098 8560 11462 8564
rect 11098 8476 11240 8560
rect 10810 8440 11000 8476
rect 10636 8436 11000 8440
tri 11000 8436 11040 8476 sw
tri 11098 8436 11138 8476 ne
rect 11138 8440 11240 8476
rect 11360 8476 11462 8560
tri 11462 8476 11550 8564 sw
tri 11560 8476 11648 8564 ne
rect 11648 8560 12012 8564
rect 11648 8476 11790 8560
rect 11360 8440 11550 8476
rect 11138 8436 11550 8440
rect 10636 8388 11040 8436
rect 10136 8338 10538 8388
rect 9616 8308 10038 8338
rect 9124 8250 9518 8308
rect 8614 8210 9026 8250
tri 9026 8210 9066 8250 sw
tri 9124 8210 9164 8250 ne
rect 9164 8210 9518 8250
tri 9518 8210 9616 8308 sw
tri 9616 8210 9714 8308 ne
rect 9714 8250 10038 8308
tri 10038 8250 10126 8338 sw
tri 10136 8250 10224 8338 ne
rect 10224 8308 10538 8338
tri 10538 8308 10618 8388 sw
tri 10636 8308 10716 8388 ne
rect 10716 8338 11040 8388
tri 11040 8338 11138 8436 sw
tri 11138 8338 11236 8436 ne
rect 11236 8388 11550 8436
tri 11550 8388 11638 8476 sw
tri 11648 8388 11736 8476 ne
rect 11736 8440 11790 8476
rect 11910 8476 12012 8560
tri 12012 8476 12100 8564 sw
tri 12110 8476 12198 8564 ne
rect 12198 8560 12562 8564
rect 12198 8476 12340 8560
rect 11910 8440 12100 8476
rect 11736 8436 12100 8440
tri 12100 8436 12140 8476 sw
tri 12198 8436 12238 8476 ne
rect 12238 8440 12340 8476
rect 12460 8476 12562 8560
tri 12562 8476 12650 8564 sw
tri 12660 8476 12748 8564 ne
rect 12748 8560 13112 8564
rect 12748 8476 12890 8560
rect 12460 8440 12650 8476
rect 12238 8436 12650 8440
rect 11736 8388 12140 8436
rect 11236 8338 11638 8388
rect 10716 8308 11138 8338
rect 10224 8250 10618 8308
rect 9714 8210 10126 8250
tri 10126 8210 10166 8250 sw
tri 10224 8210 10264 8250 ne
rect 10264 8210 10618 8250
tri 10618 8210 10716 8308 sw
tri 10716 8210 10814 8308 ne
rect 10814 8250 11138 8308
tri 11138 8250 11226 8338 sw
tri 11236 8250 11324 8338 ne
rect 11324 8308 11638 8338
tri 11638 8308 11718 8388 sw
tri 11736 8308 11816 8388 ne
rect 11816 8338 12140 8388
tri 12140 8338 12238 8436 sw
tri 12238 8338 12336 8436 ne
rect 12336 8388 12650 8436
tri 12650 8388 12738 8476 sw
tri 12748 8388 12836 8476 ne
rect 12836 8440 12890 8476
rect 13010 8476 13112 8560
tri 13112 8476 13200 8564 sw
tri 13210 8476 13298 8564 ne
rect 13298 8560 14275 8564
rect 13298 8476 13440 8560
rect 13010 8440 13200 8476
rect 12836 8436 13200 8440
tri 13200 8436 13240 8476 sw
tri 13298 8436 13338 8476 ne
rect 13338 8440 13440 8476
rect 13560 8440 14275 8560
rect 13338 8436 14275 8440
rect 12836 8388 13240 8436
rect 12336 8338 12738 8388
rect 11816 8308 12238 8338
rect 11324 8250 11718 8308
rect 10814 8210 11226 8250
tri 11226 8210 11266 8250 sw
tri 11324 8210 11364 8250 ne
rect 11364 8210 11718 8250
tri 11718 8210 11816 8308 sw
tri 11816 8210 11914 8308 ne
rect 11914 8250 12238 8308
tri 12238 8250 12326 8338 sw
tri 12336 8250 12424 8338 ne
rect 12424 8308 12738 8338
tri 12738 8308 12818 8388 sw
tri 12836 8308 12916 8388 ne
rect 12916 8338 13240 8388
tri 13240 8338 13338 8436 sw
tri 13338 8338 13436 8436 ne
rect 13436 8338 14275 8436
rect 12916 8308 13338 8338
rect 12424 8250 12818 8308
rect 11914 8210 12326 8250
tri 12326 8210 12366 8250 sw
tri 12424 8210 12464 8250 ne
rect 12464 8210 12818 8250
tri 12818 8210 12916 8308 sw
tri 12916 8210 13014 8308 ne
rect 13014 8250 13338 8308
tri 13338 8250 13426 8338 sw
tri 13436 8250 13524 8338 ne
rect 13524 8250 14275 8338
rect 13014 8210 13426 8250
tri 13426 8210 13466 8250 sw
tri 13524 8210 13564 8250 ne
rect 13564 8210 14275 8250
rect -2525 8112 -284 8210
tri -284 8112 -186 8210 sw
tri -186 8112 -88 8210 ne
rect -88 8112 266 8210
tri 266 8112 364 8210 sw
tri 364 8112 462 8210 ne
rect 462 8112 816 8210
tri 816 8112 914 8210 sw
tri 914 8112 1012 8210 ne
rect 1012 8112 1366 8210
tri 1366 8112 1464 8210 sw
tri 1464 8112 1562 8210 ne
rect 1562 8112 1916 8210
tri 1916 8112 2014 8210 sw
tri 2014 8112 2112 8210 ne
rect 2112 8112 2466 8210
tri 2466 8112 2564 8210 sw
tri 2564 8112 2662 8210 ne
rect 2662 8112 3016 8210
tri 3016 8112 3114 8210 sw
tri 3114 8112 3212 8210 ne
rect 3212 8112 3566 8210
tri 3566 8112 3664 8210 sw
tri 3664 8112 3762 8210 ne
rect 3762 8112 4116 8210
tri 4116 8112 4214 8210 sw
tri 4214 8112 4312 8210 ne
rect 4312 8112 4666 8210
tri 4666 8112 4764 8210 sw
tri 4764 8112 4862 8210 ne
rect 4862 8112 5216 8210
tri 5216 8112 5314 8210 sw
tri 5314 8112 5412 8210 ne
rect 5412 8112 5766 8210
tri 5766 8112 5864 8210 sw
tri 5864 8112 5962 8210 ne
rect 5962 8112 6316 8210
tri 6316 8112 6414 8210 sw
tri 6414 8112 6512 8210 ne
rect 6512 8112 6866 8210
tri 6866 8112 6964 8210 sw
tri 6964 8112 7062 8210 ne
rect 7062 8112 7416 8210
tri 7416 8112 7514 8210 sw
tri 7514 8112 7612 8210 ne
rect 7612 8112 7966 8210
tri 7966 8112 8064 8210 sw
tri 8064 8112 8162 8210 ne
rect 8162 8112 8516 8210
tri 8516 8112 8614 8210 sw
tri 8614 8112 8712 8210 ne
rect 8712 8112 9066 8210
tri 9066 8112 9164 8210 sw
tri 9164 8112 9262 8210 ne
rect 9262 8112 9616 8210
tri 9616 8112 9714 8210 sw
tri 9714 8112 9812 8210 ne
rect 9812 8112 10166 8210
tri 10166 8112 10264 8210 sw
tri 10264 8112 10362 8210 ne
rect 10362 8112 10716 8210
tri 10716 8112 10814 8210 sw
tri 10814 8112 10912 8210 ne
rect 10912 8112 11266 8210
tri 11266 8112 11364 8210 sw
tri 11364 8112 11462 8210 ne
rect 11462 8112 11816 8210
tri 11816 8112 11914 8210 sw
tri 11914 8112 12012 8210 ne
rect 12012 8112 12366 8210
tri 12366 8112 12464 8210 sw
tri 12464 8112 12562 8210 ne
rect 12562 8112 12916 8210
tri 12916 8112 13014 8210 sw
tri 13014 8112 13112 8210 ne
rect 13112 8112 13466 8210
tri 13466 8112 13564 8210 sw
tri 13564 8112 13662 8210 ne
rect 13662 8112 14275 8210
rect -2525 8014 -186 8112
tri -186 8014 -88 8112 sw
tri -88 8014 10 8112 ne
rect 10 8014 364 8112
tri 364 8014 462 8112 sw
tri 462 8014 560 8112 ne
rect 560 8014 914 8112
tri 914 8014 1012 8112 sw
tri 1012 8014 1110 8112 ne
rect 1110 8014 1464 8112
tri 1464 8014 1562 8112 sw
tri 1562 8014 1660 8112 ne
rect 1660 8014 2014 8112
tri 2014 8014 2112 8112 sw
tri 2112 8014 2210 8112 ne
rect 2210 8014 2564 8112
tri 2564 8014 2662 8112 sw
tri 2662 8014 2760 8112 ne
rect 2760 8014 3114 8112
tri 3114 8014 3212 8112 sw
tri 3212 8014 3310 8112 ne
rect 3310 8014 3664 8112
tri 3664 8014 3762 8112 sw
tri 3762 8014 3860 8112 ne
rect 3860 8014 4214 8112
tri 4214 8014 4312 8112 sw
tri 4312 8014 4410 8112 ne
rect 4410 8014 4764 8112
tri 4764 8014 4862 8112 sw
tri 4862 8014 4960 8112 ne
rect 4960 8014 5314 8112
tri 5314 8014 5412 8112 sw
tri 5412 8014 5510 8112 ne
rect 5510 8014 5864 8112
tri 5864 8014 5962 8112 sw
tri 5962 8014 6060 8112 ne
rect 6060 8014 6414 8112
tri 6414 8014 6512 8112 sw
tri 6512 8014 6610 8112 ne
rect 6610 8014 6964 8112
tri 6964 8014 7062 8112 sw
tri 7062 8014 7160 8112 ne
rect 7160 8014 7514 8112
tri 7514 8014 7612 8112 sw
tri 7612 8014 7710 8112 ne
rect 7710 8014 8064 8112
tri 8064 8014 8162 8112 sw
tri 8162 8014 8260 8112 ne
rect 8260 8014 8614 8112
tri 8614 8014 8712 8112 sw
tri 8712 8014 8810 8112 ne
rect 8810 8014 9164 8112
tri 9164 8014 9262 8112 sw
tri 9262 8014 9360 8112 ne
rect 9360 8014 9714 8112
tri 9714 8014 9812 8112 sw
tri 9812 8014 9910 8112 ne
rect 9910 8014 10264 8112
tri 10264 8014 10362 8112 sw
tri 10362 8014 10460 8112 ne
rect 10460 8014 10814 8112
tri 10814 8014 10912 8112 sw
tri 10912 8014 11010 8112 ne
rect 11010 8014 11364 8112
tri 11364 8014 11462 8112 sw
tri 11462 8014 11560 8112 ne
rect 11560 8014 11914 8112
tri 11914 8014 12012 8112 sw
tri 12012 8014 12110 8112 ne
rect 12110 8014 12464 8112
tri 12464 8014 12562 8112 sw
tri 12562 8014 12660 8112 ne
rect 12660 8014 13014 8112
tri 13014 8014 13112 8112 sw
tri 13112 8014 13210 8112 ne
rect 13210 8014 13564 8112
tri 13564 8014 13662 8112 sw
rect 14775 8014 15775 8662
rect -2525 8010 -88 8014
rect -2525 7890 -310 8010
rect -190 7926 -88 8010
tri -88 7926 0 8014 sw
tri 10 7926 98 8014 ne
rect 98 8010 462 8014
rect 98 7926 240 8010
rect -190 7890 0 7926
rect -2525 7886 0 7890
rect -2525 7238 -1525 7886
tri -412 7788 -314 7886 ne
rect -314 7838 0 7886
tri 0 7838 88 7926 sw
tri 98 7838 186 7926 ne
rect 186 7890 240 7926
rect 360 7926 462 8010
tri 462 7926 550 8014 sw
tri 560 7926 648 8014 ne
rect 648 8010 1012 8014
rect 648 7926 790 8010
rect 360 7890 550 7926
rect 186 7886 550 7890
tri 550 7886 590 7926 sw
tri 648 7886 688 7926 ne
rect 688 7890 790 7926
rect 910 7926 1012 8010
tri 1012 7926 1100 8014 sw
tri 1110 7926 1198 8014 ne
rect 1198 8010 1562 8014
rect 1198 7926 1340 8010
rect 910 7890 1100 7926
rect 688 7886 1100 7890
rect 186 7838 590 7886
rect -314 7788 88 7838
rect -1025 7700 -412 7788
tri -412 7700 -324 7788 sw
tri -314 7700 -226 7788 ne
rect -226 7758 88 7788
tri 88 7758 168 7838 sw
tri 186 7758 266 7838 ne
rect 266 7788 590 7838
tri 590 7788 688 7886 sw
tri 688 7788 786 7886 ne
rect 786 7838 1100 7886
tri 1100 7838 1188 7926 sw
tri 1198 7838 1286 7926 ne
rect 1286 7890 1340 7926
rect 1460 7926 1562 8010
tri 1562 7926 1650 8014 sw
tri 1660 7926 1748 8014 ne
rect 1748 8010 2112 8014
rect 1748 7926 1890 8010
rect 1460 7890 1650 7926
rect 1286 7886 1650 7890
tri 1650 7886 1690 7926 sw
tri 1748 7886 1788 7926 ne
rect 1788 7890 1890 7926
rect 2010 7926 2112 8010
tri 2112 7926 2200 8014 sw
tri 2210 7926 2298 8014 ne
rect 2298 8010 2662 8014
rect 2298 7926 2440 8010
rect 2010 7890 2200 7926
rect 1788 7886 2200 7890
rect 1286 7838 1690 7886
rect 786 7788 1188 7838
rect 266 7758 688 7788
rect -226 7700 168 7758
rect -1025 7660 -324 7700
tri -324 7660 -284 7700 sw
tri -226 7660 -186 7700 ne
rect -186 7660 168 7700
tri 168 7660 266 7758 sw
tri 266 7660 364 7758 ne
rect 364 7700 688 7758
tri 688 7700 776 7788 sw
tri 786 7700 874 7788 ne
rect 874 7758 1188 7788
tri 1188 7758 1268 7838 sw
tri 1286 7758 1366 7838 ne
rect 1366 7788 1690 7838
tri 1690 7788 1788 7886 sw
tri 1788 7788 1886 7886 ne
rect 1886 7838 2200 7886
tri 2200 7838 2288 7926 sw
tri 2298 7838 2386 7926 ne
rect 2386 7890 2440 7926
rect 2560 7926 2662 8010
tri 2662 7926 2750 8014 sw
tri 2760 7926 2848 8014 ne
rect 2848 8010 3212 8014
rect 2848 7926 2990 8010
rect 2560 7890 2750 7926
rect 2386 7886 2750 7890
tri 2750 7886 2790 7926 sw
tri 2848 7886 2888 7926 ne
rect 2888 7890 2990 7926
rect 3110 7926 3212 8010
tri 3212 7926 3300 8014 sw
tri 3310 7926 3398 8014 ne
rect 3398 8010 3762 8014
rect 3398 7926 3540 8010
rect 3110 7890 3300 7926
rect 2888 7886 3300 7890
rect 2386 7838 2790 7886
rect 1886 7788 2288 7838
rect 1366 7758 1788 7788
rect 874 7700 1268 7758
rect 364 7660 776 7700
tri 776 7660 816 7700 sw
tri 874 7660 914 7700 ne
rect 914 7660 1268 7700
tri 1268 7660 1366 7758 sw
tri 1366 7660 1464 7758 ne
rect 1464 7700 1788 7758
tri 1788 7700 1876 7788 sw
tri 1886 7700 1974 7788 ne
rect 1974 7758 2288 7788
tri 2288 7758 2368 7838 sw
tri 2386 7758 2466 7838 ne
rect 2466 7788 2790 7838
tri 2790 7788 2888 7886 sw
tri 2888 7788 2986 7886 ne
rect 2986 7838 3300 7886
tri 3300 7838 3388 7926 sw
tri 3398 7838 3486 7926 ne
rect 3486 7890 3540 7926
rect 3660 7926 3762 8010
tri 3762 7926 3850 8014 sw
tri 3860 7926 3948 8014 ne
rect 3948 8010 4312 8014
rect 3948 7926 4090 8010
rect 3660 7890 3850 7926
rect 3486 7886 3850 7890
tri 3850 7886 3890 7926 sw
tri 3948 7886 3988 7926 ne
rect 3988 7890 4090 7926
rect 4210 7926 4312 8010
tri 4312 7926 4400 8014 sw
tri 4410 7926 4498 8014 ne
rect 4498 8010 4862 8014
rect 4498 7926 4640 8010
rect 4210 7890 4400 7926
rect 3988 7886 4400 7890
rect 3486 7838 3890 7886
rect 2986 7788 3388 7838
rect 2466 7758 2888 7788
rect 1974 7700 2368 7758
rect 1464 7660 1876 7700
tri 1876 7660 1916 7700 sw
tri 1974 7660 2014 7700 ne
rect 2014 7660 2368 7700
tri 2368 7660 2466 7758 sw
tri 2466 7660 2564 7758 ne
rect 2564 7700 2888 7758
tri 2888 7700 2976 7788 sw
tri 2986 7700 3074 7788 ne
rect 3074 7758 3388 7788
tri 3388 7758 3468 7838 sw
tri 3486 7758 3566 7838 ne
rect 3566 7788 3890 7838
tri 3890 7788 3988 7886 sw
tri 3988 7788 4086 7886 ne
rect 4086 7838 4400 7886
tri 4400 7838 4488 7926 sw
tri 4498 7838 4586 7926 ne
rect 4586 7890 4640 7926
rect 4760 7926 4862 8010
tri 4862 7926 4950 8014 sw
tri 4960 7926 5048 8014 ne
rect 5048 8010 5412 8014
rect 5048 7926 5190 8010
rect 4760 7890 4950 7926
rect 4586 7886 4950 7890
tri 4950 7886 4990 7926 sw
tri 5048 7886 5088 7926 ne
rect 5088 7890 5190 7926
rect 5310 7926 5412 8010
tri 5412 7926 5500 8014 sw
tri 5510 7926 5598 8014 ne
rect 5598 8010 5962 8014
rect 5598 7926 5740 8010
rect 5310 7890 5500 7926
rect 5088 7886 5500 7890
rect 4586 7838 4990 7886
rect 4086 7788 4488 7838
rect 3566 7758 3988 7788
rect 3074 7700 3468 7758
rect 2564 7660 2976 7700
tri 2976 7660 3016 7700 sw
tri 3074 7660 3114 7700 ne
rect 3114 7660 3468 7700
tri 3468 7660 3566 7758 sw
tri 3566 7660 3664 7758 ne
rect 3664 7700 3988 7758
tri 3988 7700 4076 7788 sw
tri 4086 7700 4174 7788 ne
rect 4174 7758 4488 7788
tri 4488 7758 4568 7838 sw
tri 4586 7758 4666 7838 ne
rect 4666 7788 4990 7838
tri 4990 7788 5088 7886 sw
tri 5088 7788 5186 7886 ne
rect 5186 7838 5500 7886
tri 5500 7838 5588 7926 sw
tri 5598 7838 5686 7926 ne
rect 5686 7890 5740 7926
rect 5860 7926 5962 8010
tri 5962 7926 6050 8014 sw
tri 6060 7926 6148 8014 ne
rect 6148 8010 6512 8014
rect 6148 7926 6290 8010
rect 5860 7890 6050 7926
rect 5686 7886 6050 7890
tri 6050 7886 6090 7926 sw
tri 6148 7886 6188 7926 ne
rect 6188 7890 6290 7926
rect 6410 7926 6512 8010
tri 6512 7926 6600 8014 sw
tri 6610 7926 6698 8014 ne
rect 6698 8010 7062 8014
rect 6698 7926 6840 8010
rect 6410 7890 6600 7926
rect 6188 7886 6600 7890
rect 5686 7838 6090 7886
rect 5186 7788 5588 7838
rect 4666 7758 5088 7788
rect 4174 7700 4568 7758
rect 3664 7660 4076 7700
tri 4076 7660 4116 7700 sw
tri 4174 7660 4214 7700 ne
rect 4214 7660 4568 7700
tri 4568 7660 4666 7758 sw
tri 4666 7660 4764 7758 ne
rect 4764 7700 5088 7758
tri 5088 7700 5176 7788 sw
tri 5186 7700 5274 7788 ne
rect 5274 7758 5588 7788
tri 5588 7758 5668 7838 sw
tri 5686 7758 5766 7838 ne
rect 5766 7788 6090 7838
tri 6090 7788 6188 7886 sw
tri 6188 7788 6286 7886 ne
rect 6286 7838 6600 7886
tri 6600 7838 6688 7926 sw
tri 6698 7838 6786 7926 ne
rect 6786 7890 6840 7926
rect 6960 7926 7062 8010
tri 7062 7926 7150 8014 sw
tri 7160 7926 7248 8014 ne
rect 7248 8010 7612 8014
rect 7248 7926 7390 8010
rect 6960 7890 7150 7926
rect 6786 7886 7150 7890
tri 7150 7886 7190 7926 sw
tri 7248 7886 7288 7926 ne
rect 7288 7890 7390 7926
rect 7510 7926 7612 8010
tri 7612 7926 7700 8014 sw
tri 7710 7926 7798 8014 ne
rect 7798 8010 8162 8014
rect 7798 7926 7940 8010
rect 7510 7890 7700 7926
rect 7288 7886 7700 7890
rect 6786 7838 7190 7886
rect 6286 7788 6688 7838
rect 5766 7758 6188 7788
rect 5274 7700 5668 7758
rect 4764 7660 5176 7700
tri 5176 7660 5216 7700 sw
tri 5274 7660 5314 7700 ne
rect 5314 7660 5668 7700
tri 5668 7660 5766 7758 sw
tri 5766 7660 5864 7758 ne
rect 5864 7700 6188 7758
tri 6188 7700 6276 7788 sw
tri 6286 7700 6374 7788 ne
rect 6374 7758 6688 7788
tri 6688 7758 6768 7838 sw
tri 6786 7758 6866 7838 ne
rect 6866 7788 7190 7838
tri 7190 7788 7288 7886 sw
tri 7288 7788 7386 7886 ne
rect 7386 7838 7700 7886
tri 7700 7838 7788 7926 sw
tri 7798 7838 7886 7926 ne
rect 7886 7890 7940 7926
rect 8060 7926 8162 8010
tri 8162 7926 8250 8014 sw
tri 8260 7926 8348 8014 ne
rect 8348 8010 8712 8014
rect 8348 7926 8490 8010
rect 8060 7890 8250 7926
rect 7886 7886 8250 7890
tri 8250 7886 8290 7926 sw
tri 8348 7886 8388 7926 ne
rect 8388 7890 8490 7926
rect 8610 7926 8712 8010
tri 8712 7926 8800 8014 sw
tri 8810 7926 8898 8014 ne
rect 8898 8010 9262 8014
rect 8898 7926 9040 8010
rect 8610 7890 8800 7926
rect 8388 7886 8800 7890
rect 7886 7838 8290 7886
rect 7386 7788 7788 7838
rect 6866 7758 7288 7788
rect 6374 7700 6768 7758
rect 5864 7660 6276 7700
tri 6276 7660 6316 7700 sw
tri 6374 7660 6414 7700 ne
rect 6414 7660 6768 7700
tri 6768 7660 6866 7758 sw
tri 6866 7660 6964 7758 ne
rect 6964 7700 7288 7758
tri 7288 7700 7376 7788 sw
tri 7386 7700 7474 7788 ne
rect 7474 7758 7788 7788
tri 7788 7758 7868 7838 sw
tri 7886 7758 7966 7838 ne
rect 7966 7788 8290 7838
tri 8290 7788 8388 7886 sw
tri 8388 7788 8486 7886 ne
rect 8486 7838 8800 7886
tri 8800 7838 8888 7926 sw
tri 8898 7838 8986 7926 ne
rect 8986 7890 9040 7926
rect 9160 7926 9262 8010
tri 9262 7926 9350 8014 sw
tri 9360 7926 9448 8014 ne
rect 9448 8010 9812 8014
rect 9448 7926 9590 8010
rect 9160 7890 9350 7926
rect 8986 7886 9350 7890
tri 9350 7886 9390 7926 sw
tri 9448 7886 9488 7926 ne
rect 9488 7890 9590 7926
rect 9710 7926 9812 8010
tri 9812 7926 9900 8014 sw
tri 9910 7926 9998 8014 ne
rect 9998 8010 10362 8014
rect 9998 7926 10140 8010
rect 9710 7890 9900 7926
rect 9488 7886 9900 7890
rect 8986 7838 9390 7886
rect 8486 7788 8888 7838
rect 7966 7758 8388 7788
rect 7474 7700 7868 7758
rect 6964 7660 7376 7700
tri 7376 7660 7416 7700 sw
tri 7474 7660 7514 7700 ne
rect 7514 7660 7868 7700
tri 7868 7660 7966 7758 sw
tri 7966 7660 8064 7758 ne
rect 8064 7700 8388 7758
tri 8388 7700 8476 7788 sw
tri 8486 7700 8574 7788 ne
rect 8574 7758 8888 7788
tri 8888 7758 8968 7838 sw
tri 8986 7758 9066 7838 ne
rect 9066 7788 9390 7838
tri 9390 7788 9488 7886 sw
tri 9488 7788 9586 7886 ne
rect 9586 7838 9900 7886
tri 9900 7838 9988 7926 sw
tri 9998 7838 10086 7926 ne
rect 10086 7890 10140 7926
rect 10260 7926 10362 8010
tri 10362 7926 10450 8014 sw
tri 10460 7926 10548 8014 ne
rect 10548 8010 10912 8014
rect 10548 7926 10690 8010
rect 10260 7890 10450 7926
rect 10086 7886 10450 7890
tri 10450 7886 10490 7926 sw
tri 10548 7886 10588 7926 ne
rect 10588 7890 10690 7926
rect 10810 7926 10912 8010
tri 10912 7926 11000 8014 sw
tri 11010 7926 11098 8014 ne
rect 11098 8010 11462 8014
rect 11098 7926 11240 8010
rect 10810 7890 11000 7926
rect 10588 7886 11000 7890
rect 10086 7838 10490 7886
rect 9586 7788 9988 7838
rect 9066 7758 9488 7788
rect 8574 7700 8968 7758
rect 8064 7660 8476 7700
tri 8476 7660 8516 7700 sw
tri 8574 7660 8614 7700 ne
rect 8614 7660 8968 7700
tri 8968 7660 9066 7758 sw
tri 9066 7660 9164 7758 ne
rect 9164 7700 9488 7758
tri 9488 7700 9576 7788 sw
tri 9586 7700 9674 7788 ne
rect 9674 7758 9988 7788
tri 9988 7758 10068 7838 sw
tri 10086 7758 10166 7838 ne
rect 10166 7788 10490 7838
tri 10490 7788 10588 7886 sw
tri 10588 7788 10686 7886 ne
rect 10686 7838 11000 7886
tri 11000 7838 11088 7926 sw
tri 11098 7838 11186 7926 ne
rect 11186 7890 11240 7926
rect 11360 7926 11462 8010
tri 11462 7926 11550 8014 sw
tri 11560 7926 11648 8014 ne
rect 11648 8010 12012 8014
rect 11648 7926 11790 8010
rect 11360 7890 11550 7926
rect 11186 7886 11550 7890
tri 11550 7886 11590 7926 sw
tri 11648 7886 11688 7926 ne
rect 11688 7890 11790 7926
rect 11910 7926 12012 8010
tri 12012 7926 12100 8014 sw
tri 12110 7926 12198 8014 ne
rect 12198 8010 12562 8014
rect 12198 7926 12340 8010
rect 11910 7890 12100 7926
rect 11688 7886 12100 7890
rect 11186 7838 11590 7886
rect 10686 7788 11088 7838
rect 10166 7758 10588 7788
rect 9674 7700 10068 7758
rect 9164 7660 9576 7700
tri 9576 7660 9616 7700 sw
tri 9674 7660 9714 7700 ne
rect 9714 7660 10068 7700
tri 10068 7660 10166 7758 sw
tri 10166 7660 10264 7758 ne
rect 10264 7700 10588 7758
tri 10588 7700 10676 7788 sw
tri 10686 7700 10774 7788 ne
rect 10774 7758 11088 7788
tri 11088 7758 11168 7838 sw
tri 11186 7758 11266 7838 ne
rect 11266 7788 11590 7838
tri 11590 7788 11688 7886 sw
tri 11688 7788 11786 7886 ne
rect 11786 7838 12100 7886
tri 12100 7838 12188 7926 sw
tri 12198 7838 12286 7926 ne
rect 12286 7890 12340 7926
rect 12460 7926 12562 8010
tri 12562 7926 12650 8014 sw
tri 12660 7926 12748 8014 ne
rect 12748 8010 13112 8014
rect 12748 7926 12890 8010
rect 12460 7890 12650 7926
rect 12286 7886 12650 7890
tri 12650 7886 12690 7926 sw
tri 12748 7886 12788 7926 ne
rect 12788 7890 12890 7926
rect 13010 7926 13112 8010
tri 13112 7926 13200 8014 sw
tri 13210 7926 13298 8014 ne
rect 13298 8010 15775 8014
rect 13298 7926 13440 8010
rect 13010 7890 13200 7926
rect 12788 7886 13200 7890
rect 12286 7838 12690 7886
rect 11786 7788 12188 7838
rect 11266 7758 11688 7788
rect 10774 7700 11168 7758
rect 10264 7660 10676 7700
tri 10676 7660 10716 7700 sw
tri 10774 7660 10814 7700 ne
rect 10814 7660 11168 7700
tri 11168 7660 11266 7758 sw
tri 11266 7660 11364 7758 ne
rect 11364 7700 11688 7758
tri 11688 7700 11776 7788 sw
tri 11786 7700 11874 7788 ne
rect 11874 7758 12188 7788
tri 12188 7758 12268 7838 sw
tri 12286 7758 12366 7838 ne
rect 12366 7788 12690 7838
tri 12690 7788 12788 7886 sw
tri 12788 7788 12886 7886 ne
rect 12886 7838 13200 7886
tri 13200 7838 13288 7926 sw
tri 13298 7838 13386 7926 ne
rect 13386 7890 13440 7926
rect 13560 7890 15775 8010
rect 13386 7838 15775 7890
rect 12886 7788 13288 7838
rect 12366 7758 12788 7788
rect 11874 7700 12268 7758
rect 11364 7660 11776 7700
tri 11776 7660 11816 7700 sw
tri 11874 7660 11914 7700 ne
rect 11914 7660 12268 7700
tri 12268 7660 12366 7758 sw
tri 12366 7660 12464 7758 ne
rect 12464 7700 12788 7758
tri 12788 7700 12876 7788 sw
tri 12886 7700 12974 7788 ne
rect 12974 7758 13288 7788
tri 13288 7758 13368 7838 sw
tri 13386 7758 13466 7838 ne
rect 13466 7758 14075 7838
rect 12974 7700 13368 7758
rect 12464 7660 12876 7700
tri 12876 7660 12916 7700 sw
tri 12974 7660 13014 7700 ne
rect 13014 7660 13368 7700
tri 13368 7660 13466 7758 sw
tri 13466 7660 13564 7758 ne
rect 13564 7738 14075 7758
rect 14175 7738 15775 7838
rect 13564 7660 15775 7738
rect -1025 7612 -284 7660
rect -1025 7512 -925 7612
rect -825 7562 -284 7612
tri -284 7562 -186 7660 sw
tri -186 7562 -88 7660 ne
rect -88 7562 266 7660
tri 266 7562 364 7660 sw
tri 364 7562 462 7660 ne
rect 462 7562 816 7660
tri 816 7562 914 7660 sw
tri 914 7562 1012 7660 ne
rect 1012 7562 1366 7660
tri 1366 7562 1464 7660 sw
tri 1464 7562 1562 7660 ne
rect 1562 7562 1916 7660
tri 1916 7562 2014 7660 sw
tri 2014 7562 2112 7660 ne
rect 2112 7562 2466 7660
tri 2466 7562 2564 7660 sw
tri 2564 7562 2662 7660 ne
rect 2662 7562 3016 7660
tri 3016 7562 3114 7660 sw
tri 3114 7562 3212 7660 ne
rect 3212 7562 3566 7660
tri 3566 7562 3664 7660 sw
tri 3664 7562 3762 7660 ne
rect 3762 7562 4116 7660
tri 4116 7562 4214 7660 sw
tri 4214 7562 4312 7660 ne
rect 4312 7562 4666 7660
tri 4666 7562 4764 7660 sw
tri 4764 7562 4862 7660 ne
rect 4862 7562 5216 7660
tri 5216 7562 5314 7660 sw
tri 5314 7562 5412 7660 ne
rect 5412 7562 5766 7660
tri 5766 7562 5864 7660 sw
tri 5864 7562 5962 7660 ne
rect 5962 7562 6316 7660
tri 6316 7562 6414 7660 sw
tri 6414 7562 6512 7660 ne
rect 6512 7562 6866 7660
tri 6866 7562 6964 7660 sw
tri 6964 7562 7062 7660 ne
rect 7062 7562 7416 7660
tri 7416 7562 7514 7660 sw
tri 7514 7562 7612 7660 ne
rect 7612 7562 7966 7660
tri 7966 7562 8064 7660 sw
tri 8064 7562 8162 7660 ne
rect 8162 7562 8516 7660
tri 8516 7562 8614 7660 sw
tri 8614 7562 8712 7660 ne
rect 8712 7562 9066 7660
tri 9066 7562 9164 7660 sw
tri 9164 7562 9262 7660 ne
rect 9262 7562 9616 7660
tri 9616 7562 9714 7660 sw
tri 9714 7562 9812 7660 ne
rect 9812 7562 10166 7660
tri 10166 7562 10264 7660 sw
tri 10264 7562 10362 7660 ne
rect 10362 7562 10716 7660
tri 10716 7562 10814 7660 sw
tri 10814 7562 10912 7660 ne
rect 10912 7562 11266 7660
tri 11266 7562 11364 7660 sw
tri 11364 7562 11462 7660 ne
rect 11462 7562 11816 7660
tri 11816 7562 11914 7660 sw
tri 11914 7562 12012 7660 ne
rect 12012 7562 12366 7660
tri 12366 7562 12464 7660 sw
tri 12464 7562 12562 7660 ne
rect 12562 7562 12916 7660
tri 12916 7562 13014 7660 sw
tri 13014 7562 13112 7660 ne
rect 13112 7562 13466 7660
tri 13466 7562 13564 7660 sw
tri 13564 7562 13662 7660 ne
rect 13662 7562 15775 7660
rect -825 7512 -186 7562
rect -1025 7464 -186 7512
tri -186 7464 -88 7562 sw
tri -88 7464 10 7562 ne
rect 10 7464 364 7562
tri 364 7464 462 7562 sw
tri 462 7464 560 7562 ne
rect 560 7464 914 7562
tri 914 7464 1012 7562 sw
tri 1012 7464 1110 7562 ne
rect 1110 7464 1464 7562
tri 1464 7464 1562 7562 sw
tri 1562 7464 1660 7562 ne
rect 1660 7464 2014 7562
tri 2014 7464 2112 7562 sw
tri 2112 7464 2210 7562 ne
rect 2210 7464 2564 7562
tri 2564 7464 2662 7562 sw
tri 2662 7464 2760 7562 ne
rect 2760 7464 3114 7562
tri 3114 7464 3212 7562 sw
tri 3212 7464 3310 7562 ne
rect 3310 7464 3664 7562
tri 3664 7464 3762 7562 sw
tri 3762 7464 3860 7562 ne
rect 3860 7464 4214 7562
tri 4214 7464 4312 7562 sw
tri 4312 7464 4410 7562 ne
rect 4410 7464 4764 7562
tri 4764 7464 4862 7562 sw
tri 4862 7464 4960 7562 ne
rect 4960 7464 5314 7562
tri 5314 7464 5412 7562 sw
tri 5412 7464 5510 7562 ne
rect 5510 7464 5864 7562
tri 5864 7464 5962 7562 sw
tri 5962 7464 6060 7562 ne
rect 6060 7464 6414 7562
tri 6414 7464 6512 7562 sw
tri 6512 7464 6610 7562 ne
rect 6610 7464 6964 7562
tri 6964 7464 7062 7562 sw
tri 7062 7464 7160 7562 ne
rect 7160 7464 7514 7562
tri 7514 7464 7612 7562 sw
tri 7612 7464 7710 7562 ne
rect 7710 7464 8064 7562
tri 8064 7464 8162 7562 sw
tri 8162 7464 8260 7562 ne
rect 8260 7464 8614 7562
tri 8614 7464 8712 7562 sw
tri 8712 7464 8810 7562 ne
rect 8810 7464 9164 7562
tri 9164 7464 9262 7562 sw
tri 9262 7464 9360 7562 ne
rect 9360 7464 9714 7562
tri 9714 7464 9812 7562 sw
tri 9812 7464 9910 7562 ne
rect 9910 7464 10264 7562
tri 10264 7464 10362 7562 sw
tri 10362 7464 10460 7562 ne
rect 10460 7464 10814 7562
tri 10814 7464 10912 7562 sw
tri 10912 7464 11010 7562 ne
rect 11010 7464 11364 7562
tri 11364 7464 11462 7562 sw
tri 11462 7464 11560 7562 ne
rect 11560 7464 11914 7562
tri 11914 7464 12012 7562 sw
tri 12012 7464 12110 7562 ne
rect 12110 7464 12464 7562
tri 12464 7464 12562 7562 sw
tri 12562 7464 12660 7562 ne
rect 12660 7464 13014 7562
tri 13014 7464 13112 7562 sw
tri 13112 7464 13210 7562 ne
rect 13210 7464 13564 7562
tri 13564 7464 13662 7562 sw
rect -1025 7460 -88 7464
rect -1025 7340 -310 7460
rect -190 7376 -88 7460
tri -88 7376 0 7464 sw
tri 10 7376 98 7464 ne
rect 98 7460 462 7464
rect 98 7376 240 7460
rect -190 7340 0 7376
rect -1025 7336 0 7340
tri 0 7336 40 7376 sw
tri 98 7336 138 7376 ne
rect 138 7340 240 7376
rect 360 7376 462 7460
tri 462 7376 550 7464 sw
tri 560 7376 648 7464 ne
rect 648 7460 1012 7464
rect 648 7376 790 7460
rect 360 7340 550 7376
rect 138 7336 550 7340
tri -412 7238 -314 7336 ne
rect -314 7238 40 7336
tri 40 7238 138 7336 sw
tri 138 7238 236 7336 ne
rect 236 7288 550 7336
tri 550 7288 638 7376 sw
tri 648 7288 736 7376 ne
rect 736 7340 790 7376
rect 910 7376 1012 7460
tri 1012 7376 1100 7464 sw
tri 1110 7376 1198 7464 ne
rect 1198 7460 1562 7464
rect 1198 7376 1340 7460
rect 910 7340 1100 7376
rect 736 7336 1100 7340
tri 1100 7336 1140 7376 sw
tri 1198 7336 1238 7376 ne
rect 1238 7340 1340 7376
rect 1460 7376 1562 7460
tri 1562 7376 1650 7464 sw
tri 1660 7376 1748 7464 ne
rect 1748 7460 2112 7464
rect 1748 7376 1890 7460
rect 1460 7340 1650 7376
rect 1238 7336 1650 7340
rect 736 7288 1140 7336
rect 236 7238 638 7288
rect -2525 7150 -412 7238
tri -412 7150 -324 7238 sw
tri -314 7150 -226 7238 ne
rect -226 7150 138 7238
tri 138 7150 226 7238 sw
tri 236 7150 324 7238 ne
rect 324 7208 638 7238
tri 638 7208 718 7288 sw
tri 736 7208 816 7288 ne
rect 816 7238 1140 7288
tri 1140 7238 1238 7336 sw
tri 1238 7238 1336 7336 ne
rect 1336 7288 1650 7336
tri 1650 7288 1738 7376 sw
tri 1748 7288 1836 7376 ne
rect 1836 7340 1890 7376
rect 2010 7376 2112 7460
tri 2112 7376 2200 7464 sw
tri 2210 7376 2298 7464 ne
rect 2298 7460 2662 7464
rect 2298 7376 2440 7460
rect 2010 7340 2200 7376
rect 1836 7336 2200 7340
tri 2200 7336 2240 7376 sw
tri 2298 7336 2338 7376 ne
rect 2338 7340 2440 7376
rect 2560 7376 2662 7460
tri 2662 7376 2750 7464 sw
tri 2760 7376 2848 7464 ne
rect 2848 7460 3212 7464
rect 2848 7376 2990 7460
rect 2560 7340 2750 7376
rect 2338 7336 2750 7340
rect 1836 7288 2240 7336
rect 1336 7238 1738 7288
rect 816 7208 1238 7238
rect 324 7150 718 7208
rect -2525 7110 -324 7150
tri -324 7110 -284 7150 sw
tri -226 7110 -186 7150 ne
rect -186 7110 226 7150
tri 226 7110 266 7150 sw
tri 324 7110 364 7150 ne
rect 364 7110 718 7150
tri 718 7110 816 7208 sw
tri 816 7110 914 7208 ne
rect 914 7150 1238 7208
tri 1238 7150 1326 7238 sw
tri 1336 7150 1424 7238 ne
rect 1424 7208 1738 7238
tri 1738 7208 1818 7288 sw
tri 1836 7208 1916 7288 ne
rect 1916 7238 2240 7288
tri 2240 7238 2338 7336 sw
tri 2338 7238 2436 7336 ne
rect 2436 7288 2750 7336
tri 2750 7288 2838 7376 sw
tri 2848 7288 2936 7376 ne
rect 2936 7340 2990 7376
rect 3110 7376 3212 7460
tri 3212 7376 3300 7464 sw
tri 3310 7376 3398 7464 ne
rect 3398 7460 3762 7464
rect 3398 7376 3540 7460
rect 3110 7340 3300 7376
rect 2936 7336 3300 7340
tri 3300 7336 3340 7376 sw
tri 3398 7336 3438 7376 ne
rect 3438 7340 3540 7376
rect 3660 7376 3762 7460
tri 3762 7376 3850 7464 sw
tri 3860 7376 3948 7464 ne
rect 3948 7460 4312 7464
rect 3948 7376 4090 7460
rect 3660 7340 3850 7376
rect 3438 7336 3850 7340
rect 2936 7288 3340 7336
rect 2436 7238 2838 7288
rect 1916 7208 2338 7238
rect 1424 7150 1818 7208
rect 914 7110 1326 7150
tri 1326 7110 1366 7150 sw
tri 1424 7110 1464 7150 ne
rect 1464 7110 1818 7150
tri 1818 7110 1916 7208 sw
tri 1916 7110 2014 7208 ne
rect 2014 7150 2338 7208
tri 2338 7150 2426 7238 sw
tri 2436 7150 2524 7238 ne
rect 2524 7208 2838 7238
tri 2838 7208 2918 7288 sw
tri 2936 7208 3016 7288 ne
rect 3016 7238 3340 7288
tri 3340 7238 3438 7336 sw
tri 3438 7238 3536 7336 ne
rect 3536 7288 3850 7336
tri 3850 7288 3938 7376 sw
tri 3948 7288 4036 7376 ne
rect 4036 7340 4090 7376
rect 4210 7376 4312 7460
tri 4312 7376 4400 7464 sw
tri 4410 7376 4498 7464 ne
rect 4498 7460 4862 7464
rect 4498 7376 4640 7460
rect 4210 7340 4400 7376
rect 4036 7336 4400 7340
tri 4400 7336 4440 7376 sw
tri 4498 7336 4538 7376 ne
rect 4538 7340 4640 7376
rect 4760 7376 4862 7460
tri 4862 7376 4950 7464 sw
tri 4960 7376 5048 7464 ne
rect 5048 7460 5412 7464
rect 5048 7376 5190 7460
rect 4760 7340 4950 7376
rect 4538 7336 4950 7340
rect 4036 7288 4440 7336
rect 3536 7238 3938 7288
rect 3016 7208 3438 7238
rect 2524 7150 2918 7208
rect 2014 7110 2426 7150
tri 2426 7110 2466 7150 sw
tri 2524 7110 2564 7150 ne
rect 2564 7110 2918 7150
tri 2918 7110 3016 7208 sw
tri 3016 7110 3114 7208 ne
rect 3114 7150 3438 7208
tri 3438 7150 3526 7238 sw
tri 3536 7150 3624 7238 ne
rect 3624 7208 3938 7238
tri 3938 7208 4018 7288 sw
tri 4036 7208 4116 7288 ne
rect 4116 7238 4440 7288
tri 4440 7238 4538 7336 sw
tri 4538 7238 4636 7336 ne
rect 4636 7288 4950 7336
tri 4950 7288 5038 7376 sw
tri 5048 7288 5136 7376 ne
rect 5136 7340 5190 7376
rect 5310 7376 5412 7460
tri 5412 7376 5500 7464 sw
tri 5510 7376 5598 7464 ne
rect 5598 7460 5962 7464
rect 5598 7376 5740 7460
rect 5310 7340 5500 7376
rect 5136 7336 5500 7340
tri 5500 7336 5540 7376 sw
tri 5598 7336 5638 7376 ne
rect 5638 7340 5740 7376
rect 5860 7376 5962 7460
tri 5962 7376 6050 7464 sw
tri 6060 7376 6148 7464 ne
rect 6148 7460 6512 7464
rect 6148 7376 6290 7460
rect 5860 7340 6050 7376
rect 5638 7336 6050 7340
rect 5136 7288 5540 7336
rect 4636 7238 5038 7288
rect 4116 7208 4538 7238
rect 3624 7150 4018 7208
rect 3114 7110 3526 7150
tri 3526 7110 3566 7150 sw
tri 3624 7110 3664 7150 ne
rect 3664 7110 4018 7150
tri 4018 7110 4116 7208 sw
tri 4116 7110 4214 7208 ne
rect 4214 7150 4538 7208
tri 4538 7150 4626 7238 sw
tri 4636 7150 4724 7238 ne
rect 4724 7208 5038 7238
tri 5038 7208 5118 7288 sw
tri 5136 7208 5216 7288 ne
rect 5216 7238 5540 7288
tri 5540 7238 5638 7336 sw
tri 5638 7238 5736 7336 ne
rect 5736 7288 6050 7336
tri 6050 7288 6138 7376 sw
tri 6148 7288 6236 7376 ne
rect 6236 7340 6290 7376
rect 6410 7376 6512 7460
tri 6512 7376 6600 7464 sw
tri 6610 7376 6698 7464 ne
rect 6698 7460 7062 7464
rect 6698 7376 6840 7460
rect 6410 7340 6600 7376
rect 6236 7336 6600 7340
tri 6600 7336 6640 7376 sw
tri 6698 7336 6738 7376 ne
rect 6738 7340 6840 7376
rect 6960 7376 7062 7460
tri 7062 7376 7150 7464 sw
tri 7160 7376 7248 7464 ne
rect 7248 7460 7612 7464
rect 7248 7376 7390 7460
rect 6960 7340 7150 7376
rect 6738 7336 7150 7340
rect 6236 7288 6640 7336
rect 5736 7238 6138 7288
rect 5216 7208 5638 7238
rect 4724 7150 5118 7208
rect 4214 7110 4626 7150
tri 4626 7110 4666 7150 sw
tri 4724 7110 4764 7150 ne
rect 4764 7110 5118 7150
tri 5118 7110 5216 7208 sw
tri 5216 7110 5314 7208 ne
rect 5314 7150 5638 7208
tri 5638 7150 5726 7238 sw
tri 5736 7150 5824 7238 ne
rect 5824 7208 6138 7238
tri 6138 7208 6218 7288 sw
tri 6236 7208 6316 7288 ne
rect 6316 7238 6640 7288
tri 6640 7238 6738 7336 sw
tri 6738 7238 6836 7336 ne
rect 6836 7288 7150 7336
tri 7150 7288 7238 7376 sw
tri 7248 7288 7336 7376 ne
rect 7336 7340 7390 7376
rect 7510 7376 7612 7460
tri 7612 7376 7700 7464 sw
tri 7710 7376 7798 7464 ne
rect 7798 7460 8162 7464
rect 7798 7376 7940 7460
rect 7510 7340 7700 7376
rect 7336 7336 7700 7340
tri 7700 7336 7740 7376 sw
tri 7798 7336 7838 7376 ne
rect 7838 7340 7940 7376
rect 8060 7376 8162 7460
tri 8162 7376 8250 7464 sw
tri 8260 7376 8348 7464 ne
rect 8348 7460 8712 7464
rect 8348 7376 8490 7460
rect 8060 7340 8250 7376
rect 7838 7336 8250 7340
rect 7336 7288 7740 7336
rect 6836 7238 7238 7288
rect 6316 7208 6738 7238
rect 5824 7150 6218 7208
rect 5314 7110 5726 7150
tri 5726 7110 5766 7150 sw
tri 5824 7110 5864 7150 ne
rect 5864 7110 6218 7150
tri 6218 7110 6316 7208 sw
tri 6316 7110 6414 7208 ne
rect 6414 7150 6738 7208
tri 6738 7150 6826 7238 sw
tri 6836 7150 6924 7238 ne
rect 6924 7208 7238 7238
tri 7238 7208 7318 7288 sw
tri 7336 7208 7416 7288 ne
rect 7416 7238 7740 7288
tri 7740 7238 7838 7336 sw
tri 7838 7238 7936 7336 ne
rect 7936 7288 8250 7336
tri 8250 7288 8338 7376 sw
tri 8348 7288 8436 7376 ne
rect 8436 7340 8490 7376
rect 8610 7376 8712 7460
tri 8712 7376 8800 7464 sw
tri 8810 7376 8898 7464 ne
rect 8898 7460 9262 7464
rect 8898 7376 9040 7460
rect 8610 7340 8800 7376
rect 8436 7336 8800 7340
tri 8800 7336 8840 7376 sw
tri 8898 7336 8938 7376 ne
rect 8938 7340 9040 7376
rect 9160 7376 9262 7460
tri 9262 7376 9350 7464 sw
tri 9360 7376 9448 7464 ne
rect 9448 7460 9812 7464
rect 9448 7376 9590 7460
rect 9160 7340 9350 7376
rect 8938 7336 9350 7340
rect 8436 7288 8840 7336
rect 7936 7238 8338 7288
rect 7416 7208 7838 7238
rect 6924 7150 7318 7208
rect 6414 7110 6826 7150
tri 6826 7110 6866 7150 sw
tri 6924 7110 6964 7150 ne
rect 6964 7110 7318 7150
tri 7318 7110 7416 7208 sw
tri 7416 7110 7514 7208 ne
rect 7514 7150 7838 7208
tri 7838 7150 7926 7238 sw
tri 7936 7150 8024 7238 ne
rect 8024 7208 8338 7238
tri 8338 7208 8418 7288 sw
tri 8436 7208 8516 7288 ne
rect 8516 7238 8840 7288
tri 8840 7238 8938 7336 sw
tri 8938 7238 9036 7336 ne
rect 9036 7288 9350 7336
tri 9350 7288 9438 7376 sw
tri 9448 7288 9536 7376 ne
rect 9536 7340 9590 7376
rect 9710 7376 9812 7460
tri 9812 7376 9900 7464 sw
tri 9910 7376 9998 7464 ne
rect 9998 7460 10362 7464
rect 9998 7376 10140 7460
rect 9710 7340 9900 7376
rect 9536 7336 9900 7340
tri 9900 7336 9940 7376 sw
tri 9998 7336 10038 7376 ne
rect 10038 7340 10140 7376
rect 10260 7376 10362 7460
tri 10362 7376 10450 7464 sw
tri 10460 7376 10548 7464 ne
rect 10548 7460 10912 7464
rect 10548 7376 10690 7460
rect 10260 7340 10450 7376
rect 10038 7336 10450 7340
rect 9536 7288 9940 7336
rect 9036 7238 9438 7288
rect 8516 7208 8938 7238
rect 8024 7150 8418 7208
rect 7514 7110 7926 7150
tri 7926 7110 7966 7150 sw
tri 8024 7110 8064 7150 ne
rect 8064 7110 8418 7150
tri 8418 7110 8516 7208 sw
tri 8516 7110 8614 7208 ne
rect 8614 7150 8938 7208
tri 8938 7150 9026 7238 sw
tri 9036 7150 9124 7238 ne
rect 9124 7208 9438 7238
tri 9438 7208 9518 7288 sw
tri 9536 7208 9616 7288 ne
rect 9616 7238 9940 7288
tri 9940 7238 10038 7336 sw
tri 10038 7238 10136 7336 ne
rect 10136 7288 10450 7336
tri 10450 7288 10538 7376 sw
tri 10548 7288 10636 7376 ne
rect 10636 7340 10690 7376
rect 10810 7376 10912 7460
tri 10912 7376 11000 7464 sw
tri 11010 7376 11098 7464 ne
rect 11098 7460 11462 7464
rect 11098 7376 11240 7460
rect 10810 7340 11000 7376
rect 10636 7336 11000 7340
tri 11000 7336 11040 7376 sw
tri 11098 7336 11138 7376 ne
rect 11138 7340 11240 7376
rect 11360 7376 11462 7460
tri 11462 7376 11550 7464 sw
tri 11560 7376 11648 7464 ne
rect 11648 7460 12012 7464
rect 11648 7376 11790 7460
rect 11360 7340 11550 7376
rect 11138 7336 11550 7340
rect 10636 7288 11040 7336
rect 10136 7238 10538 7288
rect 9616 7208 10038 7238
rect 9124 7150 9518 7208
rect 8614 7110 9026 7150
tri 9026 7110 9066 7150 sw
tri 9124 7110 9164 7150 ne
rect 9164 7110 9518 7150
tri 9518 7110 9616 7208 sw
tri 9616 7110 9714 7208 ne
rect 9714 7150 10038 7208
tri 10038 7150 10126 7238 sw
tri 10136 7150 10224 7238 ne
rect 10224 7208 10538 7238
tri 10538 7208 10618 7288 sw
tri 10636 7208 10716 7288 ne
rect 10716 7238 11040 7288
tri 11040 7238 11138 7336 sw
tri 11138 7238 11236 7336 ne
rect 11236 7288 11550 7336
tri 11550 7288 11638 7376 sw
tri 11648 7288 11736 7376 ne
rect 11736 7340 11790 7376
rect 11910 7376 12012 7460
tri 12012 7376 12100 7464 sw
tri 12110 7376 12198 7464 ne
rect 12198 7460 12562 7464
rect 12198 7376 12340 7460
rect 11910 7340 12100 7376
rect 11736 7336 12100 7340
tri 12100 7336 12140 7376 sw
tri 12198 7336 12238 7376 ne
rect 12238 7340 12340 7376
rect 12460 7376 12562 7460
tri 12562 7376 12650 7464 sw
tri 12660 7376 12748 7464 ne
rect 12748 7460 13112 7464
rect 12748 7376 12890 7460
rect 12460 7340 12650 7376
rect 12238 7336 12650 7340
rect 11736 7288 12140 7336
rect 11236 7238 11638 7288
rect 10716 7208 11138 7238
rect 10224 7150 10618 7208
rect 9714 7110 10126 7150
tri 10126 7110 10166 7150 sw
tri 10224 7110 10264 7150 ne
rect 10264 7110 10618 7150
tri 10618 7110 10716 7208 sw
tri 10716 7110 10814 7208 ne
rect 10814 7150 11138 7208
tri 11138 7150 11226 7238 sw
tri 11236 7150 11324 7238 ne
rect 11324 7208 11638 7238
tri 11638 7208 11718 7288 sw
tri 11736 7208 11816 7288 ne
rect 11816 7238 12140 7288
tri 12140 7238 12238 7336 sw
tri 12238 7238 12336 7336 ne
rect 12336 7288 12650 7336
tri 12650 7288 12738 7376 sw
tri 12748 7288 12836 7376 ne
rect 12836 7340 12890 7376
rect 13010 7376 13112 7460
tri 13112 7376 13200 7464 sw
tri 13210 7376 13298 7464 ne
rect 13298 7460 14275 7464
rect 13298 7376 13440 7460
rect 13010 7340 13200 7376
rect 12836 7336 13200 7340
tri 13200 7336 13240 7376 sw
tri 13298 7336 13338 7376 ne
rect 13338 7340 13440 7376
rect 13560 7340 14275 7460
rect 13338 7336 14275 7340
rect 12836 7288 13240 7336
rect 12336 7238 12738 7288
rect 11816 7208 12238 7238
rect 11324 7150 11718 7208
rect 10814 7110 11226 7150
tri 11226 7110 11266 7150 sw
tri 11324 7110 11364 7150 ne
rect 11364 7110 11718 7150
tri 11718 7110 11816 7208 sw
tri 11816 7110 11914 7208 ne
rect 11914 7150 12238 7208
tri 12238 7150 12326 7238 sw
tri 12336 7150 12424 7238 ne
rect 12424 7208 12738 7238
tri 12738 7208 12818 7288 sw
tri 12836 7208 12916 7288 ne
rect 12916 7238 13240 7288
tri 13240 7238 13338 7336 sw
tri 13338 7238 13436 7336 ne
rect 13436 7238 14275 7336
rect 12916 7208 13338 7238
rect 12424 7150 12818 7208
rect 11914 7110 12326 7150
tri 12326 7110 12366 7150 sw
tri 12424 7110 12464 7150 ne
rect 12464 7110 12818 7150
tri 12818 7110 12916 7208 sw
tri 12916 7110 13014 7208 ne
rect 13014 7150 13338 7208
tri 13338 7150 13426 7238 sw
tri 13436 7150 13524 7238 ne
rect 13524 7150 14275 7238
rect 13014 7110 13426 7150
tri 13426 7110 13466 7150 sw
tri 13524 7110 13564 7150 ne
rect 13564 7110 14275 7150
rect -2525 7012 -284 7110
tri -284 7012 -186 7110 sw
tri -186 7012 -88 7110 ne
rect -88 7012 266 7110
tri 266 7012 364 7110 sw
tri 364 7012 462 7110 ne
rect 462 7012 816 7110
tri 816 7012 914 7110 sw
tri 914 7012 1012 7110 ne
rect 1012 7012 1366 7110
tri 1366 7012 1464 7110 sw
tri 1464 7012 1562 7110 ne
rect 1562 7012 1916 7110
tri 1916 7012 2014 7110 sw
tri 2014 7012 2112 7110 ne
rect 2112 7012 2466 7110
tri 2466 7012 2564 7110 sw
tri 2564 7012 2662 7110 ne
rect 2662 7012 3016 7110
tri 3016 7012 3114 7110 sw
tri 3114 7012 3212 7110 ne
rect 3212 7012 3566 7110
tri 3566 7012 3664 7110 sw
tri 3664 7012 3762 7110 ne
rect 3762 7012 4116 7110
tri 4116 7012 4214 7110 sw
tri 4214 7012 4312 7110 ne
rect 4312 7012 4666 7110
tri 4666 7012 4764 7110 sw
tri 4764 7012 4862 7110 ne
rect 4862 7012 5216 7110
tri 5216 7012 5314 7110 sw
tri 5314 7012 5412 7110 ne
rect 5412 7012 5766 7110
tri 5766 7012 5864 7110 sw
tri 5864 7012 5962 7110 ne
rect 5962 7012 6316 7110
tri 6316 7012 6414 7110 sw
tri 6414 7012 6512 7110 ne
rect 6512 7012 6866 7110
tri 6866 7012 6964 7110 sw
tri 6964 7012 7062 7110 ne
rect 7062 7012 7416 7110
tri 7416 7012 7514 7110 sw
tri 7514 7012 7612 7110 ne
rect 7612 7012 7966 7110
tri 7966 7012 8064 7110 sw
tri 8064 7012 8162 7110 ne
rect 8162 7012 8516 7110
tri 8516 7012 8614 7110 sw
tri 8614 7012 8712 7110 ne
rect 8712 7012 9066 7110
tri 9066 7012 9164 7110 sw
tri 9164 7012 9262 7110 ne
rect 9262 7012 9616 7110
tri 9616 7012 9714 7110 sw
tri 9714 7012 9812 7110 ne
rect 9812 7012 10166 7110
tri 10166 7012 10264 7110 sw
tri 10264 7012 10362 7110 ne
rect 10362 7012 10716 7110
tri 10716 7012 10814 7110 sw
tri 10814 7012 10912 7110 ne
rect 10912 7012 11266 7110
tri 11266 7012 11364 7110 sw
tri 11364 7012 11462 7110 ne
rect 11462 7012 11816 7110
tri 11816 7012 11914 7110 sw
tri 11914 7012 12012 7110 ne
rect 12012 7012 12366 7110
tri 12366 7012 12464 7110 sw
tri 12464 7012 12562 7110 ne
rect 12562 7012 12916 7110
tri 12916 7012 13014 7110 sw
tri 13014 7012 13112 7110 ne
rect 13112 7012 13466 7110
tri 13466 7012 13564 7110 sw
tri 13564 7012 13662 7110 ne
rect 13662 7012 14275 7110
rect -2525 6914 -186 7012
tri -186 6914 -88 7012 sw
tri -88 6914 10 7012 ne
rect 10 6914 364 7012
tri 364 6914 462 7012 sw
tri 462 6914 560 7012 ne
rect 560 6914 914 7012
tri 914 6914 1012 7012 sw
tri 1012 6914 1110 7012 ne
rect 1110 6914 1464 7012
tri 1464 6914 1562 7012 sw
tri 1562 6914 1660 7012 ne
rect 1660 6914 2014 7012
tri 2014 6914 2112 7012 sw
tri 2112 6914 2210 7012 ne
rect 2210 6914 2564 7012
tri 2564 6914 2662 7012 sw
tri 2662 6914 2760 7012 ne
rect 2760 6914 3114 7012
tri 3114 6914 3212 7012 sw
tri 3212 6914 3310 7012 ne
rect 3310 6914 3664 7012
tri 3664 6914 3762 7012 sw
tri 3762 6914 3860 7012 ne
rect 3860 6914 4214 7012
tri 4214 6914 4312 7012 sw
tri 4312 6914 4410 7012 ne
rect 4410 6914 4764 7012
tri 4764 6914 4862 7012 sw
tri 4862 6914 4960 7012 ne
rect 4960 6914 5314 7012
tri 5314 6914 5412 7012 sw
tri 5412 6914 5510 7012 ne
rect 5510 6914 5864 7012
tri 5864 6914 5962 7012 sw
tri 5962 6914 6060 7012 ne
rect 6060 6914 6414 7012
tri 6414 6914 6512 7012 sw
tri 6512 6914 6610 7012 ne
rect 6610 6914 6964 7012
tri 6964 6914 7062 7012 sw
tri 7062 6914 7160 7012 ne
rect 7160 6914 7514 7012
tri 7514 6914 7612 7012 sw
tri 7612 6914 7710 7012 ne
rect 7710 6914 8064 7012
tri 8064 6914 8162 7012 sw
tri 8162 6914 8260 7012 ne
rect 8260 6914 8614 7012
tri 8614 6914 8712 7012 sw
tri 8712 6914 8810 7012 ne
rect 8810 6914 9164 7012
tri 9164 6914 9262 7012 sw
tri 9262 6914 9360 7012 ne
rect 9360 6914 9714 7012
tri 9714 6914 9812 7012 sw
tri 9812 6914 9910 7012 ne
rect 9910 6914 10264 7012
tri 10264 6914 10362 7012 sw
tri 10362 6914 10460 7012 ne
rect 10460 6914 10814 7012
tri 10814 6914 10912 7012 sw
tri 10912 6914 11010 7012 ne
rect 11010 6914 11364 7012
tri 11364 6914 11462 7012 sw
tri 11462 6914 11560 7012 ne
rect 11560 6914 11914 7012
tri 11914 6914 12012 7012 sw
tri 12012 6914 12110 7012 ne
rect 12110 6914 12464 7012
tri 12464 6914 12562 7012 sw
tri 12562 6914 12660 7012 ne
rect 12660 6914 13014 7012
tri 13014 6914 13112 7012 sw
tri 13112 6914 13210 7012 ne
rect 13210 6914 13564 7012
tri 13564 6914 13662 7012 sw
rect 14775 6914 15775 7562
rect -2525 6910 -88 6914
rect -2525 6790 -310 6910
rect -190 6826 -88 6910
tri -88 6826 0 6914 sw
tri 10 6826 98 6914 ne
rect 98 6910 462 6914
rect 98 6826 240 6910
rect -190 6790 0 6826
rect -2525 6786 0 6790
rect -2525 6138 -1525 6786
tri -412 6688 -314 6786 ne
rect -314 6738 0 6786
tri 0 6738 88 6826 sw
tri 98 6738 186 6826 ne
rect 186 6790 240 6826
rect 360 6826 462 6910
tri 462 6826 550 6914 sw
tri 560 6826 648 6914 ne
rect 648 6910 1012 6914
rect 648 6826 790 6910
rect 360 6790 550 6826
rect 186 6786 550 6790
tri 550 6786 590 6826 sw
tri 648 6786 688 6826 ne
rect 688 6790 790 6826
rect 910 6826 1012 6910
tri 1012 6826 1100 6914 sw
tri 1110 6826 1198 6914 ne
rect 1198 6910 1562 6914
rect 1198 6826 1340 6910
rect 910 6790 1100 6826
rect 688 6786 1100 6790
rect 186 6738 590 6786
rect -314 6688 88 6738
rect -1025 6600 -412 6688
tri -412 6600 -324 6688 sw
tri -314 6600 -226 6688 ne
rect -226 6658 88 6688
tri 88 6658 168 6738 sw
tri 186 6658 266 6738 ne
rect 266 6688 590 6738
tri 590 6688 688 6786 sw
tri 688 6688 786 6786 ne
rect 786 6738 1100 6786
tri 1100 6738 1188 6826 sw
tri 1198 6738 1286 6826 ne
rect 1286 6790 1340 6826
rect 1460 6826 1562 6910
tri 1562 6826 1650 6914 sw
tri 1660 6826 1748 6914 ne
rect 1748 6910 2112 6914
rect 1748 6826 1890 6910
rect 1460 6790 1650 6826
rect 1286 6786 1650 6790
tri 1650 6786 1690 6826 sw
tri 1748 6786 1788 6826 ne
rect 1788 6790 1890 6826
rect 2010 6826 2112 6910
tri 2112 6826 2200 6914 sw
tri 2210 6826 2298 6914 ne
rect 2298 6910 2662 6914
rect 2298 6826 2440 6910
rect 2010 6790 2200 6826
rect 1788 6786 2200 6790
rect 1286 6738 1690 6786
rect 786 6688 1188 6738
rect 266 6658 688 6688
rect -226 6600 168 6658
rect -1025 6560 -324 6600
tri -324 6560 -284 6600 sw
tri -226 6560 -186 6600 ne
rect -186 6560 168 6600
tri 168 6560 266 6658 sw
tri 266 6560 364 6658 ne
rect 364 6600 688 6658
tri 688 6600 776 6688 sw
tri 786 6600 874 6688 ne
rect 874 6658 1188 6688
tri 1188 6658 1268 6738 sw
tri 1286 6658 1366 6738 ne
rect 1366 6688 1690 6738
tri 1690 6688 1788 6786 sw
tri 1788 6688 1886 6786 ne
rect 1886 6738 2200 6786
tri 2200 6738 2288 6826 sw
tri 2298 6738 2386 6826 ne
rect 2386 6790 2440 6826
rect 2560 6826 2662 6910
tri 2662 6826 2750 6914 sw
tri 2760 6826 2848 6914 ne
rect 2848 6910 3212 6914
rect 2848 6826 2990 6910
rect 2560 6790 2750 6826
rect 2386 6786 2750 6790
tri 2750 6786 2790 6826 sw
tri 2848 6786 2888 6826 ne
rect 2888 6790 2990 6826
rect 3110 6826 3212 6910
tri 3212 6826 3300 6914 sw
tri 3310 6826 3398 6914 ne
rect 3398 6910 3762 6914
rect 3398 6826 3540 6910
rect 3110 6790 3300 6826
rect 2888 6786 3300 6790
rect 2386 6738 2790 6786
rect 1886 6688 2288 6738
rect 1366 6658 1788 6688
rect 874 6600 1268 6658
rect 364 6560 776 6600
tri 776 6560 816 6600 sw
tri 874 6560 914 6600 ne
rect 914 6560 1268 6600
tri 1268 6560 1366 6658 sw
tri 1366 6560 1464 6658 ne
rect 1464 6600 1788 6658
tri 1788 6600 1876 6688 sw
tri 1886 6600 1974 6688 ne
rect 1974 6658 2288 6688
tri 2288 6658 2368 6738 sw
tri 2386 6658 2466 6738 ne
rect 2466 6688 2790 6738
tri 2790 6688 2888 6786 sw
tri 2888 6688 2986 6786 ne
rect 2986 6738 3300 6786
tri 3300 6738 3388 6826 sw
tri 3398 6738 3486 6826 ne
rect 3486 6790 3540 6826
rect 3660 6826 3762 6910
tri 3762 6826 3850 6914 sw
tri 3860 6826 3948 6914 ne
rect 3948 6910 4312 6914
rect 3948 6826 4090 6910
rect 3660 6790 3850 6826
rect 3486 6786 3850 6790
tri 3850 6786 3890 6826 sw
tri 3948 6786 3988 6826 ne
rect 3988 6790 4090 6826
rect 4210 6826 4312 6910
tri 4312 6826 4400 6914 sw
tri 4410 6826 4498 6914 ne
rect 4498 6910 4862 6914
rect 4498 6826 4640 6910
rect 4210 6790 4400 6826
rect 3988 6786 4400 6790
rect 3486 6738 3890 6786
rect 2986 6688 3388 6738
rect 2466 6658 2888 6688
rect 1974 6600 2368 6658
rect 1464 6560 1876 6600
tri 1876 6560 1916 6600 sw
tri 1974 6560 2014 6600 ne
rect 2014 6560 2368 6600
tri 2368 6560 2466 6658 sw
tri 2466 6560 2564 6658 ne
rect 2564 6600 2888 6658
tri 2888 6600 2976 6688 sw
tri 2986 6600 3074 6688 ne
rect 3074 6658 3388 6688
tri 3388 6658 3468 6738 sw
tri 3486 6658 3566 6738 ne
rect 3566 6688 3890 6738
tri 3890 6688 3988 6786 sw
tri 3988 6688 4086 6786 ne
rect 4086 6738 4400 6786
tri 4400 6738 4488 6826 sw
tri 4498 6738 4586 6826 ne
rect 4586 6790 4640 6826
rect 4760 6826 4862 6910
tri 4862 6826 4950 6914 sw
tri 4960 6826 5048 6914 ne
rect 5048 6910 5412 6914
rect 5048 6826 5190 6910
rect 4760 6790 4950 6826
rect 4586 6786 4950 6790
tri 4950 6786 4990 6826 sw
tri 5048 6786 5088 6826 ne
rect 5088 6790 5190 6826
rect 5310 6826 5412 6910
tri 5412 6826 5500 6914 sw
tri 5510 6826 5598 6914 ne
rect 5598 6910 5962 6914
rect 5598 6826 5740 6910
rect 5310 6790 5500 6826
rect 5088 6786 5500 6790
rect 4586 6738 4990 6786
rect 4086 6688 4488 6738
rect 3566 6658 3988 6688
rect 3074 6600 3468 6658
rect 2564 6560 2976 6600
tri 2976 6560 3016 6600 sw
tri 3074 6560 3114 6600 ne
rect 3114 6560 3468 6600
tri 3468 6560 3566 6658 sw
tri 3566 6560 3664 6658 ne
rect 3664 6600 3988 6658
tri 3988 6600 4076 6688 sw
tri 4086 6600 4174 6688 ne
rect 4174 6658 4488 6688
tri 4488 6658 4568 6738 sw
tri 4586 6658 4666 6738 ne
rect 4666 6688 4990 6738
tri 4990 6688 5088 6786 sw
tri 5088 6688 5186 6786 ne
rect 5186 6738 5500 6786
tri 5500 6738 5588 6826 sw
tri 5598 6738 5686 6826 ne
rect 5686 6790 5740 6826
rect 5860 6826 5962 6910
tri 5962 6826 6050 6914 sw
tri 6060 6826 6148 6914 ne
rect 6148 6910 6512 6914
rect 6148 6826 6290 6910
rect 5860 6790 6050 6826
rect 5686 6786 6050 6790
tri 6050 6786 6090 6826 sw
tri 6148 6786 6188 6826 ne
rect 6188 6790 6290 6826
rect 6410 6826 6512 6910
tri 6512 6826 6600 6914 sw
tri 6610 6826 6698 6914 ne
rect 6698 6910 7062 6914
rect 6698 6826 6840 6910
rect 6410 6790 6600 6826
rect 6188 6786 6600 6790
rect 5686 6738 6090 6786
rect 5186 6688 5588 6738
rect 4666 6658 5088 6688
rect 4174 6600 4568 6658
rect 3664 6560 4076 6600
tri 4076 6560 4116 6600 sw
tri 4174 6560 4214 6600 ne
rect 4214 6560 4568 6600
tri 4568 6560 4666 6658 sw
tri 4666 6560 4764 6658 ne
rect 4764 6600 5088 6658
tri 5088 6600 5176 6688 sw
tri 5186 6600 5274 6688 ne
rect 5274 6658 5588 6688
tri 5588 6658 5668 6738 sw
tri 5686 6658 5766 6738 ne
rect 5766 6688 6090 6738
tri 6090 6688 6188 6786 sw
tri 6188 6688 6286 6786 ne
rect 6286 6738 6600 6786
tri 6600 6738 6688 6826 sw
tri 6698 6738 6786 6826 ne
rect 6786 6790 6840 6826
rect 6960 6826 7062 6910
tri 7062 6826 7150 6914 sw
tri 7160 6826 7248 6914 ne
rect 7248 6910 7612 6914
rect 7248 6826 7390 6910
rect 6960 6790 7150 6826
rect 6786 6786 7150 6790
tri 7150 6786 7190 6826 sw
tri 7248 6786 7288 6826 ne
rect 7288 6790 7390 6826
rect 7510 6826 7612 6910
tri 7612 6826 7700 6914 sw
tri 7710 6826 7798 6914 ne
rect 7798 6910 8162 6914
rect 7798 6826 7940 6910
rect 7510 6790 7700 6826
rect 7288 6786 7700 6790
rect 6786 6738 7190 6786
rect 6286 6688 6688 6738
rect 5766 6658 6188 6688
rect 5274 6600 5668 6658
rect 4764 6560 5176 6600
tri 5176 6560 5216 6600 sw
tri 5274 6560 5314 6600 ne
rect 5314 6560 5668 6600
tri 5668 6560 5766 6658 sw
tri 5766 6560 5864 6658 ne
rect 5864 6600 6188 6658
tri 6188 6600 6276 6688 sw
tri 6286 6600 6374 6688 ne
rect 6374 6658 6688 6688
tri 6688 6658 6768 6738 sw
tri 6786 6658 6866 6738 ne
rect 6866 6688 7190 6738
tri 7190 6688 7288 6786 sw
tri 7288 6688 7386 6786 ne
rect 7386 6738 7700 6786
tri 7700 6738 7788 6826 sw
tri 7798 6738 7886 6826 ne
rect 7886 6790 7940 6826
rect 8060 6826 8162 6910
tri 8162 6826 8250 6914 sw
tri 8260 6826 8348 6914 ne
rect 8348 6910 8712 6914
rect 8348 6826 8490 6910
rect 8060 6790 8250 6826
rect 7886 6786 8250 6790
tri 8250 6786 8290 6826 sw
tri 8348 6786 8388 6826 ne
rect 8388 6790 8490 6826
rect 8610 6826 8712 6910
tri 8712 6826 8800 6914 sw
tri 8810 6826 8898 6914 ne
rect 8898 6910 9262 6914
rect 8898 6826 9040 6910
rect 8610 6790 8800 6826
rect 8388 6786 8800 6790
rect 7886 6738 8290 6786
rect 7386 6688 7788 6738
rect 6866 6658 7288 6688
rect 6374 6600 6768 6658
rect 5864 6560 6276 6600
tri 6276 6560 6316 6600 sw
tri 6374 6560 6414 6600 ne
rect 6414 6560 6768 6600
tri 6768 6560 6866 6658 sw
tri 6866 6560 6964 6658 ne
rect 6964 6600 7288 6658
tri 7288 6600 7376 6688 sw
tri 7386 6600 7474 6688 ne
rect 7474 6658 7788 6688
tri 7788 6658 7868 6738 sw
tri 7886 6658 7966 6738 ne
rect 7966 6688 8290 6738
tri 8290 6688 8388 6786 sw
tri 8388 6688 8486 6786 ne
rect 8486 6738 8800 6786
tri 8800 6738 8888 6826 sw
tri 8898 6738 8986 6826 ne
rect 8986 6790 9040 6826
rect 9160 6826 9262 6910
tri 9262 6826 9350 6914 sw
tri 9360 6826 9448 6914 ne
rect 9448 6910 9812 6914
rect 9448 6826 9590 6910
rect 9160 6790 9350 6826
rect 8986 6786 9350 6790
tri 9350 6786 9390 6826 sw
tri 9448 6786 9488 6826 ne
rect 9488 6790 9590 6826
rect 9710 6826 9812 6910
tri 9812 6826 9900 6914 sw
tri 9910 6826 9998 6914 ne
rect 9998 6910 10362 6914
rect 9998 6826 10140 6910
rect 9710 6790 9900 6826
rect 9488 6786 9900 6790
rect 8986 6738 9390 6786
rect 8486 6688 8888 6738
rect 7966 6658 8388 6688
rect 7474 6600 7868 6658
rect 6964 6560 7376 6600
tri 7376 6560 7416 6600 sw
tri 7474 6560 7514 6600 ne
rect 7514 6560 7868 6600
tri 7868 6560 7966 6658 sw
tri 7966 6560 8064 6658 ne
rect 8064 6600 8388 6658
tri 8388 6600 8476 6688 sw
tri 8486 6600 8574 6688 ne
rect 8574 6658 8888 6688
tri 8888 6658 8968 6738 sw
tri 8986 6658 9066 6738 ne
rect 9066 6688 9390 6738
tri 9390 6688 9488 6786 sw
tri 9488 6688 9586 6786 ne
rect 9586 6738 9900 6786
tri 9900 6738 9988 6826 sw
tri 9998 6738 10086 6826 ne
rect 10086 6790 10140 6826
rect 10260 6826 10362 6910
tri 10362 6826 10450 6914 sw
tri 10460 6826 10548 6914 ne
rect 10548 6910 10912 6914
rect 10548 6826 10690 6910
rect 10260 6790 10450 6826
rect 10086 6786 10450 6790
tri 10450 6786 10490 6826 sw
tri 10548 6786 10588 6826 ne
rect 10588 6790 10690 6826
rect 10810 6826 10912 6910
tri 10912 6826 11000 6914 sw
tri 11010 6826 11098 6914 ne
rect 11098 6910 11462 6914
rect 11098 6826 11240 6910
rect 10810 6790 11000 6826
rect 10588 6786 11000 6790
rect 10086 6738 10490 6786
rect 9586 6688 9988 6738
rect 9066 6658 9488 6688
rect 8574 6600 8968 6658
rect 8064 6560 8476 6600
tri 8476 6560 8516 6600 sw
tri 8574 6560 8614 6600 ne
rect 8614 6560 8968 6600
tri 8968 6560 9066 6658 sw
tri 9066 6560 9164 6658 ne
rect 9164 6600 9488 6658
tri 9488 6600 9576 6688 sw
tri 9586 6600 9674 6688 ne
rect 9674 6658 9988 6688
tri 9988 6658 10068 6738 sw
tri 10086 6658 10166 6738 ne
rect 10166 6688 10490 6738
tri 10490 6688 10588 6786 sw
tri 10588 6688 10686 6786 ne
rect 10686 6738 11000 6786
tri 11000 6738 11088 6826 sw
tri 11098 6738 11186 6826 ne
rect 11186 6790 11240 6826
rect 11360 6826 11462 6910
tri 11462 6826 11550 6914 sw
tri 11560 6826 11648 6914 ne
rect 11648 6910 12012 6914
rect 11648 6826 11790 6910
rect 11360 6790 11550 6826
rect 11186 6786 11550 6790
tri 11550 6786 11590 6826 sw
tri 11648 6786 11688 6826 ne
rect 11688 6790 11790 6826
rect 11910 6826 12012 6910
tri 12012 6826 12100 6914 sw
tri 12110 6826 12198 6914 ne
rect 12198 6910 12562 6914
rect 12198 6826 12340 6910
rect 11910 6790 12100 6826
rect 11688 6786 12100 6790
rect 11186 6738 11590 6786
rect 10686 6688 11088 6738
rect 10166 6658 10588 6688
rect 9674 6600 10068 6658
rect 9164 6560 9576 6600
tri 9576 6560 9616 6600 sw
tri 9674 6560 9714 6600 ne
rect 9714 6560 10068 6600
tri 10068 6560 10166 6658 sw
tri 10166 6560 10264 6658 ne
rect 10264 6600 10588 6658
tri 10588 6600 10676 6688 sw
tri 10686 6600 10774 6688 ne
rect 10774 6658 11088 6688
tri 11088 6658 11168 6738 sw
tri 11186 6658 11266 6738 ne
rect 11266 6688 11590 6738
tri 11590 6688 11688 6786 sw
tri 11688 6688 11786 6786 ne
rect 11786 6738 12100 6786
tri 12100 6738 12188 6826 sw
tri 12198 6738 12286 6826 ne
rect 12286 6790 12340 6826
rect 12460 6826 12562 6910
tri 12562 6826 12650 6914 sw
tri 12660 6826 12748 6914 ne
rect 12748 6910 13112 6914
rect 12748 6826 12890 6910
rect 12460 6790 12650 6826
rect 12286 6786 12650 6790
tri 12650 6786 12690 6826 sw
tri 12748 6786 12788 6826 ne
rect 12788 6790 12890 6826
rect 13010 6826 13112 6910
tri 13112 6826 13200 6914 sw
tri 13210 6826 13298 6914 ne
rect 13298 6910 15775 6914
rect 13298 6826 13440 6910
rect 13010 6790 13200 6826
rect 12788 6786 13200 6790
rect 12286 6738 12690 6786
rect 11786 6688 12188 6738
rect 11266 6658 11688 6688
rect 10774 6600 11168 6658
rect 10264 6560 10676 6600
tri 10676 6560 10716 6600 sw
tri 10774 6560 10814 6600 ne
rect 10814 6560 11168 6600
tri 11168 6560 11266 6658 sw
tri 11266 6560 11364 6658 ne
rect 11364 6600 11688 6658
tri 11688 6600 11776 6688 sw
tri 11786 6600 11874 6688 ne
rect 11874 6658 12188 6688
tri 12188 6658 12268 6738 sw
tri 12286 6658 12366 6738 ne
rect 12366 6688 12690 6738
tri 12690 6688 12788 6786 sw
tri 12788 6688 12886 6786 ne
rect 12886 6738 13200 6786
tri 13200 6738 13288 6826 sw
tri 13298 6738 13386 6826 ne
rect 13386 6790 13440 6826
rect 13560 6790 15775 6910
rect 13386 6738 15775 6790
rect 12886 6688 13288 6738
rect 12366 6658 12788 6688
rect 11874 6600 12268 6658
rect 11364 6560 11776 6600
tri 11776 6560 11816 6600 sw
tri 11874 6560 11914 6600 ne
rect 11914 6560 12268 6600
tri 12268 6560 12366 6658 sw
tri 12366 6560 12464 6658 ne
rect 12464 6600 12788 6658
tri 12788 6600 12876 6688 sw
tri 12886 6600 12974 6688 ne
rect 12974 6658 13288 6688
tri 13288 6658 13368 6738 sw
tri 13386 6658 13466 6738 ne
rect 13466 6658 14075 6738
rect 12974 6600 13368 6658
rect 12464 6560 12876 6600
tri 12876 6560 12916 6600 sw
tri 12974 6560 13014 6600 ne
rect 13014 6560 13368 6600
tri 13368 6560 13466 6658 sw
tri 13466 6560 13564 6658 ne
rect 13564 6638 14075 6658
rect 14175 6638 15775 6738
rect 13564 6560 15775 6638
rect -1025 6512 -284 6560
rect -1025 6412 -925 6512
rect -825 6462 -284 6512
tri -284 6462 -186 6560 sw
tri -186 6462 -88 6560 ne
rect -88 6462 266 6560
tri 266 6462 364 6560 sw
tri 364 6462 462 6560 ne
rect 462 6462 816 6560
tri 816 6462 914 6560 sw
tri 914 6462 1012 6560 ne
rect 1012 6462 1366 6560
tri 1366 6462 1464 6560 sw
tri 1464 6462 1562 6560 ne
rect 1562 6462 1916 6560
tri 1916 6462 2014 6560 sw
tri 2014 6462 2112 6560 ne
rect 2112 6462 2466 6560
tri 2466 6462 2564 6560 sw
tri 2564 6462 2662 6560 ne
rect 2662 6462 3016 6560
tri 3016 6462 3114 6560 sw
tri 3114 6462 3212 6560 ne
rect 3212 6462 3566 6560
tri 3566 6462 3664 6560 sw
tri 3664 6462 3762 6560 ne
rect 3762 6462 4116 6560
tri 4116 6462 4214 6560 sw
tri 4214 6462 4312 6560 ne
rect 4312 6462 4666 6560
tri 4666 6462 4764 6560 sw
tri 4764 6462 4862 6560 ne
rect 4862 6462 5216 6560
tri 5216 6462 5314 6560 sw
tri 5314 6462 5412 6560 ne
rect 5412 6462 5766 6560
tri 5766 6462 5864 6560 sw
tri 5864 6462 5962 6560 ne
rect 5962 6462 6316 6560
tri 6316 6462 6414 6560 sw
tri 6414 6462 6512 6560 ne
rect 6512 6462 6866 6560
tri 6866 6462 6964 6560 sw
tri 6964 6462 7062 6560 ne
rect 7062 6462 7416 6560
tri 7416 6462 7514 6560 sw
tri 7514 6462 7612 6560 ne
rect 7612 6462 7966 6560
tri 7966 6462 8064 6560 sw
tri 8064 6462 8162 6560 ne
rect 8162 6462 8516 6560
tri 8516 6462 8614 6560 sw
tri 8614 6462 8712 6560 ne
rect 8712 6462 9066 6560
tri 9066 6462 9164 6560 sw
tri 9164 6462 9262 6560 ne
rect 9262 6462 9616 6560
tri 9616 6462 9714 6560 sw
tri 9714 6462 9812 6560 ne
rect 9812 6462 10166 6560
tri 10166 6462 10264 6560 sw
tri 10264 6462 10362 6560 ne
rect 10362 6462 10716 6560
tri 10716 6462 10814 6560 sw
tri 10814 6462 10912 6560 ne
rect 10912 6462 11266 6560
tri 11266 6462 11364 6560 sw
tri 11364 6462 11462 6560 ne
rect 11462 6462 11816 6560
tri 11816 6462 11914 6560 sw
tri 11914 6462 12012 6560 ne
rect 12012 6462 12366 6560
tri 12366 6462 12464 6560 sw
tri 12464 6462 12562 6560 ne
rect 12562 6462 12916 6560
tri 12916 6462 13014 6560 sw
tri 13014 6462 13112 6560 ne
rect 13112 6462 13466 6560
tri 13466 6462 13564 6560 sw
tri 13564 6462 13662 6560 ne
rect 13662 6462 15775 6560
rect -825 6412 -186 6462
rect -1025 6364 -186 6412
tri -186 6364 -88 6462 sw
tri -88 6364 10 6462 ne
rect 10 6364 364 6462
tri 364 6364 462 6462 sw
tri 462 6364 560 6462 ne
rect 560 6364 914 6462
tri 914 6364 1012 6462 sw
tri 1012 6364 1110 6462 ne
rect 1110 6364 1464 6462
tri 1464 6364 1562 6462 sw
tri 1562 6364 1660 6462 ne
rect 1660 6364 2014 6462
tri 2014 6364 2112 6462 sw
tri 2112 6364 2210 6462 ne
rect 2210 6364 2564 6462
tri 2564 6364 2662 6462 sw
tri 2662 6364 2760 6462 ne
rect 2760 6364 3114 6462
tri 3114 6364 3212 6462 sw
tri 3212 6364 3310 6462 ne
rect 3310 6364 3664 6462
tri 3664 6364 3762 6462 sw
tri 3762 6364 3860 6462 ne
rect 3860 6364 4214 6462
tri 4214 6364 4312 6462 sw
tri 4312 6364 4410 6462 ne
rect 4410 6364 4764 6462
tri 4764 6364 4862 6462 sw
tri 4862 6364 4960 6462 ne
rect 4960 6364 5314 6462
tri 5314 6364 5412 6462 sw
tri 5412 6364 5510 6462 ne
rect 5510 6364 5864 6462
tri 5864 6364 5962 6462 sw
tri 5962 6364 6060 6462 ne
rect 6060 6364 6414 6462
tri 6414 6364 6512 6462 sw
tri 6512 6364 6610 6462 ne
rect 6610 6364 6964 6462
tri 6964 6364 7062 6462 sw
tri 7062 6364 7160 6462 ne
rect 7160 6364 7514 6462
tri 7514 6364 7612 6462 sw
tri 7612 6364 7710 6462 ne
rect 7710 6364 8064 6462
tri 8064 6364 8162 6462 sw
tri 8162 6364 8260 6462 ne
rect 8260 6364 8614 6462
tri 8614 6364 8712 6462 sw
tri 8712 6364 8810 6462 ne
rect 8810 6364 9164 6462
tri 9164 6364 9262 6462 sw
tri 9262 6364 9360 6462 ne
rect 9360 6364 9714 6462
tri 9714 6364 9812 6462 sw
tri 9812 6364 9910 6462 ne
rect 9910 6364 10264 6462
tri 10264 6364 10362 6462 sw
tri 10362 6364 10460 6462 ne
rect 10460 6364 10814 6462
tri 10814 6364 10912 6462 sw
tri 10912 6364 11010 6462 ne
rect 11010 6364 11364 6462
tri 11364 6364 11462 6462 sw
tri 11462 6364 11560 6462 ne
rect 11560 6364 11914 6462
tri 11914 6364 12012 6462 sw
tri 12012 6364 12110 6462 ne
rect 12110 6364 12464 6462
tri 12464 6364 12562 6462 sw
tri 12562 6364 12660 6462 ne
rect 12660 6364 13014 6462
tri 13014 6364 13112 6462 sw
tri 13112 6364 13210 6462 ne
rect 13210 6364 13564 6462
tri 13564 6364 13662 6462 sw
rect -1025 6360 -88 6364
rect -1025 6240 -310 6360
rect -190 6276 -88 6360
tri -88 6276 0 6364 sw
tri 10 6276 98 6364 ne
rect 98 6360 462 6364
rect 98 6276 240 6360
rect -190 6240 0 6276
rect -1025 6236 0 6240
tri 0 6236 40 6276 sw
tri 98 6236 138 6276 ne
rect 138 6240 240 6276
rect 360 6276 462 6360
tri 462 6276 550 6364 sw
tri 560 6276 648 6364 ne
rect 648 6360 1012 6364
rect 648 6276 790 6360
rect 360 6240 550 6276
rect 138 6236 550 6240
tri -412 6138 -314 6236 ne
rect -314 6138 40 6236
tri 40 6138 138 6236 sw
tri 138 6138 236 6236 ne
rect 236 6188 550 6236
tri 550 6188 638 6276 sw
tri 648 6188 736 6276 ne
rect 736 6240 790 6276
rect 910 6276 1012 6360
tri 1012 6276 1100 6364 sw
tri 1110 6276 1198 6364 ne
rect 1198 6360 1562 6364
rect 1198 6276 1340 6360
rect 910 6240 1100 6276
rect 736 6236 1100 6240
tri 1100 6236 1140 6276 sw
tri 1198 6236 1238 6276 ne
rect 1238 6240 1340 6276
rect 1460 6276 1562 6360
tri 1562 6276 1650 6364 sw
tri 1660 6276 1748 6364 ne
rect 1748 6360 2112 6364
rect 1748 6276 1890 6360
rect 1460 6240 1650 6276
rect 1238 6236 1650 6240
rect 736 6188 1140 6236
rect 236 6138 638 6188
rect -2525 6050 -412 6138
tri -412 6050 -324 6138 sw
tri -314 6050 -226 6138 ne
rect -226 6050 138 6138
tri 138 6050 226 6138 sw
tri 236 6050 324 6138 ne
rect 324 6108 638 6138
tri 638 6108 718 6188 sw
tri 736 6108 816 6188 ne
rect 816 6138 1140 6188
tri 1140 6138 1238 6236 sw
tri 1238 6138 1336 6236 ne
rect 1336 6188 1650 6236
tri 1650 6188 1738 6276 sw
tri 1748 6188 1836 6276 ne
rect 1836 6240 1890 6276
rect 2010 6276 2112 6360
tri 2112 6276 2200 6364 sw
tri 2210 6276 2298 6364 ne
rect 2298 6360 2662 6364
rect 2298 6276 2440 6360
rect 2010 6240 2200 6276
rect 1836 6236 2200 6240
tri 2200 6236 2240 6276 sw
tri 2298 6236 2338 6276 ne
rect 2338 6240 2440 6276
rect 2560 6276 2662 6360
tri 2662 6276 2750 6364 sw
tri 2760 6276 2848 6364 ne
rect 2848 6360 3212 6364
rect 2848 6276 2990 6360
rect 2560 6240 2750 6276
rect 2338 6236 2750 6240
rect 1836 6188 2240 6236
rect 1336 6138 1738 6188
rect 816 6108 1238 6138
rect 324 6050 718 6108
rect -2525 6010 -324 6050
tri -324 6010 -284 6050 sw
tri -226 6010 -186 6050 ne
rect -186 6010 226 6050
tri 226 6010 266 6050 sw
tri 324 6010 364 6050 ne
rect 364 6010 718 6050
tri 718 6010 816 6108 sw
tri 816 6010 914 6108 ne
rect 914 6050 1238 6108
tri 1238 6050 1326 6138 sw
tri 1336 6050 1424 6138 ne
rect 1424 6108 1738 6138
tri 1738 6108 1818 6188 sw
tri 1836 6108 1916 6188 ne
rect 1916 6138 2240 6188
tri 2240 6138 2338 6236 sw
tri 2338 6138 2436 6236 ne
rect 2436 6188 2750 6236
tri 2750 6188 2838 6276 sw
tri 2848 6188 2936 6276 ne
rect 2936 6240 2990 6276
rect 3110 6276 3212 6360
tri 3212 6276 3300 6364 sw
tri 3310 6276 3398 6364 ne
rect 3398 6360 3762 6364
rect 3398 6276 3540 6360
rect 3110 6240 3300 6276
rect 2936 6236 3300 6240
tri 3300 6236 3340 6276 sw
tri 3398 6236 3438 6276 ne
rect 3438 6240 3540 6276
rect 3660 6276 3762 6360
tri 3762 6276 3850 6364 sw
tri 3860 6276 3948 6364 ne
rect 3948 6360 4312 6364
rect 3948 6276 4090 6360
rect 3660 6240 3850 6276
rect 3438 6236 3850 6240
rect 2936 6188 3340 6236
rect 2436 6138 2838 6188
rect 1916 6108 2338 6138
rect 1424 6050 1818 6108
rect 914 6010 1326 6050
tri 1326 6010 1366 6050 sw
tri 1424 6010 1464 6050 ne
rect 1464 6010 1818 6050
tri 1818 6010 1916 6108 sw
tri 1916 6010 2014 6108 ne
rect 2014 6050 2338 6108
tri 2338 6050 2426 6138 sw
tri 2436 6050 2524 6138 ne
rect 2524 6108 2838 6138
tri 2838 6108 2918 6188 sw
tri 2936 6108 3016 6188 ne
rect 3016 6138 3340 6188
tri 3340 6138 3438 6236 sw
tri 3438 6138 3536 6236 ne
rect 3536 6188 3850 6236
tri 3850 6188 3938 6276 sw
tri 3948 6188 4036 6276 ne
rect 4036 6240 4090 6276
rect 4210 6276 4312 6360
tri 4312 6276 4400 6364 sw
tri 4410 6276 4498 6364 ne
rect 4498 6360 4862 6364
rect 4498 6276 4640 6360
rect 4210 6240 4400 6276
rect 4036 6236 4400 6240
tri 4400 6236 4440 6276 sw
tri 4498 6236 4538 6276 ne
rect 4538 6240 4640 6276
rect 4760 6276 4862 6360
tri 4862 6276 4950 6364 sw
tri 4960 6276 5048 6364 ne
rect 5048 6360 5412 6364
rect 5048 6276 5190 6360
rect 4760 6240 4950 6276
rect 4538 6236 4950 6240
rect 4036 6188 4440 6236
rect 3536 6138 3938 6188
rect 3016 6108 3438 6138
rect 2524 6050 2918 6108
rect 2014 6010 2426 6050
tri 2426 6010 2466 6050 sw
tri 2524 6010 2564 6050 ne
rect 2564 6010 2918 6050
tri 2918 6010 3016 6108 sw
tri 3016 6010 3114 6108 ne
rect 3114 6050 3438 6108
tri 3438 6050 3526 6138 sw
tri 3536 6050 3624 6138 ne
rect 3624 6108 3938 6138
tri 3938 6108 4018 6188 sw
tri 4036 6108 4116 6188 ne
rect 4116 6138 4440 6188
tri 4440 6138 4538 6236 sw
tri 4538 6138 4636 6236 ne
rect 4636 6188 4950 6236
tri 4950 6188 5038 6276 sw
tri 5048 6188 5136 6276 ne
rect 5136 6240 5190 6276
rect 5310 6276 5412 6360
tri 5412 6276 5500 6364 sw
tri 5510 6276 5598 6364 ne
rect 5598 6360 5962 6364
rect 5598 6276 5740 6360
rect 5310 6240 5500 6276
rect 5136 6236 5500 6240
tri 5500 6236 5540 6276 sw
tri 5598 6236 5638 6276 ne
rect 5638 6240 5740 6276
rect 5860 6276 5962 6360
tri 5962 6276 6050 6364 sw
tri 6060 6276 6148 6364 ne
rect 6148 6360 6512 6364
rect 6148 6276 6290 6360
rect 5860 6240 6050 6276
rect 5638 6236 6050 6240
rect 5136 6188 5540 6236
rect 4636 6138 5038 6188
rect 4116 6108 4538 6138
rect 3624 6050 4018 6108
rect 3114 6010 3526 6050
tri 3526 6010 3566 6050 sw
tri 3624 6010 3664 6050 ne
rect 3664 6010 4018 6050
tri 4018 6010 4116 6108 sw
tri 4116 6010 4214 6108 ne
rect 4214 6050 4538 6108
tri 4538 6050 4626 6138 sw
tri 4636 6050 4724 6138 ne
rect 4724 6108 5038 6138
tri 5038 6108 5118 6188 sw
tri 5136 6108 5216 6188 ne
rect 5216 6138 5540 6188
tri 5540 6138 5638 6236 sw
tri 5638 6138 5736 6236 ne
rect 5736 6188 6050 6236
tri 6050 6188 6138 6276 sw
tri 6148 6188 6236 6276 ne
rect 6236 6240 6290 6276
rect 6410 6276 6512 6360
tri 6512 6276 6600 6364 sw
tri 6610 6276 6698 6364 ne
rect 6698 6360 7062 6364
rect 6698 6276 6840 6360
rect 6410 6240 6600 6276
rect 6236 6236 6600 6240
tri 6600 6236 6640 6276 sw
tri 6698 6236 6738 6276 ne
rect 6738 6240 6840 6276
rect 6960 6276 7062 6360
tri 7062 6276 7150 6364 sw
tri 7160 6276 7248 6364 ne
rect 7248 6360 7612 6364
rect 7248 6276 7390 6360
rect 6960 6240 7150 6276
rect 6738 6236 7150 6240
rect 6236 6188 6640 6236
rect 5736 6138 6138 6188
rect 5216 6108 5638 6138
rect 4724 6050 5118 6108
rect 4214 6010 4626 6050
tri 4626 6010 4666 6050 sw
tri 4724 6010 4764 6050 ne
rect 4764 6010 5118 6050
tri 5118 6010 5216 6108 sw
tri 5216 6010 5314 6108 ne
rect 5314 6050 5638 6108
tri 5638 6050 5726 6138 sw
tri 5736 6050 5824 6138 ne
rect 5824 6108 6138 6138
tri 6138 6108 6218 6188 sw
tri 6236 6108 6316 6188 ne
rect 6316 6138 6640 6188
tri 6640 6138 6738 6236 sw
tri 6738 6138 6836 6236 ne
rect 6836 6188 7150 6236
tri 7150 6188 7238 6276 sw
tri 7248 6188 7336 6276 ne
rect 7336 6240 7390 6276
rect 7510 6276 7612 6360
tri 7612 6276 7700 6364 sw
tri 7710 6276 7798 6364 ne
rect 7798 6360 8162 6364
rect 7798 6276 7940 6360
rect 7510 6240 7700 6276
rect 7336 6236 7700 6240
tri 7700 6236 7740 6276 sw
tri 7798 6236 7838 6276 ne
rect 7838 6240 7940 6276
rect 8060 6276 8162 6360
tri 8162 6276 8250 6364 sw
tri 8260 6276 8348 6364 ne
rect 8348 6360 8712 6364
rect 8348 6276 8490 6360
rect 8060 6240 8250 6276
rect 7838 6236 8250 6240
rect 7336 6188 7740 6236
rect 6836 6138 7238 6188
rect 6316 6108 6738 6138
rect 5824 6050 6218 6108
rect 5314 6010 5726 6050
tri 5726 6010 5766 6050 sw
tri 5824 6010 5864 6050 ne
rect 5864 6010 6218 6050
tri 6218 6010 6316 6108 sw
tri 6316 6010 6414 6108 ne
rect 6414 6050 6738 6108
tri 6738 6050 6826 6138 sw
tri 6836 6050 6924 6138 ne
rect 6924 6108 7238 6138
tri 7238 6108 7318 6188 sw
tri 7336 6108 7416 6188 ne
rect 7416 6138 7740 6188
tri 7740 6138 7838 6236 sw
tri 7838 6138 7936 6236 ne
rect 7936 6188 8250 6236
tri 8250 6188 8338 6276 sw
tri 8348 6188 8436 6276 ne
rect 8436 6240 8490 6276
rect 8610 6276 8712 6360
tri 8712 6276 8800 6364 sw
tri 8810 6276 8898 6364 ne
rect 8898 6360 9262 6364
rect 8898 6276 9040 6360
rect 8610 6240 8800 6276
rect 8436 6236 8800 6240
tri 8800 6236 8840 6276 sw
tri 8898 6236 8938 6276 ne
rect 8938 6240 9040 6276
rect 9160 6276 9262 6360
tri 9262 6276 9350 6364 sw
tri 9360 6276 9448 6364 ne
rect 9448 6360 9812 6364
rect 9448 6276 9590 6360
rect 9160 6240 9350 6276
rect 8938 6236 9350 6240
rect 8436 6188 8840 6236
rect 7936 6138 8338 6188
rect 7416 6108 7838 6138
rect 6924 6050 7318 6108
rect 6414 6010 6826 6050
tri 6826 6010 6866 6050 sw
tri 6924 6010 6964 6050 ne
rect 6964 6010 7318 6050
tri 7318 6010 7416 6108 sw
tri 7416 6010 7514 6108 ne
rect 7514 6050 7838 6108
tri 7838 6050 7926 6138 sw
tri 7936 6050 8024 6138 ne
rect 8024 6108 8338 6138
tri 8338 6108 8418 6188 sw
tri 8436 6108 8516 6188 ne
rect 8516 6138 8840 6188
tri 8840 6138 8938 6236 sw
tri 8938 6138 9036 6236 ne
rect 9036 6188 9350 6236
tri 9350 6188 9438 6276 sw
tri 9448 6188 9536 6276 ne
rect 9536 6240 9590 6276
rect 9710 6276 9812 6360
tri 9812 6276 9900 6364 sw
tri 9910 6276 9998 6364 ne
rect 9998 6360 10362 6364
rect 9998 6276 10140 6360
rect 9710 6240 9900 6276
rect 9536 6236 9900 6240
tri 9900 6236 9940 6276 sw
tri 9998 6236 10038 6276 ne
rect 10038 6240 10140 6276
rect 10260 6276 10362 6360
tri 10362 6276 10450 6364 sw
tri 10460 6276 10548 6364 ne
rect 10548 6360 10912 6364
rect 10548 6276 10690 6360
rect 10260 6240 10450 6276
rect 10038 6236 10450 6240
rect 9536 6188 9940 6236
rect 9036 6138 9438 6188
rect 8516 6108 8938 6138
rect 8024 6050 8418 6108
rect 7514 6010 7926 6050
tri 7926 6010 7966 6050 sw
tri 8024 6010 8064 6050 ne
rect 8064 6010 8418 6050
tri 8418 6010 8516 6108 sw
tri 8516 6010 8614 6108 ne
rect 8614 6050 8938 6108
tri 8938 6050 9026 6138 sw
tri 9036 6050 9124 6138 ne
rect 9124 6108 9438 6138
tri 9438 6108 9518 6188 sw
tri 9536 6108 9616 6188 ne
rect 9616 6138 9940 6188
tri 9940 6138 10038 6236 sw
tri 10038 6138 10136 6236 ne
rect 10136 6188 10450 6236
tri 10450 6188 10538 6276 sw
tri 10548 6188 10636 6276 ne
rect 10636 6240 10690 6276
rect 10810 6276 10912 6360
tri 10912 6276 11000 6364 sw
tri 11010 6276 11098 6364 ne
rect 11098 6360 11462 6364
rect 11098 6276 11240 6360
rect 10810 6240 11000 6276
rect 10636 6236 11000 6240
tri 11000 6236 11040 6276 sw
tri 11098 6236 11138 6276 ne
rect 11138 6240 11240 6276
rect 11360 6276 11462 6360
tri 11462 6276 11550 6364 sw
tri 11560 6276 11648 6364 ne
rect 11648 6360 12012 6364
rect 11648 6276 11790 6360
rect 11360 6240 11550 6276
rect 11138 6236 11550 6240
rect 10636 6188 11040 6236
rect 10136 6138 10538 6188
rect 9616 6108 10038 6138
rect 9124 6050 9518 6108
rect 8614 6010 9026 6050
tri 9026 6010 9066 6050 sw
tri 9124 6010 9164 6050 ne
rect 9164 6010 9518 6050
tri 9518 6010 9616 6108 sw
tri 9616 6010 9714 6108 ne
rect 9714 6050 10038 6108
tri 10038 6050 10126 6138 sw
tri 10136 6050 10224 6138 ne
rect 10224 6108 10538 6138
tri 10538 6108 10618 6188 sw
tri 10636 6108 10716 6188 ne
rect 10716 6138 11040 6188
tri 11040 6138 11138 6236 sw
tri 11138 6138 11236 6236 ne
rect 11236 6188 11550 6236
tri 11550 6188 11638 6276 sw
tri 11648 6188 11736 6276 ne
rect 11736 6240 11790 6276
rect 11910 6276 12012 6360
tri 12012 6276 12100 6364 sw
tri 12110 6276 12198 6364 ne
rect 12198 6360 12562 6364
rect 12198 6276 12340 6360
rect 11910 6240 12100 6276
rect 11736 6236 12100 6240
tri 12100 6236 12140 6276 sw
tri 12198 6236 12238 6276 ne
rect 12238 6240 12340 6276
rect 12460 6276 12562 6360
tri 12562 6276 12650 6364 sw
tri 12660 6276 12748 6364 ne
rect 12748 6360 13112 6364
rect 12748 6276 12890 6360
rect 12460 6240 12650 6276
rect 12238 6236 12650 6240
rect 11736 6188 12140 6236
rect 11236 6138 11638 6188
rect 10716 6108 11138 6138
rect 10224 6050 10618 6108
rect 9714 6010 10126 6050
tri 10126 6010 10166 6050 sw
tri 10224 6010 10264 6050 ne
rect 10264 6010 10618 6050
tri 10618 6010 10716 6108 sw
tri 10716 6010 10814 6108 ne
rect 10814 6050 11138 6108
tri 11138 6050 11226 6138 sw
tri 11236 6050 11324 6138 ne
rect 11324 6108 11638 6138
tri 11638 6108 11718 6188 sw
tri 11736 6108 11816 6188 ne
rect 11816 6138 12140 6188
tri 12140 6138 12238 6236 sw
tri 12238 6138 12336 6236 ne
rect 12336 6188 12650 6236
tri 12650 6188 12738 6276 sw
tri 12748 6188 12836 6276 ne
rect 12836 6240 12890 6276
rect 13010 6276 13112 6360
tri 13112 6276 13200 6364 sw
tri 13210 6276 13298 6364 ne
rect 13298 6360 14275 6364
rect 13298 6276 13440 6360
rect 13010 6240 13200 6276
rect 12836 6236 13200 6240
tri 13200 6236 13240 6276 sw
tri 13298 6236 13338 6276 ne
rect 13338 6240 13440 6276
rect 13560 6240 14275 6360
rect 13338 6236 14275 6240
rect 12836 6188 13240 6236
rect 12336 6138 12738 6188
rect 11816 6108 12238 6138
rect 11324 6050 11718 6108
rect 10814 6010 11226 6050
tri 11226 6010 11266 6050 sw
tri 11324 6010 11364 6050 ne
rect 11364 6010 11718 6050
tri 11718 6010 11816 6108 sw
tri 11816 6010 11914 6108 ne
rect 11914 6050 12238 6108
tri 12238 6050 12326 6138 sw
tri 12336 6050 12424 6138 ne
rect 12424 6108 12738 6138
tri 12738 6108 12818 6188 sw
tri 12836 6108 12916 6188 ne
rect 12916 6138 13240 6188
tri 13240 6138 13338 6236 sw
tri 13338 6138 13436 6236 ne
rect 13436 6138 14275 6236
rect 12916 6108 13338 6138
rect 12424 6050 12818 6108
rect 11914 6010 12326 6050
tri 12326 6010 12366 6050 sw
tri 12424 6010 12464 6050 ne
rect 12464 6010 12818 6050
tri 12818 6010 12916 6108 sw
tri 12916 6010 13014 6108 ne
rect 13014 6050 13338 6108
tri 13338 6050 13426 6138 sw
tri 13436 6050 13524 6138 ne
rect 13524 6050 14275 6138
rect 13014 6010 13426 6050
tri 13426 6010 13466 6050 sw
tri 13524 6010 13564 6050 ne
rect 13564 6010 14275 6050
rect -2525 5912 -284 6010
tri -284 5912 -186 6010 sw
tri -186 5912 -88 6010 ne
rect -88 5912 266 6010
tri 266 5912 364 6010 sw
tri 364 5912 462 6010 ne
rect 462 5912 816 6010
tri 816 5912 914 6010 sw
tri 914 5912 1012 6010 ne
rect 1012 5912 1366 6010
tri 1366 5912 1464 6010 sw
tri 1464 5912 1562 6010 ne
rect 1562 5912 1916 6010
tri 1916 5912 2014 6010 sw
tri 2014 5912 2112 6010 ne
rect 2112 5912 2466 6010
tri 2466 5912 2564 6010 sw
tri 2564 5912 2662 6010 ne
rect 2662 5912 3016 6010
tri 3016 5912 3114 6010 sw
tri 3114 5912 3212 6010 ne
rect 3212 5912 3566 6010
tri 3566 5912 3664 6010 sw
tri 3664 5912 3762 6010 ne
rect 3762 5912 4116 6010
tri 4116 5912 4214 6010 sw
tri 4214 5912 4312 6010 ne
rect 4312 5912 4666 6010
tri 4666 5912 4764 6010 sw
tri 4764 5912 4862 6010 ne
rect 4862 5912 5216 6010
tri 5216 5912 5314 6010 sw
tri 5314 5912 5412 6010 ne
rect 5412 5912 5766 6010
tri 5766 5912 5864 6010 sw
tri 5864 5912 5962 6010 ne
rect 5962 5912 6316 6010
tri 6316 5912 6414 6010 sw
tri 6414 5912 6512 6010 ne
rect 6512 5912 6866 6010
tri 6866 5912 6964 6010 sw
tri 6964 5912 7062 6010 ne
rect 7062 5912 7416 6010
tri 7416 5912 7514 6010 sw
tri 7514 5912 7612 6010 ne
rect 7612 5912 7966 6010
tri 7966 5912 8064 6010 sw
tri 8064 5912 8162 6010 ne
rect 8162 5912 8516 6010
tri 8516 5912 8614 6010 sw
tri 8614 5912 8712 6010 ne
rect 8712 5912 9066 6010
tri 9066 5912 9164 6010 sw
tri 9164 5912 9262 6010 ne
rect 9262 5912 9616 6010
tri 9616 5912 9714 6010 sw
tri 9714 5912 9812 6010 ne
rect 9812 5912 10166 6010
tri 10166 5912 10264 6010 sw
tri 10264 5912 10362 6010 ne
rect 10362 5912 10716 6010
tri 10716 5912 10814 6010 sw
tri 10814 5912 10912 6010 ne
rect 10912 5912 11266 6010
tri 11266 5912 11364 6010 sw
tri 11364 5912 11462 6010 ne
rect 11462 5912 11816 6010
tri 11816 5912 11914 6010 sw
tri 11914 5912 12012 6010 ne
rect 12012 5912 12366 6010
tri 12366 5912 12464 6010 sw
tri 12464 5912 12562 6010 ne
rect 12562 5912 12916 6010
tri 12916 5912 13014 6010 sw
tri 13014 5912 13112 6010 ne
rect 13112 5912 13466 6010
tri 13466 5912 13564 6010 sw
tri 13564 5912 13662 6010 ne
rect 13662 5912 14275 6010
rect -2525 5814 -186 5912
tri -186 5814 -88 5912 sw
tri -88 5814 10 5912 ne
rect 10 5814 364 5912
tri 364 5814 462 5912 sw
tri 462 5814 560 5912 ne
rect 560 5814 914 5912
tri 914 5814 1012 5912 sw
tri 1012 5814 1110 5912 ne
rect 1110 5814 1464 5912
tri 1464 5814 1562 5912 sw
tri 1562 5814 1660 5912 ne
rect 1660 5814 2014 5912
tri 2014 5814 2112 5912 sw
tri 2112 5814 2210 5912 ne
rect 2210 5814 2564 5912
tri 2564 5814 2662 5912 sw
tri 2662 5814 2760 5912 ne
rect 2760 5814 3114 5912
tri 3114 5814 3212 5912 sw
tri 3212 5814 3310 5912 ne
rect 3310 5814 3664 5912
tri 3664 5814 3762 5912 sw
tri 3762 5814 3860 5912 ne
rect 3860 5814 4214 5912
tri 4214 5814 4312 5912 sw
tri 4312 5814 4410 5912 ne
rect 4410 5814 4764 5912
tri 4764 5814 4862 5912 sw
tri 4862 5814 4960 5912 ne
rect 4960 5814 5314 5912
tri 5314 5814 5412 5912 sw
tri 5412 5814 5510 5912 ne
rect 5510 5814 5864 5912
tri 5864 5814 5962 5912 sw
tri 5962 5814 6060 5912 ne
rect 6060 5814 6414 5912
tri 6414 5814 6512 5912 sw
tri 6512 5814 6610 5912 ne
rect 6610 5814 6964 5912
tri 6964 5814 7062 5912 sw
tri 7062 5814 7160 5912 ne
rect 7160 5814 7514 5912
tri 7514 5814 7612 5912 sw
tri 7612 5814 7710 5912 ne
rect 7710 5814 8064 5912
tri 8064 5814 8162 5912 sw
tri 8162 5814 8260 5912 ne
rect 8260 5814 8614 5912
tri 8614 5814 8712 5912 sw
tri 8712 5814 8810 5912 ne
rect 8810 5814 9164 5912
tri 9164 5814 9262 5912 sw
tri 9262 5814 9360 5912 ne
rect 9360 5814 9714 5912
tri 9714 5814 9812 5912 sw
tri 9812 5814 9910 5912 ne
rect 9910 5814 10264 5912
tri 10264 5814 10362 5912 sw
tri 10362 5814 10460 5912 ne
rect 10460 5814 10814 5912
tri 10814 5814 10912 5912 sw
tri 10912 5814 11010 5912 ne
rect 11010 5814 11364 5912
tri 11364 5814 11462 5912 sw
tri 11462 5814 11560 5912 ne
rect 11560 5814 11914 5912
tri 11914 5814 12012 5912 sw
tri 12012 5814 12110 5912 ne
rect 12110 5814 12464 5912
tri 12464 5814 12562 5912 sw
tri 12562 5814 12660 5912 ne
rect 12660 5814 13014 5912
tri 13014 5814 13112 5912 sw
tri 13112 5814 13210 5912 ne
rect 13210 5814 13564 5912
tri 13564 5814 13662 5912 sw
rect 14775 5814 15775 6462
rect -2525 5810 -88 5814
rect -2525 5690 -310 5810
rect -190 5726 -88 5810
tri -88 5726 0 5814 sw
tri 10 5726 98 5814 ne
rect 98 5810 462 5814
rect 98 5726 240 5810
rect -190 5690 0 5726
rect -2525 5686 0 5690
rect -2525 5038 -1525 5686
tri -412 5588 -314 5686 ne
rect -314 5638 0 5686
tri 0 5638 88 5726 sw
tri 98 5638 186 5726 ne
rect 186 5690 240 5726
rect 360 5726 462 5810
tri 462 5726 550 5814 sw
tri 560 5726 648 5814 ne
rect 648 5810 1012 5814
rect 648 5726 790 5810
rect 360 5690 550 5726
rect 186 5686 550 5690
tri 550 5686 590 5726 sw
tri 648 5686 688 5726 ne
rect 688 5690 790 5726
rect 910 5726 1012 5810
tri 1012 5726 1100 5814 sw
tri 1110 5726 1198 5814 ne
rect 1198 5810 1562 5814
rect 1198 5726 1340 5810
rect 910 5690 1100 5726
rect 688 5686 1100 5690
rect 186 5638 590 5686
rect -314 5588 88 5638
rect -1025 5500 -412 5588
tri -412 5500 -324 5588 sw
tri -314 5500 -226 5588 ne
rect -226 5558 88 5588
tri 88 5558 168 5638 sw
tri 186 5558 266 5638 ne
rect 266 5588 590 5638
tri 590 5588 688 5686 sw
tri 688 5588 786 5686 ne
rect 786 5638 1100 5686
tri 1100 5638 1188 5726 sw
tri 1198 5638 1286 5726 ne
rect 1286 5690 1340 5726
rect 1460 5726 1562 5810
tri 1562 5726 1650 5814 sw
tri 1660 5726 1748 5814 ne
rect 1748 5810 2112 5814
rect 1748 5726 1890 5810
rect 1460 5690 1650 5726
rect 1286 5686 1650 5690
tri 1650 5686 1690 5726 sw
tri 1748 5686 1788 5726 ne
rect 1788 5690 1890 5726
rect 2010 5726 2112 5810
tri 2112 5726 2200 5814 sw
tri 2210 5726 2298 5814 ne
rect 2298 5810 2662 5814
rect 2298 5726 2440 5810
rect 2010 5690 2200 5726
rect 1788 5686 2200 5690
rect 1286 5638 1690 5686
rect 786 5588 1188 5638
rect 266 5558 688 5588
rect -226 5500 168 5558
rect -1025 5460 -324 5500
tri -324 5460 -284 5500 sw
tri -226 5460 -186 5500 ne
rect -186 5460 168 5500
tri 168 5460 266 5558 sw
tri 266 5460 364 5558 ne
rect 364 5500 688 5558
tri 688 5500 776 5588 sw
tri 786 5500 874 5588 ne
rect 874 5558 1188 5588
tri 1188 5558 1268 5638 sw
tri 1286 5558 1366 5638 ne
rect 1366 5588 1690 5638
tri 1690 5588 1788 5686 sw
tri 1788 5588 1886 5686 ne
rect 1886 5638 2200 5686
tri 2200 5638 2288 5726 sw
tri 2298 5638 2386 5726 ne
rect 2386 5690 2440 5726
rect 2560 5726 2662 5810
tri 2662 5726 2750 5814 sw
tri 2760 5726 2848 5814 ne
rect 2848 5810 3212 5814
rect 2848 5726 2990 5810
rect 2560 5690 2750 5726
rect 2386 5686 2750 5690
tri 2750 5686 2790 5726 sw
tri 2848 5686 2888 5726 ne
rect 2888 5690 2990 5726
rect 3110 5726 3212 5810
tri 3212 5726 3300 5814 sw
tri 3310 5726 3398 5814 ne
rect 3398 5810 3762 5814
rect 3398 5726 3540 5810
rect 3110 5690 3300 5726
rect 2888 5686 3300 5690
rect 2386 5638 2790 5686
rect 1886 5588 2288 5638
rect 1366 5558 1788 5588
rect 874 5500 1268 5558
rect 364 5460 776 5500
tri 776 5460 816 5500 sw
tri 874 5460 914 5500 ne
rect 914 5460 1268 5500
tri 1268 5460 1366 5558 sw
tri 1366 5460 1464 5558 ne
rect 1464 5500 1788 5558
tri 1788 5500 1876 5588 sw
tri 1886 5500 1974 5588 ne
rect 1974 5558 2288 5588
tri 2288 5558 2368 5638 sw
tri 2386 5558 2466 5638 ne
rect 2466 5588 2790 5638
tri 2790 5588 2888 5686 sw
tri 2888 5588 2986 5686 ne
rect 2986 5638 3300 5686
tri 3300 5638 3388 5726 sw
tri 3398 5638 3486 5726 ne
rect 3486 5690 3540 5726
rect 3660 5726 3762 5810
tri 3762 5726 3850 5814 sw
tri 3860 5726 3948 5814 ne
rect 3948 5810 4312 5814
rect 3948 5726 4090 5810
rect 3660 5690 3850 5726
rect 3486 5686 3850 5690
tri 3850 5686 3890 5726 sw
tri 3948 5686 3988 5726 ne
rect 3988 5690 4090 5726
rect 4210 5726 4312 5810
tri 4312 5726 4400 5814 sw
tri 4410 5726 4498 5814 ne
rect 4498 5810 4862 5814
rect 4498 5726 4640 5810
rect 4210 5690 4400 5726
rect 3988 5686 4400 5690
rect 3486 5638 3890 5686
rect 2986 5588 3388 5638
rect 2466 5558 2888 5588
rect 1974 5500 2368 5558
rect 1464 5460 1876 5500
tri 1876 5460 1916 5500 sw
tri 1974 5460 2014 5500 ne
rect 2014 5460 2368 5500
tri 2368 5460 2466 5558 sw
tri 2466 5460 2564 5558 ne
rect 2564 5500 2888 5558
tri 2888 5500 2976 5588 sw
tri 2986 5500 3074 5588 ne
rect 3074 5558 3388 5588
tri 3388 5558 3468 5638 sw
tri 3486 5558 3566 5638 ne
rect 3566 5588 3890 5638
tri 3890 5588 3988 5686 sw
tri 3988 5588 4086 5686 ne
rect 4086 5638 4400 5686
tri 4400 5638 4488 5726 sw
tri 4498 5638 4586 5726 ne
rect 4586 5690 4640 5726
rect 4760 5726 4862 5810
tri 4862 5726 4950 5814 sw
tri 4960 5726 5048 5814 ne
rect 5048 5810 5412 5814
rect 5048 5726 5190 5810
rect 4760 5690 4950 5726
rect 4586 5686 4950 5690
tri 4950 5686 4990 5726 sw
tri 5048 5686 5088 5726 ne
rect 5088 5690 5190 5726
rect 5310 5726 5412 5810
tri 5412 5726 5500 5814 sw
tri 5510 5726 5598 5814 ne
rect 5598 5810 5962 5814
rect 5598 5726 5740 5810
rect 5310 5690 5500 5726
rect 5088 5686 5500 5690
rect 4586 5638 4990 5686
rect 4086 5588 4488 5638
rect 3566 5558 3988 5588
rect 3074 5500 3468 5558
rect 2564 5460 2976 5500
tri 2976 5460 3016 5500 sw
tri 3074 5460 3114 5500 ne
rect 3114 5460 3468 5500
tri 3468 5460 3566 5558 sw
tri 3566 5460 3664 5558 ne
rect 3664 5500 3988 5558
tri 3988 5500 4076 5588 sw
tri 4086 5500 4174 5588 ne
rect 4174 5558 4488 5588
tri 4488 5558 4568 5638 sw
tri 4586 5558 4666 5638 ne
rect 4666 5588 4990 5638
tri 4990 5588 5088 5686 sw
tri 5088 5588 5186 5686 ne
rect 5186 5638 5500 5686
tri 5500 5638 5588 5726 sw
tri 5598 5638 5686 5726 ne
rect 5686 5690 5740 5726
rect 5860 5726 5962 5810
tri 5962 5726 6050 5814 sw
tri 6060 5726 6148 5814 ne
rect 6148 5810 6512 5814
rect 6148 5726 6290 5810
rect 5860 5690 6050 5726
rect 5686 5686 6050 5690
tri 6050 5686 6090 5726 sw
tri 6148 5686 6188 5726 ne
rect 6188 5690 6290 5726
rect 6410 5726 6512 5810
tri 6512 5726 6600 5814 sw
tri 6610 5726 6698 5814 ne
rect 6698 5810 7062 5814
rect 6698 5726 6840 5810
rect 6410 5690 6600 5726
rect 6188 5686 6600 5690
rect 5686 5638 6090 5686
rect 5186 5588 5588 5638
rect 4666 5558 5088 5588
rect 4174 5500 4568 5558
rect 3664 5460 4076 5500
tri 4076 5460 4116 5500 sw
tri 4174 5460 4214 5500 ne
rect 4214 5460 4568 5500
tri 4568 5460 4666 5558 sw
tri 4666 5460 4764 5558 ne
rect 4764 5500 5088 5558
tri 5088 5500 5176 5588 sw
tri 5186 5500 5274 5588 ne
rect 5274 5558 5588 5588
tri 5588 5558 5668 5638 sw
tri 5686 5558 5766 5638 ne
rect 5766 5588 6090 5638
tri 6090 5588 6188 5686 sw
tri 6188 5588 6286 5686 ne
rect 6286 5638 6600 5686
tri 6600 5638 6688 5726 sw
tri 6698 5638 6786 5726 ne
rect 6786 5690 6840 5726
rect 6960 5726 7062 5810
tri 7062 5726 7150 5814 sw
tri 7160 5726 7248 5814 ne
rect 7248 5810 7612 5814
rect 7248 5726 7390 5810
rect 6960 5690 7150 5726
rect 6786 5686 7150 5690
tri 7150 5686 7190 5726 sw
tri 7248 5686 7288 5726 ne
rect 7288 5690 7390 5726
rect 7510 5726 7612 5810
tri 7612 5726 7700 5814 sw
tri 7710 5726 7798 5814 ne
rect 7798 5810 8162 5814
rect 7798 5726 7940 5810
rect 7510 5690 7700 5726
rect 7288 5686 7700 5690
rect 6786 5638 7190 5686
rect 6286 5588 6688 5638
rect 5766 5558 6188 5588
rect 5274 5500 5668 5558
rect 4764 5460 5176 5500
tri 5176 5460 5216 5500 sw
tri 5274 5460 5314 5500 ne
rect 5314 5460 5668 5500
tri 5668 5460 5766 5558 sw
tri 5766 5460 5864 5558 ne
rect 5864 5500 6188 5558
tri 6188 5500 6276 5588 sw
tri 6286 5500 6374 5588 ne
rect 6374 5558 6688 5588
tri 6688 5558 6768 5638 sw
tri 6786 5558 6866 5638 ne
rect 6866 5588 7190 5638
tri 7190 5588 7288 5686 sw
tri 7288 5588 7386 5686 ne
rect 7386 5638 7700 5686
tri 7700 5638 7788 5726 sw
tri 7798 5638 7886 5726 ne
rect 7886 5690 7940 5726
rect 8060 5726 8162 5810
tri 8162 5726 8250 5814 sw
tri 8260 5726 8348 5814 ne
rect 8348 5810 8712 5814
rect 8348 5726 8490 5810
rect 8060 5690 8250 5726
rect 7886 5686 8250 5690
tri 8250 5686 8290 5726 sw
tri 8348 5686 8388 5726 ne
rect 8388 5690 8490 5726
rect 8610 5726 8712 5810
tri 8712 5726 8800 5814 sw
tri 8810 5726 8898 5814 ne
rect 8898 5810 9262 5814
rect 8898 5726 9040 5810
rect 8610 5690 8800 5726
rect 8388 5686 8800 5690
rect 7886 5638 8290 5686
rect 7386 5588 7788 5638
rect 6866 5558 7288 5588
rect 6374 5500 6768 5558
rect 5864 5460 6276 5500
tri 6276 5460 6316 5500 sw
tri 6374 5460 6414 5500 ne
rect 6414 5460 6768 5500
tri 6768 5460 6866 5558 sw
tri 6866 5460 6964 5558 ne
rect 6964 5500 7288 5558
tri 7288 5500 7376 5588 sw
tri 7386 5500 7474 5588 ne
rect 7474 5558 7788 5588
tri 7788 5558 7868 5638 sw
tri 7886 5558 7966 5638 ne
rect 7966 5588 8290 5638
tri 8290 5588 8388 5686 sw
tri 8388 5588 8486 5686 ne
rect 8486 5638 8800 5686
tri 8800 5638 8888 5726 sw
tri 8898 5638 8986 5726 ne
rect 8986 5690 9040 5726
rect 9160 5726 9262 5810
tri 9262 5726 9350 5814 sw
tri 9360 5726 9448 5814 ne
rect 9448 5810 9812 5814
rect 9448 5726 9590 5810
rect 9160 5690 9350 5726
rect 8986 5686 9350 5690
tri 9350 5686 9390 5726 sw
tri 9448 5686 9488 5726 ne
rect 9488 5690 9590 5726
rect 9710 5726 9812 5810
tri 9812 5726 9900 5814 sw
tri 9910 5726 9998 5814 ne
rect 9998 5810 10362 5814
rect 9998 5726 10140 5810
rect 9710 5690 9900 5726
rect 9488 5686 9900 5690
rect 8986 5638 9390 5686
rect 8486 5588 8888 5638
rect 7966 5558 8388 5588
rect 7474 5500 7868 5558
rect 6964 5460 7376 5500
tri 7376 5460 7416 5500 sw
tri 7474 5460 7514 5500 ne
rect 7514 5460 7868 5500
tri 7868 5460 7966 5558 sw
tri 7966 5460 8064 5558 ne
rect 8064 5500 8388 5558
tri 8388 5500 8476 5588 sw
tri 8486 5500 8574 5588 ne
rect 8574 5558 8888 5588
tri 8888 5558 8968 5638 sw
tri 8986 5558 9066 5638 ne
rect 9066 5588 9390 5638
tri 9390 5588 9488 5686 sw
tri 9488 5588 9586 5686 ne
rect 9586 5638 9900 5686
tri 9900 5638 9988 5726 sw
tri 9998 5638 10086 5726 ne
rect 10086 5690 10140 5726
rect 10260 5726 10362 5810
tri 10362 5726 10450 5814 sw
tri 10460 5726 10548 5814 ne
rect 10548 5810 10912 5814
rect 10548 5726 10690 5810
rect 10260 5690 10450 5726
rect 10086 5686 10450 5690
tri 10450 5686 10490 5726 sw
tri 10548 5686 10588 5726 ne
rect 10588 5690 10690 5726
rect 10810 5726 10912 5810
tri 10912 5726 11000 5814 sw
tri 11010 5726 11098 5814 ne
rect 11098 5810 11462 5814
rect 11098 5726 11240 5810
rect 10810 5690 11000 5726
rect 10588 5686 11000 5690
rect 10086 5638 10490 5686
rect 9586 5588 9988 5638
rect 9066 5558 9488 5588
rect 8574 5500 8968 5558
rect 8064 5460 8476 5500
tri 8476 5460 8516 5500 sw
tri 8574 5460 8614 5500 ne
rect 8614 5460 8968 5500
tri 8968 5460 9066 5558 sw
tri 9066 5460 9164 5558 ne
rect 9164 5500 9488 5558
tri 9488 5500 9576 5588 sw
tri 9586 5500 9674 5588 ne
rect 9674 5558 9988 5588
tri 9988 5558 10068 5638 sw
tri 10086 5558 10166 5638 ne
rect 10166 5588 10490 5638
tri 10490 5588 10588 5686 sw
tri 10588 5588 10686 5686 ne
rect 10686 5638 11000 5686
tri 11000 5638 11088 5726 sw
tri 11098 5638 11186 5726 ne
rect 11186 5690 11240 5726
rect 11360 5726 11462 5810
tri 11462 5726 11550 5814 sw
tri 11560 5726 11648 5814 ne
rect 11648 5810 12012 5814
rect 11648 5726 11790 5810
rect 11360 5690 11550 5726
rect 11186 5686 11550 5690
tri 11550 5686 11590 5726 sw
tri 11648 5686 11688 5726 ne
rect 11688 5690 11790 5726
rect 11910 5726 12012 5810
tri 12012 5726 12100 5814 sw
tri 12110 5726 12198 5814 ne
rect 12198 5810 12562 5814
rect 12198 5726 12340 5810
rect 11910 5690 12100 5726
rect 11688 5686 12100 5690
rect 11186 5638 11590 5686
rect 10686 5588 11088 5638
rect 10166 5558 10588 5588
rect 9674 5500 10068 5558
rect 9164 5460 9576 5500
tri 9576 5460 9616 5500 sw
tri 9674 5460 9714 5500 ne
rect 9714 5460 10068 5500
tri 10068 5460 10166 5558 sw
tri 10166 5460 10264 5558 ne
rect 10264 5500 10588 5558
tri 10588 5500 10676 5588 sw
tri 10686 5500 10774 5588 ne
rect 10774 5558 11088 5588
tri 11088 5558 11168 5638 sw
tri 11186 5558 11266 5638 ne
rect 11266 5588 11590 5638
tri 11590 5588 11688 5686 sw
tri 11688 5588 11786 5686 ne
rect 11786 5638 12100 5686
tri 12100 5638 12188 5726 sw
tri 12198 5638 12286 5726 ne
rect 12286 5690 12340 5726
rect 12460 5726 12562 5810
tri 12562 5726 12650 5814 sw
tri 12660 5726 12748 5814 ne
rect 12748 5810 13112 5814
rect 12748 5726 12890 5810
rect 12460 5690 12650 5726
rect 12286 5686 12650 5690
tri 12650 5686 12690 5726 sw
tri 12748 5686 12788 5726 ne
rect 12788 5690 12890 5726
rect 13010 5726 13112 5810
tri 13112 5726 13200 5814 sw
tri 13210 5726 13298 5814 ne
rect 13298 5810 15775 5814
rect 13298 5726 13440 5810
rect 13010 5690 13200 5726
rect 12788 5686 13200 5690
rect 12286 5638 12690 5686
rect 11786 5588 12188 5638
rect 11266 5558 11688 5588
rect 10774 5500 11168 5558
rect 10264 5460 10676 5500
tri 10676 5460 10716 5500 sw
tri 10774 5460 10814 5500 ne
rect 10814 5460 11168 5500
tri 11168 5460 11266 5558 sw
tri 11266 5460 11364 5558 ne
rect 11364 5500 11688 5558
tri 11688 5500 11776 5588 sw
tri 11786 5500 11874 5588 ne
rect 11874 5558 12188 5588
tri 12188 5558 12268 5638 sw
tri 12286 5558 12366 5638 ne
rect 12366 5588 12690 5638
tri 12690 5588 12788 5686 sw
tri 12788 5588 12886 5686 ne
rect 12886 5638 13200 5686
tri 13200 5638 13288 5726 sw
tri 13298 5638 13386 5726 ne
rect 13386 5690 13440 5726
rect 13560 5690 15775 5810
rect 13386 5638 15775 5690
rect 12886 5588 13288 5638
rect 12366 5558 12788 5588
rect 11874 5500 12268 5558
rect 11364 5460 11776 5500
tri 11776 5460 11816 5500 sw
tri 11874 5460 11914 5500 ne
rect 11914 5460 12268 5500
tri 12268 5460 12366 5558 sw
tri 12366 5460 12464 5558 ne
rect 12464 5500 12788 5558
tri 12788 5500 12876 5588 sw
tri 12886 5500 12974 5588 ne
rect 12974 5558 13288 5588
tri 13288 5558 13368 5638 sw
tri 13386 5558 13466 5638 ne
rect 13466 5558 14075 5638
rect 12974 5500 13368 5558
rect 12464 5460 12876 5500
tri 12876 5460 12916 5500 sw
tri 12974 5460 13014 5500 ne
rect 13014 5460 13368 5500
tri 13368 5460 13466 5558 sw
tri 13466 5460 13564 5558 ne
rect 13564 5538 14075 5558
rect 14175 5538 15775 5638
rect 13564 5460 15775 5538
rect -1025 5412 -284 5460
rect -1025 5312 -925 5412
rect -825 5362 -284 5412
tri -284 5362 -186 5460 sw
tri -186 5362 -88 5460 ne
rect -88 5362 266 5460
tri 266 5362 364 5460 sw
tri 364 5362 462 5460 ne
rect 462 5362 816 5460
tri 816 5362 914 5460 sw
tri 914 5362 1012 5460 ne
rect 1012 5362 1366 5460
tri 1366 5362 1464 5460 sw
tri 1464 5362 1562 5460 ne
rect 1562 5362 1916 5460
tri 1916 5362 2014 5460 sw
tri 2014 5362 2112 5460 ne
rect 2112 5362 2466 5460
tri 2466 5362 2564 5460 sw
tri 2564 5362 2662 5460 ne
rect 2662 5362 3016 5460
tri 3016 5362 3114 5460 sw
tri 3114 5362 3212 5460 ne
rect 3212 5362 3566 5460
tri 3566 5362 3664 5460 sw
tri 3664 5362 3762 5460 ne
rect 3762 5362 4116 5460
tri 4116 5362 4214 5460 sw
tri 4214 5362 4312 5460 ne
rect 4312 5362 4666 5460
tri 4666 5362 4764 5460 sw
tri 4764 5362 4862 5460 ne
rect 4862 5362 5216 5460
tri 5216 5362 5314 5460 sw
tri 5314 5362 5412 5460 ne
rect 5412 5362 5766 5460
tri 5766 5362 5864 5460 sw
tri 5864 5362 5962 5460 ne
rect 5962 5362 6316 5460
tri 6316 5362 6414 5460 sw
tri 6414 5362 6512 5460 ne
rect 6512 5362 6866 5460
tri 6866 5362 6964 5460 sw
tri 6964 5362 7062 5460 ne
rect 7062 5362 7416 5460
tri 7416 5362 7514 5460 sw
tri 7514 5362 7612 5460 ne
rect 7612 5362 7966 5460
tri 7966 5362 8064 5460 sw
tri 8064 5362 8162 5460 ne
rect 8162 5362 8516 5460
tri 8516 5362 8614 5460 sw
tri 8614 5362 8712 5460 ne
rect 8712 5362 9066 5460
tri 9066 5362 9164 5460 sw
tri 9164 5362 9262 5460 ne
rect 9262 5362 9616 5460
tri 9616 5362 9714 5460 sw
tri 9714 5362 9812 5460 ne
rect 9812 5362 10166 5460
tri 10166 5362 10264 5460 sw
tri 10264 5362 10362 5460 ne
rect 10362 5362 10716 5460
tri 10716 5362 10814 5460 sw
tri 10814 5362 10912 5460 ne
rect 10912 5362 11266 5460
tri 11266 5362 11364 5460 sw
tri 11364 5362 11462 5460 ne
rect 11462 5362 11816 5460
tri 11816 5362 11914 5460 sw
tri 11914 5362 12012 5460 ne
rect 12012 5362 12366 5460
tri 12366 5362 12464 5460 sw
tri 12464 5362 12562 5460 ne
rect 12562 5362 12916 5460
tri 12916 5362 13014 5460 sw
tri 13014 5362 13112 5460 ne
rect 13112 5362 13466 5460
tri 13466 5362 13564 5460 sw
tri 13564 5362 13662 5460 ne
rect 13662 5362 15775 5460
rect -825 5312 -186 5362
rect -1025 5264 -186 5312
tri -186 5264 -88 5362 sw
tri -88 5264 10 5362 ne
rect 10 5264 364 5362
tri 364 5264 462 5362 sw
tri 462 5264 560 5362 ne
rect 560 5264 914 5362
tri 914 5264 1012 5362 sw
tri 1012 5264 1110 5362 ne
rect 1110 5264 1464 5362
tri 1464 5264 1562 5362 sw
tri 1562 5264 1660 5362 ne
rect 1660 5264 2014 5362
tri 2014 5264 2112 5362 sw
tri 2112 5264 2210 5362 ne
rect 2210 5264 2564 5362
tri 2564 5264 2662 5362 sw
tri 2662 5264 2760 5362 ne
rect 2760 5264 3114 5362
tri 3114 5264 3212 5362 sw
tri 3212 5264 3310 5362 ne
rect 3310 5264 3664 5362
tri 3664 5264 3762 5362 sw
tri 3762 5264 3860 5362 ne
rect 3860 5264 4214 5362
tri 4214 5264 4312 5362 sw
tri 4312 5264 4410 5362 ne
rect 4410 5264 4764 5362
tri 4764 5264 4862 5362 sw
tri 4862 5264 4960 5362 ne
rect 4960 5264 5314 5362
tri 5314 5264 5412 5362 sw
tri 5412 5264 5510 5362 ne
rect 5510 5264 5864 5362
tri 5864 5264 5962 5362 sw
tri 5962 5264 6060 5362 ne
rect 6060 5264 6414 5362
tri 6414 5264 6512 5362 sw
tri 6512 5264 6610 5362 ne
rect 6610 5264 6964 5362
tri 6964 5264 7062 5362 sw
tri 7062 5264 7160 5362 ne
rect 7160 5264 7514 5362
tri 7514 5264 7612 5362 sw
tri 7612 5264 7710 5362 ne
rect 7710 5264 8064 5362
tri 8064 5264 8162 5362 sw
tri 8162 5264 8260 5362 ne
rect 8260 5264 8614 5362
tri 8614 5264 8712 5362 sw
tri 8712 5264 8810 5362 ne
rect 8810 5264 9164 5362
tri 9164 5264 9262 5362 sw
tri 9262 5264 9360 5362 ne
rect 9360 5264 9714 5362
tri 9714 5264 9812 5362 sw
tri 9812 5264 9910 5362 ne
rect 9910 5264 10264 5362
tri 10264 5264 10362 5362 sw
tri 10362 5264 10460 5362 ne
rect 10460 5264 10814 5362
tri 10814 5264 10912 5362 sw
tri 10912 5264 11010 5362 ne
rect 11010 5264 11364 5362
tri 11364 5264 11462 5362 sw
tri 11462 5264 11560 5362 ne
rect 11560 5264 11914 5362
tri 11914 5264 12012 5362 sw
tri 12012 5264 12110 5362 ne
rect 12110 5264 12464 5362
tri 12464 5264 12562 5362 sw
tri 12562 5264 12660 5362 ne
rect 12660 5264 13014 5362
tri 13014 5264 13112 5362 sw
tri 13112 5264 13210 5362 ne
rect 13210 5264 13564 5362
tri 13564 5264 13662 5362 sw
rect -1025 5260 -88 5264
rect -1025 5140 -310 5260
rect -190 5176 -88 5260
tri -88 5176 0 5264 sw
tri 10 5176 98 5264 ne
rect 98 5260 462 5264
rect 98 5176 240 5260
rect -190 5140 0 5176
rect -1025 5136 0 5140
tri 0 5136 40 5176 sw
tri 98 5136 138 5176 ne
rect 138 5140 240 5176
rect 360 5176 462 5260
tri 462 5176 550 5264 sw
tri 560 5176 648 5264 ne
rect 648 5260 1012 5264
rect 648 5176 790 5260
rect 360 5140 550 5176
rect 138 5136 550 5140
tri -412 5038 -314 5136 ne
rect -314 5038 40 5136
tri 40 5038 138 5136 sw
tri 138 5038 236 5136 ne
rect 236 5088 550 5136
tri 550 5088 638 5176 sw
tri 648 5088 736 5176 ne
rect 736 5140 790 5176
rect 910 5176 1012 5260
tri 1012 5176 1100 5264 sw
tri 1110 5176 1198 5264 ne
rect 1198 5260 1562 5264
rect 1198 5176 1340 5260
rect 910 5140 1100 5176
rect 736 5136 1100 5140
tri 1100 5136 1140 5176 sw
tri 1198 5136 1238 5176 ne
rect 1238 5140 1340 5176
rect 1460 5176 1562 5260
tri 1562 5176 1650 5264 sw
tri 1660 5176 1748 5264 ne
rect 1748 5260 2112 5264
rect 1748 5176 1890 5260
rect 1460 5140 1650 5176
rect 1238 5136 1650 5140
rect 736 5088 1140 5136
rect 236 5038 638 5088
rect -2525 4950 -412 5038
tri -412 4950 -324 5038 sw
tri -314 4950 -226 5038 ne
rect -226 4950 138 5038
tri 138 4950 226 5038 sw
tri 236 4950 324 5038 ne
rect 324 5008 638 5038
tri 638 5008 718 5088 sw
tri 736 5008 816 5088 ne
rect 816 5038 1140 5088
tri 1140 5038 1238 5136 sw
tri 1238 5038 1336 5136 ne
rect 1336 5088 1650 5136
tri 1650 5088 1738 5176 sw
tri 1748 5088 1836 5176 ne
rect 1836 5140 1890 5176
rect 2010 5176 2112 5260
tri 2112 5176 2200 5264 sw
tri 2210 5176 2298 5264 ne
rect 2298 5260 2662 5264
rect 2298 5176 2440 5260
rect 2010 5140 2200 5176
rect 1836 5136 2200 5140
tri 2200 5136 2240 5176 sw
tri 2298 5136 2338 5176 ne
rect 2338 5140 2440 5176
rect 2560 5176 2662 5260
tri 2662 5176 2750 5264 sw
tri 2760 5176 2848 5264 ne
rect 2848 5260 3212 5264
rect 2848 5176 2990 5260
rect 2560 5140 2750 5176
rect 2338 5136 2750 5140
rect 1836 5088 2240 5136
rect 1336 5038 1738 5088
rect 816 5008 1238 5038
rect 324 4950 718 5008
rect -2525 4910 -324 4950
tri -324 4910 -284 4950 sw
tri -226 4910 -186 4950 ne
rect -186 4910 226 4950
tri 226 4910 266 4950 sw
tri 324 4910 364 4950 ne
rect 364 4910 718 4950
tri 718 4910 816 5008 sw
tri 816 4910 914 5008 ne
rect 914 4950 1238 5008
tri 1238 4950 1326 5038 sw
tri 1336 4950 1424 5038 ne
rect 1424 5008 1738 5038
tri 1738 5008 1818 5088 sw
tri 1836 5008 1916 5088 ne
rect 1916 5038 2240 5088
tri 2240 5038 2338 5136 sw
tri 2338 5038 2436 5136 ne
rect 2436 5088 2750 5136
tri 2750 5088 2838 5176 sw
tri 2848 5088 2936 5176 ne
rect 2936 5140 2990 5176
rect 3110 5176 3212 5260
tri 3212 5176 3300 5264 sw
tri 3310 5176 3398 5264 ne
rect 3398 5260 3762 5264
rect 3398 5176 3540 5260
rect 3110 5140 3300 5176
rect 2936 5136 3300 5140
tri 3300 5136 3340 5176 sw
tri 3398 5136 3438 5176 ne
rect 3438 5140 3540 5176
rect 3660 5176 3762 5260
tri 3762 5176 3850 5264 sw
tri 3860 5176 3948 5264 ne
rect 3948 5260 4312 5264
rect 3948 5176 4090 5260
rect 3660 5140 3850 5176
rect 3438 5136 3850 5140
rect 2936 5088 3340 5136
rect 2436 5038 2838 5088
rect 1916 5008 2338 5038
rect 1424 4950 1818 5008
rect 914 4910 1326 4950
tri 1326 4910 1366 4950 sw
tri 1424 4910 1464 4950 ne
rect 1464 4910 1818 4950
tri 1818 4910 1916 5008 sw
tri 1916 4910 2014 5008 ne
rect 2014 4950 2338 5008
tri 2338 4950 2426 5038 sw
tri 2436 4950 2524 5038 ne
rect 2524 5008 2838 5038
tri 2838 5008 2918 5088 sw
tri 2936 5008 3016 5088 ne
rect 3016 5038 3340 5088
tri 3340 5038 3438 5136 sw
tri 3438 5038 3536 5136 ne
rect 3536 5088 3850 5136
tri 3850 5088 3938 5176 sw
tri 3948 5088 4036 5176 ne
rect 4036 5140 4090 5176
rect 4210 5176 4312 5260
tri 4312 5176 4400 5264 sw
tri 4410 5176 4498 5264 ne
rect 4498 5260 4862 5264
rect 4498 5176 4640 5260
rect 4210 5140 4400 5176
rect 4036 5136 4400 5140
tri 4400 5136 4440 5176 sw
tri 4498 5136 4538 5176 ne
rect 4538 5140 4640 5176
rect 4760 5176 4862 5260
tri 4862 5176 4950 5264 sw
tri 4960 5176 5048 5264 ne
rect 5048 5260 5412 5264
rect 5048 5176 5190 5260
rect 4760 5140 4950 5176
rect 4538 5136 4950 5140
rect 4036 5088 4440 5136
rect 3536 5038 3938 5088
rect 3016 5008 3438 5038
rect 2524 4950 2918 5008
rect 2014 4910 2426 4950
tri 2426 4910 2466 4950 sw
tri 2524 4910 2564 4950 ne
rect 2564 4910 2918 4950
tri 2918 4910 3016 5008 sw
tri 3016 4910 3114 5008 ne
rect 3114 4950 3438 5008
tri 3438 4950 3526 5038 sw
tri 3536 4950 3624 5038 ne
rect 3624 5008 3938 5038
tri 3938 5008 4018 5088 sw
tri 4036 5008 4116 5088 ne
rect 4116 5038 4440 5088
tri 4440 5038 4538 5136 sw
tri 4538 5038 4636 5136 ne
rect 4636 5088 4950 5136
tri 4950 5088 5038 5176 sw
tri 5048 5088 5136 5176 ne
rect 5136 5140 5190 5176
rect 5310 5176 5412 5260
tri 5412 5176 5500 5264 sw
tri 5510 5176 5598 5264 ne
rect 5598 5260 5962 5264
rect 5598 5176 5740 5260
rect 5310 5140 5500 5176
rect 5136 5136 5500 5140
tri 5500 5136 5540 5176 sw
tri 5598 5136 5638 5176 ne
rect 5638 5140 5740 5176
rect 5860 5176 5962 5260
tri 5962 5176 6050 5264 sw
tri 6060 5176 6148 5264 ne
rect 6148 5260 6512 5264
rect 6148 5176 6290 5260
rect 5860 5140 6050 5176
rect 5638 5136 6050 5140
rect 5136 5088 5540 5136
rect 4636 5038 5038 5088
rect 4116 5008 4538 5038
rect 3624 4950 4018 5008
rect 3114 4910 3526 4950
tri 3526 4910 3566 4950 sw
tri 3624 4910 3664 4950 ne
rect 3664 4910 4018 4950
tri 4018 4910 4116 5008 sw
tri 4116 4910 4214 5008 ne
rect 4214 4950 4538 5008
tri 4538 4950 4626 5038 sw
tri 4636 4950 4724 5038 ne
rect 4724 5008 5038 5038
tri 5038 5008 5118 5088 sw
tri 5136 5008 5216 5088 ne
rect 5216 5038 5540 5088
tri 5540 5038 5638 5136 sw
tri 5638 5038 5736 5136 ne
rect 5736 5088 6050 5136
tri 6050 5088 6138 5176 sw
tri 6148 5088 6236 5176 ne
rect 6236 5140 6290 5176
rect 6410 5176 6512 5260
tri 6512 5176 6600 5264 sw
tri 6610 5176 6698 5264 ne
rect 6698 5260 7062 5264
rect 6698 5176 6840 5260
rect 6410 5140 6600 5176
rect 6236 5136 6600 5140
tri 6600 5136 6640 5176 sw
tri 6698 5136 6738 5176 ne
rect 6738 5140 6840 5176
rect 6960 5176 7062 5260
tri 7062 5176 7150 5264 sw
tri 7160 5176 7248 5264 ne
rect 7248 5260 7612 5264
rect 7248 5176 7390 5260
rect 6960 5140 7150 5176
rect 6738 5136 7150 5140
rect 6236 5088 6640 5136
rect 5736 5038 6138 5088
rect 5216 5008 5638 5038
rect 4724 4950 5118 5008
rect 4214 4910 4626 4950
tri 4626 4910 4666 4950 sw
tri 4724 4910 4764 4950 ne
rect 4764 4910 5118 4950
tri 5118 4910 5216 5008 sw
tri 5216 4910 5314 5008 ne
rect 5314 4950 5638 5008
tri 5638 4950 5726 5038 sw
tri 5736 4950 5824 5038 ne
rect 5824 5008 6138 5038
tri 6138 5008 6218 5088 sw
tri 6236 5008 6316 5088 ne
rect 6316 5038 6640 5088
tri 6640 5038 6738 5136 sw
tri 6738 5038 6836 5136 ne
rect 6836 5088 7150 5136
tri 7150 5088 7238 5176 sw
tri 7248 5088 7336 5176 ne
rect 7336 5140 7390 5176
rect 7510 5176 7612 5260
tri 7612 5176 7700 5264 sw
tri 7710 5176 7798 5264 ne
rect 7798 5260 8162 5264
rect 7798 5176 7940 5260
rect 7510 5140 7700 5176
rect 7336 5136 7700 5140
tri 7700 5136 7740 5176 sw
tri 7798 5136 7838 5176 ne
rect 7838 5140 7940 5176
rect 8060 5176 8162 5260
tri 8162 5176 8250 5264 sw
tri 8260 5176 8348 5264 ne
rect 8348 5260 8712 5264
rect 8348 5176 8490 5260
rect 8060 5140 8250 5176
rect 7838 5136 8250 5140
rect 7336 5088 7740 5136
rect 6836 5038 7238 5088
rect 6316 5008 6738 5038
rect 5824 4950 6218 5008
rect 5314 4910 5726 4950
tri 5726 4910 5766 4950 sw
tri 5824 4910 5864 4950 ne
rect 5864 4910 6218 4950
tri 6218 4910 6316 5008 sw
tri 6316 4910 6414 5008 ne
rect 6414 4950 6738 5008
tri 6738 4950 6826 5038 sw
tri 6836 4950 6924 5038 ne
rect 6924 5008 7238 5038
tri 7238 5008 7318 5088 sw
tri 7336 5008 7416 5088 ne
rect 7416 5038 7740 5088
tri 7740 5038 7838 5136 sw
tri 7838 5038 7936 5136 ne
rect 7936 5088 8250 5136
tri 8250 5088 8338 5176 sw
tri 8348 5088 8436 5176 ne
rect 8436 5140 8490 5176
rect 8610 5176 8712 5260
tri 8712 5176 8800 5264 sw
tri 8810 5176 8898 5264 ne
rect 8898 5260 9262 5264
rect 8898 5176 9040 5260
rect 8610 5140 8800 5176
rect 8436 5136 8800 5140
tri 8800 5136 8840 5176 sw
tri 8898 5136 8938 5176 ne
rect 8938 5140 9040 5176
rect 9160 5176 9262 5260
tri 9262 5176 9350 5264 sw
tri 9360 5176 9448 5264 ne
rect 9448 5260 9812 5264
rect 9448 5176 9590 5260
rect 9160 5140 9350 5176
rect 8938 5136 9350 5140
rect 8436 5088 8840 5136
rect 7936 5038 8338 5088
rect 7416 5008 7838 5038
rect 6924 4950 7318 5008
rect 6414 4910 6826 4950
tri 6826 4910 6866 4950 sw
tri 6924 4910 6964 4950 ne
rect 6964 4910 7318 4950
tri 7318 4910 7416 5008 sw
tri 7416 4910 7514 5008 ne
rect 7514 4950 7838 5008
tri 7838 4950 7926 5038 sw
tri 7936 4950 8024 5038 ne
rect 8024 5008 8338 5038
tri 8338 5008 8418 5088 sw
tri 8436 5008 8516 5088 ne
rect 8516 5038 8840 5088
tri 8840 5038 8938 5136 sw
tri 8938 5038 9036 5136 ne
rect 9036 5088 9350 5136
tri 9350 5088 9438 5176 sw
tri 9448 5088 9536 5176 ne
rect 9536 5140 9590 5176
rect 9710 5176 9812 5260
tri 9812 5176 9900 5264 sw
tri 9910 5176 9998 5264 ne
rect 9998 5260 10362 5264
rect 9998 5176 10140 5260
rect 9710 5140 9900 5176
rect 9536 5136 9900 5140
tri 9900 5136 9940 5176 sw
tri 9998 5136 10038 5176 ne
rect 10038 5140 10140 5176
rect 10260 5176 10362 5260
tri 10362 5176 10450 5264 sw
tri 10460 5176 10548 5264 ne
rect 10548 5260 10912 5264
rect 10548 5176 10690 5260
rect 10260 5140 10450 5176
rect 10038 5136 10450 5140
rect 9536 5088 9940 5136
rect 9036 5038 9438 5088
rect 8516 5008 8938 5038
rect 8024 4950 8418 5008
rect 7514 4910 7926 4950
tri 7926 4910 7966 4950 sw
tri 8024 4910 8064 4950 ne
rect 8064 4910 8418 4950
tri 8418 4910 8516 5008 sw
tri 8516 4910 8614 5008 ne
rect 8614 4950 8938 5008
tri 8938 4950 9026 5038 sw
tri 9036 4950 9124 5038 ne
rect 9124 5008 9438 5038
tri 9438 5008 9518 5088 sw
tri 9536 5008 9616 5088 ne
rect 9616 5038 9940 5088
tri 9940 5038 10038 5136 sw
tri 10038 5038 10136 5136 ne
rect 10136 5088 10450 5136
tri 10450 5088 10538 5176 sw
tri 10548 5088 10636 5176 ne
rect 10636 5140 10690 5176
rect 10810 5176 10912 5260
tri 10912 5176 11000 5264 sw
tri 11010 5176 11098 5264 ne
rect 11098 5260 11462 5264
rect 11098 5176 11240 5260
rect 10810 5140 11000 5176
rect 10636 5136 11000 5140
tri 11000 5136 11040 5176 sw
tri 11098 5136 11138 5176 ne
rect 11138 5140 11240 5176
rect 11360 5176 11462 5260
tri 11462 5176 11550 5264 sw
tri 11560 5176 11648 5264 ne
rect 11648 5260 12012 5264
rect 11648 5176 11790 5260
rect 11360 5140 11550 5176
rect 11138 5136 11550 5140
rect 10636 5088 11040 5136
rect 10136 5038 10538 5088
rect 9616 5008 10038 5038
rect 9124 4950 9518 5008
rect 8614 4910 9026 4950
tri 9026 4910 9066 4950 sw
tri 9124 4910 9164 4950 ne
rect 9164 4910 9518 4950
tri 9518 4910 9616 5008 sw
tri 9616 4910 9714 5008 ne
rect 9714 4950 10038 5008
tri 10038 4950 10126 5038 sw
tri 10136 4950 10224 5038 ne
rect 10224 5008 10538 5038
tri 10538 5008 10618 5088 sw
tri 10636 5008 10716 5088 ne
rect 10716 5038 11040 5088
tri 11040 5038 11138 5136 sw
tri 11138 5038 11236 5136 ne
rect 11236 5088 11550 5136
tri 11550 5088 11638 5176 sw
tri 11648 5088 11736 5176 ne
rect 11736 5140 11790 5176
rect 11910 5176 12012 5260
tri 12012 5176 12100 5264 sw
tri 12110 5176 12198 5264 ne
rect 12198 5260 12562 5264
rect 12198 5176 12340 5260
rect 11910 5140 12100 5176
rect 11736 5136 12100 5140
tri 12100 5136 12140 5176 sw
tri 12198 5136 12238 5176 ne
rect 12238 5140 12340 5176
rect 12460 5176 12562 5260
tri 12562 5176 12650 5264 sw
tri 12660 5176 12748 5264 ne
rect 12748 5260 13112 5264
rect 12748 5176 12890 5260
rect 12460 5140 12650 5176
rect 12238 5136 12650 5140
rect 11736 5088 12140 5136
rect 11236 5038 11638 5088
rect 10716 5008 11138 5038
rect 10224 4950 10618 5008
rect 9714 4910 10126 4950
tri 10126 4910 10166 4950 sw
tri 10224 4910 10264 4950 ne
rect 10264 4910 10618 4950
tri 10618 4910 10716 5008 sw
tri 10716 4910 10814 5008 ne
rect 10814 4950 11138 5008
tri 11138 4950 11226 5038 sw
tri 11236 4950 11324 5038 ne
rect 11324 5008 11638 5038
tri 11638 5008 11718 5088 sw
tri 11736 5008 11816 5088 ne
rect 11816 5038 12140 5088
tri 12140 5038 12238 5136 sw
tri 12238 5038 12336 5136 ne
rect 12336 5088 12650 5136
tri 12650 5088 12738 5176 sw
tri 12748 5088 12836 5176 ne
rect 12836 5140 12890 5176
rect 13010 5176 13112 5260
tri 13112 5176 13200 5264 sw
tri 13210 5176 13298 5264 ne
rect 13298 5260 14275 5264
rect 13298 5176 13440 5260
rect 13010 5140 13200 5176
rect 12836 5136 13200 5140
tri 13200 5136 13240 5176 sw
tri 13298 5136 13338 5176 ne
rect 13338 5140 13440 5176
rect 13560 5140 14275 5260
rect 13338 5136 14275 5140
rect 12836 5088 13240 5136
rect 12336 5038 12738 5088
rect 11816 5008 12238 5038
rect 11324 4950 11718 5008
rect 10814 4910 11226 4950
tri 11226 4910 11266 4950 sw
tri 11324 4910 11364 4950 ne
rect 11364 4910 11718 4950
tri 11718 4910 11816 5008 sw
tri 11816 4910 11914 5008 ne
rect 11914 4950 12238 5008
tri 12238 4950 12326 5038 sw
tri 12336 4950 12424 5038 ne
rect 12424 5008 12738 5038
tri 12738 5008 12818 5088 sw
tri 12836 5008 12916 5088 ne
rect 12916 5038 13240 5088
tri 13240 5038 13338 5136 sw
tri 13338 5038 13436 5136 ne
rect 13436 5038 14275 5136
rect 12916 5008 13338 5038
rect 12424 4950 12818 5008
rect 11914 4910 12326 4950
tri 12326 4910 12366 4950 sw
tri 12424 4910 12464 4950 ne
rect 12464 4910 12818 4950
tri 12818 4910 12916 5008 sw
tri 12916 4910 13014 5008 ne
rect 13014 4950 13338 5008
tri 13338 4950 13426 5038 sw
tri 13436 4950 13524 5038 ne
rect 13524 4950 14275 5038
rect 13014 4910 13426 4950
tri 13426 4910 13466 4950 sw
tri 13524 4910 13564 4950 ne
rect 13564 4910 14275 4950
rect -2525 4812 -284 4910
tri -284 4812 -186 4910 sw
tri -186 4812 -88 4910 ne
rect -88 4812 266 4910
tri 266 4812 364 4910 sw
tri 364 4812 462 4910 ne
rect 462 4812 816 4910
tri 816 4812 914 4910 sw
tri 914 4812 1012 4910 ne
rect 1012 4812 1366 4910
tri 1366 4812 1464 4910 sw
tri 1464 4812 1562 4910 ne
rect 1562 4812 1916 4910
tri 1916 4812 2014 4910 sw
tri 2014 4812 2112 4910 ne
rect 2112 4812 2466 4910
tri 2466 4812 2564 4910 sw
tri 2564 4812 2662 4910 ne
rect 2662 4812 3016 4910
tri 3016 4812 3114 4910 sw
tri 3114 4812 3212 4910 ne
rect 3212 4812 3566 4910
tri 3566 4812 3664 4910 sw
tri 3664 4812 3762 4910 ne
rect 3762 4812 4116 4910
tri 4116 4812 4214 4910 sw
tri 4214 4812 4312 4910 ne
rect 4312 4812 4666 4910
tri 4666 4812 4764 4910 sw
tri 4764 4812 4862 4910 ne
rect 4862 4812 5216 4910
tri 5216 4812 5314 4910 sw
tri 5314 4812 5412 4910 ne
rect 5412 4812 5766 4910
tri 5766 4812 5864 4910 sw
tri 5864 4812 5962 4910 ne
rect 5962 4812 6316 4910
tri 6316 4812 6414 4910 sw
tri 6414 4812 6512 4910 ne
rect 6512 4812 6866 4910
tri 6866 4812 6964 4910 sw
tri 6964 4812 7062 4910 ne
rect 7062 4812 7416 4910
tri 7416 4812 7514 4910 sw
tri 7514 4812 7612 4910 ne
rect 7612 4812 7966 4910
tri 7966 4812 8064 4910 sw
tri 8064 4812 8162 4910 ne
rect 8162 4812 8516 4910
tri 8516 4812 8614 4910 sw
tri 8614 4812 8712 4910 ne
rect 8712 4812 9066 4910
tri 9066 4812 9164 4910 sw
tri 9164 4812 9262 4910 ne
rect 9262 4812 9616 4910
tri 9616 4812 9714 4910 sw
tri 9714 4812 9812 4910 ne
rect 9812 4812 10166 4910
tri 10166 4812 10264 4910 sw
tri 10264 4812 10362 4910 ne
rect 10362 4812 10716 4910
tri 10716 4812 10814 4910 sw
tri 10814 4812 10912 4910 ne
rect 10912 4812 11266 4910
tri 11266 4812 11364 4910 sw
tri 11364 4812 11462 4910 ne
rect 11462 4812 11816 4910
tri 11816 4812 11914 4910 sw
tri 11914 4812 12012 4910 ne
rect 12012 4812 12366 4910
tri 12366 4812 12464 4910 sw
tri 12464 4812 12562 4910 ne
rect 12562 4812 12916 4910
tri 12916 4812 13014 4910 sw
tri 13014 4812 13112 4910 ne
rect 13112 4812 13466 4910
tri 13466 4812 13564 4910 sw
tri 13564 4812 13662 4910 ne
rect 13662 4812 14275 4910
rect -2525 4714 -186 4812
tri -186 4714 -88 4812 sw
tri -88 4714 10 4812 ne
rect 10 4714 364 4812
tri 364 4714 462 4812 sw
tri 462 4714 560 4812 ne
rect 560 4714 914 4812
tri 914 4714 1012 4812 sw
tri 1012 4714 1110 4812 ne
rect 1110 4714 1464 4812
tri 1464 4714 1562 4812 sw
tri 1562 4714 1660 4812 ne
rect 1660 4714 2014 4812
tri 2014 4714 2112 4812 sw
tri 2112 4714 2210 4812 ne
rect 2210 4714 2564 4812
tri 2564 4714 2662 4812 sw
tri 2662 4714 2760 4812 ne
rect 2760 4714 3114 4812
tri 3114 4714 3212 4812 sw
tri 3212 4714 3310 4812 ne
rect 3310 4714 3664 4812
tri 3664 4714 3762 4812 sw
tri 3762 4714 3860 4812 ne
rect 3860 4714 4214 4812
tri 4214 4714 4312 4812 sw
tri 4312 4714 4410 4812 ne
rect 4410 4714 4764 4812
tri 4764 4714 4862 4812 sw
tri 4862 4714 4960 4812 ne
rect 4960 4714 5314 4812
tri 5314 4714 5412 4812 sw
tri 5412 4714 5510 4812 ne
rect 5510 4714 5864 4812
tri 5864 4714 5962 4812 sw
tri 5962 4714 6060 4812 ne
rect 6060 4714 6414 4812
tri 6414 4714 6512 4812 sw
tri 6512 4714 6610 4812 ne
rect 6610 4714 6964 4812
tri 6964 4714 7062 4812 sw
tri 7062 4714 7160 4812 ne
rect 7160 4714 7514 4812
tri 7514 4714 7612 4812 sw
tri 7612 4714 7710 4812 ne
rect 7710 4714 8064 4812
tri 8064 4714 8162 4812 sw
tri 8162 4714 8260 4812 ne
rect 8260 4714 8614 4812
tri 8614 4714 8712 4812 sw
tri 8712 4714 8810 4812 ne
rect 8810 4714 9164 4812
tri 9164 4714 9262 4812 sw
tri 9262 4714 9360 4812 ne
rect 9360 4714 9714 4812
tri 9714 4714 9812 4812 sw
tri 9812 4714 9910 4812 ne
rect 9910 4714 10264 4812
tri 10264 4714 10362 4812 sw
tri 10362 4714 10460 4812 ne
rect 10460 4714 10814 4812
tri 10814 4714 10912 4812 sw
tri 10912 4714 11010 4812 ne
rect 11010 4714 11364 4812
tri 11364 4714 11462 4812 sw
tri 11462 4714 11560 4812 ne
rect 11560 4714 11914 4812
tri 11914 4714 12012 4812 sw
tri 12012 4714 12110 4812 ne
rect 12110 4714 12464 4812
tri 12464 4714 12562 4812 sw
tri 12562 4714 12660 4812 ne
rect 12660 4714 13014 4812
tri 13014 4714 13112 4812 sw
tri 13112 4714 13210 4812 ne
rect 13210 4714 13564 4812
tri 13564 4714 13662 4812 sw
rect 14775 4714 15775 5362
rect -2525 4710 -88 4714
rect -2525 4590 -310 4710
rect -190 4626 -88 4710
tri -88 4626 0 4714 sw
tri 10 4626 98 4714 ne
rect 98 4710 462 4714
rect 98 4626 240 4710
rect -190 4590 0 4626
rect -2525 4586 0 4590
rect -2525 3938 -1525 4586
tri -412 4488 -314 4586 ne
rect -314 4538 0 4586
tri 0 4538 88 4626 sw
tri 98 4538 186 4626 ne
rect 186 4590 240 4626
rect 360 4626 462 4710
tri 462 4626 550 4714 sw
tri 560 4626 648 4714 ne
rect 648 4710 1012 4714
rect 648 4626 790 4710
rect 360 4590 550 4626
rect 186 4586 550 4590
tri 550 4586 590 4626 sw
tri 648 4586 688 4626 ne
rect 688 4590 790 4626
rect 910 4626 1012 4710
tri 1012 4626 1100 4714 sw
tri 1110 4626 1198 4714 ne
rect 1198 4710 1562 4714
rect 1198 4626 1340 4710
rect 910 4590 1100 4626
rect 688 4586 1100 4590
rect 186 4538 590 4586
rect -314 4488 88 4538
rect -1025 4400 -412 4488
tri -412 4400 -324 4488 sw
tri -314 4400 -226 4488 ne
rect -226 4458 88 4488
tri 88 4458 168 4538 sw
tri 186 4458 266 4538 ne
rect 266 4488 590 4538
tri 590 4488 688 4586 sw
tri 688 4488 786 4586 ne
rect 786 4538 1100 4586
tri 1100 4538 1188 4626 sw
tri 1198 4538 1286 4626 ne
rect 1286 4590 1340 4626
rect 1460 4626 1562 4710
tri 1562 4626 1650 4714 sw
tri 1660 4626 1748 4714 ne
rect 1748 4710 2112 4714
rect 1748 4626 1890 4710
rect 1460 4590 1650 4626
rect 1286 4586 1650 4590
tri 1650 4586 1690 4626 sw
tri 1748 4586 1788 4626 ne
rect 1788 4590 1890 4626
rect 2010 4626 2112 4710
tri 2112 4626 2200 4714 sw
tri 2210 4626 2298 4714 ne
rect 2298 4710 2662 4714
rect 2298 4626 2440 4710
rect 2010 4590 2200 4626
rect 1788 4586 2200 4590
rect 1286 4538 1690 4586
rect 786 4488 1188 4538
rect 266 4458 688 4488
rect -226 4400 168 4458
rect -1025 4360 -324 4400
tri -324 4360 -284 4400 sw
tri -226 4360 -186 4400 ne
rect -186 4360 168 4400
tri 168 4360 266 4458 sw
tri 266 4360 364 4458 ne
rect 364 4400 688 4458
tri 688 4400 776 4488 sw
tri 786 4400 874 4488 ne
rect 874 4458 1188 4488
tri 1188 4458 1268 4538 sw
tri 1286 4458 1366 4538 ne
rect 1366 4488 1690 4538
tri 1690 4488 1788 4586 sw
tri 1788 4488 1886 4586 ne
rect 1886 4538 2200 4586
tri 2200 4538 2288 4626 sw
tri 2298 4538 2386 4626 ne
rect 2386 4590 2440 4626
rect 2560 4626 2662 4710
tri 2662 4626 2750 4714 sw
tri 2760 4626 2848 4714 ne
rect 2848 4710 3212 4714
rect 2848 4626 2990 4710
rect 2560 4590 2750 4626
rect 2386 4586 2750 4590
tri 2750 4586 2790 4626 sw
tri 2848 4586 2888 4626 ne
rect 2888 4590 2990 4626
rect 3110 4626 3212 4710
tri 3212 4626 3300 4714 sw
tri 3310 4626 3398 4714 ne
rect 3398 4710 3762 4714
rect 3398 4626 3540 4710
rect 3110 4590 3300 4626
rect 2888 4586 3300 4590
rect 2386 4538 2790 4586
rect 1886 4488 2288 4538
rect 1366 4458 1788 4488
rect 874 4400 1268 4458
rect 364 4360 776 4400
tri 776 4360 816 4400 sw
tri 874 4360 914 4400 ne
rect 914 4360 1268 4400
tri 1268 4360 1366 4458 sw
tri 1366 4360 1464 4458 ne
rect 1464 4400 1788 4458
tri 1788 4400 1876 4488 sw
tri 1886 4400 1974 4488 ne
rect 1974 4458 2288 4488
tri 2288 4458 2368 4538 sw
tri 2386 4458 2466 4538 ne
rect 2466 4488 2790 4538
tri 2790 4488 2888 4586 sw
tri 2888 4488 2986 4586 ne
rect 2986 4538 3300 4586
tri 3300 4538 3388 4626 sw
tri 3398 4538 3486 4626 ne
rect 3486 4590 3540 4626
rect 3660 4626 3762 4710
tri 3762 4626 3850 4714 sw
tri 3860 4626 3948 4714 ne
rect 3948 4710 4312 4714
rect 3948 4626 4090 4710
rect 3660 4590 3850 4626
rect 3486 4586 3850 4590
tri 3850 4586 3890 4626 sw
tri 3948 4586 3988 4626 ne
rect 3988 4590 4090 4626
rect 4210 4626 4312 4710
tri 4312 4626 4400 4714 sw
tri 4410 4626 4498 4714 ne
rect 4498 4710 4862 4714
rect 4498 4626 4640 4710
rect 4210 4590 4400 4626
rect 3988 4586 4400 4590
rect 3486 4538 3890 4586
rect 2986 4488 3388 4538
rect 2466 4458 2888 4488
rect 1974 4400 2368 4458
rect 1464 4360 1876 4400
tri 1876 4360 1916 4400 sw
tri 1974 4360 2014 4400 ne
rect 2014 4360 2368 4400
tri 2368 4360 2466 4458 sw
tri 2466 4360 2564 4458 ne
rect 2564 4400 2888 4458
tri 2888 4400 2976 4488 sw
tri 2986 4400 3074 4488 ne
rect 3074 4458 3388 4488
tri 3388 4458 3468 4538 sw
tri 3486 4458 3566 4538 ne
rect 3566 4488 3890 4538
tri 3890 4488 3988 4586 sw
tri 3988 4488 4086 4586 ne
rect 4086 4538 4400 4586
tri 4400 4538 4488 4626 sw
tri 4498 4538 4586 4626 ne
rect 4586 4590 4640 4626
rect 4760 4626 4862 4710
tri 4862 4626 4950 4714 sw
tri 4960 4626 5048 4714 ne
rect 5048 4710 5412 4714
rect 5048 4626 5190 4710
rect 4760 4590 4950 4626
rect 4586 4586 4950 4590
tri 4950 4586 4990 4626 sw
tri 5048 4586 5088 4626 ne
rect 5088 4590 5190 4626
rect 5310 4626 5412 4710
tri 5412 4626 5500 4714 sw
tri 5510 4626 5598 4714 ne
rect 5598 4710 5962 4714
rect 5598 4626 5740 4710
rect 5310 4590 5500 4626
rect 5088 4586 5500 4590
rect 4586 4538 4990 4586
rect 4086 4488 4488 4538
rect 3566 4458 3988 4488
rect 3074 4400 3468 4458
rect 2564 4360 2976 4400
tri 2976 4360 3016 4400 sw
tri 3074 4360 3114 4400 ne
rect 3114 4360 3468 4400
tri 3468 4360 3566 4458 sw
tri 3566 4360 3664 4458 ne
rect 3664 4400 3988 4458
tri 3988 4400 4076 4488 sw
tri 4086 4400 4174 4488 ne
rect 4174 4458 4488 4488
tri 4488 4458 4568 4538 sw
tri 4586 4458 4666 4538 ne
rect 4666 4488 4990 4538
tri 4990 4488 5088 4586 sw
tri 5088 4488 5186 4586 ne
rect 5186 4538 5500 4586
tri 5500 4538 5588 4626 sw
tri 5598 4538 5686 4626 ne
rect 5686 4590 5740 4626
rect 5860 4626 5962 4710
tri 5962 4626 6050 4714 sw
tri 6060 4626 6148 4714 ne
rect 6148 4710 6512 4714
rect 6148 4626 6290 4710
rect 5860 4590 6050 4626
rect 5686 4586 6050 4590
tri 6050 4586 6090 4626 sw
tri 6148 4586 6188 4626 ne
rect 6188 4590 6290 4626
rect 6410 4626 6512 4710
tri 6512 4626 6600 4714 sw
tri 6610 4626 6698 4714 ne
rect 6698 4710 7062 4714
rect 6698 4626 6840 4710
rect 6410 4590 6600 4626
rect 6188 4586 6600 4590
rect 5686 4538 6090 4586
rect 5186 4488 5588 4538
rect 4666 4458 5088 4488
rect 4174 4400 4568 4458
rect 3664 4360 4076 4400
tri 4076 4360 4116 4400 sw
tri 4174 4360 4214 4400 ne
rect 4214 4360 4568 4400
tri 4568 4360 4666 4458 sw
tri 4666 4360 4764 4458 ne
rect 4764 4400 5088 4458
tri 5088 4400 5176 4488 sw
tri 5186 4400 5274 4488 ne
rect 5274 4458 5588 4488
tri 5588 4458 5668 4538 sw
tri 5686 4458 5766 4538 ne
rect 5766 4488 6090 4538
tri 6090 4488 6188 4586 sw
tri 6188 4488 6286 4586 ne
rect 6286 4538 6600 4586
tri 6600 4538 6688 4626 sw
tri 6698 4538 6786 4626 ne
rect 6786 4590 6840 4626
rect 6960 4626 7062 4710
tri 7062 4626 7150 4714 sw
tri 7160 4626 7248 4714 ne
rect 7248 4710 7612 4714
rect 7248 4626 7390 4710
rect 6960 4590 7150 4626
rect 6786 4586 7150 4590
tri 7150 4586 7190 4626 sw
tri 7248 4586 7288 4626 ne
rect 7288 4590 7390 4626
rect 7510 4626 7612 4710
tri 7612 4626 7700 4714 sw
tri 7710 4626 7798 4714 ne
rect 7798 4710 8162 4714
rect 7798 4626 7940 4710
rect 7510 4590 7700 4626
rect 7288 4586 7700 4590
rect 6786 4538 7190 4586
rect 6286 4488 6688 4538
rect 5766 4458 6188 4488
rect 5274 4400 5668 4458
rect 4764 4360 5176 4400
tri 5176 4360 5216 4400 sw
tri 5274 4360 5314 4400 ne
rect 5314 4360 5668 4400
tri 5668 4360 5766 4458 sw
tri 5766 4360 5864 4458 ne
rect 5864 4400 6188 4458
tri 6188 4400 6276 4488 sw
tri 6286 4400 6374 4488 ne
rect 6374 4458 6688 4488
tri 6688 4458 6768 4538 sw
tri 6786 4458 6866 4538 ne
rect 6866 4488 7190 4538
tri 7190 4488 7288 4586 sw
tri 7288 4488 7386 4586 ne
rect 7386 4538 7700 4586
tri 7700 4538 7788 4626 sw
tri 7798 4538 7886 4626 ne
rect 7886 4590 7940 4626
rect 8060 4626 8162 4710
tri 8162 4626 8250 4714 sw
tri 8260 4626 8348 4714 ne
rect 8348 4710 8712 4714
rect 8348 4626 8490 4710
rect 8060 4590 8250 4626
rect 7886 4586 8250 4590
tri 8250 4586 8290 4626 sw
tri 8348 4586 8388 4626 ne
rect 8388 4590 8490 4626
rect 8610 4626 8712 4710
tri 8712 4626 8800 4714 sw
tri 8810 4626 8898 4714 ne
rect 8898 4710 9262 4714
rect 8898 4626 9040 4710
rect 8610 4590 8800 4626
rect 8388 4586 8800 4590
rect 7886 4538 8290 4586
rect 7386 4488 7788 4538
rect 6866 4458 7288 4488
rect 6374 4400 6768 4458
rect 5864 4360 6276 4400
tri 6276 4360 6316 4400 sw
tri 6374 4360 6414 4400 ne
rect 6414 4360 6768 4400
tri 6768 4360 6866 4458 sw
tri 6866 4360 6964 4458 ne
rect 6964 4400 7288 4458
tri 7288 4400 7376 4488 sw
tri 7386 4400 7474 4488 ne
rect 7474 4458 7788 4488
tri 7788 4458 7868 4538 sw
tri 7886 4458 7966 4538 ne
rect 7966 4488 8290 4538
tri 8290 4488 8388 4586 sw
tri 8388 4488 8486 4586 ne
rect 8486 4538 8800 4586
tri 8800 4538 8888 4626 sw
tri 8898 4538 8986 4626 ne
rect 8986 4590 9040 4626
rect 9160 4626 9262 4710
tri 9262 4626 9350 4714 sw
tri 9360 4626 9448 4714 ne
rect 9448 4710 9812 4714
rect 9448 4626 9590 4710
rect 9160 4590 9350 4626
rect 8986 4586 9350 4590
tri 9350 4586 9390 4626 sw
tri 9448 4586 9488 4626 ne
rect 9488 4590 9590 4626
rect 9710 4626 9812 4710
tri 9812 4626 9900 4714 sw
tri 9910 4626 9998 4714 ne
rect 9998 4710 10362 4714
rect 9998 4626 10140 4710
rect 9710 4590 9900 4626
rect 9488 4586 9900 4590
rect 8986 4538 9390 4586
rect 8486 4488 8888 4538
rect 7966 4458 8388 4488
rect 7474 4400 7868 4458
rect 6964 4360 7376 4400
tri 7376 4360 7416 4400 sw
tri 7474 4360 7514 4400 ne
rect 7514 4360 7868 4400
tri 7868 4360 7966 4458 sw
tri 7966 4360 8064 4458 ne
rect 8064 4400 8388 4458
tri 8388 4400 8476 4488 sw
tri 8486 4400 8574 4488 ne
rect 8574 4458 8888 4488
tri 8888 4458 8968 4538 sw
tri 8986 4458 9066 4538 ne
rect 9066 4488 9390 4538
tri 9390 4488 9488 4586 sw
tri 9488 4488 9586 4586 ne
rect 9586 4538 9900 4586
tri 9900 4538 9988 4626 sw
tri 9998 4538 10086 4626 ne
rect 10086 4590 10140 4626
rect 10260 4626 10362 4710
tri 10362 4626 10450 4714 sw
tri 10460 4626 10548 4714 ne
rect 10548 4710 10912 4714
rect 10548 4626 10690 4710
rect 10260 4590 10450 4626
rect 10086 4586 10450 4590
tri 10450 4586 10490 4626 sw
tri 10548 4586 10588 4626 ne
rect 10588 4590 10690 4626
rect 10810 4626 10912 4710
tri 10912 4626 11000 4714 sw
tri 11010 4626 11098 4714 ne
rect 11098 4710 11462 4714
rect 11098 4626 11240 4710
rect 10810 4590 11000 4626
rect 10588 4586 11000 4590
rect 10086 4538 10490 4586
rect 9586 4488 9988 4538
rect 9066 4458 9488 4488
rect 8574 4400 8968 4458
rect 8064 4360 8476 4400
tri 8476 4360 8516 4400 sw
tri 8574 4360 8614 4400 ne
rect 8614 4360 8968 4400
tri 8968 4360 9066 4458 sw
tri 9066 4360 9164 4458 ne
rect 9164 4400 9488 4458
tri 9488 4400 9576 4488 sw
tri 9586 4400 9674 4488 ne
rect 9674 4458 9988 4488
tri 9988 4458 10068 4538 sw
tri 10086 4458 10166 4538 ne
rect 10166 4488 10490 4538
tri 10490 4488 10588 4586 sw
tri 10588 4488 10686 4586 ne
rect 10686 4538 11000 4586
tri 11000 4538 11088 4626 sw
tri 11098 4538 11186 4626 ne
rect 11186 4590 11240 4626
rect 11360 4626 11462 4710
tri 11462 4626 11550 4714 sw
tri 11560 4626 11648 4714 ne
rect 11648 4710 12012 4714
rect 11648 4626 11790 4710
rect 11360 4590 11550 4626
rect 11186 4586 11550 4590
tri 11550 4586 11590 4626 sw
tri 11648 4586 11688 4626 ne
rect 11688 4590 11790 4626
rect 11910 4626 12012 4710
tri 12012 4626 12100 4714 sw
tri 12110 4626 12198 4714 ne
rect 12198 4710 12562 4714
rect 12198 4626 12340 4710
rect 11910 4590 12100 4626
rect 11688 4586 12100 4590
rect 11186 4538 11590 4586
rect 10686 4488 11088 4538
rect 10166 4458 10588 4488
rect 9674 4400 10068 4458
rect 9164 4360 9576 4400
tri 9576 4360 9616 4400 sw
tri 9674 4360 9714 4400 ne
rect 9714 4360 10068 4400
tri 10068 4360 10166 4458 sw
tri 10166 4360 10264 4458 ne
rect 10264 4400 10588 4458
tri 10588 4400 10676 4488 sw
tri 10686 4400 10774 4488 ne
rect 10774 4458 11088 4488
tri 11088 4458 11168 4538 sw
tri 11186 4458 11266 4538 ne
rect 11266 4488 11590 4538
tri 11590 4488 11688 4586 sw
tri 11688 4488 11786 4586 ne
rect 11786 4538 12100 4586
tri 12100 4538 12188 4626 sw
tri 12198 4538 12286 4626 ne
rect 12286 4590 12340 4626
rect 12460 4626 12562 4710
tri 12562 4626 12650 4714 sw
tri 12660 4626 12748 4714 ne
rect 12748 4710 13112 4714
rect 12748 4626 12890 4710
rect 12460 4590 12650 4626
rect 12286 4586 12650 4590
tri 12650 4586 12690 4626 sw
tri 12748 4586 12788 4626 ne
rect 12788 4590 12890 4626
rect 13010 4626 13112 4710
tri 13112 4626 13200 4714 sw
tri 13210 4626 13298 4714 ne
rect 13298 4710 15775 4714
rect 13298 4626 13440 4710
rect 13010 4590 13200 4626
rect 12788 4586 13200 4590
rect 12286 4538 12690 4586
rect 11786 4488 12188 4538
rect 11266 4458 11688 4488
rect 10774 4400 11168 4458
rect 10264 4360 10676 4400
tri 10676 4360 10716 4400 sw
tri 10774 4360 10814 4400 ne
rect 10814 4360 11168 4400
tri 11168 4360 11266 4458 sw
tri 11266 4360 11364 4458 ne
rect 11364 4400 11688 4458
tri 11688 4400 11776 4488 sw
tri 11786 4400 11874 4488 ne
rect 11874 4458 12188 4488
tri 12188 4458 12268 4538 sw
tri 12286 4458 12366 4538 ne
rect 12366 4488 12690 4538
tri 12690 4488 12788 4586 sw
tri 12788 4488 12886 4586 ne
rect 12886 4538 13200 4586
tri 13200 4538 13288 4626 sw
tri 13298 4538 13386 4626 ne
rect 13386 4590 13440 4626
rect 13560 4590 15775 4710
rect 13386 4538 15775 4590
rect 12886 4488 13288 4538
rect 12366 4458 12788 4488
rect 11874 4400 12268 4458
rect 11364 4360 11776 4400
tri 11776 4360 11816 4400 sw
tri 11874 4360 11914 4400 ne
rect 11914 4360 12268 4400
tri 12268 4360 12366 4458 sw
tri 12366 4360 12464 4458 ne
rect 12464 4400 12788 4458
tri 12788 4400 12876 4488 sw
tri 12886 4400 12974 4488 ne
rect 12974 4458 13288 4488
tri 13288 4458 13368 4538 sw
tri 13386 4458 13466 4538 ne
rect 13466 4458 14075 4538
rect 12974 4400 13368 4458
rect 12464 4360 12876 4400
tri 12876 4360 12916 4400 sw
tri 12974 4360 13014 4400 ne
rect 13014 4360 13368 4400
tri 13368 4360 13466 4458 sw
tri 13466 4360 13564 4458 ne
rect 13564 4438 14075 4458
rect 14175 4438 15775 4538
rect 13564 4360 15775 4438
rect -1025 4312 -284 4360
rect -1025 4212 -925 4312
rect -825 4262 -284 4312
tri -284 4262 -186 4360 sw
tri -186 4262 -88 4360 ne
rect -88 4262 266 4360
tri 266 4262 364 4360 sw
tri 364 4262 462 4360 ne
rect 462 4262 816 4360
tri 816 4262 914 4360 sw
tri 914 4262 1012 4360 ne
rect 1012 4262 1366 4360
tri 1366 4262 1464 4360 sw
tri 1464 4262 1562 4360 ne
rect 1562 4262 1916 4360
tri 1916 4262 2014 4360 sw
tri 2014 4262 2112 4360 ne
rect 2112 4262 2466 4360
tri 2466 4262 2564 4360 sw
tri 2564 4262 2662 4360 ne
rect 2662 4262 3016 4360
tri 3016 4262 3114 4360 sw
tri 3114 4262 3212 4360 ne
rect 3212 4262 3566 4360
tri 3566 4262 3664 4360 sw
tri 3664 4262 3762 4360 ne
rect 3762 4262 4116 4360
tri 4116 4262 4214 4360 sw
tri 4214 4262 4312 4360 ne
rect 4312 4262 4666 4360
tri 4666 4262 4764 4360 sw
tri 4764 4262 4862 4360 ne
rect 4862 4262 5216 4360
tri 5216 4262 5314 4360 sw
tri 5314 4262 5412 4360 ne
rect 5412 4262 5766 4360
tri 5766 4262 5864 4360 sw
tri 5864 4262 5962 4360 ne
rect 5962 4262 6316 4360
tri 6316 4262 6414 4360 sw
tri 6414 4262 6512 4360 ne
rect 6512 4262 6866 4360
tri 6866 4262 6964 4360 sw
tri 6964 4262 7062 4360 ne
rect 7062 4262 7416 4360
tri 7416 4262 7514 4360 sw
tri 7514 4262 7612 4360 ne
rect 7612 4262 7966 4360
tri 7966 4262 8064 4360 sw
tri 8064 4262 8162 4360 ne
rect 8162 4262 8516 4360
tri 8516 4262 8614 4360 sw
tri 8614 4262 8712 4360 ne
rect 8712 4262 9066 4360
tri 9066 4262 9164 4360 sw
tri 9164 4262 9262 4360 ne
rect 9262 4262 9616 4360
tri 9616 4262 9714 4360 sw
tri 9714 4262 9812 4360 ne
rect 9812 4262 10166 4360
tri 10166 4262 10264 4360 sw
tri 10264 4262 10362 4360 ne
rect 10362 4262 10716 4360
tri 10716 4262 10814 4360 sw
tri 10814 4262 10912 4360 ne
rect 10912 4262 11266 4360
tri 11266 4262 11364 4360 sw
tri 11364 4262 11462 4360 ne
rect 11462 4262 11816 4360
tri 11816 4262 11914 4360 sw
tri 11914 4262 12012 4360 ne
rect 12012 4262 12366 4360
tri 12366 4262 12464 4360 sw
tri 12464 4262 12562 4360 ne
rect 12562 4262 12916 4360
tri 12916 4262 13014 4360 sw
tri 13014 4262 13112 4360 ne
rect 13112 4262 13466 4360
tri 13466 4262 13564 4360 sw
tri 13564 4262 13662 4360 ne
rect 13662 4262 15775 4360
rect -825 4212 -186 4262
rect -1025 4164 -186 4212
tri -186 4164 -88 4262 sw
tri -88 4164 10 4262 ne
rect 10 4164 364 4262
tri 364 4164 462 4262 sw
tri 462 4164 560 4262 ne
rect 560 4164 914 4262
tri 914 4164 1012 4262 sw
tri 1012 4164 1110 4262 ne
rect 1110 4164 1464 4262
tri 1464 4164 1562 4262 sw
tri 1562 4164 1660 4262 ne
rect 1660 4164 2014 4262
tri 2014 4164 2112 4262 sw
tri 2112 4164 2210 4262 ne
rect 2210 4164 2564 4262
tri 2564 4164 2662 4262 sw
tri 2662 4164 2760 4262 ne
rect 2760 4164 3114 4262
tri 3114 4164 3212 4262 sw
tri 3212 4164 3310 4262 ne
rect 3310 4164 3664 4262
tri 3664 4164 3762 4262 sw
tri 3762 4164 3860 4262 ne
rect 3860 4164 4214 4262
tri 4214 4164 4312 4262 sw
tri 4312 4164 4410 4262 ne
rect 4410 4164 4764 4262
tri 4764 4164 4862 4262 sw
tri 4862 4164 4960 4262 ne
rect 4960 4164 5314 4262
tri 5314 4164 5412 4262 sw
tri 5412 4164 5510 4262 ne
rect 5510 4164 5864 4262
tri 5864 4164 5962 4262 sw
tri 5962 4164 6060 4262 ne
rect 6060 4164 6414 4262
tri 6414 4164 6512 4262 sw
tri 6512 4164 6610 4262 ne
rect 6610 4164 6964 4262
tri 6964 4164 7062 4262 sw
tri 7062 4164 7160 4262 ne
rect 7160 4164 7514 4262
tri 7514 4164 7612 4262 sw
tri 7612 4164 7710 4262 ne
rect 7710 4164 8064 4262
tri 8064 4164 8162 4262 sw
tri 8162 4164 8260 4262 ne
rect 8260 4164 8614 4262
tri 8614 4164 8712 4262 sw
tri 8712 4164 8810 4262 ne
rect 8810 4164 9164 4262
tri 9164 4164 9262 4262 sw
tri 9262 4164 9360 4262 ne
rect 9360 4164 9714 4262
tri 9714 4164 9812 4262 sw
tri 9812 4164 9910 4262 ne
rect 9910 4164 10264 4262
tri 10264 4164 10362 4262 sw
tri 10362 4164 10460 4262 ne
rect 10460 4164 10814 4262
tri 10814 4164 10912 4262 sw
tri 10912 4164 11010 4262 ne
rect 11010 4164 11364 4262
tri 11364 4164 11462 4262 sw
tri 11462 4164 11560 4262 ne
rect 11560 4164 11914 4262
tri 11914 4164 12012 4262 sw
tri 12012 4164 12110 4262 ne
rect 12110 4164 12464 4262
tri 12464 4164 12562 4262 sw
tri 12562 4164 12660 4262 ne
rect 12660 4164 13014 4262
tri 13014 4164 13112 4262 sw
tri 13112 4164 13210 4262 ne
rect 13210 4164 13564 4262
tri 13564 4164 13662 4262 sw
rect -1025 4160 -88 4164
rect -1025 4040 -310 4160
rect -190 4076 -88 4160
tri -88 4076 0 4164 sw
tri 10 4076 98 4164 ne
rect 98 4160 462 4164
rect 98 4076 240 4160
rect -190 4040 0 4076
rect -1025 4036 0 4040
tri 0 4036 40 4076 sw
tri 98 4036 138 4076 ne
rect 138 4040 240 4076
rect 360 4076 462 4160
tri 462 4076 550 4164 sw
tri 560 4076 648 4164 ne
rect 648 4160 1012 4164
rect 648 4076 790 4160
rect 360 4040 550 4076
rect 138 4036 550 4040
tri -412 3938 -314 4036 ne
rect -314 3938 40 4036
tri 40 3938 138 4036 sw
tri 138 3938 236 4036 ne
rect 236 3988 550 4036
tri 550 3988 638 4076 sw
tri 648 3988 736 4076 ne
rect 736 4040 790 4076
rect 910 4076 1012 4160
tri 1012 4076 1100 4164 sw
tri 1110 4076 1198 4164 ne
rect 1198 4160 1562 4164
rect 1198 4076 1340 4160
rect 910 4040 1100 4076
rect 736 4036 1100 4040
tri 1100 4036 1140 4076 sw
tri 1198 4036 1238 4076 ne
rect 1238 4040 1340 4076
rect 1460 4076 1562 4160
tri 1562 4076 1650 4164 sw
tri 1660 4076 1748 4164 ne
rect 1748 4160 2112 4164
rect 1748 4076 1890 4160
rect 1460 4040 1650 4076
rect 1238 4036 1650 4040
rect 736 3988 1140 4036
rect 236 3938 638 3988
rect -2525 3850 -412 3938
tri -412 3850 -324 3938 sw
tri -314 3850 -226 3938 ne
rect -226 3850 138 3938
tri 138 3850 226 3938 sw
tri 236 3850 324 3938 ne
rect 324 3908 638 3938
tri 638 3908 718 3988 sw
tri 736 3908 816 3988 ne
rect 816 3938 1140 3988
tri 1140 3938 1238 4036 sw
tri 1238 3938 1336 4036 ne
rect 1336 3988 1650 4036
tri 1650 3988 1738 4076 sw
tri 1748 3988 1836 4076 ne
rect 1836 4040 1890 4076
rect 2010 4076 2112 4160
tri 2112 4076 2200 4164 sw
tri 2210 4076 2298 4164 ne
rect 2298 4160 2662 4164
rect 2298 4076 2440 4160
rect 2010 4040 2200 4076
rect 1836 4036 2200 4040
tri 2200 4036 2240 4076 sw
tri 2298 4036 2338 4076 ne
rect 2338 4040 2440 4076
rect 2560 4076 2662 4160
tri 2662 4076 2750 4164 sw
tri 2760 4076 2848 4164 ne
rect 2848 4160 3212 4164
rect 2848 4076 2990 4160
rect 2560 4040 2750 4076
rect 2338 4036 2750 4040
rect 1836 3988 2240 4036
rect 1336 3938 1738 3988
rect 816 3908 1238 3938
rect 324 3850 718 3908
rect -2525 3810 -324 3850
tri -324 3810 -284 3850 sw
tri -226 3810 -186 3850 ne
rect -186 3810 226 3850
tri 226 3810 266 3850 sw
tri 324 3810 364 3850 ne
rect 364 3810 718 3850
tri 718 3810 816 3908 sw
tri 816 3810 914 3908 ne
rect 914 3850 1238 3908
tri 1238 3850 1326 3938 sw
tri 1336 3850 1424 3938 ne
rect 1424 3908 1738 3938
tri 1738 3908 1818 3988 sw
tri 1836 3908 1916 3988 ne
rect 1916 3938 2240 3988
tri 2240 3938 2338 4036 sw
tri 2338 3938 2436 4036 ne
rect 2436 3988 2750 4036
tri 2750 3988 2838 4076 sw
tri 2848 3988 2936 4076 ne
rect 2936 4040 2990 4076
rect 3110 4076 3212 4160
tri 3212 4076 3300 4164 sw
tri 3310 4076 3398 4164 ne
rect 3398 4160 3762 4164
rect 3398 4076 3540 4160
rect 3110 4040 3300 4076
rect 2936 4036 3300 4040
tri 3300 4036 3340 4076 sw
tri 3398 4036 3438 4076 ne
rect 3438 4040 3540 4076
rect 3660 4076 3762 4160
tri 3762 4076 3850 4164 sw
tri 3860 4076 3948 4164 ne
rect 3948 4160 4312 4164
rect 3948 4076 4090 4160
rect 3660 4040 3850 4076
rect 3438 4036 3850 4040
rect 2936 3988 3340 4036
rect 2436 3938 2838 3988
rect 1916 3908 2338 3938
rect 1424 3850 1818 3908
rect 914 3810 1326 3850
tri 1326 3810 1366 3850 sw
tri 1424 3810 1464 3850 ne
rect 1464 3810 1818 3850
tri 1818 3810 1916 3908 sw
tri 1916 3810 2014 3908 ne
rect 2014 3850 2338 3908
tri 2338 3850 2426 3938 sw
tri 2436 3850 2524 3938 ne
rect 2524 3908 2838 3938
tri 2838 3908 2918 3988 sw
tri 2936 3908 3016 3988 ne
rect 3016 3938 3340 3988
tri 3340 3938 3438 4036 sw
tri 3438 3938 3536 4036 ne
rect 3536 3988 3850 4036
tri 3850 3988 3938 4076 sw
tri 3948 3988 4036 4076 ne
rect 4036 4040 4090 4076
rect 4210 4076 4312 4160
tri 4312 4076 4400 4164 sw
tri 4410 4076 4498 4164 ne
rect 4498 4160 4862 4164
rect 4498 4076 4640 4160
rect 4210 4040 4400 4076
rect 4036 4036 4400 4040
tri 4400 4036 4440 4076 sw
tri 4498 4036 4538 4076 ne
rect 4538 4040 4640 4076
rect 4760 4076 4862 4160
tri 4862 4076 4950 4164 sw
tri 4960 4076 5048 4164 ne
rect 5048 4160 5412 4164
rect 5048 4076 5190 4160
rect 4760 4040 4950 4076
rect 4538 4036 4950 4040
rect 4036 3988 4440 4036
rect 3536 3938 3938 3988
rect 3016 3908 3438 3938
rect 2524 3850 2918 3908
rect 2014 3810 2426 3850
tri 2426 3810 2466 3850 sw
tri 2524 3810 2564 3850 ne
rect 2564 3810 2918 3850
tri 2918 3810 3016 3908 sw
tri 3016 3810 3114 3908 ne
rect 3114 3850 3438 3908
tri 3438 3850 3526 3938 sw
tri 3536 3850 3624 3938 ne
rect 3624 3908 3938 3938
tri 3938 3908 4018 3988 sw
tri 4036 3908 4116 3988 ne
rect 4116 3938 4440 3988
tri 4440 3938 4538 4036 sw
tri 4538 3938 4636 4036 ne
rect 4636 3988 4950 4036
tri 4950 3988 5038 4076 sw
tri 5048 3988 5136 4076 ne
rect 5136 4040 5190 4076
rect 5310 4076 5412 4160
tri 5412 4076 5500 4164 sw
tri 5510 4076 5598 4164 ne
rect 5598 4160 5962 4164
rect 5598 4076 5740 4160
rect 5310 4040 5500 4076
rect 5136 4036 5500 4040
tri 5500 4036 5540 4076 sw
tri 5598 4036 5638 4076 ne
rect 5638 4040 5740 4076
rect 5860 4076 5962 4160
tri 5962 4076 6050 4164 sw
tri 6060 4076 6148 4164 ne
rect 6148 4160 6512 4164
rect 6148 4076 6290 4160
rect 5860 4040 6050 4076
rect 5638 4036 6050 4040
rect 5136 3988 5540 4036
rect 4636 3938 5038 3988
rect 4116 3908 4538 3938
rect 3624 3850 4018 3908
rect 3114 3810 3526 3850
tri 3526 3810 3566 3850 sw
tri 3624 3810 3664 3850 ne
rect 3664 3810 4018 3850
tri 4018 3810 4116 3908 sw
tri 4116 3810 4214 3908 ne
rect 4214 3850 4538 3908
tri 4538 3850 4626 3938 sw
tri 4636 3850 4724 3938 ne
rect 4724 3908 5038 3938
tri 5038 3908 5118 3988 sw
tri 5136 3908 5216 3988 ne
rect 5216 3938 5540 3988
tri 5540 3938 5638 4036 sw
tri 5638 3938 5736 4036 ne
rect 5736 3988 6050 4036
tri 6050 3988 6138 4076 sw
tri 6148 3988 6236 4076 ne
rect 6236 4040 6290 4076
rect 6410 4076 6512 4160
tri 6512 4076 6600 4164 sw
tri 6610 4076 6698 4164 ne
rect 6698 4160 7062 4164
rect 6698 4076 6840 4160
rect 6410 4040 6600 4076
rect 6236 4036 6600 4040
tri 6600 4036 6640 4076 sw
tri 6698 4036 6738 4076 ne
rect 6738 4040 6840 4076
rect 6960 4076 7062 4160
tri 7062 4076 7150 4164 sw
tri 7160 4076 7248 4164 ne
rect 7248 4160 7612 4164
rect 7248 4076 7390 4160
rect 6960 4040 7150 4076
rect 6738 4036 7150 4040
rect 6236 3988 6640 4036
rect 5736 3938 6138 3988
rect 5216 3908 5638 3938
rect 4724 3850 5118 3908
rect 4214 3810 4626 3850
tri 4626 3810 4666 3850 sw
tri 4724 3810 4764 3850 ne
rect 4764 3810 5118 3850
tri 5118 3810 5216 3908 sw
tri 5216 3810 5314 3908 ne
rect 5314 3850 5638 3908
tri 5638 3850 5726 3938 sw
tri 5736 3850 5824 3938 ne
rect 5824 3908 6138 3938
tri 6138 3908 6218 3988 sw
tri 6236 3908 6316 3988 ne
rect 6316 3938 6640 3988
tri 6640 3938 6738 4036 sw
tri 6738 3938 6836 4036 ne
rect 6836 3988 7150 4036
tri 7150 3988 7238 4076 sw
tri 7248 3988 7336 4076 ne
rect 7336 4040 7390 4076
rect 7510 4076 7612 4160
tri 7612 4076 7700 4164 sw
tri 7710 4076 7798 4164 ne
rect 7798 4160 8162 4164
rect 7798 4076 7940 4160
rect 7510 4040 7700 4076
rect 7336 4036 7700 4040
tri 7700 4036 7740 4076 sw
tri 7798 4036 7838 4076 ne
rect 7838 4040 7940 4076
rect 8060 4076 8162 4160
tri 8162 4076 8250 4164 sw
tri 8260 4076 8348 4164 ne
rect 8348 4160 8712 4164
rect 8348 4076 8490 4160
rect 8060 4040 8250 4076
rect 7838 4036 8250 4040
rect 7336 3988 7740 4036
rect 6836 3938 7238 3988
rect 6316 3908 6738 3938
rect 5824 3850 6218 3908
rect 5314 3810 5726 3850
tri 5726 3810 5766 3850 sw
tri 5824 3810 5864 3850 ne
rect 5864 3810 6218 3850
tri 6218 3810 6316 3908 sw
tri 6316 3810 6414 3908 ne
rect 6414 3850 6738 3908
tri 6738 3850 6826 3938 sw
tri 6836 3850 6924 3938 ne
rect 6924 3908 7238 3938
tri 7238 3908 7318 3988 sw
tri 7336 3908 7416 3988 ne
rect 7416 3938 7740 3988
tri 7740 3938 7838 4036 sw
tri 7838 3938 7936 4036 ne
rect 7936 3988 8250 4036
tri 8250 3988 8338 4076 sw
tri 8348 3988 8436 4076 ne
rect 8436 4040 8490 4076
rect 8610 4076 8712 4160
tri 8712 4076 8800 4164 sw
tri 8810 4076 8898 4164 ne
rect 8898 4160 9262 4164
rect 8898 4076 9040 4160
rect 8610 4040 8800 4076
rect 8436 4036 8800 4040
tri 8800 4036 8840 4076 sw
tri 8898 4036 8938 4076 ne
rect 8938 4040 9040 4076
rect 9160 4076 9262 4160
tri 9262 4076 9350 4164 sw
tri 9360 4076 9448 4164 ne
rect 9448 4160 9812 4164
rect 9448 4076 9590 4160
rect 9160 4040 9350 4076
rect 8938 4036 9350 4040
rect 8436 3988 8840 4036
rect 7936 3938 8338 3988
rect 7416 3908 7838 3938
rect 6924 3850 7318 3908
rect 6414 3810 6826 3850
tri 6826 3810 6866 3850 sw
tri 6924 3810 6964 3850 ne
rect 6964 3810 7318 3850
tri 7318 3810 7416 3908 sw
tri 7416 3810 7514 3908 ne
rect 7514 3850 7838 3908
tri 7838 3850 7926 3938 sw
tri 7936 3850 8024 3938 ne
rect 8024 3908 8338 3938
tri 8338 3908 8418 3988 sw
tri 8436 3908 8516 3988 ne
rect 8516 3938 8840 3988
tri 8840 3938 8938 4036 sw
tri 8938 3938 9036 4036 ne
rect 9036 3988 9350 4036
tri 9350 3988 9438 4076 sw
tri 9448 3988 9536 4076 ne
rect 9536 4040 9590 4076
rect 9710 4076 9812 4160
tri 9812 4076 9900 4164 sw
tri 9910 4076 9998 4164 ne
rect 9998 4160 10362 4164
rect 9998 4076 10140 4160
rect 9710 4040 9900 4076
rect 9536 4036 9900 4040
tri 9900 4036 9940 4076 sw
tri 9998 4036 10038 4076 ne
rect 10038 4040 10140 4076
rect 10260 4076 10362 4160
tri 10362 4076 10450 4164 sw
tri 10460 4076 10548 4164 ne
rect 10548 4160 10912 4164
rect 10548 4076 10690 4160
rect 10260 4040 10450 4076
rect 10038 4036 10450 4040
rect 9536 3988 9940 4036
rect 9036 3938 9438 3988
rect 8516 3908 8938 3938
rect 8024 3850 8418 3908
rect 7514 3810 7926 3850
tri 7926 3810 7966 3850 sw
tri 8024 3810 8064 3850 ne
rect 8064 3810 8418 3850
tri 8418 3810 8516 3908 sw
tri 8516 3810 8614 3908 ne
rect 8614 3850 8938 3908
tri 8938 3850 9026 3938 sw
tri 9036 3850 9124 3938 ne
rect 9124 3908 9438 3938
tri 9438 3908 9518 3988 sw
tri 9536 3908 9616 3988 ne
rect 9616 3938 9940 3988
tri 9940 3938 10038 4036 sw
tri 10038 3938 10136 4036 ne
rect 10136 3988 10450 4036
tri 10450 3988 10538 4076 sw
tri 10548 3988 10636 4076 ne
rect 10636 4040 10690 4076
rect 10810 4076 10912 4160
tri 10912 4076 11000 4164 sw
tri 11010 4076 11098 4164 ne
rect 11098 4160 11462 4164
rect 11098 4076 11240 4160
rect 10810 4040 11000 4076
rect 10636 4036 11000 4040
tri 11000 4036 11040 4076 sw
tri 11098 4036 11138 4076 ne
rect 11138 4040 11240 4076
rect 11360 4076 11462 4160
tri 11462 4076 11550 4164 sw
tri 11560 4076 11648 4164 ne
rect 11648 4160 12012 4164
rect 11648 4076 11790 4160
rect 11360 4040 11550 4076
rect 11138 4036 11550 4040
rect 10636 3988 11040 4036
rect 10136 3938 10538 3988
rect 9616 3908 10038 3938
rect 9124 3850 9518 3908
rect 8614 3810 9026 3850
tri 9026 3810 9066 3850 sw
tri 9124 3810 9164 3850 ne
rect 9164 3810 9518 3850
tri 9518 3810 9616 3908 sw
tri 9616 3810 9714 3908 ne
rect 9714 3850 10038 3908
tri 10038 3850 10126 3938 sw
tri 10136 3850 10224 3938 ne
rect 10224 3908 10538 3938
tri 10538 3908 10618 3988 sw
tri 10636 3908 10716 3988 ne
rect 10716 3938 11040 3988
tri 11040 3938 11138 4036 sw
tri 11138 3938 11236 4036 ne
rect 11236 3988 11550 4036
tri 11550 3988 11638 4076 sw
tri 11648 3988 11736 4076 ne
rect 11736 4040 11790 4076
rect 11910 4076 12012 4160
tri 12012 4076 12100 4164 sw
tri 12110 4076 12198 4164 ne
rect 12198 4160 12562 4164
rect 12198 4076 12340 4160
rect 11910 4040 12100 4076
rect 11736 4036 12100 4040
tri 12100 4036 12140 4076 sw
tri 12198 4036 12238 4076 ne
rect 12238 4040 12340 4076
rect 12460 4076 12562 4160
tri 12562 4076 12650 4164 sw
tri 12660 4076 12748 4164 ne
rect 12748 4160 13112 4164
rect 12748 4076 12890 4160
rect 12460 4040 12650 4076
rect 12238 4036 12650 4040
rect 11736 3988 12140 4036
rect 11236 3938 11638 3988
rect 10716 3908 11138 3938
rect 10224 3850 10618 3908
rect 9714 3810 10126 3850
tri 10126 3810 10166 3850 sw
tri 10224 3810 10264 3850 ne
rect 10264 3810 10618 3850
tri 10618 3810 10716 3908 sw
tri 10716 3810 10814 3908 ne
rect 10814 3850 11138 3908
tri 11138 3850 11226 3938 sw
tri 11236 3850 11324 3938 ne
rect 11324 3908 11638 3938
tri 11638 3908 11718 3988 sw
tri 11736 3908 11816 3988 ne
rect 11816 3938 12140 3988
tri 12140 3938 12238 4036 sw
tri 12238 3938 12336 4036 ne
rect 12336 3988 12650 4036
tri 12650 3988 12738 4076 sw
tri 12748 3988 12836 4076 ne
rect 12836 4040 12890 4076
rect 13010 4076 13112 4160
tri 13112 4076 13200 4164 sw
tri 13210 4076 13298 4164 ne
rect 13298 4160 14275 4164
rect 13298 4076 13440 4160
rect 13010 4040 13200 4076
rect 12836 4036 13200 4040
tri 13200 4036 13240 4076 sw
tri 13298 4036 13338 4076 ne
rect 13338 4040 13440 4076
rect 13560 4040 14275 4160
rect 13338 4036 14275 4040
rect 12836 3988 13240 4036
rect 12336 3938 12738 3988
rect 11816 3908 12238 3938
rect 11324 3850 11718 3908
rect 10814 3810 11226 3850
tri 11226 3810 11266 3850 sw
tri 11324 3810 11364 3850 ne
rect 11364 3810 11718 3850
tri 11718 3810 11816 3908 sw
tri 11816 3810 11914 3908 ne
rect 11914 3850 12238 3908
tri 12238 3850 12326 3938 sw
tri 12336 3850 12424 3938 ne
rect 12424 3908 12738 3938
tri 12738 3908 12818 3988 sw
tri 12836 3908 12916 3988 ne
rect 12916 3938 13240 3988
tri 13240 3938 13338 4036 sw
tri 13338 3938 13436 4036 ne
rect 13436 3938 14275 4036
rect 12916 3908 13338 3938
rect 12424 3850 12818 3908
rect 11914 3810 12326 3850
tri 12326 3810 12366 3850 sw
tri 12424 3810 12464 3850 ne
rect 12464 3810 12818 3850
tri 12818 3810 12916 3908 sw
tri 12916 3810 13014 3908 ne
rect 13014 3850 13338 3908
tri 13338 3850 13426 3938 sw
tri 13436 3850 13524 3938 ne
rect 13524 3850 14275 3938
rect 13014 3810 13426 3850
tri 13426 3810 13466 3850 sw
tri 13524 3810 13564 3850 ne
rect 13564 3810 14275 3850
rect -2525 3712 -284 3810
tri -284 3712 -186 3810 sw
tri -186 3712 -88 3810 ne
rect -88 3712 266 3810
tri 266 3712 364 3810 sw
tri 364 3712 462 3810 ne
rect 462 3712 816 3810
tri 816 3712 914 3810 sw
tri 914 3712 1012 3810 ne
rect 1012 3712 1366 3810
tri 1366 3712 1464 3810 sw
tri 1464 3712 1562 3810 ne
rect 1562 3712 1916 3810
tri 1916 3712 2014 3810 sw
tri 2014 3712 2112 3810 ne
rect 2112 3712 2466 3810
tri 2466 3712 2564 3810 sw
tri 2564 3712 2662 3810 ne
rect 2662 3712 3016 3810
tri 3016 3712 3114 3810 sw
tri 3114 3712 3212 3810 ne
rect 3212 3712 3566 3810
tri 3566 3712 3664 3810 sw
tri 3664 3712 3762 3810 ne
rect 3762 3712 4116 3810
tri 4116 3712 4214 3810 sw
tri 4214 3712 4312 3810 ne
rect 4312 3712 4666 3810
tri 4666 3712 4764 3810 sw
tri 4764 3712 4862 3810 ne
rect 4862 3712 5216 3810
tri 5216 3712 5314 3810 sw
tri 5314 3712 5412 3810 ne
rect 5412 3712 5766 3810
tri 5766 3712 5864 3810 sw
tri 5864 3712 5962 3810 ne
rect 5962 3712 6316 3810
tri 6316 3712 6414 3810 sw
tri 6414 3712 6512 3810 ne
rect 6512 3712 6866 3810
tri 6866 3712 6964 3810 sw
tri 6964 3712 7062 3810 ne
rect 7062 3712 7416 3810
tri 7416 3712 7514 3810 sw
tri 7514 3712 7612 3810 ne
rect 7612 3712 7966 3810
tri 7966 3712 8064 3810 sw
tri 8064 3712 8162 3810 ne
rect 8162 3712 8516 3810
tri 8516 3712 8614 3810 sw
tri 8614 3712 8712 3810 ne
rect 8712 3712 9066 3810
tri 9066 3712 9164 3810 sw
tri 9164 3712 9262 3810 ne
rect 9262 3712 9616 3810
tri 9616 3712 9714 3810 sw
tri 9714 3712 9812 3810 ne
rect 9812 3712 10166 3810
tri 10166 3712 10264 3810 sw
tri 10264 3712 10362 3810 ne
rect 10362 3712 10716 3810
tri 10716 3712 10814 3810 sw
tri 10814 3712 10912 3810 ne
rect 10912 3712 11266 3810
tri 11266 3712 11364 3810 sw
tri 11364 3712 11462 3810 ne
rect 11462 3712 11816 3810
tri 11816 3712 11914 3810 sw
tri 11914 3712 12012 3810 ne
rect 12012 3712 12366 3810
tri 12366 3712 12464 3810 sw
tri 12464 3712 12562 3810 ne
rect 12562 3712 12916 3810
tri 12916 3712 13014 3810 sw
tri 13014 3712 13112 3810 ne
rect 13112 3712 13466 3810
tri 13466 3712 13564 3810 sw
tri 13564 3712 13662 3810 ne
rect 13662 3712 14275 3810
rect -2525 3614 -186 3712
tri -186 3614 -88 3712 sw
tri -88 3614 10 3712 ne
rect 10 3614 364 3712
tri 364 3614 462 3712 sw
tri 462 3614 560 3712 ne
rect 560 3614 914 3712
tri 914 3614 1012 3712 sw
tri 1012 3614 1110 3712 ne
rect 1110 3614 1464 3712
tri 1464 3614 1562 3712 sw
tri 1562 3614 1660 3712 ne
rect 1660 3614 2014 3712
tri 2014 3614 2112 3712 sw
tri 2112 3614 2210 3712 ne
rect 2210 3614 2564 3712
tri 2564 3614 2662 3712 sw
tri 2662 3614 2760 3712 ne
rect 2760 3614 3114 3712
tri 3114 3614 3212 3712 sw
tri 3212 3614 3310 3712 ne
rect 3310 3614 3664 3712
tri 3664 3614 3762 3712 sw
tri 3762 3614 3860 3712 ne
rect 3860 3614 4214 3712
tri 4214 3614 4312 3712 sw
tri 4312 3614 4410 3712 ne
rect 4410 3614 4764 3712
tri 4764 3614 4862 3712 sw
tri 4862 3614 4960 3712 ne
rect 4960 3614 5314 3712
tri 5314 3614 5412 3712 sw
tri 5412 3614 5510 3712 ne
rect 5510 3614 5864 3712
tri 5864 3614 5962 3712 sw
tri 5962 3614 6060 3712 ne
rect 6060 3614 6414 3712
tri 6414 3614 6512 3712 sw
tri 6512 3614 6610 3712 ne
rect 6610 3614 6964 3712
tri 6964 3614 7062 3712 sw
tri 7062 3614 7160 3712 ne
rect 7160 3614 7514 3712
tri 7514 3614 7612 3712 sw
tri 7612 3614 7710 3712 ne
rect 7710 3614 8064 3712
tri 8064 3614 8162 3712 sw
tri 8162 3614 8260 3712 ne
rect 8260 3614 8614 3712
tri 8614 3614 8712 3712 sw
tri 8712 3614 8810 3712 ne
rect 8810 3614 9164 3712
tri 9164 3614 9262 3712 sw
tri 9262 3614 9360 3712 ne
rect 9360 3614 9714 3712
tri 9714 3614 9812 3712 sw
tri 9812 3614 9910 3712 ne
rect 9910 3614 10264 3712
tri 10264 3614 10362 3712 sw
tri 10362 3614 10460 3712 ne
rect 10460 3614 10814 3712
tri 10814 3614 10912 3712 sw
tri 10912 3614 11010 3712 ne
rect 11010 3614 11364 3712
tri 11364 3614 11462 3712 sw
tri 11462 3614 11560 3712 ne
rect 11560 3614 11914 3712
tri 11914 3614 12012 3712 sw
tri 12012 3614 12110 3712 ne
rect 12110 3614 12464 3712
tri 12464 3614 12562 3712 sw
tri 12562 3614 12660 3712 ne
rect 12660 3614 13014 3712
tri 13014 3614 13112 3712 sw
tri 13112 3614 13210 3712 ne
rect 13210 3614 13564 3712
tri 13564 3614 13662 3712 sw
rect 14775 3614 15775 4262
rect -2525 3610 -88 3614
rect -2525 3490 -310 3610
rect -190 3526 -88 3610
tri -88 3526 0 3614 sw
tri 10 3526 98 3614 ne
rect 98 3610 462 3614
rect 98 3526 240 3610
rect -190 3490 0 3526
rect -2525 3486 0 3490
rect -2525 2838 -1525 3486
tri -412 3388 -314 3486 ne
rect -314 3438 0 3486
tri 0 3438 88 3526 sw
tri 98 3438 186 3526 ne
rect 186 3490 240 3526
rect 360 3526 462 3610
tri 462 3526 550 3614 sw
tri 560 3526 648 3614 ne
rect 648 3610 1012 3614
rect 648 3526 790 3610
rect 360 3490 550 3526
rect 186 3486 550 3490
tri 550 3486 590 3526 sw
tri 648 3486 688 3526 ne
rect 688 3490 790 3526
rect 910 3526 1012 3610
tri 1012 3526 1100 3614 sw
tri 1110 3526 1198 3614 ne
rect 1198 3610 1562 3614
rect 1198 3526 1340 3610
rect 910 3490 1100 3526
rect 688 3486 1100 3490
rect 186 3438 590 3486
rect -314 3388 88 3438
rect -1025 3300 -412 3388
tri -412 3300 -324 3388 sw
tri -314 3300 -226 3388 ne
rect -226 3358 88 3388
tri 88 3358 168 3438 sw
tri 186 3358 266 3438 ne
rect 266 3388 590 3438
tri 590 3388 688 3486 sw
tri 688 3388 786 3486 ne
rect 786 3438 1100 3486
tri 1100 3438 1188 3526 sw
tri 1198 3438 1286 3526 ne
rect 1286 3490 1340 3526
rect 1460 3526 1562 3610
tri 1562 3526 1650 3614 sw
tri 1660 3526 1748 3614 ne
rect 1748 3610 2112 3614
rect 1748 3526 1890 3610
rect 1460 3490 1650 3526
rect 1286 3486 1650 3490
tri 1650 3486 1690 3526 sw
tri 1748 3486 1788 3526 ne
rect 1788 3490 1890 3526
rect 2010 3526 2112 3610
tri 2112 3526 2200 3614 sw
tri 2210 3526 2298 3614 ne
rect 2298 3610 2662 3614
rect 2298 3526 2440 3610
rect 2010 3490 2200 3526
rect 1788 3486 2200 3490
rect 1286 3438 1690 3486
rect 786 3388 1188 3438
rect 266 3358 688 3388
rect -226 3300 168 3358
rect -1025 3260 -324 3300
tri -324 3260 -284 3300 sw
tri -226 3260 -186 3300 ne
rect -186 3260 168 3300
tri 168 3260 266 3358 sw
tri 266 3260 364 3358 ne
rect 364 3300 688 3358
tri 688 3300 776 3388 sw
tri 786 3300 874 3388 ne
rect 874 3358 1188 3388
tri 1188 3358 1268 3438 sw
tri 1286 3358 1366 3438 ne
rect 1366 3388 1690 3438
tri 1690 3388 1788 3486 sw
tri 1788 3388 1886 3486 ne
rect 1886 3438 2200 3486
tri 2200 3438 2288 3526 sw
tri 2298 3438 2386 3526 ne
rect 2386 3490 2440 3526
rect 2560 3526 2662 3610
tri 2662 3526 2750 3614 sw
tri 2760 3526 2848 3614 ne
rect 2848 3610 3212 3614
rect 2848 3526 2990 3610
rect 2560 3490 2750 3526
rect 2386 3486 2750 3490
tri 2750 3486 2790 3526 sw
tri 2848 3486 2888 3526 ne
rect 2888 3490 2990 3526
rect 3110 3526 3212 3610
tri 3212 3526 3300 3614 sw
tri 3310 3526 3398 3614 ne
rect 3398 3610 3762 3614
rect 3398 3526 3540 3610
rect 3110 3490 3300 3526
rect 2888 3486 3300 3490
rect 2386 3438 2790 3486
rect 1886 3388 2288 3438
rect 1366 3358 1788 3388
rect 874 3300 1268 3358
rect 364 3260 776 3300
tri 776 3260 816 3300 sw
tri 874 3260 914 3300 ne
rect 914 3260 1268 3300
tri 1268 3260 1366 3358 sw
tri 1366 3260 1464 3358 ne
rect 1464 3300 1788 3358
tri 1788 3300 1876 3388 sw
tri 1886 3300 1974 3388 ne
rect 1974 3358 2288 3388
tri 2288 3358 2368 3438 sw
tri 2386 3358 2466 3438 ne
rect 2466 3388 2790 3438
tri 2790 3388 2888 3486 sw
tri 2888 3388 2986 3486 ne
rect 2986 3438 3300 3486
tri 3300 3438 3388 3526 sw
tri 3398 3438 3486 3526 ne
rect 3486 3490 3540 3526
rect 3660 3526 3762 3610
tri 3762 3526 3850 3614 sw
tri 3860 3526 3948 3614 ne
rect 3948 3610 4312 3614
rect 3948 3526 4090 3610
rect 3660 3490 3850 3526
rect 3486 3486 3850 3490
tri 3850 3486 3890 3526 sw
tri 3948 3486 3988 3526 ne
rect 3988 3490 4090 3526
rect 4210 3526 4312 3610
tri 4312 3526 4400 3614 sw
tri 4410 3526 4498 3614 ne
rect 4498 3610 4862 3614
rect 4498 3526 4640 3610
rect 4210 3490 4400 3526
rect 3988 3486 4400 3490
rect 3486 3438 3890 3486
rect 2986 3388 3388 3438
rect 2466 3358 2888 3388
rect 1974 3300 2368 3358
rect 1464 3260 1876 3300
tri 1876 3260 1916 3300 sw
tri 1974 3260 2014 3300 ne
rect 2014 3260 2368 3300
tri 2368 3260 2466 3358 sw
tri 2466 3260 2564 3358 ne
rect 2564 3300 2888 3358
tri 2888 3300 2976 3388 sw
tri 2986 3300 3074 3388 ne
rect 3074 3358 3388 3388
tri 3388 3358 3468 3438 sw
tri 3486 3358 3566 3438 ne
rect 3566 3388 3890 3438
tri 3890 3388 3988 3486 sw
tri 3988 3388 4086 3486 ne
rect 4086 3438 4400 3486
tri 4400 3438 4488 3526 sw
tri 4498 3438 4586 3526 ne
rect 4586 3490 4640 3526
rect 4760 3526 4862 3610
tri 4862 3526 4950 3614 sw
tri 4960 3526 5048 3614 ne
rect 5048 3610 5412 3614
rect 5048 3526 5190 3610
rect 4760 3490 4950 3526
rect 4586 3486 4950 3490
tri 4950 3486 4990 3526 sw
tri 5048 3486 5088 3526 ne
rect 5088 3490 5190 3526
rect 5310 3526 5412 3610
tri 5412 3526 5500 3614 sw
tri 5510 3526 5598 3614 ne
rect 5598 3610 5962 3614
rect 5598 3526 5740 3610
rect 5310 3490 5500 3526
rect 5088 3486 5500 3490
rect 4586 3438 4990 3486
rect 4086 3388 4488 3438
rect 3566 3358 3988 3388
rect 3074 3300 3468 3358
rect 2564 3260 2976 3300
tri 2976 3260 3016 3300 sw
tri 3074 3260 3114 3300 ne
rect 3114 3260 3468 3300
tri 3468 3260 3566 3358 sw
tri 3566 3260 3664 3358 ne
rect 3664 3300 3988 3358
tri 3988 3300 4076 3388 sw
tri 4086 3300 4174 3388 ne
rect 4174 3358 4488 3388
tri 4488 3358 4568 3438 sw
tri 4586 3358 4666 3438 ne
rect 4666 3388 4990 3438
tri 4990 3388 5088 3486 sw
tri 5088 3388 5186 3486 ne
rect 5186 3438 5500 3486
tri 5500 3438 5588 3526 sw
tri 5598 3438 5686 3526 ne
rect 5686 3490 5740 3526
rect 5860 3526 5962 3610
tri 5962 3526 6050 3614 sw
tri 6060 3526 6148 3614 ne
rect 6148 3610 6512 3614
rect 6148 3526 6290 3610
rect 5860 3490 6050 3526
rect 5686 3486 6050 3490
tri 6050 3486 6090 3526 sw
tri 6148 3486 6188 3526 ne
rect 6188 3490 6290 3526
rect 6410 3526 6512 3610
tri 6512 3526 6600 3614 sw
tri 6610 3526 6698 3614 ne
rect 6698 3610 7062 3614
rect 6698 3526 6840 3610
rect 6410 3490 6600 3526
rect 6188 3486 6600 3490
rect 5686 3438 6090 3486
rect 5186 3388 5588 3438
rect 4666 3358 5088 3388
rect 4174 3300 4568 3358
rect 3664 3260 4076 3300
tri 4076 3260 4116 3300 sw
tri 4174 3260 4214 3300 ne
rect 4214 3260 4568 3300
tri 4568 3260 4666 3358 sw
tri 4666 3260 4764 3358 ne
rect 4764 3300 5088 3358
tri 5088 3300 5176 3388 sw
tri 5186 3300 5274 3388 ne
rect 5274 3358 5588 3388
tri 5588 3358 5668 3438 sw
tri 5686 3358 5766 3438 ne
rect 5766 3388 6090 3438
tri 6090 3388 6188 3486 sw
tri 6188 3388 6286 3486 ne
rect 6286 3438 6600 3486
tri 6600 3438 6688 3526 sw
tri 6698 3438 6786 3526 ne
rect 6786 3490 6840 3526
rect 6960 3526 7062 3610
tri 7062 3526 7150 3614 sw
tri 7160 3526 7248 3614 ne
rect 7248 3610 7612 3614
rect 7248 3526 7390 3610
rect 6960 3490 7150 3526
rect 6786 3486 7150 3490
tri 7150 3486 7190 3526 sw
tri 7248 3486 7288 3526 ne
rect 7288 3490 7390 3526
rect 7510 3526 7612 3610
tri 7612 3526 7700 3614 sw
tri 7710 3526 7798 3614 ne
rect 7798 3610 8162 3614
rect 7798 3526 7940 3610
rect 7510 3490 7700 3526
rect 7288 3486 7700 3490
rect 6786 3438 7190 3486
rect 6286 3388 6688 3438
rect 5766 3358 6188 3388
rect 5274 3300 5668 3358
rect 4764 3260 5176 3300
tri 5176 3260 5216 3300 sw
tri 5274 3260 5314 3300 ne
rect 5314 3260 5668 3300
tri 5668 3260 5766 3358 sw
tri 5766 3260 5864 3358 ne
rect 5864 3300 6188 3358
tri 6188 3300 6276 3388 sw
tri 6286 3300 6374 3388 ne
rect 6374 3358 6688 3388
tri 6688 3358 6768 3438 sw
tri 6786 3358 6866 3438 ne
rect 6866 3388 7190 3438
tri 7190 3388 7288 3486 sw
tri 7288 3388 7386 3486 ne
rect 7386 3438 7700 3486
tri 7700 3438 7788 3526 sw
tri 7798 3438 7886 3526 ne
rect 7886 3490 7940 3526
rect 8060 3526 8162 3610
tri 8162 3526 8250 3614 sw
tri 8260 3526 8348 3614 ne
rect 8348 3610 8712 3614
rect 8348 3526 8490 3610
rect 8060 3490 8250 3526
rect 7886 3486 8250 3490
tri 8250 3486 8290 3526 sw
tri 8348 3486 8388 3526 ne
rect 8388 3490 8490 3526
rect 8610 3526 8712 3610
tri 8712 3526 8800 3614 sw
tri 8810 3526 8898 3614 ne
rect 8898 3610 9262 3614
rect 8898 3526 9040 3610
rect 8610 3490 8800 3526
rect 8388 3486 8800 3490
rect 7886 3438 8290 3486
rect 7386 3388 7788 3438
rect 6866 3358 7288 3388
rect 6374 3300 6768 3358
rect 5864 3260 6276 3300
tri 6276 3260 6316 3300 sw
tri 6374 3260 6414 3300 ne
rect 6414 3260 6768 3300
tri 6768 3260 6866 3358 sw
tri 6866 3260 6964 3358 ne
rect 6964 3300 7288 3358
tri 7288 3300 7376 3388 sw
tri 7386 3300 7474 3388 ne
rect 7474 3358 7788 3388
tri 7788 3358 7868 3438 sw
tri 7886 3358 7966 3438 ne
rect 7966 3388 8290 3438
tri 8290 3388 8388 3486 sw
tri 8388 3388 8486 3486 ne
rect 8486 3438 8800 3486
tri 8800 3438 8888 3526 sw
tri 8898 3438 8986 3526 ne
rect 8986 3490 9040 3526
rect 9160 3526 9262 3610
tri 9262 3526 9350 3614 sw
tri 9360 3526 9448 3614 ne
rect 9448 3610 9812 3614
rect 9448 3526 9590 3610
rect 9160 3490 9350 3526
rect 8986 3486 9350 3490
tri 9350 3486 9390 3526 sw
tri 9448 3486 9488 3526 ne
rect 9488 3490 9590 3526
rect 9710 3526 9812 3610
tri 9812 3526 9900 3614 sw
tri 9910 3526 9998 3614 ne
rect 9998 3610 10362 3614
rect 9998 3526 10140 3610
rect 9710 3490 9900 3526
rect 9488 3486 9900 3490
rect 8986 3438 9390 3486
rect 8486 3388 8888 3438
rect 7966 3358 8388 3388
rect 7474 3300 7868 3358
rect 6964 3260 7376 3300
tri 7376 3260 7416 3300 sw
tri 7474 3260 7514 3300 ne
rect 7514 3260 7868 3300
tri 7868 3260 7966 3358 sw
tri 7966 3260 8064 3358 ne
rect 8064 3300 8388 3358
tri 8388 3300 8476 3388 sw
tri 8486 3300 8574 3388 ne
rect 8574 3358 8888 3388
tri 8888 3358 8968 3438 sw
tri 8986 3358 9066 3438 ne
rect 9066 3388 9390 3438
tri 9390 3388 9488 3486 sw
tri 9488 3388 9586 3486 ne
rect 9586 3438 9900 3486
tri 9900 3438 9988 3526 sw
tri 9998 3438 10086 3526 ne
rect 10086 3490 10140 3526
rect 10260 3526 10362 3610
tri 10362 3526 10450 3614 sw
tri 10460 3526 10548 3614 ne
rect 10548 3610 10912 3614
rect 10548 3526 10690 3610
rect 10260 3490 10450 3526
rect 10086 3486 10450 3490
tri 10450 3486 10490 3526 sw
tri 10548 3486 10588 3526 ne
rect 10588 3490 10690 3526
rect 10810 3526 10912 3610
tri 10912 3526 11000 3614 sw
tri 11010 3526 11098 3614 ne
rect 11098 3610 11462 3614
rect 11098 3526 11240 3610
rect 10810 3490 11000 3526
rect 10588 3486 11000 3490
rect 10086 3438 10490 3486
rect 9586 3388 9988 3438
rect 9066 3358 9488 3388
rect 8574 3300 8968 3358
rect 8064 3260 8476 3300
tri 8476 3260 8516 3300 sw
tri 8574 3260 8614 3300 ne
rect 8614 3260 8968 3300
tri 8968 3260 9066 3358 sw
tri 9066 3260 9164 3358 ne
rect 9164 3300 9488 3358
tri 9488 3300 9576 3388 sw
tri 9586 3300 9674 3388 ne
rect 9674 3358 9988 3388
tri 9988 3358 10068 3438 sw
tri 10086 3358 10166 3438 ne
rect 10166 3388 10490 3438
tri 10490 3388 10588 3486 sw
tri 10588 3388 10686 3486 ne
rect 10686 3438 11000 3486
tri 11000 3438 11088 3526 sw
tri 11098 3438 11186 3526 ne
rect 11186 3490 11240 3526
rect 11360 3526 11462 3610
tri 11462 3526 11550 3614 sw
tri 11560 3526 11648 3614 ne
rect 11648 3610 12012 3614
rect 11648 3526 11790 3610
rect 11360 3490 11550 3526
rect 11186 3486 11550 3490
tri 11550 3486 11590 3526 sw
tri 11648 3486 11688 3526 ne
rect 11688 3490 11790 3526
rect 11910 3526 12012 3610
tri 12012 3526 12100 3614 sw
tri 12110 3526 12198 3614 ne
rect 12198 3610 12562 3614
rect 12198 3526 12340 3610
rect 11910 3490 12100 3526
rect 11688 3486 12100 3490
rect 11186 3438 11590 3486
rect 10686 3388 11088 3438
rect 10166 3358 10588 3388
rect 9674 3300 10068 3358
rect 9164 3260 9576 3300
tri 9576 3260 9616 3300 sw
tri 9674 3260 9714 3300 ne
rect 9714 3260 10068 3300
tri 10068 3260 10166 3358 sw
tri 10166 3260 10264 3358 ne
rect 10264 3300 10588 3358
tri 10588 3300 10676 3388 sw
tri 10686 3300 10774 3388 ne
rect 10774 3358 11088 3388
tri 11088 3358 11168 3438 sw
tri 11186 3358 11266 3438 ne
rect 11266 3388 11590 3438
tri 11590 3388 11688 3486 sw
tri 11688 3388 11786 3486 ne
rect 11786 3438 12100 3486
tri 12100 3438 12188 3526 sw
tri 12198 3438 12286 3526 ne
rect 12286 3490 12340 3526
rect 12460 3526 12562 3610
tri 12562 3526 12650 3614 sw
tri 12660 3526 12748 3614 ne
rect 12748 3610 13112 3614
rect 12748 3526 12890 3610
rect 12460 3490 12650 3526
rect 12286 3486 12650 3490
tri 12650 3486 12690 3526 sw
tri 12748 3486 12788 3526 ne
rect 12788 3490 12890 3526
rect 13010 3526 13112 3610
tri 13112 3526 13200 3614 sw
tri 13210 3526 13298 3614 ne
rect 13298 3610 15775 3614
rect 13298 3526 13440 3610
rect 13010 3490 13200 3526
rect 12788 3486 13200 3490
rect 12286 3438 12690 3486
rect 11786 3388 12188 3438
rect 11266 3358 11688 3388
rect 10774 3300 11168 3358
rect 10264 3260 10676 3300
tri 10676 3260 10716 3300 sw
tri 10774 3260 10814 3300 ne
rect 10814 3260 11168 3300
tri 11168 3260 11266 3358 sw
tri 11266 3260 11364 3358 ne
rect 11364 3300 11688 3358
tri 11688 3300 11776 3388 sw
tri 11786 3300 11874 3388 ne
rect 11874 3358 12188 3388
tri 12188 3358 12268 3438 sw
tri 12286 3358 12366 3438 ne
rect 12366 3388 12690 3438
tri 12690 3388 12788 3486 sw
tri 12788 3388 12886 3486 ne
rect 12886 3438 13200 3486
tri 13200 3438 13288 3526 sw
tri 13298 3438 13386 3526 ne
rect 13386 3490 13440 3526
rect 13560 3490 15775 3610
rect 13386 3438 15775 3490
rect 12886 3388 13288 3438
rect 12366 3358 12788 3388
rect 11874 3300 12268 3358
rect 11364 3260 11776 3300
tri 11776 3260 11816 3300 sw
tri 11874 3260 11914 3300 ne
rect 11914 3260 12268 3300
tri 12268 3260 12366 3358 sw
tri 12366 3260 12464 3358 ne
rect 12464 3300 12788 3358
tri 12788 3300 12876 3388 sw
tri 12886 3300 12974 3388 ne
rect 12974 3358 13288 3388
tri 13288 3358 13368 3438 sw
tri 13386 3358 13466 3438 ne
rect 13466 3358 14075 3438
rect 12974 3300 13368 3358
rect 12464 3260 12876 3300
tri 12876 3260 12916 3300 sw
tri 12974 3260 13014 3300 ne
rect 13014 3260 13368 3300
tri 13368 3260 13466 3358 sw
tri 13466 3260 13564 3358 ne
rect 13564 3338 14075 3358
rect 14175 3338 15775 3438
rect 13564 3260 15775 3338
rect -1025 3212 -284 3260
rect -1025 3112 -925 3212
rect -825 3162 -284 3212
tri -284 3162 -186 3260 sw
tri -186 3162 -88 3260 ne
rect -88 3162 266 3260
tri 266 3162 364 3260 sw
tri 364 3162 462 3260 ne
rect 462 3162 816 3260
tri 816 3162 914 3260 sw
tri 914 3162 1012 3260 ne
rect 1012 3162 1366 3260
tri 1366 3162 1464 3260 sw
tri 1464 3162 1562 3260 ne
rect 1562 3162 1916 3260
tri 1916 3162 2014 3260 sw
tri 2014 3162 2112 3260 ne
rect 2112 3162 2466 3260
tri 2466 3162 2564 3260 sw
tri 2564 3162 2662 3260 ne
rect 2662 3162 3016 3260
tri 3016 3162 3114 3260 sw
tri 3114 3162 3212 3260 ne
rect 3212 3162 3566 3260
tri 3566 3162 3664 3260 sw
tri 3664 3162 3762 3260 ne
rect 3762 3162 4116 3260
tri 4116 3162 4214 3260 sw
tri 4214 3162 4312 3260 ne
rect 4312 3162 4666 3260
tri 4666 3162 4764 3260 sw
tri 4764 3162 4862 3260 ne
rect 4862 3162 5216 3260
tri 5216 3162 5314 3260 sw
tri 5314 3162 5412 3260 ne
rect 5412 3162 5766 3260
tri 5766 3162 5864 3260 sw
tri 5864 3162 5962 3260 ne
rect 5962 3162 6316 3260
tri 6316 3162 6414 3260 sw
tri 6414 3162 6512 3260 ne
rect 6512 3162 6866 3260
tri 6866 3162 6964 3260 sw
tri 6964 3162 7062 3260 ne
rect 7062 3162 7416 3260
tri 7416 3162 7514 3260 sw
tri 7514 3162 7612 3260 ne
rect 7612 3162 7966 3260
tri 7966 3162 8064 3260 sw
tri 8064 3162 8162 3260 ne
rect 8162 3162 8516 3260
tri 8516 3162 8614 3260 sw
tri 8614 3162 8712 3260 ne
rect 8712 3162 9066 3260
tri 9066 3162 9164 3260 sw
tri 9164 3162 9262 3260 ne
rect 9262 3162 9616 3260
tri 9616 3162 9714 3260 sw
tri 9714 3162 9812 3260 ne
rect 9812 3162 10166 3260
tri 10166 3162 10264 3260 sw
tri 10264 3162 10362 3260 ne
rect 10362 3162 10716 3260
tri 10716 3162 10814 3260 sw
tri 10814 3162 10912 3260 ne
rect 10912 3162 11266 3260
tri 11266 3162 11364 3260 sw
tri 11364 3162 11462 3260 ne
rect 11462 3162 11816 3260
tri 11816 3162 11914 3260 sw
tri 11914 3162 12012 3260 ne
rect 12012 3162 12366 3260
tri 12366 3162 12464 3260 sw
tri 12464 3162 12562 3260 ne
rect 12562 3162 12916 3260
tri 12916 3162 13014 3260 sw
tri 13014 3162 13112 3260 ne
rect 13112 3162 13466 3260
tri 13466 3162 13564 3260 sw
tri 13564 3162 13662 3260 ne
rect 13662 3162 15775 3260
rect -825 3112 -186 3162
rect -1025 3064 -186 3112
tri -186 3064 -88 3162 sw
tri -88 3064 10 3162 ne
rect 10 3064 364 3162
tri 364 3064 462 3162 sw
tri 462 3064 560 3162 ne
rect 560 3064 914 3162
tri 914 3064 1012 3162 sw
tri 1012 3064 1110 3162 ne
rect 1110 3064 1464 3162
tri 1464 3064 1562 3162 sw
tri 1562 3064 1660 3162 ne
rect 1660 3064 2014 3162
tri 2014 3064 2112 3162 sw
tri 2112 3064 2210 3162 ne
rect 2210 3064 2564 3162
tri 2564 3064 2662 3162 sw
tri 2662 3064 2760 3162 ne
rect 2760 3064 3114 3162
tri 3114 3064 3212 3162 sw
tri 3212 3064 3310 3162 ne
rect 3310 3064 3664 3162
tri 3664 3064 3762 3162 sw
tri 3762 3064 3860 3162 ne
rect 3860 3064 4214 3162
tri 4214 3064 4312 3162 sw
tri 4312 3064 4410 3162 ne
rect 4410 3064 4764 3162
tri 4764 3064 4862 3162 sw
tri 4862 3064 4960 3162 ne
rect 4960 3064 5314 3162
tri 5314 3064 5412 3162 sw
tri 5412 3064 5510 3162 ne
rect 5510 3064 5864 3162
tri 5864 3064 5962 3162 sw
tri 5962 3064 6060 3162 ne
rect 6060 3064 6414 3162
tri 6414 3064 6512 3162 sw
tri 6512 3064 6610 3162 ne
rect 6610 3064 6964 3162
tri 6964 3064 7062 3162 sw
tri 7062 3064 7160 3162 ne
rect 7160 3064 7514 3162
tri 7514 3064 7612 3162 sw
tri 7612 3064 7710 3162 ne
rect 7710 3064 8064 3162
tri 8064 3064 8162 3162 sw
tri 8162 3064 8260 3162 ne
rect 8260 3064 8614 3162
tri 8614 3064 8712 3162 sw
tri 8712 3064 8810 3162 ne
rect 8810 3064 9164 3162
tri 9164 3064 9262 3162 sw
tri 9262 3064 9360 3162 ne
rect 9360 3064 9714 3162
tri 9714 3064 9812 3162 sw
tri 9812 3064 9910 3162 ne
rect 9910 3064 10264 3162
tri 10264 3064 10362 3162 sw
tri 10362 3064 10460 3162 ne
rect 10460 3064 10814 3162
tri 10814 3064 10912 3162 sw
tri 10912 3064 11010 3162 ne
rect 11010 3064 11364 3162
tri 11364 3064 11462 3162 sw
tri 11462 3064 11560 3162 ne
rect 11560 3064 11914 3162
tri 11914 3064 12012 3162 sw
tri 12012 3064 12110 3162 ne
rect 12110 3064 12464 3162
tri 12464 3064 12562 3162 sw
tri 12562 3064 12660 3162 ne
rect 12660 3064 13014 3162
tri 13014 3064 13112 3162 sw
tri 13112 3064 13210 3162 ne
rect 13210 3064 13564 3162
tri 13564 3064 13662 3162 sw
rect -1025 3060 -88 3064
rect -1025 2940 -310 3060
rect -190 2976 -88 3060
tri -88 2976 0 3064 sw
tri 10 2976 98 3064 ne
rect 98 3060 462 3064
rect 98 2976 240 3060
rect -190 2940 0 2976
rect -1025 2936 0 2940
tri 0 2936 40 2976 sw
tri 98 2936 138 2976 ne
rect 138 2940 240 2976
rect 360 2976 462 3060
tri 462 2976 550 3064 sw
tri 560 2976 648 3064 ne
rect 648 3060 1012 3064
rect 648 2976 790 3060
rect 360 2940 550 2976
rect 138 2936 550 2940
tri -412 2838 -314 2936 ne
rect -314 2838 40 2936
tri 40 2838 138 2936 sw
tri 138 2838 236 2936 ne
rect 236 2888 550 2936
tri 550 2888 638 2976 sw
tri 648 2888 736 2976 ne
rect 736 2940 790 2976
rect 910 2976 1012 3060
tri 1012 2976 1100 3064 sw
tri 1110 2976 1198 3064 ne
rect 1198 3060 1562 3064
rect 1198 2976 1340 3060
rect 910 2940 1100 2976
rect 736 2936 1100 2940
tri 1100 2936 1140 2976 sw
tri 1198 2936 1238 2976 ne
rect 1238 2940 1340 2976
rect 1460 2976 1562 3060
tri 1562 2976 1650 3064 sw
tri 1660 2976 1748 3064 ne
rect 1748 3060 2112 3064
rect 1748 2976 1890 3060
rect 1460 2940 1650 2976
rect 1238 2936 1650 2940
rect 736 2888 1140 2936
rect 236 2838 638 2888
rect -2525 2750 -412 2838
tri -412 2750 -324 2838 sw
tri -314 2750 -226 2838 ne
rect -226 2750 138 2838
tri 138 2750 226 2838 sw
tri 236 2750 324 2838 ne
rect 324 2808 638 2838
tri 638 2808 718 2888 sw
tri 736 2808 816 2888 ne
rect 816 2838 1140 2888
tri 1140 2838 1238 2936 sw
tri 1238 2838 1336 2936 ne
rect 1336 2888 1650 2936
tri 1650 2888 1738 2976 sw
tri 1748 2888 1836 2976 ne
rect 1836 2940 1890 2976
rect 2010 2976 2112 3060
tri 2112 2976 2200 3064 sw
tri 2210 2976 2298 3064 ne
rect 2298 3060 2662 3064
rect 2298 2976 2440 3060
rect 2010 2940 2200 2976
rect 1836 2936 2200 2940
tri 2200 2936 2240 2976 sw
tri 2298 2936 2338 2976 ne
rect 2338 2940 2440 2976
rect 2560 2976 2662 3060
tri 2662 2976 2750 3064 sw
tri 2760 2976 2848 3064 ne
rect 2848 3060 3212 3064
rect 2848 2976 2990 3060
rect 2560 2940 2750 2976
rect 2338 2936 2750 2940
rect 1836 2888 2240 2936
rect 1336 2838 1738 2888
rect 816 2808 1238 2838
rect 324 2750 718 2808
rect -2525 2710 -324 2750
tri -324 2710 -284 2750 sw
tri -226 2710 -186 2750 ne
rect -186 2710 226 2750
tri 226 2710 266 2750 sw
tri 324 2710 364 2750 ne
rect 364 2710 718 2750
tri 718 2710 816 2808 sw
tri 816 2710 914 2808 ne
rect 914 2750 1238 2808
tri 1238 2750 1326 2838 sw
tri 1336 2750 1424 2838 ne
rect 1424 2808 1738 2838
tri 1738 2808 1818 2888 sw
tri 1836 2808 1916 2888 ne
rect 1916 2838 2240 2888
tri 2240 2838 2338 2936 sw
tri 2338 2838 2436 2936 ne
rect 2436 2888 2750 2936
tri 2750 2888 2838 2976 sw
tri 2848 2888 2936 2976 ne
rect 2936 2940 2990 2976
rect 3110 2976 3212 3060
tri 3212 2976 3300 3064 sw
tri 3310 2976 3398 3064 ne
rect 3398 3060 3762 3064
rect 3398 2976 3540 3060
rect 3110 2940 3300 2976
rect 2936 2936 3300 2940
tri 3300 2936 3340 2976 sw
tri 3398 2936 3438 2976 ne
rect 3438 2940 3540 2976
rect 3660 2976 3762 3060
tri 3762 2976 3850 3064 sw
tri 3860 2976 3948 3064 ne
rect 3948 3060 4312 3064
rect 3948 2976 4090 3060
rect 3660 2940 3850 2976
rect 3438 2936 3850 2940
rect 2936 2888 3340 2936
rect 2436 2838 2838 2888
rect 1916 2808 2338 2838
rect 1424 2750 1818 2808
rect 914 2710 1326 2750
tri 1326 2710 1366 2750 sw
tri 1424 2710 1464 2750 ne
rect 1464 2710 1818 2750
tri 1818 2710 1916 2808 sw
tri 1916 2710 2014 2808 ne
rect 2014 2750 2338 2808
tri 2338 2750 2426 2838 sw
tri 2436 2750 2524 2838 ne
rect 2524 2808 2838 2838
tri 2838 2808 2918 2888 sw
tri 2936 2808 3016 2888 ne
rect 3016 2838 3340 2888
tri 3340 2838 3438 2936 sw
tri 3438 2838 3536 2936 ne
rect 3536 2888 3850 2936
tri 3850 2888 3938 2976 sw
tri 3948 2888 4036 2976 ne
rect 4036 2940 4090 2976
rect 4210 2976 4312 3060
tri 4312 2976 4400 3064 sw
tri 4410 2976 4498 3064 ne
rect 4498 3060 4862 3064
rect 4498 2976 4640 3060
rect 4210 2940 4400 2976
rect 4036 2936 4400 2940
tri 4400 2936 4440 2976 sw
tri 4498 2936 4538 2976 ne
rect 4538 2940 4640 2976
rect 4760 2976 4862 3060
tri 4862 2976 4950 3064 sw
tri 4960 2976 5048 3064 ne
rect 5048 3060 5412 3064
rect 5048 2976 5190 3060
rect 4760 2940 4950 2976
rect 4538 2936 4950 2940
rect 4036 2888 4440 2936
rect 3536 2838 3938 2888
rect 3016 2808 3438 2838
rect 2524 2750 2918 2808
rect 2014 2710 2426 2750
tri 2426 2710 2466 2750 sw
tri 2524 2710 2564 2750 ne
rect 2564 2710 2918 2750
tri 2918 2710 3016 2808 sw
tri 3016 2710 3114 2808 ne
rect 3114 2750 3438 2808
tri 3438 2750 3526 2838 sw
tri 3536 2750 3624 2838 ne
rect 3624 2808 3938 2838
tri 3938 2808 4018 2888 sw
tri 4036 2808 4116 2888 ne
rect 4116 2838 4440 2888
tri 4440 2838 4538 2936 sw
tri 4538 2838 4636 2936 ne
rect 4636 2888 4950 2936
tri 4950 2888 5038 2976 sw
tri 5048 2888 5136 2976 ne
rect 5136 2940 5190 2976
rect 5310 2976 5412 3060
tri 5412 2976 5500 3064 sw
tri 5510 2976 5598 3064 ne
rect 5598 3060 5962 3064
rect 5598 2976 5740 3060
rect 5310 2940 5500 2976
rect 5136 2936 5500 2940
tri 5500 2936 5540 2976 sw
tri 5598 2936 5638 2976 ne
rect 5638 2940 5740 2976
rect 5860 2976 5962 3060
tri 5962 2976 6050 3064 sw
tri 6060 2976 6148 3064 ne
rect 6148 3060 6512 3064
rect 6148 2976 6290 3060
rect 5860 2940 6050 2976
rect 5638 2936 6050 2940
rect 5136 2888 5540 2936
rect 4636 2838 5038 2888
rect 4116 2808 4538 2838
rect 3624 2750 4018 2808
rect 3114 2710 3526 2750
tri 3526 2710 3566 2750 sw
tri 3624 2710 3664 2750 ne
rect 3664 2710 4018 2750
tri 4018 2710 4116 2808 sw
tri 4116 2710 4214 2808 ne
rect 4214 2750 4538 2808
tri 4538 2750 4626 2838 sw
tri 4636 2750 4724 2838 ne
rect 4724 2808 5038 2838
tri 5038 2808 5118 2888 sw
tri 5136 2808 5216 2888 ne
rect 5216 2838 5540 2888
tri 5540 2838 5638 2936 sw
tri 5638 2838 5736 2936 ne
rect 5736 2888 6050 2936
tri 6050 2888 6138 2976 sw
tri 6148 2888 6236 2976 ne
rect 6236 2940 6290 2976
rect 6410 2976 6512 3060
tri 6512 2976 6600 3064 sw
tri 6610 2976 6698 3064 ne
rect 6698 3060 7062 3064
rect 6698 2976 6840 3060
rect 6410 2940 6600 2976
rect 6236 2936 6600 2940
tri 6600 2936 6640 2976 sw
tri 6698 2936 6738 2976 ne
rect 6738 2940 6840 2976
rect 6960 2976 7062 3060
tri 7062 2976 7150 3064 sw
tri 7160 2976 7248 3064 ne
rect 7248 3060 7612 3064
rect 7248 2976 7390 3060
rect 6960 2940 7150 2976
rect 6738 2936 7150 2940
rect 6236 2888 6640 2936
rect 5736 2838 6138 2888
rect 5216 2808 5638 2838
rect 4724 2750 5118 2808
rect 4214 2710 4626 2750
tri 4626 2710 4666 2750 sw
tri 4724 2710 4764 2750 ne
rect 4764 2710 5118 2750
tri 5118 2710 5216 2808 sw
tri 5216 2710 5314 2808 ne
rect 5314 2750 5638 2808
tri 5638 2750 5726 2838 sw
tri 5736 2750 5824 2838 ne
rect 5824 2808 6138 2838
tri 6138 2808 6218 2888 sw
tri 6236 2808 6316 2888 ne
rect 6316 2838 6640 2888
tri 6640 2838 6738 2936 sw
tri 6738 2838 6836 2936 ne
rect 6836 2888 7150 2936
tri 7150 2888 7238 2976 sw
tri 7248 2888 7336 2976 ne
rect 7336 2940 7390 2976
rect 7510 2976 7612 3060
tri 7612 2976 7700 3064 sw
tri 7710 2976 7798 3064 ne
rect 7798 3060 8162 3064
rect 7798 2976 7940 3060
rect 7510 2940 7700 2976
rect 7336 2936 7700 2940
tri 7700 2936 7740 2976 sw
tri 7798 2936 7838 2976 ne
rect 7838 2940 7940 2976
rect 8060 2976 8162 3060
tri 8162 2976 8250 3064 sw
tri 8260 2976 8348 3064 ne
rect 8348 3060 8712 3064
rect 8348 2976 8490 3060
rect 8060 2940 8250 2976
rect 7838 2936 8250 2940
rect 7336 2888 7740 2936
rect 6836 2838 7238 2888
rect 6316 2808 6738 2838
rect 5824 2750 6218 2808
rect 5314 2710 5726 2750
tri 5726 2710 5766 2750 sw
tri 5824 2710 5864 2750 ne
rect 5864 2710 6218 2750
tri 6218 2710 6316 2808 sw
tri 6316 2710 6414 2808 ne
rect 6414 2750 6738 2808
tri 6738 2750 6826 2838 sw
tri 6836 2750 6924 2838 ne
rect 6924 2808 7238 2838
tri 7238 2808 7318 2888 sw
tri 7336 2808 7416 2888 ne
rect 7416 2838 7740 2888
tri 7740 2838 7838 2936 sw
tri 7838 2838 7936 2936 ne
rect 7936 2888 8250 2936
tri 8250 2888 8338 2976 sw
tri 8348 2888 8436 2976 ne
rect 8436 2940 8490 2976
rect 8610 2976 8712 3060
tri 8712 2976 8800 3064 sw
tri 8810 2976 8898 3064 ne
rect 8898 3060 9262 3064
rect 8898 2976 9040 3060
rect 8610 2940 8800 2976
rect 8436 2936 8800 2940
tri 8800 2936 8840 2976 sw
tri 8898 2936 8938 2976 ne
rect 8938 2940 9040 2976
rect 9160 2976 9262 3060
tri 9262 2976 9350 3064 sw
tri 9360 2976 9448 3064 ne
rect 9448 3060 9812 3064
rect 9448 2976 9590 3060
rect 9160 2940 9350 2976
rect 8938 2936 9350 2940
rect 8436 2888 8840 2936
rect 7936 2838 8338 2888
rect 7416 2808 7838 2838
rect 6924 2750 7318 2808
rect 6414 2710 6826 2750
tri 6826 2710 6866 2750 sw
tri 6924 2710 6964 2750 ne
rect 6964 2710 7318 2750
tri 7318 2710 7416 2808 sw
tri 7416 2710 7514 2808 ne
rect 7514 2750 7838 2808
tri 7838 2750 7926 2838 sw
tri 7936 2750 8024 2838 ne
rect 8024 2808 8338 2838
tri 8338 2808 8418 2888 sw
tri 8436 2808 8516 2888 ne
rect 8516 2838 8840 2888
tri 8840 2838 8938 2936 sw
tri 8938 2838 9036 2936 ne
rect 9036 2888 9350 2936
tri 9350 2888 9438 2976 sw
tri 9448 2888 9536 2976 ne
rect 9536 2940 9590 2976
rect 9710 2976 9812 3060
tri 9812 2976 9900 3064 sw
tri 9910 2976 9998 3064 ne
rect 9998 3060 10362 3064
rect 9998 2976 10140 3060
rect 9710 2940 9900 2976
rect 9536 2936 9900 2940
tri 9900 2936 9940 2976 sw
tri 9998 2936 10038 2976 ne
rect 10038 2940 10140 2976
rect 10260 2976 10362 3060
tri 10362 2976 10450 3064 sw
tri 10460 2976 10548 3064 ne
rect 10548 3060 10912 3064
rect 10548 2976 10690 3060
rect 10260 2940 10450 2976
rect 10038 2936 10450 2940
rect 9536 2888 9940 2936
rect 9036 2838 9438 2888
rect 8516 2808 8938 2838
rect 8024 2750 8418 2808
rect 7514 2710 7926 2750
tri 7926 2710 7966 2750 sw
tri 8024 2710 8064 2750 ne
rect 8064 2710 8418 2750
tri 8418 2710 8516 2808 sw
tri 8516 2710 8614 2808 ne
rect 8614 2750 8938 2808
tri 8938 2750 9026 2838 sw
tri 9036 2750 9124 2838 ne
rect 9124 2808 9438 2838
tri 9438 2808 9518 2888 sw
tri 9536 2808 9616 2888 ne
rect 9616 2838 9940 2888
tri 9940 2838 10038 2936 sw
tri 10038 2838 10136 2936 ne
rect 10136 2888 10450 2936
tri 10450 2888 10538 2976 sw
tri 10548 2888 10636 2976 ne
rect 10636 2940 10690 2976
rect 10810 2976 10912 3060
tri 10912 2976 11000 3064 sw
tri 11010 2976 11098 3064 ne
rect 11098 3060 11462 3064
rect 11098 2976 11240 3060
rect 10810 2940 11000 2976
rect 10636 2936 11000 2940
tri 11000 2936 11040 2976 sw
tri 11098 2936 11138 2976 ne
rect 11138 2940 11240 2976
rect 11360 2976 11462 3060
tri 11462 2976 11550 3064 sw
tri 11560 2976 11648 3064 ne
rect 11648 3060 12012 3064
rect 11648 2976 11790 3060
rect 11360 2940 11550 2976
rect 11138 2936 11550 2940
rect 10636 2888 11040 2936
rect 10136 2838 10538 2888
rect 9616 2808 10038 2838
rect 9124 2750 9518 2808
rect 8614 2710 9026 2750
tri 9026 2710 9066 2750 sw
tri 9124 2710 9164 2750 ne
rect 9164 2710 9518 2750
tri 9518 2710 9616 2808 sw
tri 9616 2710 9714 2808 ne
rect 9714 2750 10038 2808
tri 10038 2750 10126 2838 sw
tri 10136 2750 10224 2838 ne
rect 10224 2808 10538 2838
tri 10538 2808 10618 2888 sw
tri 10636 2808 10716 2888 ne
rect 10716 2838 11040 2888
tri 11040 2838 11138 2936 sw
tri 11138 2838 11236 2936 ne
rect 11236 2888 11550 2936
tri 11550 2888 11638 2976 sw
tri 11648 2888 11736 2976 ne
rect 11736 2940 11790 2976
rect 11910 2976 12012 3060
tri 12012 2976 12100 3064 sw
tri 12110 2976 12198 3064 ne
rect 12198 3060 12562 3064
rect 12198 2976 12340 3060
rect 11910 2940 12100 2976
rect 11736 2936 12100 2940
tri 12100 2936 12140 2976 sw
tri 12198 2936 12238 2976 ne
rect 12238 2940 12340 2976
rect 12460 2976 12562 3060
tri 12562 2976 12650 3064 sw
tri 12660 2976 12748 3064 ne
rect 12748 3060 13112 3064
rect 12748 2976 12890 3060
rect 12460 2940 12650 2976
rect 12238 2936 12650 2940
rect 11736 2888 12140 2936
rect 11236 2838 11638 2888
rect 10716 2808 11138 2838
rect 10224 2750 10618 2808
rect 9714 2710 10126 2750
tri 10126 2710 10166 2750 sw
tri 10224 2710 10264 2750 ne
rect 10264 2710 10618 2750
tri 10618 2710 10716 2808 sw
tri 10716 2710 10814 2808 ne
rect 10814 2750 11138 2808
tri 11138 2750 11226 2838 sw
tri 11236 2750 11324 2838 ne
rect 11324 2808 11638 2838
tri 11638 2808 11718 2888 sw
tri 11736 2808 11816 2888 ne
rect 11816 2838 12140 2888
tri 12140 2838 12238 2936 sw
tri 12238 2838 12336 2936 ne
rect 12336 2888 12650 2936
tri 12650 2888 12738 2976 sw
tri 12748 2888 12836 2976 ne
rect 12836 2940 12890 2976
rect 13010 2976 13112 3060
tri 13112 2976 13200 3064 sw
tri 13210 2976 13298 3064 ne
rect 13298 3060 14275 3064
rect 13298 2976 13440 3060
rect 13010 2940 13200 2976
rect 12836 2936 13200 2940
tri 13200 2936 13240 2976 sw
tri 13298 2936 13338 2976 ne
rect 13338 2940 13440 2976
rect 13560 2940 14275 3060
rect 13338 2936 14275 2940
rect 12836 2888 13240 2936
rect 12336 2838 12738 2888
rect 11816 2808 12238 2838
rect 11324 2750 11718 2808
rect 10814 2710 11226 2750
tri 11226 2710 11266 2750 sw
tri 11324 2710 11364 2750 ne
rect 11364 2710 11718 2750
tri 11718 2710 11816 2808 sw
tri 11816 2710 11914 2808 ne
rect 11914 2750 12238 2808
tri 12238 2750 12326 2838 sw
tri 12336 2750 12424 2838 ne
rect 12424 2808 12738 2838
tri 12738 2808 12818 2888 sw
tri 12836 2808 12916 2888 ne
rect 12916 2838 13240 2888
tri 13240 2838 13338 2936 sw
tri 13338 2838 13436 2936 ne
rect 13436 2838 14275 2936
rect 12916 2808 13338 2838
rect 12424 2750 12818 2808
rect 11914 2710 12326 2750
tri 12326 2710 12366 2750 sw
tri 12424 2710 12464 2750 ne
rect 12464 2710 12818 2750
tri 12818 2710 12916 2808 sw
tri 12916 2710 13014 2808 ne
rect 13014 2750 13338 2808
tri 13338 2750 13426 2838 sw
tri 13436 2750 13524 2838 ne
rect 13524 2750 14275 2838
rect 13014 2710 13426 2750
tri 13426 2710 13466 2750 sw
tri 13524 2710 13564 2750 ne
rect 13564 2710 14275 2750
rect -2525 2612 -284 2710
tri -284 2612 -186 2710 sw
tri -186 2612 -88 2710 ne
rect -88 2612 266 2710
tri 266 2612 364 2710 sw
tri 364 2612 462 2710 ne
rect 462 2612 816 2710
tri 816 2612 914 2710 sw
tri 914 2612 1012 2710 ne
rect 1012 2612 1366 2710
tri 1366 2612 1464 2710 sw
tri 1464 2612 1562 2710 ne
rect 1562 2612 1916 2710
tri 1916 2612 2014 2710 sw
tri 2014 2612 2112 2710 ne
rect 2112 2612 2466 2710
tri 2466 2612 2564 2710 sw
tri 2564 2612 2662 2710 ne
rect 2662 2612 3016 2710
tri 3016 2612 3114 2710 sw
tri 3114 2612 3212 2710 ne
rect 3212 2612 3566 2710
tri 3566 2612 3664 2710 sw
tri 3664 2612 3762 2710 ne
rect 3762 2612 4116 2710
tri 4116 2612 4214 2710 sw
tri 4214 2612 4312 2710 ne
rect 4312 2612 4666 2710
tri 4666 2612 4764 2710 sw
tri 4764 2612 4862 2710 ne
rect 4862 2612 5216 2710
tri 5216 2612 5314 2710 sw
tri 5314 2612 5412 2710 ne
rect 5412 2612 5766 2710
tri 5766 2612 5864 2710 sw
tri 5864 2612 5962 2710 ne
rect 5962 2612 6316 2710
tri 6316 2612 6414 2710 sw
tri 6414 2612 6512 2710 ne
rect 6512 2612 6866 2710
tri 6866 2612 6964 2710 sw
tri 6964 2612 7062 2710 ne
rect 7062 2612 7416 2710
tri 7416 2612 7514 2710 sw
tri 7514 2612 7612 2710 ne
rect 7612 2612 7966 2710
tri 7966 2612 8064 2710 sw
tri 8064 2612 8162 2710 ne
rect 8162 2612 8516 2710
tri 8516 2612 8614 2710 sw
tri 8614 2612 8712 2710 ne
rect 8712 2612 9066 2710
tri 9066 2612 9164 2710 sw
tri 9164 2612 9262 2710 ne
rect 9262 2612 9616 2710
tri 9616 2612 9714 2710 sw
tri 9714 2612 9812 2710 ne
rect 9812 2612 10166 2710
tri 10166 2612 10264 2710 sw
tri 10264 2612 10362 2710 ne
rect 10362 2612 10716 2710
tri 10716 2612 10814 2710 sw
tri 10814 2612 10912 2710 ne
rect 10912 2612 11266 2710
tri 11266 2612 11364 2710 sw
tri 11364 2612 11462 2710 ne
rect 11462 2612 11816 2710
tri 11816 2612 11914 2710 sw
tri 11914 2612 12012 2710 ne
rect 12012 2612 12366 2710
tri 12366 2612 12464 2710 sw
tri 12464 2612 12562 2710 ne
rect 12562 2612 12916 2710
tri 12916 2612 13014 2710 sw
tri 13014 2612 13112 2710 ne
rect 13112 2612 13466 2710
tri 13466 2612 13564 2710 sw
tri 13564 2612 13662 2710 ne
rect 13662 2612 14275 2710
rect -2525 2514 -186 2612
tri -186 2514 -88 2612 sw
tri -88 2514 10 2612 ne
rect 10 2514 364 2612
tri 364 2514 462 2612 sw
tri 462 2514 560 2612 ne
rect 560 2514 914 2612
tri 914 2514 1012 2612 sw
tri 1012 2514 1110 2612 ne
rect 1110 2514 1464 2612
tri 1464 2514 1562 2612 sw
tri 1562 2514 1660 2612 ne
rect 1660 2514 2014 2612
tri 2014 2514 2112 2612 sw
tri 2112 2514 2210 2612 ne
rect 2210 2514 2564 2612
tri 2564 2514 2662 2612 sw
tri 2662 2514 2760 2612 ne
rect 2760 2514 3114 2612
tri 3114 2514 3212 2612 sw
tri 3212 2514 3310 2612 ne
rect 3310 2514 3664 2612
tri 3664 2514 3762 2612 sw
tri 3762 2514 3860 2612 ne
rect 3860 2514 4214 2612
tri 4214 2514 4312 2612 sw
tri 4312 2514 4410 2612 ne
rect 4410 2514 4764 2612
tri 4764 2514 4862 2612 sw
tri 4862 2514 4960 2612 ne
rect 4960 2514 5314 2612
tri 5314 2514 5412 2612 sw
tri 5412 2514 5510 2612 ne
rect 5510 2514 5864 2612
tri 5864 2514 5962 2612 sw
tri 5962 2514 6060 2612 ne
rect 6060 2514 6414 2612
tri 6414 2514 6512 2612 sw
tri 6512 2514 6610 2612 ne
rect 6610 2514 6964 2612
tri 6964 2514 7062 2612 sw
tri 7062 2514 7160 2612 ne
rect 7160 2514 7514 2612
tri 7514 2514 7612 2612 sw
tri 7612 2514 7710 2612 ne
rect 7710 2514 8064 2612
tri 8064 2514 8162 2612 sw
tri 8162 2514 8260 2612 ne
rect 8260 2514 8614 2612
tri 8614 2514 8712 2612 sw
tri 8712 2514 8810 2612 ne
rect 8810 2514 9164 2612
tri 9164 2514 9262 2612 sw
tri 9262 2514 9360 2612 ne
rect 9360 2514 9714 2612
tri 9714 2514 9812 2612 sw
tri 9812 2514 9910 2612 ne
rect 9910 2514 10264 2612
tri 10264 2514 10362 2612 sw
tri 10362 2514 10460 2612 ne
rect 10460 2514 10814 2612
tri 10814 2514 10912 2612 sw
tri 10912 2514 11010 2612 ne
rect 11010 2514 11364 2612
tri 11364 2514 11462 2612 sw
tri 11462 2514 11560 2612 ne
rect 11560 2514 11914 2612
tri 11914 2514 12012 2612 sw
tri 12012 2514 12110 2612 ne
rect 12110 2514 12464 2612
tri 12464 2514 12562 2612 sw
tri 12562 2514 12660 2612 ne
rect 12660 2514 13014 2612
tri 13014 2514 13112 2612 sw
tri 13112 2514 13210 2612 ne
rect 13210 2514 13564 2612
tri 13564 2514 13662 2612 sw
rect 14775 2514 15775 3162
rect -2525 2510 -88 2514
rect -2525 2390 -310 2510
rect -190 2426 -88 2510
tri -88 2426 0 2514 sw
tri 10 2426 98 2514 ne
rect 98 2510 462 2514
rect 98 2426 240 2510
rect -190 2390 0 2426
rect -2525 2386 0 2390
rect -2525 1738 -1525 2386
tri -412 2288 -314 2386 ne
rect -314 2338 0 2386
tri 0 2338 88 2426 sw
tri 98 2338 186 2426 ne
rect 186 2390 240 2426
rect 360 2426 462 2510
tri 462 2426 550 2514 sw
tri 560 2426 648 2514 ne
rect 648 2510 1012 2514
rect 648 2426 790 2510
rect 360 2390 550 2426
rect 186 2386 550 2390
tri 550 2386 590 2426 sw
tri 648 2386 688 2426 ne
rect 688 2390 790 2426
rect 910 2426 1012 2510
tri 1012 2426 1100 2514 sw
tri 1110 2426 1198 2514 ne
rect 1198 2510 1562 2514
rect 1198 2426 1340 2510
rect 910 2390 1100 2426
rect 688 2386 1100 2390
rect 186 2338 590 2386
rect -314 2288 88 2338
rect -1025 2200 -412 2288
tri -412 2200 -324 2288 sw
tri -314 2200 -226 2288 ne
rect -226 2258 88 2288
tri 88 2258 168 2338 sw
tri 186 2258 266 2338 ne
rect 266 2288 590 2338
tri 590 2288 688 2386 sw
tri 688 2288 786 2386 ne
rect 786 2338 1100 2386
tri 1100 2338 1188 2426 sw
tri 1198 2338 1286 2426 ne
rect 1286 2390 1340 2426
rect 1460 2426 1562 2510
tri 1562 2426 1650 2514 sw
tri 1660 2426 1748 2514 ne
rect 1748 2510 2112 2514
rect 1748 2426 1890 2510
rect 1460 2390 1650 2426
rect 1286 2386 1650 2390
tri 1650 2386 1690 2426 sw
tri 1748 2386 1788 2426 ne
rect 1788 2390 1890 2426
rect 2010 2426 2112 2510
tri 2112 2426 2200 2514 sw
tri 2210 2426 2298 2514 ne
rect 2298 2510 2662 2514
rect 2298 2426 2440 2510
rect 2010 2390 2200 2426
rect 1788 2386 2200 2390
rect 1286 2338 1690 2386
rect 786 2288 1188 2338
rect 266 2258 688 2288
rect -226 2200 168 2258
rect -1025 2160 -324 2200
tri -324 2160 -284 2200 sw
tri -226 2160 -186 2200 ne
rect -186 2160 168 2200
tri 168 2160 266 2258 sw
tri 266 2160 364 2258 ne
rect 364 2200 688 2258
tri 688 2200 776 2288 sw
tri 786 2200 874 2288 ne
rect 874 2258 1188 2288
tri 1188 2258 1268 2338 sw
tri 1286 2258 1366 2338 ne
rect 1366 2288 1690 2338
tri 1690 2288 1788 2386 sw
tri 1788 2288 1886 2386 ne
rect 1886 2338 2200 2386
tri 2200 2338 2288 2426 sw
tri 2298 2338 2386 2426 ne
rect 2386 2390 2440 2426
rect 2560 2426 2662 2510
tri 2662 2426 2750 2514 sw
tri 2760 2426 2848 2514 ne
rect 2848 2510 3212 2514
rect 2848 2426 2990 2510
rect 2560 2390 2750 2426
rect 2386 2386 2750 2390
tri 2750 2386 2790 2426 sw
tri 2848 2386 2888 2426 ne
rect 2888 2390 2990 2426
rect 3110 2426 3212 2510
tri 3212 2426 3300 2514 sw
tri 3310 2426 3398 2514 ne
rect 3398 2510 3762 2514
rect 3398 2426 3540 2510
rect 3110 2390 3300 2426
rect 2888 2386 3300 2390
rect 2386 2338 2790 2386
rect 1886 2288 2288 2338
rect 1366 2258 1788 2288
rect 874 2200 1268 2258
rect 364 2160 776 2200
tri 776 2160 816 2200 sw
tri 874 2160 914 2200 ne
rect 914 2160 1268 2200
tri 1268 2160 1366 2258 sw
tri 1366 2160 1464 2258 ne
rect 1464 2200 1788 2258
tri 1788 2200 1876 2288 sw
tri 1886 2200 1974 2288 ne
rect 1974 2258 2288 2288
tri 2288 2258 2368 2338 sw
tri 2386 2258 2466 2338 ne
rect 2466 2288 2790 2338
tri 2790 2288 2888 2386 sw
tri 2888 2288 2986 2386 ne
rect 2986 2338 3300 2386
tri 3300 2338 3388 2426 sw
tri 3398 2338 3486 2426 ne
rect 3486 2390 3540 2426
rect 3660 2426 3762 2510
tri 3762 2426 3850 2514 sw
tri 3860 2426 3948 2514 ne
rect 3948 2510 4312 2514
rect 3948 2426 4090 2510
rect 3660 2390 3850 2426
rect 3486 2386 3850 2390
tri 3850 2386 3890 2426 sw
tri 3948 2386 3988 2426 ne
rect 3988 2390 4090 2426
rect 4210 2426 4312 2510
tri 4312 2426 4400 2514 sw
tri 4410 2426 4498 2514 ne
rect 4498 2510 4862 2514
rect 4498 2426 4640 2510
rect 4210 2390 4400 2426
rect 3988 2386 4400 2390
rect 3486 2338 3890 2386
rect 2986 2288 3388 2338
rect 2466 2258 2888 2288
rect 1974 2200 2368 2258
rect 1464 2160 1876 2200
tri 1876 2160 1916 2200 sw
tri 1974 2160 2014 2200 ne
rect 2014 2160 2368 2200
tri 2368 2160 2466 2258 sw
tri 2466 2160 2564 2258 ne
rect 2564 2200 2888 2258
tri 2888 2200 2976 2288 sw
tri 2986 2200 3074 2288 ne
rect 3074 2258 3388 2288
tri 3388 2258 3468 2338 sw
tri 3486 2258 3566 2338 ne
rect 3566 2288 3890 2338
tri 3890 2288 3988 2386 sw
tri 3988 2288 4086 2386 ne
rect 4086 2338 4400 2386
tri 4400 2338 4488 2426 sw
tri 4498 2338 4586 2426 ne
rect 4586 2390 4640 2426
rect 4760 2426 4862 2510
tri 4862 2426 4950 2514 sw
tri 4960 2426 5048 2514 ne
rect 5048 2510 5412 2514
rect 5048 2426 5190 2510
rect 4760 2390 4950 2426
rect 4586 2386 4950 2390
tri 4950 2386 4990 2426 sw
tri 5048 2386 5088 2426 ne
rect 5088 2390 5190 2426
rect 5310 2426 5412 2510
tri 5412 2426 5500 2514 sw
tri 5510 2426 5598 2514 ne
rect 5598 2510 5962 2514
rect 5598 2426 5740 2510
rect 5310 2390 5500 2426
rect 5088 2386 5500 2390
rect 4586 2338 4990 2386
rect 4086 2288 4488 2338
rect 3566 2258 3988 2288
rect 3074 2200 3468 2258
rect 2564 2160 2976 2200
tri 2976 2160 3016 2200 sw
tri 3074 2160 3114 2200 ne
rect 3114 2160 3468 2200
tri 3468 2160 3566 2258 sw
tri 3566 2160 3664 2258 ne
rect 3664 2200 3988 2258
tri 3988 2200 4076 2288 sw
tri 4086 2200 4174 2288 ne
rect 4174 2258 4488 2288
tri 4488 2258 4568 2338 sw
tri 4586 2258 4666 2338 ne
rect 4666 2288 4990 2338
tri 4990 2288 5088 2386 sw
tri 5088 2288 5186 2386 ne
rect 5186 2338 5500 2386
tri 5500 2338 5588 2426 sw
tri 5598 2338 5686 2426 ne
rect 5686 2390 5740 2426
rect 5860 2426 5962 2510
tri 5962 2426 6050 2514 sw
tri 6060 2426 6148 2514 ne
rect 6148 2510 6512 2514
rect 6148 2426 6290 2510
rect 5860 2390 6050 2426
rect 5686 2386 6050 2390
tri 6050 2386 6090 2426 sw
tri 6148 2386 6188 2426 ne
rect 6188 2390 6290 2426
rect 6410 2426 6512 2510
tri 6512 2426 6600 2514 sw
tri 6610 2426 6698 2514 ne
rect 6698 2510 7062 2514
rect 6698 2426 6840 2510
rect 6410 2390 6600 2426
rect 6188 2386 6600 2390
rect 5686 2338 6090 2386
rect 5186 2288 5588 2338
rect 4666 2258 5088 2288
rect 4174 2200 4568 2258
rect 3664 2160 4076 2200
tri 4076 2160 4116 2200 sw
tri 4174 2160 4214 2200 ne
rect 4214 2160 4568 2200
tri 4568 2160 4666 2258 sw
tri 4666 2160 4764 2258 ne
rect 4764 2200 5088 2258
tri 5088 2200 5176 2288 sw
tri 5186 2200 5274 2288 ne
rect 5274 2258 5588 2288
tri 5588 2258 5668 2338 sw
tri 5686 2258 5766 2338 ne
rect 5766 2288 6090 2338
tri 6090 2288 6188 2386 sw
tri 6188 2288 6286 2386 ne
rect 6286 2338 6600 2386
tri 6600 2338 6688 2426 sw
tri 6698 2338 6786 2426 ne
rect 6786 2390 6840 2426
rect 6960 2426 7062 2510
tri 7062 2426 7150 2514 sw
tri 7160 2426 7248 2514 ne
rect 7248 2510 7612 2514
rect 7248 2426 7390 2510
rect 6960 2390 7150 2426
rect 6786 2386 7150 2390
tri 7150 2386 7190 2426 sw
tri 7248 2386 7288 2426 ne
rect 7288 2390 7390 2426
rect 7510 2426 7612 2510
tri 7612 2426 7700 2514 sw
tri 7710 2426 7798 2514 ne
rect 7798 2510 8162 2514
rect 7798 2426 7940 2510
rect 7510 2390 7700 2426
rect 7288 2386 7700 2390
rect 6786 2338 7190 2386
rect 6286 2288 6688 2338
rect 5766 2258 6188 2288
rect 5274 2200 5668 2258
rect 4764 2160 5176 2200
tri 5176 2160 5216 2200 sw
tri 5274 2160 5314 2200 ne
rect 5314 2160 5668 2200
tri 5668 2160 5766 2258 sw
tri 5766 2160 5864 2258 ne
rect 5864 2200 6188 2258
tri 6188 2200 6276 2288 sw
tri 6286 2200 6374 2288 ne
rect 6374 2258 6688 2288
tri 6688 2258 6768 2338 sw
tri 6786 2258 6866 2338 ne
rect 6866 2288 7190 2338
tri 7190 2288 7288 2386 sw
tri 7288 2288 7386 2386 ne
rect 7386 2338 7700 2386
tri 7700 2338 7788 2426 sw
tri 7798 2338 7886 2426 ne
rect 7886 2390 7940 2426
rect 8060 2426 8162 2510
tri 8162 2426 8250 2514 sw
tri 8260 2426 8348 2514 ne
rect 8348 2510 8712 2514
rect 8348 2426 8490 2510
rect 8060 2390 8250 2426
rect 7886 2386 8250 2390
tri 8250 2386 8290 2426 sw
tri 8348 2386 8388 2426 ne
rect 8388 2390 8490 2426
rect 8610 2426 8712 2510
tri 8712 2426 8800 2514 sw
tri 8810 2426 8898 2514 ne
rect 8898 2510 9262 2514
rect 8898 2426 9040 2510
rect 8610 2390 8800 2426
rect 8388 2386 8800 2390
rect 7886 2338 8290 2386
rect 7386 2288 7788 2338
rect 6866 2258 7288 2288
rect 6374 2200 6768 2258
rect 5864 2160 6276 2200
tri 6276 2160 6316 2200 sw
tri 6374 2160 6414 2200 ne
rect 6414 2160 6768 2200
tri 6768 2160 6866 2258 sw
tri 6866 2160 6964 2258 ne
rect 6964 2200 7288 2258
tri 7288 2200 7376 2288 sw
tri 7386 2200 7474 2288 ne
rect 7474 2258 7788 2288
tri 7788 2258 7868 2338 sw
tri 7886 2258 7966 2338 ne
rect 7966 2288 8290 2338
tri 8290 2288 8388 2386 sw
tri 8388 2288 8486 2386 ne
rect 8486 2338 8800 2386
tri 8800 2338 8888 2426 sw
tri 8898 2338 8986 2426 ne
rect 8986 2390 9040 2426
rect 9160 2426 9262 2510
tri 9262 2426 9350 2514 sw
tri 9360 2426 9448 2514 ne
rect 9448 2510 9812 2514
rect 9448 2426 9590 2510
rect 9160 2390 9350 2426
rect 8986 2386 9350 2390
tri 9350 2386 9390 2426 sw
tri 9448 2386 9488 2426 ne
rect 9488 2390 9590 2426
rect 9710 2426 9812 2510
tri 9812 2426 9900 2514 sw
tri 9910 2426 9998 2514 ne
rect 9998 2510 10362 2514
rect 9998 2426 10140 2510
rect 9710 2390 9900 2426
rect 9488 2386 9900 2390
rect 8986 2338 9390 2386
rect 8486 2288 8888 2338
rect 7966 2258 8388 2288
rect 7474 2200 7868 2258
rect 6964 2160 7376 2200
tri 7376 2160 7416 2200 sw
tri 7474 2160 7514 2200 ne
rect 7514 2160 7868 2200
tri 7868 2160 7966 2258 sw
tri 7966 2160 8064 2258 ne
rect 8064 2200 8388 2258
tri 8388 2200 8476 2288 sw
tri 8486 2200 8574 2288 ne
rect 8574 2258 8888 2288
tri 8888 2258 8968 2338 sw
tri 8986 2258 9066 2338 ne
rect 9066 2288 9390 2338
tri 9390 2288 9488 2386 sw
tri 9488 2288 9586 2386 ne
rect 9586 2338 9900 2386
tri 9900 2338 9988 2426 sw
tri 9998 2338 10086 2426 ne
rect 10086 2390 10140 2426
rect 10260 2426 10362 2510
tri 10362 2426 10450 2514 sw
tri 10460 2426 10548 2514 ne
rect 10548 2510 10912 2514
rect 10548 2426 10690 2510
rect 10260 2390 10450 2426
rect 10086 2386 10450 2390
tri 10450 2386 10490 2426 sw
tri 10548 2386 10588 2426 ne
rect 10588 2390 10690 2426
rect 10810 2426 10912 2510
tri 10912 2426 11000 2514 sw
tri 11010 2426 11098 2514 ne
rect 11098 2510 11462 2514
rect 11098 2426 11240 2510
rect 10810 2390 11000 2426
rect 10588 2386 11000 2390
rect 10086 2338 10490 2386
rect 9586 2288 9988 2338
rect 9066 2258 9488 2288
rect 8574 2200 8968 2258
rect 8064 2160 8476 2200
tri 8476 2160 8516 2200 sw
tri 8574 2160 8614 2200 ne
rect 8614 2160 8968 2200
tri 8968 2160 9066 2258 sw
tri 9066 2160 9164 2258 ne
rect 9164 2200 9488 2258
tri 9488 2200 9576 2288 sw
tri 9586 2200 9674 2288 ne
rect 9674 2258 9988 2288
tri 9988 2258 10068 2338 sw
tri 10086 2258 10166 2338 ne
rect 10166 2288 10490 2338
tri 10490 2288 10588 2386 sw
tri 10588 2288 10686 2386 ne
rect 10686 2338 11000 2386
tri 11000 2338 11088 2426 sw
tri 11098 2338 11186 2426 ne
rect 11186 2390 11240 2426
rect 11360 2426 11462 2510
tri 11462 2426 11550 2514 sw
tri 11560 2426 11648 2514 ne
rect 11648 2510 12012 2514
rect 11648 2426 11790 2510
rect 11360 2390 11550 2426
rect 11186 2386 11550 2390
tri 11550 2386 11590 2426 sw
tri 11648 2386 11688 2426 ne
rect 11688 2390 11790 2426
rect 11910 2426 12012 2510
tri 12012 2426 12100 2514 sw
tri 12110 2426 12198 2514 ne
rect 12198 2510 12562 2514
rect 12198 2426 12340 2510
rect 11910 2390 12100 2426
rect 11688 2386 12100 2390
rect 11186 2338 11590 2386
rect 10686 2288 11088 2338
rect 10166 2258 10588 2288
rect 9674 2200 10068 2258
rect 9164 2160 9576 2200
tri 9576 2160 9616 2200 sw
tri 9674 2160 9714 2200 ne
rect 9714 2160 10068 2200
tri 10068 2160 10166 2258 sw
tri 10166 2160 10264 2258 ne
rect 10264 2200 10588 2258
tri 10588 2200 10676 2288 sw
tri 10686 2200 10774 2288 ne
rect 10774 2258 11088 2288
tri 11088 2258 11168 2338 sw
tri 11186 2258 11266 2338 ne
rect 11266 2288 11590 2338
tri 11590 2288 11688 2386 sw
tri 11688 2288 11786 2386 ne
rect 11786 2338 12100 2386
tri 12100 2338 12188 2426 sw
tri 12198 2338 12286 2426 ne
rect 12286 2390 12340 2426
rect 12460 2426 12562 2510
tri 12562 2426 12650 2514 sw
tri 12660 2426 12748 2514 ne
rect 12748 2510 13112 2514
rect 12748 2426 12890 2510
rect 12460 2390 12650 2426
rect 12286 2386 12650 2390
tri 12650 2386 12690 2426 sw
tri 12748 2386 12788 2426 ne
rect 12788 2390 12890 2426
rect 13010 2426 13112 2510
tri 13112 2426 13200 2514 sw
tri 13210 2426 13298 2514 ne
rect 13298 2510 15775 2514
rect 13298 2426 13440 2510
rect 13010 2390 13200 2426
rect 12788 2386 13200 2390
rect 12286 2338 12690 2386
rect 11786 2288 12188 2338
rect 11266 2258 11688 2288
rect 10774 2200 11168 2258
rect 10264 2160 10676 2200
tri 10676 2160 10716 2200 sw
tri 10774 2160 10814 2200 ne
rect 10814 2160 11168 2200
tri 11168 2160 11266 2258 sw
tri 11266 2160 11364 2258 ne
rect 11364 2200 11688 2258
tri 11688 2200 11776 2288 sw
tri 11786 2200 11874 2288 ne
rect 11874 2258 12188 2288
tri 12188 2258 12268 2338 sw
tri 12286 2258 12366 2338 ne
rect 12366 2288 12690 2338
tri 12690 2288 12788 2386 sw
tri 12788 2288 12886 2386 ne
rect 12886 2338 13200 2386
tri 13200 2338 13288 2426 sw
tri 13298 2338 13386 2426 ne
rect 13386 2390 13440 2426
rect 13560 2390 15775 2510
rect 13386 2338 15775 2390
rect 12886 2288 13288 2338
rect 12366 2258 12788 2288
rect 11874 2200 12268 2258
rect 11364 2160 11776 2200
tri 11776 2160 11816 2200 sw
tri 11874 2160 11914 2200 ne
rect 11914 2160 12268 2200
tri 12268 2160 12366 2258 sw
tri 12366 2160 12464 2258 ne
rect 12464 2200 12788 2258
tri 12788 2200 12876 2288 sw
tri 12886 2200 12974 2288 ne
rect 12974 2258 13288 2288
tri 13288 2258 13368 2338 sw
tri 13386 2258 13466 2338 ne
rect 13466 2258 14075 2338
rect 12974 2200 13368 2258
rect 12464 2160 12876 2200
tri 12876 2160 12916 2200 sw
tri 12974 2160 13014 2200 ne
rect 13014 2160 13368 2200
tri 13368 2160 13466 2258 sw
tri 13466 2160 13564 2258 ne
rect 13564 2238 14075 2258
rect 14175 2238 15775 2338
rect 13564 2160 15775 2238
rect -1025 2112 -284 2160
rect -1025 2012 -925 2112
rect -825 2062 -284 2112
tri -284 2062 -186 2160 sw
tri -186 2062 -88 2160 ne
rect -88 2062 266 2160
tri 266 2062 364 2160 sw
tri 364 2062 462 2160 ne
rect 462 2062 816 2160
tri 816 2062 914 2160 sw
tri 914 2062 1012 2160 ne
rect 1012 2062 1366 2160
tri 1366 2062 1464 2160 sw
tri 1464 2062 1562 2160 ne
rect 1562 2062 1916 2160
tri 1916 2062 2014 2160 sw
tri 2014 2062 2112 2160 ne
rect 2112 2062 2466 2160
tri 2466 2062 2564 2160 sw
tri 2564 2062 2662 2160 ne
rect 2662 2062 3016 2160
tri 3016 2062 3114 2160 sw
tri 3114 2062 3212 2160 ne
rect 3212 2062 3566 2160
tri 3566 2062 3664 2160 sw
tri 3664 2062 3762 2160 ne
rect 3762 2062 4116 2160
tri 4116 2062 4214 2160 sw
tri 4214 2062 4312 2160 ne
rect 4312 2062 4666 2160
tri 4666 2062 4764 2160 sw
tri 4764 2062 4862 2160 ne
rect 4862 2062 5216 2160
tri 5216 2062 5314 2160 sw
tri 5314 2062 5412 2160 ne
rect 5412 2062 5766 2160
tri 5766 2062 5864 2160 sw
tri 5864 2062 5962 2160 ne
rect 5962 2062 6316 2160
tri 6316 2062 6414 2160 sw
tri 6414 2062 6512 2160 ne
rect 6512 2062 6866 2160
tri 6866 2062 6964 2160 sw
tri 6964 2062 7062 2160 ne
rect 7062 2062 7416 2160
tri 7416 2062 7514 2160 sw
tri 7514 2062 7612 2160 ne
rect 7612 2062 7966 2160
tri 7966 2062 8064 2160 sw
tri 8064 2062 8162 2160 ne
rect 8162 2062 8516 2160
tri 8516 2062 8614 2160 sw
tri 8614 2062 8712 2160 ne
rect 8712 2062 9066 2160
tri 9066 2062 9164 2160 sw
tri 9164 2062 9262 2160 ne
rect 9262 2062 9616 2160
tri 9616 2062 9714 2160 sw
tri 9714 2062 9812 2160 ne
rect 9812 2062 10166 2160
tri 10166 2062 10264 2160 sw
tri 10264 2062 10362 2160 ne
rect 10362 2062 10716 2160
tri 10716 2062 10814 2160 sw
tri 10814 2062 10912 2160 ne
rect 10912 2062 11266 2160
tri 11266 2062 11364 2160 sw
tri 11364 2062 11462 2160 ne
rect 11462 2062 11816 2160
tri 11816 2062 11914 2160 sw
tri 11914 2062 12012 2160 ne
rect 12012 2062 12366 2160
tri 12366 2062 12464 2160 sw
tri 12464 2062 12562 2160 ne
rect 12562 2062 12916 2160
tri 12916 2062 13014 2160 sw
tri 13014 2062 13112 2160 ne
rect 13112 2062 13466 2160
tri 13466 2062 13564 2160 sw
tri 13564 2062 13662 2160 ne
rect 13662 2062 15775 2160
rect -825 2012 -186 2062
rect -1025 1964 -186 2012
tri -186 1964 -88 2062 sw
tri -88 1964 10 2062 ne
rect 10 1964 364 2062
tri 364 1964 462 2062 sw
tri 462 1964 560 2062 ne
rect 560 1964 914 2062
tri 914 1964 1012 2062 sw
tri 1012 1964 1110 2062 ne
rect 1110 1964 1464 2062
tri 1464 1964 1562 2062 sw
tri 1562 1964 1660 2062 ne
rect 1660 1964 2014 2062
tri 2014 1964 2112 2062 sw
tri 2112 1964 2210 2062 ne
rect 2210 1964 2564 2062
tri 2564 1964 2662 2062 sw
tri 2662 1964 2760 2062 ne
rect 2760 1964 3114 2062
tri 3114 1964 3212 2062 sw
tri 3212 1964 3310 2062 ne
rect 3310 1964 3664 2062
tri 3664 1964 3762 2062 sw
tri 3762 1964 3860 2062 ne
rect 3860 1964 4214 2062
tri 4214 1964 4312 2062 sw
tri 4312 1964 4410 2062 ne
rect 4410 1964 4764 2062
tri 4764 1964 4862 2062 sw
tri 4862 1964 4960 2062 ne
rect 4960 1964 5314 2062
tri 5314 1964 5412 2062 sw
tri 5412 1964 5510 2062 ne
rect 5510 1964 5864 2062
tri 5864 1964 5962 2062 sw
tri 5962 1964 6060 2062 ne
rect 6060 1964 6414 2062
tri 6414 1964 6512 2062 sw
tri 6512 1964 6610 2062 ne
rect 6610 1964 6964 2062
tri 6964 1964 7062 2062 sw
tri 7062 1964 7160 2062 ne
rect 7160 1964 7514 2062
tri 7514 1964 7612 2062 sw
tri 7612 1964 7710 2062 ne
rect 7710 1964 8064 2062
tri 8064 1964 8162 2062 sw
tri 8162 1964 8260 2062 ne
rect 8260 1964 8614 2062
tri 8614 1964 8712 2062 sw
tri 8712 1964 8810 2062 ne
rect 8810 1964 9164 2062
tri 9164 1964 9262 2062 sw
tri 9262 1964 9360 2062 ne
rect 9360 1964 9714 2062
tri 9714 1964 9812 2062 sw
tri 9812 1964 9910 2062 ne
rect 9910 1964 10264 2062
tri 10264 1964 10362 2062 sw
tri 10362 1964 10460 2062 ne
rect 10460 1964 10814 2062
tri 10814 1964 10912 2062 sw
tri 10912 1964 11010 2062 ne
rect 11010 1964 11364 2062
tri 11364 1964 11462 2062 sw
tri 11462 1964 11560 2062 ne
rect 11560 1964 11914 2062
tri 11914 1964 12012 2062 sw
tri 12012 1964 12110 2062 ne
rect 12110 1964 12464 2062
tri 12464 1964 12562 2062 sw
tri 12562 1964 12660 2062 ne
rect 12660 1964 13014 2062
tri 13014 1964 13112 2062 sw
tri 13112 1964 13210 2062 ne
rect 13210 1964 13564 2062
tri 13564 1964 13662 2062 sw
rect -1025 1960 -88 1964
rect -1025 1840 -310 1960
rect -190 1876 -88 1960
tri -88 1876 0 1964 sw
tri 10 1876 98 1964 ne
rect 98 1960 462 1964
rect 98 1876 240 1960
rect -190 1840 0 1876
rect -1025 1836 0 1840
tri 0 1836 40 1876 sw
tri 98 1836 138 1876 ne
rect 138 1840 240 1876
rect 360 1876 462 1960
tri 462 1876 550 1964 sw
tri 560 1876 648 1964 ne
rect 648 1960 1012 1964
rect 648 1876 790 1960
rect 360 1840 550 1876
rect 138 1836 550 1840
tri -412 1738 -314 1836 ne
rect -314 1738 40 1836
tri 40 1738 138 1836 sw
tri 138 1738 236 1836 ne
rect 236 1788 550 1836
tri 550 1788 638 1876 sw
tri 648 1788 736 1876 ne
rect 736 1840 790 1876
rect 910 1876 1012 1960
tri 1012 1876 1100 1964 sw
tri 1110 1876 1198 1964 ne
rect 1198 1960 1562 1964
rect 1198 1876 1340 1960
rect 910 1840 1100 1876
rect 736 1836 1100 1840
tri 1100 1836 1140 1876 sw
tri 1198 1836 1238 1876 ne
rect 1238 1840 1340 1876
rect 1460 1876 1562 1960
tri 1562 1876 1650 1964 sw
tri 1660 1876 1748 1964 ne
rect 1748 1960 2112 1964
rect 1748 1876 1890 1960
rect 1460 1840 1650 1876
rect 1238 1836 1650 1840
rect 736 1788 1140 1836
rect 236 1738 638 1788
rect -2525 1650 -412 1738
tri -412 1650 -324 1738 sw
tri -314 1650 -226 1738 ne
rect -226 1650 138 1738
tri 138 1650 226 1738 sw
tri 236 1650 324 1738 ne
rect 324 1708 638 1738
tri 638 1708 718 1788 sw
tri 736 1708 816 1788 ne
rect 816 1738 1140 1788
tri 1140 1738 1238 1836 sw
tri 1238 1738 1336 1836 ne
rect 1336 1788 1650 1836
tri 1650 1788 1738 1876 sw
tri 1748 1788 1836 1876 ne
rect 1836 1840 1890 1876
rect 2010 1876 2112 1960
tri 2112 1876 2200 1964 sw
tri 2210 1876 2298 1964 ne
rect 2298 1960 2662 1964
rect 2298 1876 2440 1960
rect 2010 1840 2200 1876
rect 1836 1836 2200 1840
tri 2200 1836 2240 1876 sw
tri 2298 1836 2338 1876 ne
rect 2338 1840 2440 1876
rect 2560 1876 2662 1960
tri 2662 1876 2750 1964 sw
tri 2760 1876 2848 1964 ne
rect 2848 1960 3212 1964
rect 2848 1876 2990 1960
rect 2560 1840 2750 1876
rect 2338 1836 2750 1840
rect 1836 1788 2240 1836
rect 1336 1738 1738 1788
rect 816 1708 1238 1738
rect 324 1650 718 1708
rect -2525 1610 -324 1650
tri -324 1610 -284 1650 sw
tri -226 1610 -186 1650 ne
rect -186 1610 226 1650
tri 226 1610 266 1650 sw
tri 324 1610 364 1650 ne
rect 364 1610 718 1650
tri 718 1610 816 1708 sw
tri 816 1610 914 1708 ne
rect 914 1650 1238 1708
tri 1238 1650 1326 1738 sw
tri 1336 1650 1424 1738 ne
rect 1424 1708 1738 1738
tri 1738 1708 1818 1788 sw
tri 1836 1708 1916 1788 ne
rect 1916 1738 2240 1788
tri 2240 1738 2338 1836 sw
tri 2338 1738 2436 1836 ne
rect 2436 1788 2750 1836
tri 2750 1788 2838 1876 sw
tri 2848 1788 2936 1876 ne
rect 2936 1840 2990 1876
rect 3110 1876 3212 1960
tri 3212 1876 3300 1964 sw
tri 3310 1876 3398 1964 ne
rect 3398 1960 3762 1964
rect 3398 1876 3540 1960
rect 3110 1840 3300 1876
rect 2936 1836 3300 1840
tri 3300 1836 3340 1876 sw
tri 3398 1836 3438 1876 ne
rect 3438 1840 3540 1876
rect 3660 1876 3762 1960
tri 3762 1876 3850 1964 sw
tri 3860 1876 3948 1964 ne
rect 3948 1960 4312 1964
rect 3948 1876 4090 1960
rect 3660 1840 3850 1876
rect 3438 1836 3850 1840
rect 2936 1788 3340 1836
rect 2436 1738 2838 1788
rect 1916 1708 2338 1738
rect 1424 1650 1818 1708
rect 914 1610 1326 1650
tri 1326 1610 1366 1650 sw
tri 1424 1610 1464 1650 ne
rect 1464 1610 1818 1650
tri 1818 1610 1916 1708 sw
tri 1916 1610 2014 1708 ne
rect 2014 1650 2338 1708
tri 2338 1650 2426 1738 sw
tri 2436 1650 2524 1738 ne
rect 2524 1708 2838 1738
tri 2838 1708 2918 1788 sw
tri 2936 1708 3016 1788 ne
rect 3016 1738 3340 1788
tri 3340 1738 3438 1836 sw
tri 3438 1738 3536 1836 ne
rect 3536 1788 3850 1836
tri 3850 1788 3938 1876 sw
tri 3948 1788 4036 1876 ne
rect 4036 1840 4090 1876
rect 4210 1876 4312 1960
tri 4312 1876 4400 1964 sw
tri 4410 1876 4498 1964 ne
rect 4498 1960 4862 1964
rect 4498 1876 4640 1960
rect 4210 1840 4400 1876
rect 4036 1836 4400 1840
tri 4400 1836 4440 1876 sw
tri 4498 1836 4538 1876 ne
rect 4538 1840 4640 1876
rect 4760 1876 4862 1960
tri 4862 1876 4950 1964 sw
tri 4960 1876 5048 1964 ne
rect 5048 1960 5412 1964
rect 5048 1876 5190 1960
rect 4760 1840 4950 1876
rect 4538 1836 4950 1840
rect 4036 1788 4440 1836
rect 3536 1738 3938 1788
rect 3016 1708 3438 1738
rect 2524 1650 2918 1708
rect 2014 1610 2426 1650
tri 2426 1610 2466 1650 sw
tri 2524 1610 2564 1650 ne
rect 2564 1610 2918 1650
tri 2918 1610 3016 1708 sw
tri 3016 1610 3114 1708 ne
rect 3114 1650 3438 1708
tri 3438 1650 3526 1738 sw
tri 3536 1650 3624 1738 ne
rect 3624 1708 3938 1738
tri 3938 1708 4018 1788 sw
tri 4036 1708 4116 1788 ne
rect 4116 1738 4440 1788
tri 4440 1738 4538 1836 sw
tri 4538 1738 4636 1836 ne
rect 4636 1788 4950 1836
tri 4950 1788 5038 1876 sw
tri 5048 1788 5136 1876 ne
rect 5136 1840 5190 1876
rect 5310 1876 5412 1960
tri 5412 1876 5500 1964 sw
tri 5510 1876 5598 1964 ne
rect 5598 1960 5962 1964
rect 5598 1876 5740 1960
rect 5310 1840 5500 1876
rect 5136 1836 5500 1840
tri 5500 1836 5540 1876 sw
tri 5598 1836 5638 1876 ne
rect 5638 1840 5740 1876
rect 5860 1876 5962 1960
tri 5962 1876 6050 1964 sw
tri 6060 1876 6148 1964 ne
rect 6148 1960 6512 1964
rect 6148 1876 6290 1960
rect 5860 1840 6050 1876
rect 5638 1836 6050 1840
rect 5136 1788 5540 1836
rect 4636 1738 5038 1788
rect 4116 1708 4538 1738
rect 3624 1650 4018 1708
rect 3114 1610 3526 1650
tri 3526 1610 3566 1650 sw
tri 3624 1610 3664 1650 ne
rect 3664 1610 4018 1650
tri 4018 1610 4116 1708 sw
tri 4116 1610 4214 1708 ne
rect 4214 1650 4538 1708
tri 4538 1650 4626 1738 sw
tri 4636 1650 4724 1738 ne
rect 4724 1708 5038 1738
tri 5038 1708 5118 1788 sw
tri 5136 1708 5216 1788 ne
rect 5216 1738 5540 1788
tri 5540 1738 5638 1836 sw
tri 5638 1738 5736 1836 ne
rect 5736 1788 6050 1836
tri 6050 1788 6138 1876 sw
tri 6148 1788 6236 1876 ne
rect 6236 1840 6290 1876
rect 6410 1876 6512 1960
tri 6512 1876 6600 1964 sw
tri 6610 1876 6698 1964 ne
rect 6698 1960 7062 1964
rect 6698 1876 6840 1960
rect 6410 1840 6600 1876
rect 6236 1836 6600 1840
tri 6600 1836 6640 1876 sw
tri 6698 1836 6738 1876 ne
rect 6738 1840 6840 1876
rect 6960 1876 7062 1960
tri 7062 1876 7150 1964 sw
tri 7160 1876 7248 1964 ne
rect 7248 1960 7612 1964
rect 7248 1876 7390 1960
rect 6960 1840 7150 1876
rect 6738 1836 7150 1840
rect 6236 1788 6640 1836
rect 5736 1738 6138 1788
rect 5216 1708 5638 1738
rect 4724 1650 5118 1708
rect 4214 1610 4626 1650
tri 4626 1610 4666 1650 sw
tri 4724 1610 4764 1650 ne
rect 4764 1610 5118 1650
tri 5118 1610 5216 1708 sw
tri 5216 1610 5314 1708 ne
rect 5314 1650 5638 1708
tri 5638 1650 5726 1738 sw
tri 5736 1650 5824 1738 ne
rect 5824 1708 6138 1738
tri 6138 1708 6218 1788 sw
tri 6236 1708 6316 1788 ne
rect 6316 1738 6640 1788
tri 6640 1738 6738 1836 sw
tri 6738 1738 6836 1836 ne
rect 6836 1788 7150 1836
tri 7150 1788 7238 1876 sw
tri 7248 1788 7336 1876 ne
rect 7336 1840 7390 1876
rect 7510 1876 7612 1960
tri 7612 1876 7700 1964 sw
tri 7710 1876 7798 1964 ne
rect 7798 1960 8162 1964
rect 7798 1876 7940 1960
rect 7510 1840 7700 1876
rect 7336 1836 7700 1840
tri 7700 1836 7740 1876 sw
tri 7798 1836 7838 1876 ne
rect 7838 1840 7940 1876
rect 8060 1876 8162 1960
tri 8162 1876 8250 1964 sw
tri 8260 1876 8348 1964 ne
rect 8348 1960 8712 1964
rect 8348 1876 8490 1960
rect 8060 1840 8250 1876
rect 7838 1836 8250 1840
rect 7336 1788 7740 1836
rect 6836 1738 7238 1788
rect 6316 1708 6738 1738
rect 5824 1650 6218 1708
rect 5314 1610 5726 1650
tri 5726 1610 5766 1650 sw
tri 5824 1610 5864 1650 ne
rect 5864 1610 6218 1650
tri 6218 1610 6316 1708 sw
tri 6316 1610 6414 1708 ne
rect 6414 1650 6738 1708
tri 6738 1650 6826 1738 sw
tri 6836 1650 6924 1738 ne
rect 6924 1708 7238 1738
tri 7238 1708 7318 1788 sw
tri 7336 1708 7416 1788 ne
rect 7416 1738 7740 1788
tri 7740 1738 7838 1836 sw
tri 7838 1738 7936 1836 ne
rect 7936 1788 8250 1836
tri 8250 1788 8338 1876 sw
tri 8348 1788 8436 1876 ne
rect 8436 1840 8490 1876
rect 8610 1876 8712 1960
tri 8712 1876 8800 1964 sw
tri 8810 1876 8898 1964 ne
rect 8898 1960 9262 1964
rect 8898 1876 9040 1960
rect 8610 1840 8800 1876
rect 8436 1836 8800 1840
tri 8800 1836 8840 1876 sw
tri 8898 1836 8938 1876 ne
rect 8938 1840 9040 1876
rect 9160 1876 9262 1960
tri 9262 1876 9350 1964 sw
tri 9360 1876 9448 1964 ne
rect 9448 1960 9812 1964
rect 9448 1876 9590 1960
rect 9160 1840 9350 1876
rect 8938 1836 9350 1840
rect 8436 1788 8840 1836
rect 7936 1738 8338 1788
rect 7416 1708 7838 1738
rect 6924 1650 7318 1708
rect 6414 1610 6826 1650
tri 6826 1610 6866 1650 sw
tri 6924 1610 6964 1650 ne
rect 6964 1610 7318 1650
tri 7318 1610 7416 1708 sw
tri 7416 1610 7514 1708 ne
rect 7514 1650 7838 1708
tri 7838 1650 7926 1738 sw
tri 7936 1650 8024 1738 ne
rect 8024 1708 8338 1738
tri 8338 1708 8418 1788 sw
tri 8436 1708 8516 1788 ne
rect 8516 1738 8840 1788
tri 8840 1738 8938 1836 sw
tri 8938 1738 9036 1836 ne
rect 9036 1788 9350 1836
tri 9350 1788 9438 1876 sw
tri 9448 1788 9536 1876 ne
rect 9536 1840 9590 1876
rect 9710 1876 9812 1960
tri 9812 1876 9900 1964 sw
tri 9910 1876 9998 1964 ne
rect 9998 1960 10362 1964
rect 9998 1876 10140 1960
rect 9710 1840 9900 1876
rect 9536 1836 9900 1840
tri 9900 1836 9940 1876 sw
tri 9998 1836 10038 1876 ne
rect 10038 1840 10140 1876
rect 10260 1876 10362 1960
tri 10362 1876 10450 1964 sw
tri 10460 1876 10548 1964 ne
rect 10548 1960 10912 1964
rect 10548 1876 10690 1960
rect 10260 1840 10450 1876
rect 10038 1836 10450 1840
rect 9536 1788 9940 1836
rect 9036 1738 9438 1788
rect 8516 1708 8938 1738
rect 8024 1650 8418 1708
rect 7514 1610 7926 1650
tri 7926 1610 7966 1650 sw
tri 8024 1610 8064 1650 ne
rect 8064 1610 8418 1650
tri 8418 1610 8516 1708 sw
tri 8516 1610 8614 1708 ne
rect 8614 1650 8938 1708
tri 8938 1650 9026 1738 sw
tri 9036 1650 9124 1738 ne
rect 9124 1708 9438 1738
tri 9438 1708 9518 1788 sw
tri 9536 1708 9616 1788 ne
rect 9616 1738 9940 1788
tri 9940 1738 10038 1836 sw
tri 10038 1738 10136 1836 ne
rect 10136 1788 10450 1836
tri 10450 1788 10538 1876 sw
tri 10548 1788 10636 1876 ne
rect 10636 1840 10690 1876
rect 10810 1876 10912 1960
tri 10912 1876 11000 1964 sw
tri 11010 1876 11098 1964 ne
rect 11098 1960 11462 1964
rect 11098 1876 11240 1960
rect 10810 1840 11000 1876
rect 10636 1836 11000 1840
tri 11000 1836 11040 1876 sw
tri 11098 1836 11138 1876 ne
rect 11138 1840 11240 1876
rect 11360 1876 11462 1960
tri 11462 1876 11550 1964 sw
tri 11560 1876 11648 1964 ne
rect 11648 1960 12012 1964
rect 11648 1876 11790 1960
rect 11360 1840 11550 1876
rect 11138 1836 11550 1840
rect 10636 1788 11040 1836
rect 10136 1738 10538 1788
rect 9616 1708 10038 1738
rect 9124 1650 9518 1708
rect 8614 1610 9026 1650
tri 9026 1610 9066 1650 sw
tri 9124 1610 9164 1650 ne
rect 9164 1610 9518 1650
tri 9518 1610 9616 1708 sw
tri 9616 1610 9714 1708 ne
rect 9714 1650 10038 1708
tri 10038 1650 10126 1738 sw
tri 10136 1650 10224 1738 ne
rect 10224 1708 10538 1738
tri 10538 1708 10618 1788 sw
tri 10636 1708 10716 1788 ne
rect 10716 1738 11040 1788
tri 11040 1738 11138 1836 sw
tri 11138 1738 11236 1836 ne
rect 11236 1788 11550 1836
tri 11550 1788 11638 1876 sw
tri 11648 1788 11736 1876 ne
rect 11736 1840 11790 1876
rect 11910 1876 12012 1960
tri 12012 1876 12100 1964 sw
tri 12110 1876 12198 1964 ne
rect 12198 1960 12562 1964
rect 12198 1876 12340 1960
rect 11910 1840 12100 1876
rect 11736 1836 12100 1840
tri 12100 1836 12140 1876 sw
tri 12198 1836 12238 1876 ne
rect 12238 1840 12340 1876
rect 12460 1876 12562 1960
tri 12562 1876 12650 1964 sw
tri 12660 1876 12748 1964 ne
rect 12748 1960 13112 1964
rect 12748 1876 12890 1960
rect 12460 1840 12650 1876
rect 12238 1836 12650 1840
rect 11736 1788 12140 1836
rect 11236 1738 11638 1788
rect 10716 1708 11138 1738
rect 10224 1650 10618 1708
rect 9714 1610 10126 1650
tri 10126 1610 10166 1650 sw
tri 10224 1610 10264 1650 ne
rect 10264 1610 10618 1650
tri 10618 1610 10716 1708 sw
tri 10716 1610 10814 1708 ne
rect 10814 1650 11138 1708
tri 11138 1650 11226 1738 sw
tri 11236 1650 11324 1738 ne
rect 11324 1708 11638 1738
tri 11638 1708 11718 1788 sw
tri 11736 1708 11816 1788 ne
rect 11816 1738 12140 1788
tri 12140 1738 12238 1836 sw
tri 12238 1738 12336 1836 ne
rect 12336 1788 12650 1836
tri 12650 1788 12738 1876 sw
tri 12748 1788 12836 1876 ne
rect 12836 1840 12890 1876
rect 13010 1876 13112 1960
tri 13112 1876 13200 1964 sw
tri 13210 1876 13298 1964 ne
rect 13298 1960 14275 1964
rect 13298 1876 13440 1960
rect 13010 1840 13200 1876
rect 12836 1836 13200 1840
tri 13200 1836 13240 1876 sw
tri 13298 1836 13338 1876 ne
rect 13338 1840 13440 1876
rect 13560 1840 14275 1960
rect 13338 1836 14275 1840
rect 12836 1788 13240 1836
rect 12336 1738 12738 1788
rect 11816 1708 12238 1738
rect 11324 1650 11718 1708
rect 10814 1610 11226 1650
tri 11226 1610 11266 1650 sw
tri 11324 1610 11364 1650 ne
rect 11364 1610 11718 1650
tri 11718 1610 11816 1708 sw
tri 11816 1610 11914 1708 ne
rect 11914 1650 12238 1708
tri 12238 1650 12326 1738 sw
tri 12336 1650 12424 1738 ne
rect 12424 1708 12738 1738
tri 12738 1708 12818 1788 sw
tri 12836 1708 12916 1788 ne
rect 12916 1738 13240 1788
tri 13240 1738 13338 1836 sw
tri 13338 1738 13436 1836 ne
rect 13436 1738 14275 1836
rect 12916 1708 13338 1738
rect 12424 1650 12818 1708
rect 11914 1610 12326 1650
tri 12326 1610 12366 1650 sw
tri 12424 1610 12464 1650 ne
rect 12464 1610 12818 1650
tri 12818 1610 12916 1708 sw
tri 12916 1610 13014 1708 ne
rect 13014 1650 13338 1708
tri 13338 1650 13426 1738 sw
tri 13436 1650 13524 1738 ne
rect 13524 1650 14275 1738
rect 13014 1610 13426 1650
tri 13426 1610 13466 1650 sw
tri 13524 1610 13564 1650 ne
rect 13564 1610 14275 1650
rect -2525 1512 -284 1610
tri -284 1512 -186 1610 sw
tri -186 1512 -88 1610 ne
rect -88 1512 266 1610
tri 266 1512 364 1610 sw
tri 364 1512 462 1610 ne
rect 462 1512 816 1610
tri 816 1512 914 1610 sw
tri 914 1512 1012 1610 ne
rect 1012 1512 1366 1610
tri 1366 1512 1464 1610 sw
tri 1464 1512 1562 1610 ne
rect 1562 1512 1916 1610
tri 1916 1512 2014 1610 sw
tri 2014 1512 2112 1610 ne
rect 2112 1512 2466 1610
tri 2466 1512 2564 1610 sw
tri 2564 1512 2662 1610 ne
rect 2662 1512 3016 1610
tri 3016 1512 3114 1610 sw
tri 3114 1512 3212 1610 ne
rect 3212 1512 3566 1610
tri 3566 1512 3664 1610 sw
tri 3664 1512 3762 1610 ne
rect 3762 1512 4116 1610
tri 4116 1512 4214 1610 sw
tri 4214 1512 4312 1610 ne
rect 4312 1512 4666 1610
tri 4666 1512 4764 1610 sw
tri 4764 1512 4862 1610 ne
rect 4862 1512 5216 1610
tri 5216 1512 5314 1610 sw
tri 5314 1512 5412 1610 ne
rect 5412 1512 5766 1610
tri 5766 1512 5864 1610 sw
tri 5864 1512 5962 1610 ne
rect 5962 1512 6316 1610
tri 6316 1512 6414 1610 sw
tri 6414 1512 6512 1610 ne
rect 6512 1512 6866 1610
tri 6866 1512 6964 1610 sw
tri 6964 1512 7062 1610 ne
rect 7062 1512 7416 1610
tri 7416 1512 7514 1610 sw
tri 7514 1512 7612 1610 ne
rect 7612 1512 7966 1610
tri 7966 1512 8064 1610 sw
tri 8064 1512 8162 1610 ne
rect 8162 1512 8516 1610
tri 8516 1512 8614 1610 sw
tri 8614 1512 8712 1610 ne
rect 8712 1512 9066 1610
tri 9066 1512 9164 1610 sw
tri 9164 1512 9262 1610 ne
rect 9262 1512 9616 1610
tri 9616 1512 9714 1610 sw
tri 9714 1512 9812 1610 ne
rect 9812 1512 10166 1610
tri 10166 1512 10264 1610 sw
tri 10264 1512 10362 1610 ne
rect 10362 1512 10716 1610
tri 10716 1512 10814 1610 sw
tri 10814 1512 10912 1610 ne
rect 10912 1512 11266 1610
tri 11266 1512 11364 1610 sw
tri 11364 1512 11462 1610 ne
rect 11462 1512 11816 1610
tri 11816 1512 11914 1610 sw
tri 11914 1512 12012 1610 ne
rect 12012 1512 12366 1610
tri 12366 1512 12464 1610 sw
tri 12464 1512 12562 1610 ne
rect 12562 1512 12916 1610
tri 12916 1512 13014 1610 sw
tri 13014 1512 13112 1610 ne
rect 13112 1512 13466 1610
tri 13466 1512 13564 1610 sw
tri 13564 1512 13662 1610 ne
rect 13662 1512 14275 1610
rect -2525 1414 -186 1512
tri -186 1414 -88 1512 sw
tri -88 1414 10 1512 ne
rect 10 1414 364 1512
tri 364 1414 462 1512 sw
tri 462 1414 560 1512 ne
rect 560 1414 914 1512
tri 914 1414 1012 1512 sw
tri 1012 1414 1110 1512 ne
rect 1110 1414 1464 1512
tri 1464 1414 1562 1512 sw
tri 1562 1414 1660 1512 ne
rect 1660 1414 2014 1512
tri 2014 1414 2112 1512 sw
tri 2112 1414 2210 1512 ne
rect 2210 1414 2564 1512
tri 2564 1414 2662 1512 sw
tri 2662 1414 2760 1512 ne
rect 2760 1414 3114 1512
tri 3114 1414 3212 1512 sw
tri 3212 1414 3310 1512 ne
rect 3310 1414 3664 1512
tri 3664 1414 3762 1512 sw
tri 3762 1414 3860 1512 ne
rect 3860 1414 4214 1512
tri 4214 1414 4312 1512 sw
tri 4312 1414 4410 1512 ne
rect 4410 1414 4764 1512
tri 4764 1414 4862 1512 sw
tri 4862 1414 4960 1512 ne
rect 4960 1414 5314 1512
tri 5314 1414 5412 1512 sw
tri 5412 1414 5510 1512 ne
rect 5510 1414 5864 1512
tri 5864 1414 5962 1512 sw
tri 5962 1414 6060 1512 ne
rect 6060 1414 6414 1512
tri 6414 1414 6512 1512 sw
tri 6512 1414 6610 1512 ne
rect 6610 1414 6964 1512
tri 6964 1414 7062 1512 sw
tri 7062 1414 7160 1512 ne
rect 7160 1414 7514 1512
tri 7514 1414 7612 1512 sw
tri 7612 1414 7710 1512 ne
rect 7710 1414 8064 1512
tri 8064 1414 8162 1512 sw
tri 8162 1414 8260 1512 ne
rect 8260 1414 8614 1512
tri 8614 1414 8712 1512 sw
tri 8712 1414 8810 1512 ne
rect 8810 1414 9164 1512
tri 9164 1414 9262 1512 sw
tri 9262 1414 9360 1512 ne
rect 9360 1414 9714 1512
tri 9714 1414 9812 1512 sw
tri 9812 1414 9910 1512 ne
rect 9910 1414 10264 1512
tri 10264 1414 10362 1512 sw
tri 10362 1414 10460 1512 ne
rect 10460 1414 10814 1512
tri 10814 1414 10912 1512 sw
tri 10912 1414 11010 1512 ne
rect 11010 1414 11364 1512
tri 11364 1414 11462 1512 sw
tri 11462 1414 11560 1512 ne
rect 11560 1414 11914 1512
tri 11914 1414 12012 1512 sw
tri 12012 1414 12110 1512 ne
rect 12110 1414 12464 1512
tri 12464 1414 12562 1512 sw
tri 12562 1414 12660 1512 ne
rect 12660 1414 13014 1512
tri 13014 1414 13112 1512 sw
tri 13112 1414 13210 1512 ne
rect 13210 1414 13564 1512
tri 13564 1414 13662 1512 sw
rect 14775 1414 15775 2062
rect -2525 1410 -88 1414
rect -2525 1290 -310 1410
rect -190 1326 -88 1410
tri -88 1326 0 1414 sw
tri 10 1326 98 1414 ne
rect 98 1410 462 1414
rect 98 1326 240 1410
rect -190 1290 0 1326
rect -2525 1286 0 1290
rect -2525 638 -1525 1286
tri -412 1188 -314 1286 ne
rect -314 1238 0 1286
tri 0 1238 88 1326 sw
tri 98 1238 186 1326 ne
rect 186 1290 240 1326
rect 360 1326 462 1410
tri 462 1326 550 1414 sw
tri 560 1326 648 1414 ne
rect 648 1410 1012 1414
rect 648 1326 790 1410
rect 360 1290 550 1326
rect 186 1286 550 1290
tri 550 1286 590 1326 sw
tri 648 1286 688 1326 ne
rect 688 1290 790 1326
rect 910 1326 1012 1410
tri 1012 1326 1100 1414 sw
tri 1110 1326 1198 1414 ne
rect 1198 1410 1562 1414
rect 1198 1326 1340 1410
rect 910 1290 1100 1326
rect 688 1286 1100 1290
rect 186 1238 590 1286
rect -314 1188 88 1238
rect -1025 1100 -412 1188
tri -412 1100 -324 1188 sw
tri -314 1100 -226 1188 ne
rect -226 1158 88 1188
tri 88 1158 168 1238 sw
tri 186 1158 266 1238 ne
rect 266 1188 590 1238
tri 590 1188 688 1286 sw
tri 688 1188 786 1286 ne
rect 786 1238 1100 1286
tri 1100 1238 1188 1326 sw
tri 1198 1238 1286 1326 ne
rect 1286 1290 1340 1326
rect 1460 1326 1562 1410
tri 1562 1326 1650 1414 sw
tri 1660 1326 1748 1414 ne
rect 1748 1410 2112 1414
rect 1748 1326 1890 1410
rect 1460 1290 1650 1326
rect 1286 1286 1650 1290
tri 1650 1286 1690 1326 sw
tri 1748 1286 1788 1326 ne
rect 1788 1290 1890 1326
rect 2010 1326 2112 1410
tri 2112 1326 2200 1414 sw
tri 2210 1326 2298 1414 ne
rect 2298 1410 2662 1414
rect 2298 1326 2440 1410
rect 2010 1290 2200 1326
rect 1788 1286 2200 1290
rect 1286 1238 1690 1286
rect 786 1188 1188 1238
rect 266 1158 688 1188
rect -226 1100 168 1158
rect -1025 1060 -324 1100
tri -324 1060 -284 1100 sw
tri -226 1060 -186 1100 ne
rect -186 1060 168 1100
tri 168 1060 266 1158 sw
tri 266 1060 364 1158 ne
rect 364 1100 688 1158
tri 688 1100 776 1188 sw
tri 786 1100 874 1188 ne
rect 874 1158 1188 1188
tri 1188 1158 1268 1238 sw
tri 1286 1158 1366 1238 ne
rect 1366 1188 1690 1238
tri 1690 1188 1788 1286 sw
tri 1788 1188 1886 1286 ne
rect 1886 1238 2200 1286
tri 2200 1238 2288 1326 sw
tri 2298 1238 2386 1326 ne
rect 2386 1290 2440 1326
rect 2560 1326 2662 1410
tri 2662 1326 2750 1414 sw
tri 2760 1326 2848 1414 ne
rect 2848 1410 3212 1414
rect 2848 1326 2990 1410
rect 2560 1290 2750 1326
rect 2386 1286 2750 1290
tri 2750 1286 2790 1326 sw
tri 2848 1286 2888 1326 ne
rect 2888 1290 2990 1326
rect 3110 1326 3212 1410
tri 3212 1326 3300 1414 sw
tri 3310 1326 3398 1414 ne
rect 3398 1410 3762 1414
rect 3398 1326 3540 1410
rect 3110 1290 3300 1326
rect 2888 1286 3300 1290
rect 2386 1238 2790 1286
rect 1886 1188 2288 1238
rect 1366 1158 1788 1188
rect 874 1100 1268 1158
rect 364 1060 776 1100
tri 776 1060 816 1100 sw
tri 874 1060 914 1100 ne
rect 914 1060 1268 1100
tri 1268 1060 1366 1158 sw
tri 1366 1060 1464 1158 ne
rect 1464 1100 1788 1158
tri 1788 1100 1876 1188 sw
tri 1886 1100 1974 1188 ne
rect 1974 1158 2288 1188
tri 2288 1158 2368 1238 sw
tri 2386 1158 2466 1238 ne
rect 2466 1188 2790 1238
tri 2790 1188 2888 1286 sw
tri 2888 1188 2986 1286 ne
rect 2986 1238 3300 1286
tri 3300 1238 3388 1326 sw
tri 3398 1238 3486 1326 ne
rect 3486 1290 3540 1326
rect 3660 1326 3762 1410
tri 3762 1326 3850 1414 sw
tri 3860 1326 3948 1414 ne
rect 3948 1410 4312 1414
rect 3948 1326 4090 1410
rect 3660 1290 3850 1326
rect 3486 1286 3850 1290
tri 3850 1286 3890 1326 sw
tri 3948 1286 3988 1326 ne
rect 3988 1290 4090 1326
rect 4210 1326 4312 1410
tri 4312 1326 4400 1414 sw
tri 4410 1326 4498 1414 ne
rect 4498 1410 4862 1414
rect 4498 1326 4640 1410
rect 4210 1290 4400 1326
rect 3988 1286 4400 1290
rect 3486 1238 3890 1286
rect 2986 1188 3388 1238
rect 2466 1158 2888 1188
rect 1974 1100 2368 1158
rect 1464 1060 1876 1100
tri 1876 1060 1916 1100 sw
tri 1974 1060 2014 1100 ne
rect 2014 1060 2368 1100
tri 2368 1060 2466 1158 sw
tri 2466 1060 2564 1158 ne
rect 2564 1100 2888 1158
tri 2888 1100 2976 1188 sw
tri 2986 1100 3074 1188 ne
rect 3074 1158 3388 1188
tri 3388 1158 3468 1238 sw
tri 3486 1158 3566 1238 ne
rect 3566 1188 3890 1238
tri 3890 1188 3988 1286 sw
tri 3988 1188 4086 1286 ne
rect 4086 1238 4400 1286
tri 4400 1238 4488 1326 sw
tri 4498 1238 4586 1326 ne
rect 4586 1290 4640 1326
rect 4760 1326 4862 1410
tri 4862 1326 4950 1414 sw
tri 4960 1326 5048 1414 ne
rect 5048 1410 5412 1414
rect 5048 1326 5190 1410
rect 4760 1290 4950 1326
rect 4586 1286 4950 1290
tri 4950 1286 4990 1326 sw
tri 5048 1286 5088 1326 ne
rect 5088 1290 5190 1326
rect 5310 1326 5412 1410
tri 5412 1326 5500 1414 sw
tri 5510 1326 5598 1414 ne
rect 5598 1410 5962 1414
rect 5598 1326 5740 1410
rect 5310 1290 5500 1326
rect 5088 1286 5500 1290
rect 4586 1238 4990 1286
rect 4086 1188 4488 1238
rect 3566 1158 3988 1188
rect 3074 1100 3468 1158
rect 2564 1060 2976 1100
tri 2976 1060 3016 1100 sw
tri 3074 1060 3114 1100 ne
rect 3114 1060 3468 1100
tri 3468 1060 3566 1158 sw
tri 3566 1060 3664 1158 ne
rect 3664 1100 3988 1158
tri 3988 1100 4076 1188 sw
tri 4086 1100 4174 1188 ne
rect 4174 1158 4488 1188
tri 4488 1158 4568 1238 sw
tri 4586 1158 4666 1238 ne
rect 4666 1188 4990 1238
tri 4990 1188 5088 1286 sw
tri 5088 1188 5186 1286 ne
rect 5186 1238 5500 1286
tri 5500 1238 5588 1326 sw
tri 5598 1238 5686 1326 ne
rect 5686 1290 5740 1326
rect 5860 1326 5962 1410
tri 5962 1326 6050 1414 sw
tri 6060 1326 6148 1414 ne
rect 6148 1410 6512 1414
rect 6148 1326 6290 1410
rect 5860 1290 6050 1326
rect 5686 1286 6050 1290
tri 6050 1286 6090 1326 sw
tri 6148 1286 6188 1326 ne
rect 6188 1290 6290 1326
rect 6410 1326 6512 1410
tri 6512 1326 6600 1414 sw
tri 6610 1326 6698 1414 ne
rect 6698 1410 7062 1414
rect 6698 1326 6840 1410
rect 6410 1290 6600 1326
rect 6188 1286 6600 1290
rect 5686 1238 6090 1286
rect 5186 1188 5588 1238
rect 4666 1158 5088 1188
rect 4174 1100 4568 1158
rect 3664 1060 4076 1100
tri 4076 1060 4116 1100 sw
tri 4174 1060 4214 1100 ne
rect 4214 1060 4568 1100
tri 4568 1060 4666 1158 sw
tri 4666 1060 4764 1158 ne
rect 4764 1100 5088 1158
tri 5088 1100 5176 1188 sw
tri 5186 1100 5274 1188 ne
rect 5274 1158 5588 1188
tri 5588 1158 5668 1238 sw
tri 5686 1158 5766 1238 ne
rect 5766 1188 6090 1238
tri 6090 1188 6188 1286 sw
tri 6188 1188 6286 1286 ne
rect 6286 1238 6600 1286
tri 6600 1238 6688 1326 sw
tri 6698 1238 6786 1326 ne
rect 6786 1290 6840 1326
rect 6960 1326 7062 1410
tri 7062 1326 7150 1414 sw
tri 7160 1326 7248 1414 ne
rect 7248 1410 7612 1414
rect 7248 1326 7390 1410
rect 6960 1290 7150 1326
rect 6786 1286 7150 1290
tri 7150 1286 7190 1326 sw
tri 7248 1286 7288 1326 ne
rect 7288 1290 7390 1326
rect 7510 1326 7612 1410
tri 7612 1326 7700 1414 sw
tri 7710 1326 7798 1414 ne
rect 7798 1410 8162 1414
rect 7798 1326 7940 1410
rect 7510 1290 7700 1326
rect 7288 1286 7700 1290
rect 6786 1238 7190 1286
rect 6286 1188 6688 1238
rect 5766 1158 6188 1188
rect 5274 1100 5668 1158
rect 4764 1060 5176 1100
tri 5176 1060 5216 1100 sw
tri 5274 1060 5314 1100 ne
rect 5314 1060 5668 1100
tri 5668 1060 5766 1158 sw
tri 5766 1060 5864 1158 ne
rect 5864 1100 6188 1158
tri 6188 1100 6276 1188 sw
tri 6286 1100 6374 1188 ne
rect 6374 1158 6688 1188
tri 6688 1158 6768 1238 sw
tri 6786 1158 6866 1238 ne
rect 6866 1188 7190 1238
tri 7190 1188 7288 1286 sw
tri 7288 1188 7386 1286 ne
rect 7386 1238 7700 1286
tri 7700 1238 7788 1326 sw
tri 7798 1238 7886 1326 ne
rect 7886 1290 7940 1326
rect 8060 1326 8162 1410
tri 8162 1326 8250 1414 sw
tri 8260 1326 8348 1414 ne
rect 8348 1410 8712 1414
rect 8348 1326 8490 1410
rect 8060 1290 8250 1326
rect 7886 1286 8250 1290
tri 8250 1286 8290 1326 sw
tri 8348 1286 8388 1326 ne
rect 8388 1290 8490 1326
rect 8610 1326 8712 1410
tri 8712 1326 8800 1414 sw
tri 8810 1326 8898 1414 ne
rect 8898 1410 9262 1414
rect 8898 1326 9040 1410
rect 8610 1290 8800 1326
rect 8388 1286 8800 1290
rect 7886 1238 8290 1286
rect 7386 1188 7788 1238
rect 6866 1158 7288 1188
rect 6374 1100 6768 1158
rect 5864 1060 6276 1100
tri 6276 1060 6316 1100 sw
tri 6374 1060 6414 1100 ne
rect 6414 1060 6768 1100
tri 6768 1060 6866 1158 sw
tri 6866 1060 6964 1158 ne
rect 6964 1100 7288 1158
tri 7288 1100 7376 1188 sw
tri 7386 1100 7474 1188 ne
rect 7474 1158 7788 1188
tri 7788 1158 7868 1238 sw
tri 7886 1158 7966 1238 ne
rect 7966 1188 8290 1238
tri 8290 1188 8388 1286 sw
tri 8388 1188 8486 1286 ne
rect 8486 1238 8800 1286
tri 8800 1238 8888 1326 sw
tri 8898 1238 8986 1326 ne
rect 8986 1290 9040 1326
rect 9160 1326 9262 1410
tri 9262 1326 9350 1414 sw
tri 9360 1326 9448 1414 ne
rect 9448 1410 9812 1414
rect 9448 1326 9590 1410
rect 9160 1290 9350 1326
rect 8986 1286 9350 1290
tri 9350 1286 9390 1326 sw
tri 9448 1286 9488 1326 ne
rect 9488 1290 9590 1326
rect 9710 1326 9812 1410
tri 9812 1326 9900 1414 sw
tri 9910 1326 9998 1414 ne
rect 9998 1410 10362 1414
rect 9998 1326 10140 1410
rect 9710 1290 9900 1326
rect 9488 1286 9900 1290
rect 8986 1238 9390 1286
rect 8486 1188 8888 1238
rect 7966 1158 8388 1188
rect 7474 1100 7868 1158
rect 6964 1060 7376 1100
tri 7376 1060 7416 1100 sw
tri 7474 1060 7514 1100 ne
rect 7514 1060 7868 1100
tri 7868 1060 7966 1158 sw
tri 7966 1060 8064 1158 ne
rect 8064 1100 8388 1158
tri 8388 1100 8476 1188 sw
tri 8486 1100 8574 1188 ne
rect 8574 1158 8888 1188
tri 8888 1158 8968 1238 sw
tri 8986 1158 9066 1238 ne
rect 9066 1188 9390 1238
tri 9390 1188 9488 1286 sw
tri 9488 1188 9586 1286 ne
rect 9586 1238 9900 1286
tri 9900 1238 9988 1326 sw
tri 9998 1238 10086 1326 ne
rect 10086 1290 10140 1326
rect 10260 1326 10362 1410
tri 10362 1326 10450 1414 sw
tri 10460 1326 10548 1414 ne
rect 10548 1410 10912 1414
rect 10548 1326 10690 1410
rect 10260 1290 10450 1326
rect 10086 1286 10450 1290
tri 10450 1286 10490 1326 sw
tri 10548 1286 10588 1326 ne
rect 10588 1290 10690 1326
rect 10810 1326 10912 1410
tri 10912 1326 11000 1414 sw
tri 11010 1326 11098 1414 ne
rect 11098 1410 11462 1414
rect 11098 1326 11240 1410
rect 10810 1290 11000 1326
rect 10588 1286 11000 1290
rect 10086 1238 10490 1286
rect 9586 1188 9988 1238
rect 9066 1158 9488 1188
rect 8574 1100 8968 1158
rect 8064 1060 8476 1100
tri 8476 1060 8516 1100 sw
tri 8574 1060 8614 1100 ne
rect 8614 1060 8968 1100
tri 8968 1060 9066 1158 sw
tri 9066 1060 9164 1158 ne
rect 9164 1100 9488 1158
tri 9488 1100 9576 1188 sw
tri 9586 1100 9674 1188 ne
rect 9674 1158 9988 1188
tri 9988 1158 10068 1238 sw
tri 10086 1158 10166 1238 ne
rect 10166 1188 10490 1238
tri 10490 1188 10588 1286 sw
tri 10588 1188 10686 1286 ne
rect 10686 1238 11000 1286
tri 11000 1238 11088 1326 sw
tri 11098 1238 11186 1326 ne
rect 11186 1290 11240 1326
rect 11360 1326 11462 1410
tri 11462 1326 11550 1414 sw
tri 11560 1326 11648 1414 ne
rect 11648 1410 12012 1414
rect 11648 1326 11790 1410
rect 11360 1290 11550 1326
rect 11186 1286 11550 1290
tri 11550 1286 11590 1326 sw
tri 11648 1286 11688 1326 ne
rect 11688 1290 11790 1326
rect 11910 1326 12012 1410
tri 12012 1326 12100 1414 sw
tri 12110 1326 12198 1414 ne
rect 12198 1410 12562 1414
rect 12198 1326 12340 1410
rect 11910 1290 12100 1326
rect 11688 1286 12100 1290
rect 11186 1238 11590 1286
rect 10686 1188 11088 1238
rect 10166 1158 10588 1188
rect 9674 1100 10068 1158
rect 9164 1060 9576 1100
tri 9576 1060 9616 1100 sw
tri 9674 1060 9714 1100 ne
rect 9714 1060 10068 1100
tri 10068 1060 10166 1158 sw
tri 10166 1060 10264 1158 ne
rect 10264 1100 10588 1158
tri 10588 1100 10676 1188 sw
tri 10686 1100 10774 1188 ne
rect 10774 1158 11088 1188
tri 11088 1158 11168 1238 sw
tri 11186 1158 11266 1238 ne
rect 11266 1188 11590 1238
tri 11590 1188 11688 1286 sw
tri 11688 1188 11786 1286 ne
rect 11786 1238 12100 1286
tri 12100 1238 12188 1326 sw
tri 12198 1238 12286 1326 ne
rect 12286 1290 12340 1326
rect 12460 1326 12562 1410
tri 12562 1326 12650 1414 sw
tri 12660 1326 12748 1414 ne
rect 12748 1410 13112 1414
rect 12748 1326 12890 1410
rect 12460 1290 12650 1326
rect 12286 1286 12650 1290
tri 12650 1286 12690 1326 sw
tri 12748 1286 12788 1326 ne
rect 12788 1290 12890 1326
rect 13010 1326 13112 1410
tri 13112 1326 13200 1414 sw
tri 13210 1326 13298 1414 ne
rect 13298 1410 15775 1414
rect 13298 1326 13440 1410
rect 13010 1290 13200 1326
rect 12788 1286 13200 1290
rect 12286 1238 12690 1286
rect 11786 1188 12188 1238
rect 11266 1158 11688 1188
rect 10774 1100 11168 1158
rect 10264 1060 10676 1100
tri 10676 1060 10716 1100 sw
tri 10774 1060 10814 1100 ne
rect 10814 1060 11168 1100
tri 11168 1060 11266 1158 sw
tri 11266 1060 11364 1158 ne
rect 11364 1100 11688 1158
tri 11688 1100 11776 1188 sw
tri 11786 1100 11874 1188 ne
rect 11874 1158 12188 1188
tri 12188 1158 12268 1238 sw
tri 12286 1158 12366 1238 ne
rect 12366 1188 12690 1238
tri 12690 1188 12788 1286 sw
tri 12788 1188 12886 1286 ne
rect 12886 1238 13200 1286
tri 13200 1238 13288 1326 sw
tri 13298 1238 13386 1326 ne
rect 13386 1290 13440 1326
rect 13560 1290 15775 1410
rect 13386 1238 15775 1290
rect 12886 1188 13288 1238
rect 12366 1158 12788 1188
rect 11874 1100 12268 1158
rect 11364 1060 11776 1100
tri 11776 1060 11816 1100 sw
tri 11874 1060 11914 1100 ne
rect 11914 1060 12268 1100
tri 12268 1060 12366 1158 sw
tri 12366 1060 12464 1158 ne
rect 12464 1100 12788 1158
tri 12788 1100 12876 1188 sw
tri 12886 1100 12974 1188 ne
rect 12974 1158 13288 1188
tri 13288 1158 13368 1238 sw
tri 13386 1158 13466 1238 ne
rect 13466 1158 14075 1238
rect 12974 1100 13368 1158
rect 12464 1060 12876 1100
tri 12876 1060 12916 1100 sw
tri 12974 1060 13014 1100 ne
rect 13014 1060 13368 1100
tri 13368 1060 13466 1158 sw
tri 13466 1060 13564 1158 ne
rect 13564 1138 14075 1158
rect 14175 1138 15775 1238
rect 13564 1060 15775 1138
rect -1025 1012 -284 1060
rect -1025 912 -925 1012
rect -825 962 -284 1012
tri -284 962 -186 1060 sw
tri -186 962 -88 1060 ne
rect -88 962 266 1060
tri 266 962 364 1060 sw
tri 364 962 462 1060 ne
rect 462 962 816 1060
tri 816 962 914 1060 sw
tri 914 962 1012 1060 ne
rect 1012 962 1366 1060
tri 1366 962 1464 1060 sw
tri 1464 962 1562 1060 ne
rect 1562 962 1916 1060
tri 1916 962 2014 1060 sw
tri 2014 962 2112 1060 ne
rect 2112 962 2466 1060
tri 2466 962 2564 1060 sw
tri 2564 962 2662 1060 ne
rect 2662 962 3016 1060
tri 3016 962 3114 1060 sw
tri 3114 962 3212 1060 ne
rect 3212 962 3566 1060
tri 3566 962 3664 1060 sw
tri 3664 962 3762 1060 ne
rect 3762 962 4116 1060
tri 4116 962 4214 1060 sw
tri 4214 962 4312 1060 ne
rect 4312 962 4666 1060
tri 4666 962 4764 1060 sw
tri 4764 962 4862 1060 ne
rect 4862 962 5216 1060
tri 5216 962 5314 1060 sw
tri 5314 962 5412 1060 ne
rect 5412 962 5766 1060
tri 5766 962 5864 1060 sw
tri 5864 962 5962 1060 ne
rect 5962 962 6316 1060
tri 6316 962 6414 1060 sw
tri 6414 962 6512 1060 ne
rect 6512 962 6866 1060
tri 6866 962 6964 1060 sw
tri 6964 962 7062 1060 ne
rect 7062 962 7416 1060
tri 7416 962 7514 1060 sw
tri 7514 962 7612 1060 ne
rect 7612 962 7966 1060
tri 7966 962 8064 1060 sw
tri 8064 962 8162 1060 ne
rect 8162 962 8516 1060
tri 8516 962 8614 1060 sw
tri 8614 962 8712 1060 ne
rect 8712 962 9066 1060
tri 9066 962 9164 1060 sw
tri 9164 962 9262 1060 ne
rect 9262 962 9616 1060
tri 9616 962 9714 1060 sw
tri 9714 962 9812 1060 ne
rect 9812 962 10166 1060
tri 10166 962 10264 1060 sw
tri 10264 962 10362 1060 ne
rect 10362 962 10716 1060
tri 10716 962 10814 1060 sw
tri 10814 962 10912 1060 ne
rect 10912 962 11266 1060
tri 11266 962 11364 1060 sw
tri 11364 962 11462 1060 ne
rect 11462 962 11816 1060
tri 11816 962 11914 1060 sw
tri 11914 962 12012 1060 ne
rect 12012 962 12366 1060
tri 12366 962 12464 1060 sw
tri 12464 962 12562 1060 ne
rect 12562 962 12916 1060
tri 12916 962 13014 1060 sw
tri 13014 962 13112 1060 ne
rect 13112 962 13466 1060
tri 13466 962 13564 1060 sw
tri 13564 962 13662 1060 ne
rect 13662 962 15775 1060
rect -825 912 -186 962
rect -1025 864 -186 912
tri -186 864 -88 962 sw
tri -88 864 10 962 ne
rect 10 864 364 962
tri 364 864 462 962 sw
tri 462 864 560 962 ne
rect 560 864 914 962
tri 914 864 1012 962 sw
tri 1012 864 1110 962 ne
rect 1110 864 1464 962
tri 1464 864 1562 962 sw
tri 1562 864 1660 962 ne
rect 1660 864 2014 962
tri 2014 864 2112 962 sw
tri 2112 864 2210 962 ne
rect 2210 864 2564 962
tri 2564 864 2662 962 sw
tri 2662 864 2760 962 ne
rect 2760 864 3114 962
tri 3114 864 3212 962 sw
tri 3212 864 3310 962 ne
rect 3310 864 3664 962
tri 3664 864 3762 962 sw
tri 3762 864 3860 962 ne
rect 3860 864 4214 962
tri 4214 864 4312 962 sw
tri 4312 864 4410 962 ne
rect 4410 864 4764 962
tri 4764 864 4862 962 sw
tri 4862 864 4960 962 ne
rect 4960 864 5314 962
tri 5314 864 5412 962 sw
tri 5412 864 5510 962 ne
rect 5510 864 5864 962
tri 5864 864 5962 962 sw
tri 5962 864 6060 962 ne
rect 6060 864 6414 962
tri 6414 864 6512 962 sw
tri 6512 864 6610 962 ne
rect 6610 864 6964 962
tri 6964 864 7062 962 sw
tri 7062 864 7160 962 ne
rect 7160 864 7514 962
tri 7514 864 7612 962 sw
tri 7612 864 7710 962 ne
rect 7710 864 8064 962
tri 8064 864 8162 962 sw
tri 8162 864 8260 962 ne
rect 8260 864 8614 962
tri 8614 864 8712 962 sw
tri 8712 864 8810 962 ne
rect 8810 864 9164 962
tri 9164 864 9262 962 sw
tri 9262 864 9360 962 ne
rect 9360 864 9714 962
tri 9714 864 9812 962 sw
tri 9812 864 9910 962 ne
rect 9910 864 10264 962
tri 10264 864 10362 962 sw
tri 10362 864 10460 962 ne
rect 10460 864 10814 962
tri 10814 864 10912 962 sw
tri 10912 864 11010 962 ne
rect 11010 864 11364 962
tri 11364 864 11462 962 sw
tri 11462 864 11560 962 ne
rect 11560 864 11914 962
tri 11914 864 12012 962 sw
tri 12012 864 12110 962 ne
rect 12110 864 12464 962
tri 12464 864 12562 962 sw
tri 12562 864 12660 962 ne
rect 12660 864 13014 962
tri 13014 864 13112 962 sw
tri 13112 864 13210 962 ne
rect 13210 864 13564 962
tri 13564 864 13662 962 sw
rect -1025 860 -88 864
rect -1025 740 -310 860
rect -190 776 -88 860
tri -88 776 0 864 sw
tri 10 776 98 864 ne
rect 98 860 462 864
rect 98 776 240 860
rect -190 740 0 776
rect -1025 736 0 740
tri 0 736 40 776 sw
tri 98 736 138 776 ne
rect 138 740 240 776
rect 360 776 462 860
tri 462 776 550 864 sw
tri 560 776 648 864 ne
rect 648 860 1012 864
rect 648 776 790 860
rect 360 740 550 776
rect 138 736 550 740
tri -412 638 -314 736 ne
rect -314 638 40 736
tri 40 638 138 736 sw
tri 138 638 236 736 ne
rect 236 688 550 736
tri 550 688 638 776 sw
tri 648 688 736 776 ne
rect 736 740 790 776
rect 910 776 1012 860
tri 1012 776 1100 864 sw
tri 1110 776 1198 864 ne
rect 1198 860 1562 864
rect 1198 776 1340 860
rect 910 740 1100 776
rect 736 736 1100 740
tri 1100 736 1140 776 sw
tri 1198 736 1238 776 ne
rect 1238 740 1340 776
rect 1460 776 1562 860
tri 1562 776 1650 864 sw
tri 1660 776 1748 864 ne
rect 1748 860 2112 864
rect 1748 776 1890 860
rect 1460 740 1650 776
rect 1238 736 1650 740
rect 736 688 1140 736
rect 236 638 638 688
rect -2525 550 -412 638
tri -412 550 -324 638 sw
tri -314 550 -226 638 ne
rect -226 550 138 638
tri 138 550 226 638 sw
tri 236 550 324 638 ne
rect 324 608 638 638
tri 638 608 718 688 sw
tri 736 608 816 688 ne
rect 816 638 1140 688
tri 1140 638 1238 736 sw
tri 1238 638 1336 736 ne
rect 1336 688 1650 736
tri 1650 688 1738 776 sw
tri 1748 688 1836 776 ne
rect 1836 740 1890 776
rect 2010 776 2112 860
tri 2112 776 2200 864 sw
tri 2210 776 2298 864 ne
rect 2298 860 2662 864
rect 2298 776 2440 860
rect 2010 740 2200 776
rect 1836 736 2200 740
tri 2200 736 2240 776 sw
tri 2298 736 2338 776 ne
rect 2338 740 2440 776
rect 2560 776 2662 860
tri 2662 776 2750 864 sw
tri 2760 776 2848 864 ne
rect 2848 860 3212 864
rect 2848 776 2990 860
rect 2560 740 2750 776
rect 2338 736 2750 740
rect 1836 688 2240 736
rect 1336 638 1738 688
rect 816 608 1238 638
rect 324 550 718 608
rect -2525 510 -324 550
tri -324 510 -284 550 sw
tri -226 510 -186 550 ne
rect -186 510 226 550
tri 226 510 266 550 sw
tri 324 510 364 550 ne
rect 364 510 718 550
tri 718 510 816 608 sw
tri 816 510 914 608 ne
rect 914 550 1238 608
tri 1238 550 1326 638 sw
tri 1336 550 1424 638 ne
rect 1424 608 1738 638
tri 1738 608 1818 688 sw
tri 1836 608 1916 688 ne
rect 1916 638 2240 688
tri 2240 638 2338 736 sw
tri 2338 638 2436 736 ne
rect 2436 688 2750 736
tri 2750 688 2838 776 sw
tri 2848 688 2936 776 ne
rect 2936 740 2990 776
rect 3110 776 3212 860
tri 3212 776 3300 864 sw
tri 3310 776 3398 864 ne
rect 3398 860 3762 864
rect 3398 776 3540 860
rect 3110 740 3300 776
rect 2936 736 3300 740
tri 3300 736 3340 776 sw
tri 3398 736 3438 776 ne
rect 3438 740 3540 776
rect 3660 776 3762 860
tri 3762 776 3850 864 sw
tri 3860 776 3948 864 ne
rect 3948 860 4312 864
rect 3948 776 4090 860
rect 3660 740 3850 776
rect 3438 736 3850 740
rect 2936 688 3340 736
rect 2436 638 2838 688
rect 1916 608 2338 638
rect 1424 550 1818 608
rect 914 510 1326 550
tri 1326 510 1366 550 sw
tri 1424 510 1464 550 ne
rect 1464 510 1818 550
tri 1818 510 1916 608 sw
tri 1916 510 2014 608 ne
rect 2014 550 2338 608
tri 2338 550 2426 638 sw
tri 2436 550 2524 638 ne
rect 2524 608 2838 638
tri 2838 608 2918 688 sw
tri 2936 608 3016 688 ne
rect 3016 638 3340 688
tri 3340 638 3438 736 sw
tri 3438 638 3536 736 ne
rect 3536 688 3850 736
tri 3850 688 3938 776 sw
tri 3948 688 4036 776 ne
rect 4036 740 4090 776
rect 4210 776 4312 860
tri 4312 776 4400 864 sw
tri 4410 776 4498 864 ne
rect 4498 860 4862 864
rect 4498 776 4640 860
rect 4210 740 4400 776
rect 4036 736 4400 740
tri 4400 736 4440 776 sw
tri 4498 736 4538 776 ne
rect 4538 740 4640 776
rect 4760 776 4862 860
tri 4862 776 4950 864 sw
tri 4960 776 5048 864 ne
rect 5048 860 5412 864
rect 5048 776 5190 860
rect 4760 740 4950 776
rect 4538 736 4950 740
rect 4036 688 4440 736
rect 3536 638 3938 688
rect 3016 608 3438 638
rect 2524 550 2918 608
rect 2014 510 2426 550
tri 2426 510 2466 550 sw
tri 2524 510 2564 550 ne
rect 2564 510 2918 550
tri 2918 510 3016 608 sw
tri 3016 510 3114 608 ne
rect 3114 550 3438 608
tri 3438 550 3526 638 sw
tri 3536 550 3624 638 ne
rect 3624 608 3938 638
tri 3938 608 4018 688 sw
tri 4036 608 4116 688 ne
rect 4116 638 4440 688
tri 4440 638 4538 736 sw
tri 4538 638 4636 736 ne
rect 4636 688 4950 736
tri 4950 688 5038 776 sw
tri 5048 688 5136 776 ne
rect 5136 740 5190 776
rect 5310 776 5412 860
tri 5412 776 5500 864 sw
tri 5510 776 5598 864 ne
rect 5598 860 5962 864
rect 5598 776 5740 860
rect 5310 740 5500 776
rect 5136 736 5500 740
tri 5500 736 5540 776 sw
tri 5598 736 5638 776 ne
rect 5638 740 5740 776
rect 5860 776 5962 860
tri 5962 776 6050 864 sw
tri 6060 776 6148 864 ne
rect 6148 860 6512 864
rect 6148 776 6290 860
rect 5860 740 6050 776
rect 5638 736 6050 740
rect 5136 688 5540 736
rect 4636 638 5038 688
rect 4116 608 4538 638
rect 3624 550 4018 608
rect 3114 510 3526 550
tri 3526 510 3566 550 sw
tri 3624 510 3664 550 ne
rect 3664 510 4018 550
tri 4018 510 4116 608 sw
tri 4116 510 4214 608 ne
rect 4214 550 4538 608
tri 4538 550 4626 638 sw
tri 4636 550 4724 638 ne
rect 4724 608 5038 638
tri 5038 608 5118 688 sw
tri 5136 608 5216 688 ne
rect 5216 638 5540 688
tri 5540 638 5638 736 sw
tri 5638 638 5736 736 ne
rect 5736 688 6050 736
tri 6050 688 6138 776 sw
tri 6148 688 6236 776 ne
rect 6236 740 6290 776
rect 6410 776 6512 860
tri 6512 776 6600 864 sw
tri 6610 776 6698 864 ne
rect 6698 860 7062 864
rect 6698 776 6840 860
rect 6410 740 6600 776
rect 6236 736 6600 740
tri 6600 736 6640 776 sw
tri 6698 736 6738 776 ne
rect 6738 740 6840 776
rect 6960 776 7062 860
tri 7062 776 7150 864 sw
tri 7160 776 7248 864 ne
rect 7248 860 7612 864
rect 7248 776 7390 860
rect 6960 740 7150 776
rect 6738 736 7150 740
rect 6236 688 6640 736
rect 5736 638 6138 688
rect 5216 608 5638 638
rect 4724 550 5118 608
rect 4214 510 4626 550
tri 4626 510 4666 550 sw
tri 4724 510 4764 550 ne
rect 4764 510 5118 550
tri 5118 510 5216 608 sw
tri 5216 510 5314 608 ne
rect 5314 550 5638 608
tri 5638 550 5726 638 sw
tri 5736 550 5824 638 ne
rect 5824 608 6138 638
tri 6138 608 6218 688 sw
tri 6236 608 6316 688 ne
rect 6316 638 6640 688
tri 6640 638 6738 736 sw
tri 6738 638 6836 736 ne
rect 6836 688 7150 736
tri 7150 688 7238 776 sw
tri 7248 688 7336 776 ne
rect 7336 740 7390 776
rect 7510 776 7612 860
tri 7612 776 7700 864 sw
tri 7710 776 7798 864 ne
rect 7798 860 8162 864
rect 7798 776 7940 860
rect 7510 740 7700 776
rect 7336 736 7700 740
tri 7700 736 7740 776 sw
tri 7798 736 7838 776 ne
rect 7838 740 7940 776
rect 8060 776 8162 860
tri 8162 776 8250 864 sw
tri 8260 776 8348 864 ne
rect 8348 860 8712 864
rect 8348 776 8490 860
rect 8060 740 8250 776
rect 7838 736 8250 740
rect 7336 688 7740 736
rect 6836 638 7238 688
rect 6316 608 6738 638
rect 5824 550 6218 608
rect 5314 510 5726 550
tri 5726 510 5766 550 sw
tri 5824 510 5864 550 ne
rect 5864 510 6218 550
tri 6218 510 6316 608 sw
tri 6316 510 6414 608 ne
rect 6414 550 6738 608
tri 6738 550 6826 638 sw
tri 6836 550 6924 638 ne
rect 6924 608 7238 638
tri 7238 608 7318 688 sw
tri 7336 608 7416 688 ne
rect 7416 638 7740 688
tri 7740 638 7838 736 sw
tri 7838 638 7936 736 ne
rect 7936 688 8250 736
tri 8250 688 8338 776 sw
tri 8348 688 8436 776 ne
rect 8436 740 8490 776
rect 8610 776 8712 860
tri 8712 776 8800 864 sw
tri 8810 776 8898 864 ne
rect 8898 860 9262 864
rect 8898 776 9040 860
rect 8610 740 8800 776
rect 8436 736 8800 740
tri 8800 736 8840 776 sw
tri 8898 736 8938 776 ne
rect 8938 740 9040 776
rect 9160 776 9262 860
tri 9262 776 9350 864 sw
tri 9360 776 9448 864 ne
rect 9448 860 9812 864
rect 9448 776 9590 860
rect 9160 740 9350 776
rect 8938 736 9350 740
rect 8436 688 8840 736
rect 7936 638 8338 688
rect 7416 608 7838 638
rect 6924 550 7318 608
rect 6414 510 6826 550
tri 6826 510 6866 550 sw
tri 6924 510 6964 550 ne
rect 6964 510 7318 550
tri 7318 510 7416 608 sw
tri 7416 510 7514 608 ne
rect 7514 550 7838 608
tri 7838 550 7926 638 sw
tri 7936 550 8024 638 ne
rect 8024 608 8338 638
tri 8338 608 8418 688 sw
tri 8436 608 8516 688 ne
rect 8516 638 8840 688
tri 8840 638 8938 736 sw
tri 8938 638 9036 736 ne
rect 9036 688 9350 736
tri 9350 688 9438 776 sw
tri 9448 688 9536 776 ne
rect 9536 740 9590 776
rect 9710 776 9812 860
tri 9812 776 9900 864 sw
tri 9910 776 9998 864 ne
rect 9998 860 10362 864
rect 9998 776 10140 860
rect 9710 740 9900 776
rect 9536 736 9900 740
tri 9900 736 9940 776 sw
tri 9998 736 10038 776 ne
rect 10038 740 10140 776
rect 10260 776 10362 860
tri 10362 776 10450 864 sw
tri 10460 776 10548 864 ne
rect 10548 860 10912 864
rect 10548 776 10690 860
rect 10260 740 10450 776
rect 10038 736 10450 740
rect 9536 688 9940 736
rect 9036 638 9438 688
rect 8516 608 8938 638
rect 8024 550 8418 608
rect 7514 510 7926 550
tri 7926 510 7966 550 sw
tri 8024 510 8064 550 ne
rect 8064 510 8418 550
tri 8418 510 8516 608 sw
tri 8516 510 8614 608 ne
rect 8614 550 8938 608
tri 8938 550 9026 638 sw
tri 9036 550 9124 638 ne
rect 9124 608 9438 638
tri 9438 608 9518 688 sw
tri 9536 608 9616 688 ne
rect 9616 638 9940 688
tri 9940 638 10038 736 sw
tri 10038 638 10136 736 ne
rect 10136 688 10450 736
tri 10450 688 10538 776 sw
tri 10548 688 10636 776 ne
rect 10636 740 10690 776
rect 10810 776 10912 860
tri 10912 776 11000 864 sw
tri 11010 776 11098 864 ne
rect 11098 860 11462 864
rect 11098 776 11240 860
rect 10810 740 11000 776
rect 10636 736 11000 740
tri 11000 736 11040 776 sw
tri 11098 736 11138 776 ne
rect 11138 740 11240 776
rect 11360 776 11462 860
tri 11462 776 11550 864 sw
tri 11560 776 11648 864 ne
rect 11648 860 12012 864
rect 11648 776 11790 860
rect 11360 740 11550 776
rect 11138 736 11550 740
rect 10636 688 11040 736
rect 10136 638 10538 688
rect 9616 608 10038 638
rect 9124 550 9518 608
rect 8614 510 9026 550
tri 9026 510 9066 550 sw
tri 9124 510 9164 550 ne
rect 9164 510 9518 550
tri 9518 510 9616 608 sw
tri 9616 510 9714 608 ne
rect 9714 550 10038 608
tri 10038 550 10126 638 sw
tri 10136 550 10224 638 ne
rect 10224 608 10538 638
tri 10538 608 10618 688 sw
tri 10636 608 10716 688 ne
rect 10716 638 11040 688
tri 11040 638 11138 736 sw
tri 11138 638 11236 736 ne
rect 11236 688 11550 736
tri 11550 688 11638 776 sw
tri 11648 688 11736 776 ne
rect 11736 740 11790 776
rect 11910 776 12012 860
tri 12012 776 12100 864 sw
tri 12110 776 12198 864 ne
rect 12198 860 12562 864
rect 12198 776 12340 860
rect 11910 740 12100 776
rect 11736 736 12100 740
tri 12100 736 12140 776 sw
tri 12198 736 12238 776 ne
rect 12238 740 12340 776
rect 12460 776 12562 860
tri 12562 776 12650 864 sw
tri 12660 776 12748 864 ne
rect 12748 860 13112 864
rect 12748 776 12890 860
rect 12460 740 12650 776
rect 12238 736 12650 740
rect 11736 688 12140 736
rect 11236 638 11638 688
rect 10716 608 11138 638
rect 10224 550 10618 608
rect 9714 510 10126 550
tri 10126 510 10166 550 sw
tri 10224 510 10264 550 ne
rect 10264 510 10618 550
tri 10618 510 10716 608 sw
tri 10716 510 10814 608 ne
rect 10814 550 11138 608
tri 11138 550 11226 638 sw
tri 11236 550 11324 638 ne
rect 11324 608 11638 638
tri 11638 608 11718 688 sw
tri 11736 608 11816 688 ne
rect 11816 638 12140 688
tri 12140 638 12238 736 sw
tri 12238 638 12336 736 ne
rect 12336 688 12650 736
tri 12650 688 12738 776 sw
tri 12748 688 12836 776 ne
rect 12836 740 12890 776
rect 13010 776 13112 860
tri 13112 776 13200 864 sw
tri 13210 776 13298 864 ne
rect 13298 860 14275 864
rect 13298 776 13440 860
rect 13010 740 13200 776
rect 12836 736 13200 740
tri 13200 736 13240 776 sw
tri 13298 736 13338 776 ne
rect 13338 740 13440 776
rect 13560 740 14275 860
rect 13338 736 14275 740
rect 12836 688 13240 736
rect 12336 638 12738 688
rect 11816 608 12238 638
rect 11324 550 11718 608
rect 10814 510 11226 550
tri 11226 510 11266 550 sw
tri 11324 510 11364 550 ne
rect 11364 510 11718 550
tri 11718 510 11816 608 sw
tri 11816 510 11914 608 ne
rect 11914 550 12238 608
tri 12238 550 12326 638 sw
tri 12336 550 12424 638 ne
rect 12424 608 12738 638
tri 12738 608 12818 688 sw
tri 12836 608 12916 688 ne
rect 12916 638 13240 688
tri 13240 638 13338 736 sw
tri 13338 638 13436 736 ne
rect 13436 638 14275 736
rect 12916 608 13338 638
rect 12424 550 12818 608
rect 11914 510 12326 550
tri 12326 510 12366 550 sw
tri 12424 510 12464 550 ne
rect 12464 510 12818 550
tri 12818 510 12916 608 sw
tri 12916 510 13014 608 ne
rect 13014 550 13338 608
tri 13338 550 13426 638 sw
tri 13436 550 13524 638 ne
rect 13524 550 14275 638
rect 13014 510 13426 550
tri 13426 510 13466 550 sw
tri 13524 510 13564 550 ne
rect 13564 510 14275 550
rect -2525 412 -284 510
tri -284 412 -186 510 sw
tri -186 412 -88 510 ne
rect -88 412 266 510
tri 266 412 364 510 sw
tri 364 412 462 510 ne
rect 462 412 816 510
tri 816 412 914 510 sw
tri 914 412 1012 510 ne
rect 1012 412 1366 510
tri 1366 412 1464 510 sw
tri 1464 412 1562 510 ne
rect 1562 412 1916 510
tri 1916 412 2014 510 sw
tri 2014 412 2112 510 ne
rect 2112 412 2466 510
tri 2466 412 2564 510 sw
tri 2564 412 2662 510 ne
rect 2662 412 3016 510
tri 3016 412 3114 510 sw
tri 3114 412 3212 510 ne
rect 3212 412 3566 510
tri 3566 412 3664 510 sw
tri 3664 412 3762 510 ne
rect 3762 412 4116 510
tri 4116 412 4214 510 sw
tri 4214 412 4312 510 ne
rect 4312 412 4666 510
tri 4666 412 4764 510 sw
tri 4764 412 4862 510 ne
rect 4862 412 5216 510
tri 5216 412 5314 510 sw
tri 5314 412 5412 510 ne
rect 5412 412 5766 510
tri 5766 412 5864 510 sw
tri 5864 412 5962 510 ne
rect 5962 412 6316 510
tri 6316 412 6414 510 sw
tri 6414 412 6512 510 ne
rect 6512 412 6866 510
tri 6866 412 6964 510 sw
tri 6964 412 7062 510 ne
rect 7062 412 7416 510
tri 7416 412 7514 510 sw
tri 7514 412 7612 510 ne
rect 7612 412 7966 510
tri 7966 412 8064 510 sw
tri 8064 412 8162 510 ne
rect 8162 412 8516 510
tri 8516 412 8614 510 sw
tri 8614 412 8712 510 ne
rect 8712 412 9066 510
tri 9066 412 9164 510 sw
tri 9164 412 9262 510 ne
rect 9262 412 9616 510
tri 9616 412 9714 510 sw
tri 9714 412 9812 510 ne
rect 9812 412 10166 510
tri 10166 412 10264 510 sw
tri 10264 412 10362 510 ne
rect 10362 412 10716 510
tri 10716 412 10814 510 sw
tri 10814 412 10912 510 ne
rect 10912 412 11266 510
tri 11266 412 11364 510 sw
tri 11364 412 11462 510 ne
rect 11462 412 11816 510
tri 11816 412 11914 510 sw
tri 11914 412 12012 510 ne
rect 12012 412 12366 510
tri 12366 412 12464 510 sw
tri 12464 412 12562 510 ne
rect 12562 412 12916 510
tri 12916 412 13014 510 sw
tri 13014 412 13112 510 ne
rect 13112 412 13466 510
tri 13466 412 13564 510 sw
tri 13564 412 13662 510 ne
rect 13662 412 14275 510
rect -2525 314 -186 412
tri -186 314 -88 412 sw
tri -88 314 10 412 ne
rect 10 314 364 412
tri 364 314 462 412 sw
tri 462 314 560 412 ne
rect 560 314 914 412
tri 914 314 1012 412 sw
tri 1012 314 1110 412 ne
rect 1110 314 1464 412
tri 1464 314 1562 412 sw
tri 1562 314 1660 412 ne
rect 1660 314 2014 412
tri 2014 314 2112 412 sw
tri 2112 314 2210 412 ne
rect 2210 314 2564 412
tri 2564 314 2662 412 sw
tri 2662 314 2760 412 ne
rect 2760 314 3114 412
tri 3114 314 3212 412 sw
tri 3212 314 3310 412 ne
rect 3310 314 3664 412
tri 3664 314 3762 412 sw
tri 3762 314 3860 412 ne
rect 3860 314 4214 412
tri 4214 314 4312 412 sw
tri 4312 314 4410 412 ne
rect 4410 314 4764 412
tri 4764 314 4862 412 sw
tri 4862 314 4960 412 ne
rect 4960 314 5314 412
tri 5314 314 5412 412 sw
tri 5412 314 5510 412 ne
rect 5510 314 5864 412
tri 5864 314 5962 412 sw
tri 5962 314 6060 412 ne
rect 6060 314 6414 412
tri 6414 314 6512 412 sw
tri 6512 314 6610 412 ne
rect 6610 314 6964 412
tri 6964 314 7062 412 sw
tri 7062 314 7160 412 ne
rect 7160 314 7514 412
tri 7514 314 7612 412 sw
tri 7612 314 7710 412 ne
rect 7710 314 8064 412
tri 8064 314 8162 412 sw
tri 8162 314 8260 412 ne
rect 8260 314 8614 412
tri 8614 314 8712 412 sw
tri 8712 314 8810 412 ne
rect 8810 314 9164 412
tri 9164 314 9262 412 sw
tri 9262 314 9360 412 ne
rect 9360 314 9714 412
tri 9714 314 9812 412 sw
tri 9812 314 9910 412 ne
rect 9910 314 10264 412
tri 10264 314 10362 412 sw
tri 10362 314 10460 412 ne
rect 10460 314 10814 412
tri 10814 314 10912 412 sw
tri 10912 314 11010 412 ne
rect 11010 314 11364 412
tri 11364 314 11462 412 sw
tri 11462 314 11560 412 ne
rect 11560 314 11914 412
tri 11914 314 12012 412 sw
tri 12012 314 12110 412 ne
rect 12110 314 12464 412
tri 12464 314 12562 412 sw
tri 12562 314 12660 412 ne
rect 12660 314 13014 412
tri 13014 314 13112 412 sw
tri 13112 314 13210 412 ne
rect 13210 314 13564 412
tri 13564 314 13662 412 sw
rect 14775 314 15775 962
rect -2525 310 -88 314
rect -2525 190 -310 310
rect -190 226 -88 310
tri -88 226 0 314 sw
tri 10 226 98 314 ne
rect 98 310 462 314
rect 98 226 240 310
rect -190 190 0 226
rect -2525 186 0 190
rect -2525 -575 -1525 186
tri -412 88 -314 186 ne
rect -314 138 0 186
tri 0 138 88 226 sw
tri 98 138 186 226 ne
rect 186 190 240 226
rect 360 226 462 310
tri 462 226 550 314 sw
tri 560 226 648 314 ne
rect 648 310 1012 314
rect 648 226 790 310
rect 360 190 550 226
rect 186 186 550 190
tri 550 186 590 226 sw
tri 648 186 688 226 ne
rect 688 190 790 226
rect 910 226 1012 310
tri 1012 226 1100 314 sw
tri 1110 226 1198 314 ne
rect 1198 310 1562 314
rect 1198 226 1340 310
rect 910 190 1100 226
rect 688 186 1100 190
rect 186 138 590 186
rect -314 88 88 138
rect -1025 0 -412 88
tri -412 0 -324 88 sw
tri -314 0 -226 88 ne
rect -226 58 88 88
tri 88 58 168 138 sw
tri 186 58 266 138 ne
rect 266 88 590 138
tri 590 88 688 186 sw
tri 688 88 786 186 ne
rect 786 138 1100 186
tri 1100 138 1188 226 sw
tri 1198 138 1286 226 ne
rect 1286 190 1340 226
rect 1460 226 1562 310
tri 1562 226 1650 314 sw
tri 1660 226 1748 314 ne
rect 1748 310 2112 314
rect 1748 226 1890 310
rect 1460 190 1650 226
rect 1286 186 1650 190
tri 1650 186 1690 226 sw
tri 1748 186 1788 226 ne
rect 1788 190 1890 226
rect 2010 226 2112 310
tri 2112 226 2200 314 sw
tri 2210 226 2298 314 ne
rect 2298 310 2662 314
rect 2298 226 2440 310
rect 2010 190 2200 226
rect 1788 186 2200 190
rect 1286 138 1690 186
rect 786 88 1188 138
rect 266 58 688 88
rect -226 0 168 58
tri 168 0 226 58 sw
tri 266 0 324 58 ne
rect 324 0 688 58
tri 688 0 776 88 sw
tri 786 0 874 88 ne
rect 874 58 1188 88
tri 1188 58 1268 138 sw
tri 1286 58 1366 138 ne
rect 1366 88 1690 138
tri 1690 88 1788 186 sw
tri 1788 88 1886 186 ne
rect 1886 138 2200 186
tri 2200 138 2288 226 sw
tri 2298 138 2386 226 ne
rect 2386 190 2440 226
rect 2560 226 2662 310
tri 2662 226 2750 314 sw
tri 2760 226 2848 314 ne
rect 2848 310 3212 314
rect 2848 226 2990 310
rect 2560 190 2750 226
rect 2386 186 2750 190
tri 2750 186 2790 226 sw
tri 2848 186 2888 226 ne
rect 2888 190 2990 226
rect 3110 226 3212 310
tri 3212 226 3300 314 sw
tri 3310 226 3398 314 ne
rect 3398 310 3762 314
rect 3398 226 3540 310
rect 3110 190 3300 226
rect 2888 186 3300 190
rect 2386 138 2790 186
rect 1886 88 2288 138
rect 1366 58 1788 88
rect 874 0 1268 58
tri 1268 0 1326 58 sw
tri 1366 0 1424 58 ne
rect 1424 0 1788 58
tri 1788 0 1876 88 sw
tri 1886 0 1974 88 ne
rect 1974 58 2288 88
tri 2288 58 2368 138 sw
tri 2386 58 2466 138 ne
rect 2466 88 2790 138
tri 2790 88 2888 186 sw
tri 2888 88 2986 186 ne
rect 2986 138 3300 186
tri 3300 138 3388 226 sw
tri 3398 138 3486 226 ne
rect 3486 190 3540 226
rect 3660 226 3762 310
tri 3762 226 3850 314 sw
tri 3860 226 3948 314 ne
rect 3948 310 4312 314
rect 3948 226 4090 310
rect 3660 190 3850 226
rect 3486 186 3850 190
tri 3850 186 3890 226 sw
tri 3948 186 3988 226 ne
rect 3988 190 4090 226
rect 4210 226 4312 310
tri 4312 226 4400 314 sw
tri 4410 226 4498 314 ne
rect 4498 310 4862 314
rect 4498 226 4640 310
rect 4210 190 4400 226
rect 3988 186 4400 190
rect 3486 138 3890 186
rect 2986 88 3388 138
rect 2466 58 2888 88
rect 1974 0 2368 58
tri 2368 0 2426 58 sw
tri 2466 0 2524 58 ne
rect 2524 0 2888 58
tri 2888 0 2976 88 sw
tri 2986 0 3074 88 ne
rect 3074 58 3388 88
tri 3388 58 3468 138 sw
tri 3486 58 3566 138 ne
rect 3566 88 3890 138
tri 3890 88 3988 186 sw
tri 3988 88 4086 186 ne
rect 4086 138 4400 186
tri 4400 138 4488 226 sw
tri 4498 138 4586 226 ne
rect 4586 190 4640 226
rect 4760 226 4862 310
tri 4862 226 4950 314 sw
tri 4960 226 5048 314 ne
rect 5048 310 5412 314
rect 5048 226 5190 310
rect 4760 190 4950 226
rect 4586 186 4950 190
tri 4950 186 4990 226 sw
tri 5048 186 5088 226 ne
rect 5088 190 5190 226
rect 5310 226 5412 310
tri 5412 226 5500 314 sw
tri 5510 226 5598 314 ne
rect 5598 310 5962 314
rect 5598 226 5740 310
rect 5310 190 5500 226
rect 5088 186 5500 190
rect 4586 138 4990 186
rect 4086 88 4488 138
rect 3566 58 3988 88
rect 3074 0 3468 58
tri 3468 0 3526 58 sw
tri 3566 0 3624 58 ne
rect 3624 0 3988 58
tri 3988 0 4076 88 sw
tri 4086 0 4174 88 ne
rect 4174 58 4488 88
tri 4488 58 4568 138 sw
tri 4586 58 4666 138 ne
rect 4666 88 4990 138
tri 4990 88 5088 186 sw
tri 5088 88 5186 186 ne
rect 5186 138 5500 186
tri 5500 138 5588 226 sw
tri 5598 138 5686 226 ne
rect 5686 190 5740 226
rect 5860 226 5962 310
tri 5962 226 6050 314 sw
tri 6060 226 6148 314 ne
rect 6148 310 6512 314
rect 6148 226 6290 310
rect 5860 190 6050 226
rect 5686 186 6050 190
tri 6050 186 6090 226 sw
tri 6148 186 6188 226 ne
rect 6188 190 6290 226
rect 6410 226 6512 310
tri 6512 226 6600 314 sw
tri 6610 226 6698 314 ne
rect 6698 310 7062 314
rect 6698 226 6840 310
rect 6410 190 6600 226
rect 6188 186 6600 190
rect 5686 138 6090 186
rect 5186 88 5588 138
rect 4666 58 5088 88
rect 4174 0 4568 58
tri 4568 0 4626 58 sw
tri 4666 0 4724 58 ne
rect 4724 0 5088 58
tri 5088 0 5176 88 sw
tri 5186 0 5274 88 ne
rect 5274 58 5588 88
tri 5588 58 5668 138 sw
tri 5686 58 5766 138 ne
rect 5766 88 6090 138
tri 6090 88 6188 186 sw
tri 6188 88 6286 186 ne
rect 6286 138 6600 186
tri 6600 138 6688 226 sw
tri 6698 138 6786 226 ne
rect 6786 190 6840 226
rect 6960 226 7062 310
tri 7062 226 7150 314 sw
tri 7160 226 7248 314 ne
rect 7248 310 7612 314
rect 7248 226 7390 310
rect 6960 190 7150 226
rect 6786 186 7150 190
tri 7150 186 7190 226 sw
tri 7248 186 7288 226 ne
rect 7288 190 7390 226
rect 7510 226 7612 310
tri 7612 226 7700 314 sw
tri 7710 226 7798 314 ne
rect 7798 310 8162 314
rect 7798 226 7940 310
rect 7510 190 7700 226
rect 7288 186 7700 190
rect 6786 138 7190 186
rect 6286 88 6688 138
rect 5766 58 6188 88
rect 5274 0 5668 58
tri 5668 0 5726 58 sw
tri 5766 0 5824 58 ne
rect 5824 0 6188 58
tri 6188 0 6276 88 sw
tri 6286 0 6374 88 ne
rect 6374 58 6688 88
tri 6688 58 6768 138 sw
tri 6786 58 6866 138 ne
rect 6866 88 7190 138
tri 7190 88 7288 186 sw
tri 7288 88 7386 186 ne
rect 7386 138 7700 186
tri 7700 138 7788 226 sw
tri 7798 138 7886 226 ne
rect 7886 190 7940 226
rect 8060 226 8162 310
tri 8162 226 8250 314 sw
tri 8260 226 8348 314 ne
rect 8348 310 8712 314
rect 8348 226 8490 310
rect 8060 190 8250 226
rect 7886 186 8250 190
tri 8250 186 8290 226 sw
tri 8348 186 8388 226 ne
rect 8388 190 8490 226
rect 8610 226 8712 310
tri 8712 226 8800 314 sw
tri 8810 226 8898 314 ne
rect 8898 310 9262 314
rect 8898 226 9040 310
rect 8610 190 8800 226
rect 8388 186 8800 190
rect 7886 138 8290 186
rect 7386 88 7788 138
rect 6866 58 7288 88
rect 6374 0 6768 58
tri 6768 0 6826 58 sw
tri 6866 0 6924 58 ne
rect 6924 0 7288 58
tri 7288 0 7376 88 sw
tri 7386 0 7474 88 ne
rect 7474 58 7788 88
tri 7788 58 7868 138 sw
tri 7886 58 7966 138 ne
rect 7966 88 8290 138
tri 8290 88 8388 186 sw
tri 8388 88 8486 186 ne
rect 8486 138 8800 186
tri 8800 138 8888 226 sw
tri 8898 138 8986 226 ne
rect 8986 190 9040 226
rect 9160 226 9262 310
tri 9262 226 9350 314 sw
tri 9360 226 9448 314 ne
rect 9448 310 9812 314
rect 9448 226 9590 310
rect 9160 190 9350 226
rect 8986 186 9350 190
tri 9350 186 9390 226 sw
tri 9448 186 9488 226 ne
rect 9488 190 9590 226
rect 9710 226 9812 310
tri 9812 226 9900 314 sw
tri 9910 226 9998 314 ne
rect 9998 310 10362 314
rect 9998 226 10140 310
rect 9710 190 9900 226
rect 9488 186 9900 190
rect 8986 138 9390 186
rect 8486 88 8888 138
rect 7966 58 8388 88
rect 7474 0 7868 58
tri 7868 0 7926 58 sw
tri 7966 0 8024 58 ne
rect 8024 0 8388 58
tri 8388 0 8476 88 sw
tri 8486 0 8574 88 ne
rect 8574 58 8888 88
tri 8888 58 8968 138 sw
tri 8986 58 9066 138 ne
rect 9066 88 9390 138
tri 9390 88 9488 186 sw
tri 9488 88 9586 186 ne
rect 9586 138 9900 186
tri 9900 138 9988 226 sw
tri 9998 138 10086 226 ne
rect 10086 190 10140 226
rect 10260 226 10362 310
tri 10362 226 10450 314 sw
tri 10460 226 10548 314 ne
rect 10548 310 10912 314
rect 10548 226 10690 310
rect 10260 190 10450 226
rect 10086 186 10450 190
tri 10450 186 10490 226 sw
tri 10548 186 10588 226 ne
rect 10588 190 10690 226
rect 10810 226 10912 310
tri 10912 226 11000 314 sw
tri 11010 226 11098 314 ne
rect 11098 310 11462 314
rect 11098 226 11240 310
rect 10810 190 11000 226
rect 10588 186 11000 190
rect 10086 138 10490 186
rect 9586 88 9988 138
rect 9066 58 9488 88
rect 8574 0 8968 58
tri 8968 0 9026 58 sw
tri 9066 0 9124 58 ne
rect 9124 0 9488 58
tri 9488 0 9576 88 sw
tri 9586 0 9674 88 ne
rect 9674 58 9988 88
tri 9988 58 10068 138 sw
tri 10086 58 10166 138 ne
rect 10166 88 10490 138
tri 10490 88 10588 186 sw
tri 10588 88 10686 186 ne
rect 10686 138 11000 186
tri 11000 138 11088 226 sw
tri 11098 138 11186 226 ne
rect 11186 190 11240 226
rect 11360 226 11462 310
tri 11462 226 11550 314 sw
tri 11560 226 11648 314 ne
rect 11648 310 12012 314
rect 11648 226 11790 310
rect 11360 190 11550 226
rect 11186 186 11550 190
tri 11550 186 11590 226 sw
tri 11648 186 11688 226 ne
rect 11688 190 11790 226
rect 11910 226 12012 310
tri 12012 226 12100 314 sw
tri 12110 226 12198 314 ne
rect 12198 310 12562 314
rect 12198 226 12340 310
rect 11910 190 12100 226
rect 11688 186 12100 190
rect 11186 138 11590 186
rect 10686 88 11088 138
rect 10166 58 10588 88
rect 9674 0 10068 58
tri 10068 0 10126 58 sw
tri 10166 0 10224 58 ne
rect 10224 0 10588 58
tri 10588 0 10676 88 sw
tri 10686 0 10774 88 ne
rect 10774 58 11088 88
tri 11088 58 11168 138 sw
tri 11186 58 11266 138 ne
rect 11266 88 11590 138
tri 11590 88 11688 186 sw
tri 11688 88 11786 186 ne
rect 11786 138 12100 186
tri 12100 138 12188 226 sw
tri 12198 138 12286 226 ne
rect 12286 190 12340 226
rect 12460 226 12562 310
tri 12562 226 12650 314 sw
tri 12660 226 12748 314 ne
rect 12748 310 13112 314
rect 12748 226 12890 310
rect 12460 190 12650 226
rect 12286 186 12650 190
tri 12650 186 12690 226 sw
tri 12748 186 12788 226 ne
rect 12788 190 12890 226
rect 13010 226 13112 310
tri 13112 226 13200 314 sw
tri 13210 226 13298 314 ne
rect 13298 310 15775 314
rect 13298 226 13440 310
rect 13010 190 13200 226
rect 12788 186 13200 190
rect 12286 138 12690 186
rect 11786 88 12188 138
rect 11266 58 11688 88
rect 10774 0 11168 58
tri 11168 0 11226 58 sw
tri 11266 0 11324 58 ne
rect 11324 0 11688 58
tri 11688 0 11776 88 sw
tri 11786 0 11874 88 ne
rect 11874 58 12188 88
tri 12188 58 12268 138 sw
tri 12286 58 12366 138 ne
rect 12366 88 12690 138
tri 12690 88 12788 186 sw
tri 12788 88 12886 186 ne
rect 12886 138 13200 186
tri 13200 138 13288 226 sw
tri 13298 138 13386 226 ne
rect 13386 190 13440 226
rect 13560 190 15775 310
rect 13386 138 15775 190
rect 12886 88 13288 138
rect 12366 58 12788 88
rect 11874 0 12268 58
tri 12268 0 12326 58 sw
tri 12366 0 12424 58 ne
rect 12424 0 12788 58
tri 12788 0 12876 88 sw
tri 12886 0 12974 88 ne
rect 12974 58 13288 88
tri 13288 58 13368 138 sw
tri 13386 58 13466 138 ne
rect 13466 58 14075 138
rect 12974 0 13368 58
rect -1025 -40 -324 0
tri -324 -40 -284 0 sw
tri -226 -40 -186 0 ne
rect -186 -40 226 0
rect -1025 -88 -284 -40
rect -1025 -188 -925 -88
rect -825 -138 -284 -88
tri -284 -138 -186 -40 sw
tri -186 -138 -88 -40 ne
rect -88 -98 226 -40
tri 226 -98 324 0 sw
tri 324 -98 422 0 ne
rect 422 -98 776 0
tri 776 -98 874 0 sw
tri 874 -98 972 0 ne
rect 972 -98 1326 0
tri 1326 -98 1424 0 sw
tri 1424 -98 1522 0 ne
rect 1522 -98 1876 0
tri 1876 -98 1974 0 sw
tri 1974 -98 2072 0 ne
rect 2072 -98 2426 0
tri 2426 -98 2524 0 sw
tri 2524 -98 2622 0 ne
rect 2622 -98 2976 0
tri 2976 -98 3074 0 sw
tri 3074 -98 3172 0 ne
rect 3172 -98 3526 0
tri 3526 -98 3624 0 sw
tri 3624 -98 3722 0 ne
rect 3722 -98 4076 0
tri 4076 -98 4174 0 sw
tri 4174 -98 4272 0 ne
rect 4272 -98 4626 0
tri 4626 -98 4724 0 sw
tri 4724 -98 4822 0 ne
rect 4822 -98 5176 0
tri 5176 -98 5274 0 sw
tri 5274 -98 5372 0 ne
rect 5372 -98 5726 0
tri 5726 -98 5824 0 sw
tri 5824 -98 5922 0 ne
rect 5922 -98 6276 0
tri 6276 -98 6374 0 sw
tri 6374 -98 6472 0 ne
rect 6472 -98 6826 0
tri 6826 -98 6924 0 sw
tri 6924 -98 7022 0 ne
rect 7022 -98 7376 0
tri 7376 -98 7474 0 sw
tri 7474 -98 7572 0 ne
rect 7572 -98 7926 0
tri 7926 -98 8024 0 sw
tri 8024 -98 8122 0 ne
rect 8122 -98 8476 0
tri 8476 -98 8574 0 sw
tri 8574 -98 8672 0 ne
rect 8672 -98 9026 0
tri 9026 -98 9124 0 sw
tri 9124 -98 9222 0 ne
rect 9222 -98 9576 0
tri 9576 -98 9674 0 sw
tri 9674 -98 9772 0 ne
rect 9772 -98 10126 0
tri 10126 -98 10224 0 sw
tri 10224 -98 10322 0 ne
rect 10322 -98 10676 0
tri 10676 -98 10774 0 sw
tri 10774 -98 10872 0 ne
rect 10872 -98 11226 0
tri 11226 -98 11324 0 sw
tri 11324 -98 11422 0 ne
rect 11422 -98 11776 0
tri 11776 -98 11874 0 sw
tri 11874 -98 11972 0 ne
rect 11972 -98 12326 0
tri 12326 -98 12424 0 sw
tri 12424 -98 12522 0 ne
rect 12522 -98 12876 0
tri 12876 -98 12974 0 sw
tri 12974 -98 13072 0 ne
rect 13072 -40 13368 0
tri 13368 -40 13466 58 sw
tri 13466 -40 13564 58 ne
rect 13564 38 14075 58
rect 14175 38 15775 138
rect 13564 -40 15775 38
rect 13072 -98 13466 -40
rect -88 -138 324 -98
tri 324 -138 364 -98 sw
tri 422 -138 462 -98 ne
rect 462 -138 874 -98
rect -825 -188 -186 -138
rect -1025 -236 -186 -188
tri -186 -236 -88 -138 sw
tri -88 -236 10 -138 ne
rect 10 -236 364 -138
tri 364 -236 462 -138 sw
tri 462 -236 560 -138 ne
rect 560 -186 874 -138
tri 874 -186 962 -98 sw
tri 972 -186 1060 -98 ne
rect 1060 -138 1424 -98
tri 1424 -138 1464 -98 sw
tri 1522 -138 1562 -98 ne
rect 1562 -138 1974 -98
rect 1060 -186 1464 -138
rect 560 -236 962 -186
rect -1025 -240 -88 -236
rect -1025 -360 -310 -240
rect -190 -324 -88 -240
tri -88 -324 0 -236 sw
tri 10 -324 98 -236 ne
rect 98 -240 462 -236
rect 98 -324 240 -240
rect -190 -360 0 -324
rect -1025 -364 0 -360
tri 0 -364 40 -324 sw
tri 98 -364 138 -324 ne
rect 138 -360 240 -324
rect 360 -324 462 -240
tri 462 -324 550 -236 sw
tri 560 -324 648 -236 ne
rect 648 -240 962 -236
rect 648 -324 790 -240
rect 360 -360 550 -324
rect 138 -364 550 -360
tri 550 -364 590 -324 sw
tri 648 -364 688 -324 ne
rect 688 -360 790 -324
rect 910 -266 962 -240
tri 962 -266 1042 -186 sw
tri 1060 -266 1140 -186 ne
rect 1140 -236 1464 -186
tri 1464 -236 1562 -138 sw
tri 1562 -236 1660 -138 ne
rect 1660 -186 1974 -138
tri 1974 -186 2062 -98 sw
tri 2072 -186 2160 -98 ne
rect 2160 -138 2524 -98
tri 2524 -138 2564 -98 sw
tri 2622 -138 2662 -98 ne
rect 2662 -138 3074 -98
rect 2160 -186 2564 -138
rect 1660 -236 2062 -186
rect 1140 -240 1562 -236
rect 1140 -266 1340 -240
rect 910 -360 1042 -266
rect 688 -364 1042 -360
tri 1042 -364 1140 -266 sw
tri 1140 -364 1238 -266 ne
rect 1238 -360 1340 -266
rect 1460 -324 1562 -240
tri 1562 -324 1650 -236 sw
tri 1660 -324 1748 -236 ne
rect 1748 -240 2062 -236
rect 1748 -324 1890 -240
rect 1460 -360 1650 -324
rect 1238 -364 1650 -360
tri 1650 -364 1690 -324 sw
tri 1748 -364 1788 -324 ne
rect 1788 -360 1890 -324
rect 2010 -266 2062 -240
tri 2062 -266 2142 -186 sw
tri 2160 -266 2240 -186 ne
rect 2240 -236 2564 -186
tri 2564 -236 2662 -138 sw
tri 2662 -236 2760 -138 ne
rect 2760 -186 3074 -138
tri 3074 -186 3162 -98 sw
tri 3172 -186 3260 -98 ne
rect 3260 -138 3624 -98
tri 3624 -138 3664 -98 sw
tri 3722 -138 3762 -98 ne
rect 3762 -138 4174 -98
rect 3260 -186 3664 -138
rect 2760 -236 3162 -186
rect 2240 -240 2662 -236
rect 2240 -266 2440 -240
rect 2010 -360 2142 -266
rect 1788 -364 2142 -360
tri 2142 -364 2240 -266 sw
tri 2240 -324 2298 -266 ne
rect 2298 -324 2440 -266
tri 2298 -364 2338 -324 ne
rect 2338 -360 2440 -324
rect 2560 -324 2662 -240
tri 2662 -324 2750 -236 sw
tri 2760 -324 2848 -236 ne
rect 2848 -240 3162 -236
rect 2848 -324 2990 -240
rect 2560 -360 2750 -324
rect 2338 -364 2750 -360
tri 2750 -364 2790 -324 sw
tri 2848 -364 2888 -324 ne
rect 2888 -360 2990 -324
rect 3110 -266 3162 -240
tri 3162 -266 3242 -186 sw
tri 3260 -266 3340 -186 ne
rect 3340 -236 3664 -186
tri 3664 -236 3762 -138 sw
tri 3762 -236 3860 -138 ne
rect 3860 -186 4174 -138
tri 4174 -186 4262 -98 sw
tri 4272 -186 4360 -98 ne
rect 4360 -138 4724 -98
tri 4724 -138 4764 -98 sw
tri 4822 -138 4862 -98 ne
rect 4862 -138 5274 -98
rect 4360 -186 4764 -138
rect 3860 -236 4262 -186
rect 3340 -240 3762 -236
rect 3340 -266 3540 -240
rect 3110 -360 3242 -266
rect 2888 -364 3242 -360
tri 3242 -364 3340 -266 sw
tri 3340 -324 3398 -266 ne
rect 3398 -324 3540 -266
tri 3398 -364 3438 -324 ne
rect 3438 -360 3540 -324
rect 3660 -324 3762 -240
tri 3762 -324 3850 -236 sw
tri 3860 -324 3948 -236 ne
rect 3948 -240 4262 -236
rect 3948 -324 4090 -240
rect 3660 -360 3850 -324
rect 3438 -364 3850 -360
tri 3850 -364 3890 -324 sw
tri 3948 -364 3988 -324 ne
rect 3988 -360 4090 -324
rect 4210 -266 4262 -240
tri 4262 -266 4342 -186 sw
tri 4360 -266 4440 -186 ne
rect 4440 -236 4764 -186
tri 4764 -236 4862 -138 sw
tri 4862 -236 4960 -138 ne
rect 4960 -186 5274 -138
tri 5274 -186 5362 -98 sw
tri 5372 -186 5460 -98 ne
rect 5460 -138 5824 -98
tri 5824 -138 5864 -98 sw
tri 5922 -138 5962 -98 ne
rect 5962 -138 6374 -98
rect 5460 -186 5864 -138
rect 4960 -236 5362 -186
rect 4440 -240 4862 -236
rect 4440 -266 4640 -240
rect 4210 -360 4342 -266
rect 3988 -364 4342 -360
tri 4342 -364 4440 -266 sw
tri 4440 -364 4538 -266 ne
rect 4538 -360 4640 -266
rect 4760 -324 4862 -240
tri 4862 -324 4950 -236 sw
tri 4960 -324 5048 -236 ne
rect 5048 -240 5362 -236
rect 5048 -324 5190 -240
rect 4760 -360 4950 -324
rect 4538 -364 4950 -360
tri 4950 -364 4990 -324 sw
tri 5048 -364 5088 -324 ne
rect 5088 -360 5190 -324
rect 5310 -266 5362 -240
tri 5362 -266 5442 -186 sw
tri 5460 -266 5540 -186 ne
rect 5540 -236 5864 -186
tri 5864 -236 5962 -138 sw
tri 5962 -236 6060 -138 ne
rect 6060 -186 6374 -138
tri 6374 -186 6462 -98 sw
tri 6472 -186 6560 -98 ne
rect 6560 -138 6924 -98
tri 6924 -138 6964 -98 sw
tri 7022 -138 7062 -98 ne
rect 7062 -138 7474 -98
rect 6560 -186 6964 -138
rect 6060 -236 6462 -186
rect 5540 -240 5962 -236
rect 5540 -266 5740 -240
rect 5310 -360 5442 -266
rect 5088 -364 5442 -360
tri 5442 -364 5540 -266 sw
tri 5540 -324 5598 -266 ne
rect 5598 -324 5740 -266
tri 5598 -364 5638 -324 ne
rect 5638 -360 5740 -324
rect 5860 -324 5962 -240
tri 5962 -324 6050 -236 sw
tri 6060 -324 6148 -236 ne
rect 6148 -240 6462 -236
rect 6148 -324 6290 -240
rect 5860 -360 6050 -324
rect 5638 -364 6050 -360
tri 6050 -364 6090 -324 sw
tri 6148 -364 6188 -324 ne
rect 6188 -360 6290 -324
rect 6410 -266 6462 -240
tri 6462 -266 6542 -186 sw
tri 6560 -266 6640 -186 ne
rect 6640 -236 6964 -186
tri 6964 -236 7062 -138 sw
tri 7062 -236 7160 -138 ne
rect 7160 -186 7474 -138
tri 7474 -186 7562 -98 sw
tri 7572 -186 7660 -98 ne
rect 7660 -138 8024 -98
tri 8024 -138 8064 -98 sw
tri 8122 -138 8162 -98 ne
rect 8162 -138 8574 -98
rect 7660 -186 8064 -138
rect 7160 -236 7562 -186
rect 6640 -240 7062 -236
rect 6640 -266 6840 -240
rect 6410 -360 6542 -266
rect 6188 -364 6542 -360
tri 6542 -364 6640 -266 sw
tri 6640 -324 6698 -266 ne
rect 6698 -324 6840 -266
tri 6698 -364 6738 -324 ne
rect 6738 -360 6840 -324
rect 6960 -324 7062 -240
tri 7062 -324 7150 -236 sw
tri 7160 -324 7248 -236 ne
rect 7248 -240 7562 -236
rect 7248 -324 7390 -240
rect 6960 -360 7150 -324
rect 6738 -364 7150 -360
tri 7150 -364 7190 -324 sw
tri 7248 -364 7288 -324 ne
rect 7288 -360 7390 -324
rect 7510 -266 7562 -240
tri 7562 -266 7642 -186 sw
tri 7660 -266 7740 -186 ne
rect 7740 -236 8064 -186
tri 8064 -236 8162 -138 sw
tri 8162 -236 8260 -138 ne
rect 8260 -186 8574 -138
tri 8574 -186 8662 -98 sw
tri 8672 -186 8760 -98 ne
rect 8760 -138 9124 -98
tri 9124 -138 9164 -98 sw
tri 9222 -138 9262 -98 ne
rect 9262 -138 9674 -98
rect 8760 -186 9164 -138
rect 8260 -236 8662 -186
rect 7740 -240 8162 -236
rect 7740 -266 7940 -240
rect 7510 -360 7642 -266
rect 7288 -364 7642 -360
tri 7642 -364 7740 -266 sw
tri 7740 -364 7838 -266 ne
rect 7838 -360 7940 -266
rect 8060 -324 8162 -240
tri 8162 -324 8250 -236 sw
tri 8260 -324 8348 -236 ne
rect 8348 -240 8662 -236
rect 8348 -324 8490 -240
rect 8060 -360 8250 -324
rect 7838 -364 8250 -360
tri 8250 -364 8290 -324 sw
tri 8348 -364 8388 -324 ne
rect 8388 -360 8490 -324
rect 8610 -266 8662 -240
tri 8662 -266 8742 -186 sw
tri 8760 -266 8840 -186 ne
rect 8840 -236 9164 -186
tri 9164 -236 9262 -138 sw
tri 9262 -236 9360 -138 ne
rect 9360 -186 9674 -138
tri 9674 -186 9762 -98 sw
tri 9772 -186 9860 -98 ne
rect 9860 -138 10224 -98
tri 10224 -138 10264 -98 sw
tri 10322 -138 10362 -98 ne
rect 10362 -138 10774 -98
rect 9860 -186 10264 -138
rect 9360 -236 9762 -186
rect 8840 -240 9262 -236
rect 8840 -266 9040 -240
rect 8610 -360 8742 -266
rect 8388 -364 8742 -360
tri 8742 -364 8840 -266 sw
tri 8840 -324 8898 -266 ne
rect 8898 -324 9040 -266
tri 8898 -364 8938 -324 ne
rect 8938 -360 9040 -324
rect 9160 -324 9262 -240
tri 9262 -324 9350 -236 sw
tri 9360 -324 9448 -236 ne
rect 9448 -240 9762 -236
rect 9448 -324 9590 -240
rect 9160 -360 9350 -324
rect 8938 -364 9350 -360
tri 9350 -364 9390 -324 sw
tri 9448 -364 9488 -324 ne
rect 9488 -360 9590 -324
rect 9710 -266 9762 -240
tri 9762 -266 9842 -186 sw
tri 9860 -266 9940 -186 ne
rect 9940 -236 10264 -186
tri 10264 -236 10362 -138 sw
tri 10362 -236 10460 -138 ne
rect 10460 -186 10774 -138
tri 10774 -186 10862 -98 sw
tri 10872 -186 10960 -98 ne
rect 10960 -138 11324 -98
tri 11324 -138 11364 -98 sw
tri 11422 -138 11462 -98 ne
rect 11462 -138 11874 -98
rect 10960 -186 11364 -138
rect 10460 -236 10862 -186
rect 9940 -240 10362 -236
rect 9940 -266 10140 -240
rect 9710 -360 9842 -266
rect 9488 -364 9842 -360
tri 9842 -364 9940 -266 sw
tri 9940 -324 9998 -266 ne
rect 9998 -324 10140 -266
tri 9998 -364 10038 -324 ne
rect 10038 -360 10140 -324
rect 10260 -324 10362 -240
tri 10362 -324 10450 -236 sw
tri 10460 -324 10548 -236 ne
rect 10548 -240 10862 -236
rect 10548 -324 10690 -240
rect 10260 -360 10450 -324
rect 10038 -364 10450 -360
tri 10450 -364 10490 -324 sw
tri 10548 -364 10588 -324 ne
rect 10588 -360 10690 -324
rect 10810 -266 10862 -240
tri 10862 -266 10942 -186 sw
tri 10960 -266 11040 -186 ne
rect 11040 -236 11364 -186
tri 11364 -236 11462 -138 sw
tri 11462 -236 11560 -138 ne
rect 11560 -186 11874 -138
tri 11874 -186 11962 -98 sw
tri 11972 -186 12060 -98 ne
rect 12060 -138 12424 -98
tri 12424 -138 12464 -98 sw
tri 12522 -138 12562 -98 ne
rect 12562 -138 12974 -98
rect 12060 -186 12464 -138
rect 11560 -236 11962 -186
rect 11040 -240 11462 -236
rect 11040 -266 11240 -240
rect 10810 -360 10942 -266
rect 10588 -364 10942 -360
tri 10942 -364 11040 -266 sw
tri 11040 -364 11138 -266 ne
rect 11138 -360 11240 -266
rect 11360 -324 11462 -240
tri 11462 -324 11550 -236 sw
tri 11560 -324 11648 -236 ne
rect 11648 -240 11962 -236
rect 11648 -324 11790 -240
rect 11360 -360 11550 -324
rect 11138 -364 11550 -360
tri 11550 -364 11590 -324 sw
tri 11648 -364 11688 -324 ne
rect 11688 -360 11790 -324
rect 11910 -266 11962 -240
tri 11962 -266 12042 -186 sw
tri 12060 -266 12140 -186 ne
rect 12140 -236 12464 -186
tri 12464 -236 12562 -138 sw
tri 12562 -236 12660 -138 ne
rect 12660 -186 12974 -138
tri 12974 -186 13062 -98 sw
tri 13072 -186 13160 -98 ne
rect 13160 -138 13466 -98
tri 13466 -138 13564 -40 sw
tri 13564 -138 13662 -40 ne
rect 13662 -138 15775 -40
rect 13160 -186 13564 -138
rect 12660 -236 13062 -186
rect 12140 -240 12562 -236
rect 12140 -266 12340 -240
rect 11910 -360 12042 -266
rect 11688 -364 12042 -360
tri 12042 -364 12140 -266 sw
tri 12140 -324 12198 -266 ne
rect 12198 -324 12340 -266
tri 12198 -364 12238 -324 ne
rect 12238 -360 12340 -324
rect 12460 -324 12562 -240
tri 12562 -324 12650 -236 sw
tri 12660 -324 12748 -236 ne
rect 12748 -240 13062 -236
rect 12748 -324 12890 -240
rect 12460 -360 12650 -324
rect 12238 -364 12650 -360
tri 12650 -364 12690 -324 sw
tri 12748 -364 12788 -324 ne
rect 12788 -360 12890 -324
rect 13010 -266 13062 -240
tri 13062 -266 13142 -186 sw
tri 13160 -266 13240 -186 ne
rect 13240 -236 13564 -186
tri 13564 -236 13662 -138 sw
rect 13240 -240 14275 -236
rect 13240 -266 13440 -240
rect 13010 -360 13142 -266
rect 12788 -364 13142 -360
tri 13142 -364 13240 -266 sw
tri 13240 -324 13298 -266 ne
rect 13298 -324 13440 -266
tri 13298 -364 13338 -324 ne
rect 13338 -360 13440 -324
rect 13560 -360 14275 -240
rect 13338 -364 14275 -360
tri -412 -462 -314 -364 ne
rect -314 -462 40 -364
tri 40 -462 138 -364 sw
tri 138 -462 236 -364 ne
rect 236 -462 590 -364
tri 590 -462 688 -364 sw
tri 688 -462 786 -364 ne
rect 786 -462 1140 -364
tri 1140 -462 1238 -364 sw
tri 1238 -462 1336 -364 ne
rect 1336 -462 1690 -364
tri 1690 -462 1788 -364 sw
tri 1788 -462 1886 -364 ne
rect 1886 -462 2240 -364
tri 2240 -462 2338 -364 sw
tri 2338 -462 2436 -364 ne
rect 2436 -462 2790 -364
tri 2790 -462 2888 -364 sw
tri 2888 -462 2986 -364 ne
rect 2986 -462 3340 -364
tri 3340 -462 3438 -364 sw
tri 3438 -462 3536 -364 ne
rect 3536 -462 3890 -364
tri 3890 -462 3988 -364 sw
tri 3988 -462 4086 -364 ne
rect 4086 -462 4440 -364
tri 4440 -462 4538 -364 sw
tri 4538 -462 4636 -364 ne
rect 4636 -462 4990 -364
tri 4990 -462 5088 -364 sw
tri 5088 -462 5186 -364 ne
rect 5186 -462 5540 -364
tri 5540 -462 5638 -364 sw
tri 5638 -462 5736 -364 ne
rect 5736 -462 6090 -364
tri 6090 -462 6188 -364 sw
tri 6188 -462 6286 -364 ne
rect 6286 -462 6640 -364
tri 6640 -462 6738 -364 sw
tri 6738 -462 6836 -364 ne
rect 6836 -462 7190 -364
tri 7190 -462 7288 -364 sw
tri 7288 -462 7386 -364 ne
rect 7386 -462 7740 -364
tri 7740 -462 7838 -364 sw
tri 7838 -462 7936 -364 ne
rect 7936 -462 8290 -364
tri 8290 -462 8388 -364 sw
tri 8388 -462 8486 -364 ne
rect 8486 -462 8840 -364
tri 8840 -462 8938 -364 sw
tri 8938 -462 9036 -364 ne
rect 9036 -462 9390 -364
tri 9390 -462 9488 -364 sw
tri 9488 -462 9586 -364 ne
rect 9586 -462 9940 -364
tri 9940 -462 10038 -364 sw
tri 10038 -462 10136 -364 ne
rect 10136 -462 10490 -364
tri 10490 -462 10588 -364 sw
tri 10588 -462 10686 -364 ne
rect 10686 -462 11040 -364
tri 11040 -462 11138 -364 sw
tri 11138 -462 11236 -364 ne
rect 11236 -462 11590 -364
tri 11590 -462 11688 -364 sw
tri 11688 -462 11786 -364 ne
rect 11786 -462 12140 -364
tri 12140 -462 12238 -364 sw
tri 12238 -462 12336 -364 ne
rect 12336 -462 12690 -364
tri 12690 -462 12788 -364 sw
tri 12788 -462 12886 -364 ne
rect 12886 -462 13240 -364
tri 13240 -462 13338 -364 sw
tri 13338 -462 13436 -364 ne
rect -314 -875 138 -462
rect -314 -975 -138 -875
rect -38 -975 138 -875
rect -314 -1575 138 -975
rect 236 -1075 688 -462
rect 786 -875 1238 -462
rect 786 -975 962 -875
rect 1062 -975 1238 -875
rect 786 -1575 1238 -975
rect 1336 -1075 1788 -462
rect 1886 -875 2338 -462
rect 1886 -975 2062 -875
rect 2162 -975 2338 -875
rect 1886 -1575 2338 -975
rect 2436 -1075 2888 -462
rect 2986 -875 3438 -462
rect 2986 -975 3162 -875
rect 3262 -975 3438 -875
rect 2986 -1575 3438 -975
rect 3536 -1075 3988 -462
rect 4086 -875 4538 -462
rect 4086 -975 4262 -875
rect 4362 -975 4538 -875
rect 4086 -1575 4538 -975
rect 4636 -1075 5088 -462
rect 5186 -875 5638 -462
rect 5186 -975 5362 -875
rect 5462 -975 5638 -875
rect 5186 -1575 5638 -975
rect 5736 -1075 6188 -462
rect 6286 -875 6738 -462
rect 6286 -975 6462 -875
rect 6562 -975 6738 -875
rect 6286 -1575 6738 -975
rect 6836 -1075 7288 -462
rect 7386 -875 7838 -462
rect 7386 -975 7562 -875
rect 7662 -975 7838 -875
rect 7386 -1575 7838 -975
rect 7936 -1075 8388 -462
rect 8486 -875 8938 -462
rect 8486 -975 8662 -875
rect 8762 -975 8938 -875
rect 8486 -1575 8938 -975
rect 9036 -1075 9488 -462
rect 9586 -875 10038 -462
rect 9586 -975 9762 -875
rect 9862 -975 10038 -875
rect 9586 -1575 10038 -975
rect 10136 -1075 10588 -462
rect 10686 -875 11138 -462
rect 10686 -975 10862 -875
rect 10962 -975 11138 -875
rect 10686 -1575 11138 -975
rect 11236 -1075 11688 -462
rect 11786 -875 12238 -462
rect 11786 -975 11962 -875
rect 12062 -975 12238 -875
rect 11786 -1575 12238 -975
rect 12336 -1075 12788 -462
rect 12886 -875 13338 -462
rect 12886 -975 13062 -875
rect 13162 -975 13338 -875
rect 12886 -1575 13338 -975
rect 13436 -688 14275 -364
rect 13436 -1075 13888 -688
rect 14775 -1575 15775 -138
rect -525 -2575 15775 -1575
<< via4 >>
rect -310 13390 -190 13510
rect 240 13390 360 13510
rect 790 13390 910 13510
rect 1340 13390 1460 13510
rect 1890 13390 2010 13510
rect 2440 13390 2560 13510
rect 2990 13390 3110 13510
rect 3540 13390 3660 13510
rect 4090 13390 4210 13510
rect 4640 13390 4760 13510
rect 5190 13390 5310 13510
rect 5740 13390 5860 13510
rect 6290 13390 6410 13510
rect 6840 13390 6960 13510
rect 7390 13390 7510 13510
rect 7940 13390 8060 13510
rect 8490 13390 8610 13510
rect 9040 13390 9160 13510
rect 9590 13390 9710 13510
rect 10140 13390 10260 13510
rect 10690 13390 10810 13510
rect 11240 13390 11360 13510
rect 11790 13390 11910 13510
rect 12340 13390 12460 13510
rect 12890 13390 13010 13510
rect 13440 13390 13560 13510
rect -310 12840 -190 12960
rect 240 12840 360 12960
rect 790 12840 910 12960
rect 1340 12840 1460 12960
rect 1890 12840 2010 12960
rect 2440 12840 2560 12960
rect 2990 12840 3110 12960
rect 3540 12840 3660 12960
rect 4090 12840 4210 12960
rect 4640 12840 4760 12960
rect 5190 12840 5310 12960
rect 5740 12840 5860 12960
rect 6290 12840 6410 12960
rect 6840 12840 6960 12960
rect 7390 12840 7510 12960
rect 7940 12840 8060 12960
rect 8490 12840 8610 12960
rect 9040 12840 9160 12960
rect 9590 12840 9710 12960
rect 10140 12840 10260 12960
rect 10690 12840 10810 12960
rect 11240 12840 11360 12960
rect 11790 12840 11910 12960
rect 12340 12840 12460 12960
rect 12890 12840 13010 12960
rect 13440 12840 13560 12960
rect -310 12290 -190 12410
rect 240 12290 360 12410
rect 790 12290 910 12410
rect 1340 12290 1460 12410
rect 1890 12290 2010 12410
rect 2440 12290 2560 12410
rect 2990 12290 3110 12410
rect 3540 12290 3660 12410
rect 4090 12290 4210 12410
rect 4640 12290 4760 12410
rect 5190 12290 5310 12410
rect 5740 12290 5860 12410
rect 6290 12290 6410 12410
rect 6840 12290 6960 12410
rect 7390 12290 7510 12410
rect 7940 12290 8060 12410
rect 8490 12290 8610 12410
rect 9040 12290 9160 12410
rect 9590 12290 9710 12410
rect 10140 12290 10260 12410
rect 10690 12290 10810 12410
rect 11240 12290 11360 12410
rect 11790 12290 11910 12410
rect 12340 12290 12460 12410
rect 12890 12290 13010 12410
rect 13440 12290 13560 12410
rect -310 11740 -190 11860
rect 240 11740 360 11860
rect 790 11740 910 11860
rect 1340 11740 1460 11860
rect 1890 11740 2010 11860
rect 2440 11740 2560 11860
rect 2990 11740 3110 11860
rect 3540 11740 3660 11860
rect 4090 11740 4210 11860
rect 4640 11740 4760 11860
rect 5190 11740 5310 11860
rect 5740 11740 5860 11860
rect 6290 11740 6410 11860
rect 6840 11740 6960 11860
rect 7390 11740 7510 11860
rect 7940 11740 8060 11860
rect 8490 11740 8610 11860
rect 9040 11740 9160 11860
rect 9590 11740 9710 11860
rect 10140 11740 10260 11860
rect 10690 11740 10810 11860
rect 11240 11740 11360 11860
rect 11790 11740 11910 11860
rect 12340 11740 12460 11860
rect 12890 11740 13010 11860
rect 13440 11740 13560 11860
rect -310 11190 -190 11310
rect 240 11190 360 11310
rect 790 11190 910 11310
rect 1340 11190 1460 11310
rect 1890 11190 2010 11310
rect 2440 11190 2560 11310
rect 2990 11190 3110 11310
rect 3540 11190 3660 11310
rect 4090 11190 4210 11310
rect 4640 11190 4760 11310
rect 5190 11190 5310 11310
rect 5740 11190 5860 11310
rect 6290 11190 6410 11310
rect 6840 11190 6960 11310
rect 7390 11190 7510 11310
rect 7940 11190 8060 11310
rect 8490 11190 8610 11310
rect 9040 11190 9160 11310
rect 9590 11190 9710 11310
rect 10140 11190 10260 11310
rect 10690 11190 10810 11310
rect 11240 11190 11360 11310
rect 11790 11190 11910 11310
rect 12340 11190 12460 11310
rect 12890 11190 13010 11310
rect 13440 11190 13560 11310
rect -310 10640 -190 10760
rect 240 10640 360 10760
rect 790 10640 910 10760
rect 1340 10640 1460 10760
rect 1890 10640 2010 10760
rect 2440 10640 2560 10760
rect 2990 10640 3110 10760
rect 3540 10640 3660 10760
rect 4090 10640 4210 10760
rect 4640 10640 4760 10760
rect 5190 10640 5310 10760
rect 5740 10640 5860 10760
rect 6290 10640 6410 10760
rect 6840 10640 6960 10760
rect 7390 10640 7510 10760
rect 7940 10640 8060 10760
rect 8490 10640 8610 10760
rect 9040 10640 9160 10760
rect 9590 10640 9710 10760
rect 10140 10640 10260 10760
rect 10690 10640 10810 10760
rect 11240 10640 11360 10760
rect 11790 10640 11910 10760
rect 12340 10640 12460 10760
rect 12890 10640 13010 10760
rect 13440 10640 13560 10760
rect -310 10090 -190 10210
rect 240 10090 360 10210
rect 790 10090 910 10210
rect 1340 10090 1460 10210
rect 1890 10090 2010 10210
rect 2440 10090 2560 10210
rect 2990 10090 3110 10210
rect 3540 10090 3660 10210
rect 4090 10090 4210 10210
rect 4640 10090 4760 10210
rect 5190 10090 5310 10210
rect 5740 10090 5860 10210
rect 6290 10090 6410 10210
rect 6840 10090 6960 10210
rect 7390 10090 7510 10210
rect 7940 10090 8060 10210
rect 8490 10090 8610 10210
rect 9040 10090 9160 10210
rect 9590 10090 9710 10210
rect 10140 10090 10260 10210
rect 10690 10090 10810 10210
rect 11240 10090 11360 10210
rect 11790 10090 11910 10210
rect 12340 10090 12460 10210
rect 12890 10090 13010 10210
rect 13440 10090 13560 10210
rect -310 9540 -190 9660
rect 240 9540 360 9660
rect 790 9540 910 9660
rect 1340 9540 1460 9660
rect 1890 9540 2010 9660
rect 2440 9540 2560 9660
rect 2990 9540 3110 9660
rect 3540 9540 3660 9660
rect 4090 9540 4210 9660
rect 4640 9540 4760 9660
rect 5190 9540 5310 9660
rect 5740 9540 5860 9660
rect 6290 9540 6410 9660
rect 6840 9540 6960 9660
rect 7390 9540 7510 9660
rect 7940 9540 8060 9660
rect 8490 9540 8610 9660
rect 9040 9540 9160 9660
rect 9590 9540 9710 9660
rect 10140 9540 10260 9660
rect 10690 9540 10810 9660
rect 11240 9540 11360 9660
rect 11790 9540 11910 9660
rect 12340 9540 12460 9660
rect 12890 9540 13010 9660
rect 13440 9540 13560 9660
rect -310 8990 -190 9110
rect 240 8990 360 9110
rect 790 8990 910 9110
rect 1340 8990 1460 9110
rect 1890 8990 2010 9110
rect 2440 8990 2560 9110
rect 2990 8990 3110 9110
rect 3540 8990 3660 9110
rect 4090 8990 4210 9110
rect 4640 8990 4760 9110
rect 5190 8990 5310 9110
rect 5740 8990 5860 9110
rect 6290 8990 6410 9110
rect 6840 8990 6960 9110
rect 7390 8990 7510 9110
rect 7940 8990 8060 9110
rect 8490 8990 8610 9110
rect 9040 8990 9160 9110
rect 9590 8990 9710 9110
rect 10140 8990 10260 9110
rect 10690 8990 10810 9110
rect 11240 8990 11360 9110
rect 11790 8990 11910 9110
rect 12340 8990 12460 9110
rect 12890 8990 13010 9110
rect 13440 8990 13560 9110
rect -310 8440 -190 8560
rect 240 8440 360 8560
rect 790 8440 910 8560
rect 1340 8440 1460 8560
rect 1890 8440 2010 8560
rect 2440 8440 2560 8560
rect 2990 8440 3110 8560
rect 3540 8440 3660 8560
rect 4090 8440 4210 8560
rect 4640 8440 4760 8560
rect 5190 8440 5310 8560
rect 5740 8440 5860 8560
rect 6290 8440 6410 8560
rect 6840 8440 6960 8560
rect 7390 8440 7510 8560
rect 7940 8440 8060 8560
rect 8490 8440 8610 8560
rect 9040 8440 9160 8560
rect 9590 8440 9710 8560
rect 10140 8440 10260 8560
rect 10690 8440 10810 8560
rect 11240 8440 11360 8560
rect 11790 8440 11910 8560
rect 12340 8440 12460 8560
rect 12890 8440 13010 8560
rect 13440 8440 13560 8560
rect -310 7890 -190 8010
rect 240 7890 360 8010
rect 790 7890 910 8010
rect 1340 7890 1460 8010
rect 1890 7890 2010 8010
rect 2440 7890 2560 8010
rect 2990 7890 3110 8010
rect 3540 7890 3660 8010
rect 4090 7890 4210 8010
rect 4640 7890 4760 8010
rect 5190 7890 5310 8010
rect 5740 7890 5860 8010
rect 6290 7890 6410 8010
rect 6840 7890 6960 8010
rect 7390 7890 7510 8010
rect 7940 7890 8060 8010
rect 8490 7890 8610 8010
rect 9040 7890 9160 8010
rect 9590 7890 9710 8010
rect 10140 7890 10260 8010
rect 10690 7890 10810 8010
rect 11240 7890 11360 8010
rect 11790 7890 11910 8010
rect 12340 7890 12460 8010
rect 12890 7890 13010 8010
rect 13440 7890 13560 8010
rect -310 7340 -190 7460
rect 240 7340 360 7460
rect 790 7340 910 7460
rect 1340 7340 1460 7460
rect 1890 7340 2010 7460
rect 2440 7340 2560 7460
rect 2990 7340 3110 7460
rect 3540 7340 3660 7460
rect 4090 7340 4210 7460
rect 4640 7340 4760 7460
rect 5190 7340 5310 7460
rect 5740 7340 5860 7460
rect 6290 7340 6410 7460
rect 6840 7340 6960 7460
rect 7390 7340 7510 7460
rect 7940 7340 8060 7460
rect 8490 7340 8610 7460
rect 9040 7340 9160 7460
rect 9590 7340 9710 7460
rect 10140 7340 10260 7460
rect 10690 7340 10810 7460
rect 11240 7340 11360 7460
rect 11790 7340 11910 7460
rect 12340 7340 12460 7460
rect 12890 7340 13010 7460
rect 13440 7340 13560 7460
rect -310 6790 -190 6910
rect 240 6790 360 6910
rect 790 6790 910 6910
rect 1340 6790 1460 6910
rect 1890 6790 2010 6910
rect 2440 6790 2560 6910
rect 2990 6790 3110 6910
rect 3540 6790 3660 6910
rect 4090 6790 4210 6910
rect 4640 6790 4760 6910
rect 5190 6790 5310 6910
rect 5740 6790 5860 6910
rect 6290 6790 6410 6910
rect 6840 6790 6960 6910
rect 7390 6790 7510 6910
rect 7940 6790 8060 6910
rect 8490 6790 8610 6910
rect 9040 6790 9160 6910
rect 9590 6790 9710 6910
rect 10140 6790 10260 6910
rect 10690 6790 10810 6910
rect 11240 6790 11360 6910
rect 11790 6790 11910 6910
rect 12340 6790 12460 6910
rect 12890 6790 13010 6910
rect 13440 6790 13560 6910
rect -310 6240 -190 6360
rect 240 6240 360 6360
rect 790 6240 910 6360
rect 1340 6240 1460 6360
rect 1890 6240 2010 6360
rect 2440 6240 2560 6360
rect 2990 6240 3110 6360
rect 3540 6240 3660 6360
rect 4090 6240 4210 6360
rect 4640 6240 4760 6360
rect 5190 6240 5310 6360
rect 5740 6240 5860 6360
rect 6290 6240 6410 6360
rect 6840 6240 6960 6360
rect 7390 6240 7510 6360
rect 7940 6240 8060 6360
rect 8490 6240 8610 6360
rect 9040 6240 9160 6360
rect 9590 6240 9710 6360
rect 10140 6240 10260 6360
rect 10690 6240 10810 6360
rect 11240 6240 11360 6360
rect 11790 6240 11910 6360
rect 12340 6240 12460 6360
rect 12890 6240 13010 6360
rect 13440 6240 13560 6360
rect -310 5690 -190 5810
rect 240 5690 360 5810
rect 790 5690 910 5810
rect 1340 5690 1460 5810
rect 1890 5690 2010 5810
rect 2440 5690 2560 5810
rect 2990 5690 3110 5810
rect 3540 5690 3660 5810
rect 4090 5690 4210 5810
rect 4640 5690 4760 5810
rect 5190 5690 5310 5810
rect 5740 5690 5860 5810
rect 6290 5690 6410 5810
rect 6840 5690 6960 5810
rect 7390 5690 7510 5810
rect 7940 5690 8060 5810
rect 8490 5690 8610 5810
rect 9040 5690 9160 5810
rect 9590 5690 9710 5810
rect 10140 5690 10260 5810
rect 10690 5690 10810 5810
rect 11240 5690 11360 5810
rect 11790 5690 11910 5810
rect 12340 5690 12460 5810
rect 12890 5690 13010 5810
rect 13440 5690 13560 5810
rect -310 5140 -190 5260
rect 240 5140 360 5260
rect 790 5140 910 5260
rect 1340 5140 1460 5260
rect 1890 5140 2010 5260
rect 2440 5140 2560 5260
rect 2990 5140 3110 5260
rect 3540 5140 3660 5260
rect 4090 5140 4210 5260
rect 4640 5140 4760 5260
rect 5190 5140 5310 5260
rect 5740 5140 5860 5260
rect 6290 5140 6410 5260
rect 6840 5140 6960 5260
rect 7390 5140 7510 5260
rect 7940 5140 8060 5260
rect 8490 5140 8610 5260
rect 9040 5140 9160 5260
rect 9590 5140 9710 5260
rect 10140 5140 10260 5260
rect 10690 5140 10810 5260
rect 11240 5140 11360 5260
rect 11790 5140 11910 5260
rect 12340 5140 12460 5260
rect 12890 5140 13010 5260
rect 13440 5140 13560 5260
rect -310 4590 -190 4710
rect 240 4590 360 4710
rect 790 4590 910 4710
rect 1340 4590 1460 4710
rect 1890 4590 2010 4710
rect 2440 4590 2560 4710
rect 2990 4590 3110 4710
rect 3540 4590 3660 4710
rect 4090 4590 4210 4710
rect 4640 4590 4760 4710
rect 5190 4590 5310 4710
rect 5740 4590 5860 4710
rect 6290 4590 6410 4710
rect 6840 4590 6960 4710
rect 7390 4590 7510 4710
rect 7940 4590 8060 4710
rect 8490 4590 8610 4710
rect 9040 4590 9160 4710
rect 9590 4590 9710 4710
rect 10140 4590 10260 4710
rect 10690 4590 10810 4710
rect 11240 4590 11360 4710
rect 11790 4590 11910 4710
rect 12340 4590 12460 4710
rect 12890 4590 13010 4710
rect 13440 4590 13560 4710
rect -310 4040 -190 4160
rect 240 4040 360 4160
rect 790 4040 910 4160
rect 1340 4040 1460 4160
rect 1890 4040 2010 4160
rect 2440 4040 2560 4160
rect 2990 4040 3110 4160
rect 3540 4040 3660 4160
rect 4090 4040 4210 4160
rect 4640 4040 4760 4160
rect 5190 4040 5310 4160
rect 5740 4040 5860 4160
rect 6290 4040 6410 4160
rect 6840 4040 6960 4160
rect 7390 4040 7510 4160
rect 7940 4040 8060 4160
rect 8490 4040 8610 4160
rect 9040 4040 9160 4160
rect 9590 4040 9710 4160
rect 10140 4040 10260 4160
rect 10690 4040 10810 4160
rect 11240 4040 11360 4160
rect 11790 4040 11910 4160
rect 12340 4040 12460 4160
rect 12890 4040 13010 4160
rect 13440 4040 13560 4160
rect -310 3490 -190 3610
rect 240 3490 360 3610
rect 790 3490 910 3610
rect 1340 3490 1460 3610
rect 1890 3490 2010 3610
rect 2440 3490 2560 3610
rect 2990 3490 3110 3610
rect 3540 3490 3660 3610
rect 4090 3490 4210 3610
rect 4640 3490 4760 3610
rect 5190 3490 5310 3610
rect 5740 3490 5860 3610
rect 6290 3490 6410 3610
rect 6840 3490 6960 3610
rect 7390 3490 7510 3610
rect 7940 3490 8060 3610
rect 8490 3490 8610 3610
rect 9040 3490 9160 3610
rect 9590 3490 9710 3610
rect 10140 3490 10260 3610
rect 10690 3490 10810 3610
rect 11240 3490 11360 3610
rect 11790 3490 11910 3610
rect 12340 3490 12460 3610
rect 12890 3490 13010 3610
rect 13440 3490 13560 3610
rect -310 2940 -190 3060
rect 240 2940 360 3060
rect 790 2940 910 3060
rect 1340 2940 1460 3060
rect 1890 2940 2010 3060
rect 2440 2940 2560 3060
rect 2990 2940 3110 3060
rect 3540 2940 3660 3060
rect 4090 2940 4210 3060
rect 4640 2940 4760 3060
rect 5190 2940 5310 3060
rect 5740 2940 5860 3060
rect 6290 2940 6410 3060
rect 6840 2940 6960 3060
rect 7390 2940 7510 3060
rect 7940 2940 8060 3060
rect 8490 2940 8610 3060
rect 9040 2940 9160 3060
rect 9590 2940 9710 3060
rect 10140 2940 10260 3060
rect 10690 2940 10810 3060
rect 11240 2940 11360 3060
rect 11790 2940 11910 3060
rect 12340 2940 12460 3060
rect 12890 2940 13010 3060
rect 13440 2940 13560 3060
rect -310 2390 -190 2510
rect 240 2390 360 2510
rect 790 2390 910 2510
rect 1340 2390 1460 2510
rect 1890 2390 2010 2510
rect 2440 2390 2560 2510
rect 2990 2390 3110 2510
rect 3540 2390 3660 2510
rect 4090 2390 4210 2510
rect 4640 2390 4760 2510
rect 5190 2390 5310 2510
rect 5740 2390 5860 2510
rect 6290 2390 6410 2510
rect 6840 2390 6960 2510
rect 7390 2390 7510 2510
rect 7940 2390 8060 2510
rect 8490 2390 8610 2510
rect 9040 2390 9160 2510
rect 9590 2390 9710 2510
rect 10140 2390 10260 2510
rect 10690 2390 10810 2510
rect 11240 2390 11360 2510
rect 11790 2390 11910 2510
rect 12340 2390 12460 2510
rect 12890 2390 13010 2510
rect 13440 2390 13560 2510
rect -310 1840 -190 1960
rect 240 1840 360 1960
rect 790 1840 910 1960
rect 1340 1840 1460 1960
rect 1890 1840 2010 1960
rect 2440 1840 2560 1960
rect 2990 1840 3110 1960
rect 3540 1840 3660 1960
rect 4090 1840 4210 1960
rect 4640 1840 4760 1960
rect 5190 1840 5310 1960
rect 5740 1840 5860 1960
rect 6290 1840 6410 1960
rect 6840 1840 6960 1960
rect 7390 1840 7510 1960
rect 7940 1840 8060 1960
rect 8490 1840 8610 1960
rect 9040 1840 9160 1960
rect 9590 1840 9710 1960
rect 10140 1840 10260 1960
rect 10690 1840 10810 1960
rect 11240 1840 11360 1960
rect 11790 1840 11910 1960
rect 12340 1840 12460 1960
rect 12890 1840 13010 1960
rect 13440 1840 13560 1960
rect -310 1290 -190 1410
rect 240 1290 360 1410
rect 790 1290 910 1410
rect 1340 1290 1460 1410
rect 1890 1290 2010 1410
rect 2440 1290 2560 1410
rect 2990 1290 3110 1410
rect 3540 1290 3660 1410
rect 4090 1290 4210 1410
rect 4640 1290 4760 1410
rect 5190 1290 5310 1410
rect 5740 1290 5860 1410
rect 6290 1290 6410 1410
rect 6840 1290 6960 1410
rect 7390 1290 7510 1410
rect 7940 1290 8060 1410
rect 8490 1290 8610 1410
rect 9040 1290 9160 1410
rect 9590 1290 9710 1410
rect 10140 1290 10260 1410
rect 10690 1290 10810 1410
rect 11240 1290 11360 1410
rect 11790 1290 11910 1410
rect 12340 1290 12460 1410
rect 12890 1290 13010 1410
rect 13440 1290 13560 1410
rect -310 740 -190 860
rect 240 740 360 860
rect 790 740 910 860
rect 1340 740 1460 860
rect 1890 740 2010 860
rect 2440 740 2560 860
rect 2990 740 3110 860
rect 3540 740 3660 860
rect 4090 740 4210 860
rect 4640 740 4760 860
rect 5190 740 5310 860
rect 5740 740 5860 860
rect 6290 740 6410 860
rect 6840 740 6960 860
rect 7390 740 7510 860
rect 7940 740 8060 860
rect 8490 740 8610 860
rect 9040 740 9160 860
rect 9590 740 9710 860
rect 10140 740 10260 860
rect 10690 740 10810 860
rect 11240 740 11360 860
rect 11790 740 11910 860
rect 12340 740 12460 860
rect 12890 740 13010 860
rect 13440 740 13560 860
rect -310 190 -190 310
rect 240 190 360 310
rect 790 190 910 310
rect 1340 190 1460 310
rect 1890 190 2010 310
rect 2440 190 2560 310
rect 2990 190 3110 310
rect 3540 190 3660 310
rect 4090 190 4210 310
rect 4640 190 4760 310
rect 5190 190 5310 310
rect 5740 190 5860 310
rect 6290 190 6410 310
rect 6840 190 6960 310
rect 7390 190 7510 310
rect 7940 190 8060 310
rect 8490 190 8610 310
rect 9040 190 9160 310
rect 9590 190 9710 310
rect 10140 190 10260 310
rect 10690 190 10810 310
rect 11240 190 11360 310
rect 11790 190 11910 310
rect 12340 190 12460 310
rect 12890 190 13010 310
rect 13440 190 13560 310
rect -310 -360 -190 -240
rect 240 -360 360 -240
rect 790 -360 910 -240
rect 1340 -360 1460 -240
rect 1890 -360 2010 -240
rect 2440 -360 2560 -240
rect 2990 -360 3110 -240
rect 3540 -360 3660 -240
rect 4090 -360 4210 -240
rect 4640 -360 4760 -240
rect 5190 -360 5310 -240
rect 5740 -360 5860 -240
rect 6290 -360 6410 -240
rect 6840 -360 6960 -240
rect 7390 -360 7510 -240
rect 7940 -360 8060 -240
rect 8490 -360 8610 -240
rect 9040 -360 9160 -240
rect 9590 -360 9710 -240
rect 10140 -360 10260 -240
rect 10690 -360 10810 -240
rect 11240 -360 11360 -240
rect 11790 -360 11910 -240
rect 12340 -360 12460 -240
rect 12890 -360 13010 -240
rect 13440 -360 13560 -240
<< metal5 >>
rect -2525 14725 13775 15725
rect -2525 13803 -1525 14725
rect -603 13803 -292 14725
rect -2525 13510 -292 13803
tri -292 13510 -154 13648 sw
rect -53 13647 258 14225
tri -53 13510 84 13647 ne
rect 84 13546 258 13647
tri 258 13546 360 13648 sw
rect 497 13647 808 14725
tri 497 13546 598 13647 ne
rect 598 13546 808 13647
tri 808 13546 910 13648 sw
rect 1047 13647 1358 14225
tri 1047 13546 1148 13647 ne
rect 1148 13546 1358 13647
tri 1358 13546 1460 13648 sw
rect 1597 13647 1908 14725
tri 1597 13546 1698 13647 ne
rect 1698 13546 1908 13647
tri 1908 13546 2010 13648 sw
rect 2147 13647 2458 14225
tri 2147 13546 2248 13647 ne
rect 2248 13546 2458 13647
tri 2458 13546 2560 13648 sw
rect 2697 13647 3008 14725
tri 2697 13546 2798 13647 ne
rect 2798 13546 3008 13647
tri 3008 13546 3110 13648 sw
rect 3247 13647 3558 14225
tri 3247 13546 3348 13647 ne
rect 3348 13546 3558 13647
tri 3558 13546 3660 13648 sw
rect 3797 13647 4108 14725
tri 3797 13546 3898 13647 ne
rect 3898 13546 4108 13647
tri 4108 13546 4210 13648 sw
rect 4347 13647 4658 14225
tri 4347 13546 4448 13647 ne
rect 4448 13546 4658 13647
tri 4658 13546 4760 13648 sw
rect 4897 13647 5208 14725
tri 4897 13546 4998 13647 ne
rect 4998 13546 5208 13647
tri 5208 13546 5310 13648 sw
rect 5447 13647 5758 14225
tri 5447 13546 5548 13647 ne
rect 5548 13546 5758 13647
tri 5758 13546 5860 13648 sw
rect 5997 13647 6308 14725
tri 5997 13546 6098 13647 ne
rect 6098 13546 6308 13647
tri 6308 13546 6410 13648 sw
rect 6547 13647 6858 14225
tri 6547 13546 6648 13647 ne
rect 6648 13546 6858 13647
tri 6858 13546 6960 13648 sw
rect 7097 13647 7408 14725
tri 7097 13546 7198 13647 ne
rect 7198 13546 7408 13647
tri 7408 13546 7510 13648 sw
rect 7647 13647 7958 14225
tri 7647 13546 7748 13647 ne
rect 7748 13546 7958 13647
tri 7958 13546 8060 13648 sw
rect 8197 13647 8508 14725
tri 8197 13546 8298 13647 ne
rect 8298 13546 8508 13647
tri 8508 13546 8610 13648 sw
rect 8747 13647 9058 14225
tri 8747 13546 8848 13647 ne
rect 8848 13546 9058 13647
tri 9058 13546 9160 13648 sw
rect 9297 13647 9608 14725
tri 9297 13546 9398 13647 ne
rect 9398 13546 9608 13647
tri 9608 13546 9710 13648 sw
rect 9847 13647 10158 14225
tri 9847 13546 9948 13647 ne
rect 9948 13546 10158 13647
tri 10158 13546 10260 13648 sw
rect 10397 13647 10708 14725
tri 10397 13546 10498 13647 ne
rect 10498 13546 10708 13647
tri 10708 13546 10810 13648 sw
rect 10947 13647 11258 14225
tri 10947 13546 11048 13647 ne
rect 11048 13546 11258 13647
tri 11258 13546 11360 13648 sw
rect 11497 13647 11808 14725
tri 11497 13546 11598 13647 ne
rect 11598 13546 11808 13647
tri 11808 13546 11910 13648 sw
rect 12047 13647 12358 14225
tri 12047 13546 12148 13647 ne
rect 12148 13546 12358 13647
tri 12358 13546 12460 13648 sw
rect 12597 13647 12908 14725
tri 12597 13546 12698 13647 ne
rect 12698 13546 12908 13647
tri 12908 13546 13010 13648 sw
rect 13147 13647 13458 14225
tri 13147 13546 13248 13647 ne
rect 13248 13546 13458 13647
rect 84 13510 360 13546
rect -2525 13492 -310 13510
rect -2525 12703 -1525 13492
tri -448 13356 -312 13492 ne
rect -312 13390 -310 13492
rect -190 13390 -154 13510
rect -312 13356 -154 13390
tri -154 13356 0 13510 sw
tri 84 13356 238 13510 ne
rect 238 13390 240 13510
rect 238 13356 360 13390
tri 360 13356 550 13546 sw
tri 598 13356 788 13546 ne
rect 788 13510 910 13546
rect 788 13390 790 13510
rect 788 13356 910 13390
tri 910 13356 1100 13546 sw
tri 1148 13356 1338 13546 ne
rect 1338 13510 1460 13546
rect 1338 13390 1340 13510
rect 1338 13356 1460 13390
tri 1460 13356 1650 13546 sw
tri 1698 13356 1888 13546 ne
rect 1888 13510 2010 13546
rect 1888 13390 1890 13510
rect 1888 13356 2010 13390
tri 2010 13356 2200 13546 sw
tri 2248 13356 2438 13546 ne
rect 2438 13510 2560 13546
rect 2438 13390 2440 13510
rect 2438 13356 2560 13390
tri 2560 13356 2750 13546 sw
tri 2798 13356 2988 13546 ne
rect 2988 13510 3110 13546
rect 2988 13390 2990 13510
rect 2988 13356 3110 13390
tri 3110 13356 3300 13546 sw
tri 3348 13356 3538 13546 ne
rect 3538 13510 3660 13546
rect 3538 13390 3540 13510
rect 3538 13356 3660 13390
tri 3660 13356 3850 13546 sw
tri 3898 13356 4088 13546 ne
rect 4088 13510 4210 13546
rect 4088 13390 4090 13510
rect 4088 13356 4210 13390
tri 4210 13356 4400 13546 sw
tri 4448 13356 4638 13546 ne
rect 4638 13510 4760 13546
rect 4638 13390 4640 13510
rect 4638 13356 4760 13390
tri 4760 13356 4950 13546 sw
tri 4998 13356 5188 13546 ne
rect 5188 13510 5310 13546
rect 5188 13390 5190 13510
rect 5188 13356 5310 13390
tri 5310 13356 5500 13546 sw
tri 5548 13356 5738 13546 ne
rect 5738 13510 5860 13546
rect 5738 13390 5740 13510
rect 5738 13356 5860 13390
tri 5860 13356 6050 13546 sw
tri 6098 13356 6288 13546 ne
rect 6288 13510 6410 13546
rect 6288 13390 6290 13510
rect 6288 13356 6410 13390
tri 6410 13356 6600 13546 sw
tri 6648 13356 6838 13546 ne
rect 6838 13510 6960 13546
rect 6838 13390 6840 13510
rect 6838 13356 6960 13390
tri 6960 13356 7150 13546 sw
tri 7198 13356 7388 13546 ne
rect 7388 13510 7510 13546
rect 7388 13390 7390 13510
rect 7388 13356 7510 13390
tri 7510 13356 7700 13546 sw
tri 7748 13356 7938 13546 ne
rect 7938 13510 8060 13546
rect 7938 13390 7940 13510
rect 7938 13356 8060 13390
tri 8060 13356 8250 13546 sw
tri 8298 13356 8488 13546 ne
rect 8488 13510 8610 13546
rect 8488 13390 8490 13510
rect 8488 13356 8610 13390
tri 8610 13356 8800 13546 sw
tri 8848 13356 9038 13546 ne
rect 9038 13510 9160 13546
rect 9038 13390 9040 13510
rect 9038 13356 9160 13390
tri 9160 13356 9350 13546 sw
tri 9398 13356 9588 13546 ne
rect 9588 13510 9710 13546
rect 9588 13390 9590 13510
rect 9588 13356 9710 13390
tri 9710 13356 9900 13546 sw
tri 9948 13356 10138 13546 ne
rect 10138 13510 10260 13546
rect 10138 13390 10140 13510
rect 10138 13356 10260 13390
tri 10260 13356 10450 13546 sw
tri 10498 13356 10688 13546 ne
rect 10688 13510 10810 13546
rect 10688 13390 10690 13510
rect 10688 13356 10810 13390
tri 10810 13356 11000 13546 sw
tri 11048 13356 11238 13546 ne
rect 11238 13510 11360 13546
rect 11238 13390 11240 13510
rect 11238 13356 11360 13390
tri 11360 13356 11550 13546 sw
tri 11598 13356 11788 13546 ne
rect 11788 13510 11910 13546
rect 11788 13390 11790 13510
rect 11788 13356 11910 13390
tri 11910 13356 12100 13546 sw
tri 12148 13356 12338 13546 ne
rect 12338 13510 12460 13546
rect 12338 13390 12340 13510
rect 12338 13356 12460 13390
tri 12460 13356 12650 13546 sw
tri 12698 13356 12888 13546 ne
rect 12888 13510 13010 13546
rect 12888 13390 12890 13510
rect 12888 13356 13010 13390
tri 13010 13356 13200 13546 sw
tri 13248 13356 13438 13546 ne
rect 13438 13510 13458 13546
tri 13458 13510 13596 13648 sw
rect 13438 13390 13440 13510
rect 13560 13408 13596 13510
tri 13596 13408 13698 13510 sw
rect 14775 13408 15775 13725
rect 13560 13390 15775 13408
rect 13438 13356 15775 13390
rect -1025 13200 -447 13253
tri -447 13200 -394 13253 sw
tri -312 13200 -156 13356 ne
rect -156 13200 0 13356
tri 0 13200 156 13356 sw
tri 238 13200 394 13356 ne
rect 394 13200 550 13356
tri 550 13200 706 13356 sw
tri 788 13200 944 13356 ne
rect 944 13200 1100 13356
tri 1100 13200 1256 13356 sw
tri 1338 13200 1494 13356 ne
rect 1494 13200 1650 13356
tri 1650 13200 1806 13356 sw
tri 1888 13200 2044 13356 ne
rect 2044 13200 2200 13356
tri 2200 13200 2356 13356 sw
tri 2438 13200 2594 13356 ne
rect 2594 13200 2750 13356
tri 2750 13200 2906 13356 sw
tri 2988 13200 3144 13356 ne
rect 3144 13200 3300 13356
tri 3300 13200 3456 13356 sw
tri 3538 13200 3694 13356 ne
rect 3694 13200 3850 13356
tri 3850 13200 4006 13356 sw
tri 4088 13200 4244 13356 ne
rect 4244 13200 4400 13356
tri 4400 13200 4556 13356 sw
tri 4638 13200 4794 13356 ne
rect 4794 13200 4950 13356
tri 4950 13200 5106 13356 sw
tri 5188 13200 5344 13356 ne
rect 5344 13200 5500 13356
tri 5500 13200 5656 13356 sw
tri 5738 13200 5894 13356 ne
rect 5894 13200 6050 13356
tri 6050 13200 6206 13356 sw
tri 6288 13200 6444 13356 ne
rect 6444 13200 6600 13356
tri 6600 13200 6756 13356 sw
tri 6838 13200 6994 13356 ne
rect 6994 13200 7150 13356
tri 7150 13200 7306 13356 sw
tri 7388 13200 7544 13356 ne
rect 7544 13200 7700 13356
tri 7700 13200 7856 13356 sw
tri 7938 13200 8094 13356 ne
rect 8094 13200 8250 13356
tri 8250 13200 8406 13356 sw
tri 8488 13200 8644 13356 ne
rect 8644 13200 8800 13356
tri 8800 13200 8956 13356 sw
tri 9038 13200 9194 13356 ne
rect 9194 13200 9350 13356
tri 9350 13200 9506 13356 sw
tri 9588 13200 9744 13356 ne
rect 9744 13200 9900 13356
tri 9900 13200 10056 13356 sw
tri 10138 13200 10294 13356 ne
rect 10294 13200 10450 13356
tri 10450 13200 10606 13356 sw
tri 10688 13200 10844 13356 ne
rect 10844 13200 11000 13356
tri 11000 13200 11156 13356 sw
tri 11238 13200 11394 13356 ne
rect 11394 13200 11550 13356
tri 11550 13200 11706 13356 sw
tri 11788 13200 11944 13356 ne
rect 11944 13200 12100 13356
tri 12100 13200 12256 13356 sw
tri 12338 13200 12494 13356 ne
rect 12494 13200 12650 13356
tri 12650 13200 12806 13356 sw
tri 12888 13200 13044 13356 ne
rect 13044 13200 13200 13356
tri 13200 13200 13356 13356 sw
tri 13438 13200 13594 13356 ne
rect 13594 13200 15775 13356
rect -1025 13097 -394 13200
tri -394 13097 -291 13200 sw
tri -156 13097 -53 13200 ne
rect -53 13097 156 13200
tri 156 13097 259 13200 sw
tri 394 13097 497 13200 ne
rect 497 13097 706 13200
tri 706 13097 809 13200 sw
tri 944 13097 1047 13200 ne
rect 1047 13097 1256 13200
tri 1256 13097 1359 13200 sw
tri 1494 13097 1597 13200 ne
rect 1597 13097 1806 13200
tri 1806 13097 1909 13200 sw
tri 2044 13097 2147 13200 ne
rect 2147 13097 2356 13200
tri 2356 13097 2459 13200 sw
tri 2594 13097 2697 13200 ne
rect 2697 13097 2906 13200
tri 2906 13097 3009 13200 sw
tri 3144 13097 3247 13200 ne
rect 3247 13097 3456 13200
tri 3456 13097 3559 13200 sw
tri 3694 13097 3797 13200 ne
rect 3797 13097 4006 13200
tri 4006 13097 4109 13200 sw
tri 4244 13097 4347 13200 ne
rect 4347 13097 4556 13200
tri 4556 13097 4659 13200 sw
tri 4794 13097 4897 13200 ne
rect 4897 13097 5106 13200
tri 5106 13097 5209 13200 sw
tri 5344 13097 5447 13200 ne
rect 5447 13097 5656 13200
tri 5656 13097 5759 13200 sw
tri 5894 13097 5997 13200 ne
rect 5997 13097 6206 13200
tri 6206 13097 6309 13200 sw
tri 6444 13097 6547 13200 ne
rect 6547 13097 6756 13200
tri 6756 13097 6859 13200 sw
tri 6994 13097 7097 13200 ne
rect 7097 13097 7306 13200
tri 7306 13097 7409 13200 sw
tri 7544 13097 7647 13200 ne
rect 7647 13097 7856 13200
tri 7856 13097 7959 13200 sw
tri 8094 13097 8197 13200 ne
rect 8197 13097 8406 13200
tri 8406 13097 8509 13200 sw
tri 8644 13097 8747 13200 ne
rect 8747 13097 8956 13200
tri 8956 13097 9059 13200 sw
tri 9194 13097 9297 13200 ne
rect 9297 13097 9506 13200
tri 9506 13097 9609 13200 sw
tri 9744 13097 9847 13200 ne
rect 9847 13097 10056 13200
tri 10056 13097 10159 13200 sw
tri 10294 13097 10397 13200 ne
rect 10397 13097 10606 13200
tri 10606 13097 10709 13200 sw
tri 10844 13097 10947 13200 ne
rect 10947 13097 11156 13200
tri 11156 13097 11259 13200 sw
tri 11394 13097 11497 13200 ne
rect 11497 13097 11706 13200
tri 11706 13097 11809 13200 sw
tri 11944 13097 12047 13200 ne
rect 12047 13097 12256 13200
tri 12256 13097 12359 13200 sw
tri 12494 13097 12597 13200 ne
rect 12597 13097 12806 13200
tri 12806 13097 12909 13200 sw
tri 13044 13097 13147 13200 ne
rect 13147 13097 13356 13200
tri 13356 13097 13459 13200 sw
tri 13594 13097 13697 13200 ne
rect 13697 13097 15775 13200
rect -1025 12960 -291 13097
tri -291 12960 -154 13097 sw
tri -53 12960 84 13097 ne
rect 84 12960 259 13097
tri 259 12960 396 13097 sw
tri 497 12960 634 13097 ne
rect 634 12960 809 13097
tri 809 12960 946 13097 sw
tri 1047 12960 1184 13097 ne
rect 1184 12960 1359 13097
tri 1359 12960 1496 13097 sw
tri 1597 12960 1734 13097 ne
rect 1734 12960 1909 13097
tri 1909 12960 2046 13097 sw
tri 2147 12960 2284 13097 ne
rect 2284 12960 2459 13097
tri 2459 12960 2596 13097 sw
tri 2697 12960 2834 13097 ne
rect 2834 12960 3009 13097
tri 3009 12960 3146 13097 sw
tri 3247 12960 3384 13097 ne
rect 3384 12960 3559 13097
tri 3559 12960 3696 13097 sw
tri 3797 12960 3934 13097 ne
rect 3934 12960 4109 13097
tri 4109 12960 4246 13097 sw
tri 4347 12960 4484 13097 ne
rect 4484 12960 4659 13097
tri 4659 12960 4796 13097 sw
tri 4897 12960 5034 13097 ne
rect 5034 12960 5209 13097
tri 5209 12960 5346 13097 sw
tri 5447 12960 5584 13097 ne
rect 5584 12960 5759 13097
tri 5759 12960 5896 13097 sw
tri 5997 12960 6134 13097 ne
rect 6134 12960 6309 13097
tri 6309 12960 6446 13097 sw
tri 6547 12960 6684 13097 ne
rect 6684 12960 6859 13097
tri 6859 12960 6996 13097 sw
tri 7097 12960 7234 13097 ne
rect 7234 12960 7409 13097
tri 7409 12960 7546 13097 sw
tri 7647 12960 7784 13097 ne
rect 7784 12960 7959 13097
tri 7959 12960 8096 13097 sw
tri 8197 12960 8334 13097 ne
rect 8334 12960 8509 13097
tri 8509 12960 8646 13097 sw
tri 8747 12960 8884 13097 ne
rect 8884 12960 9059 13097
tri 9059 12960 9196 13097 sw
tri 9297 12960 9434 13097 ne
rect 9434 12960 9609 13097
tri 9609 12960 9746 13097 sw
tri 9847 12960 9984 13097 ne
rect 9984 12960 10159 13097
tri 10159 12960 10296 13097 sw
tri 10397 12960 10534 13097 ne
rect 10534 12960 10709 13097
tri 10709 12960 10846 13097 sw
tri 10947 12960 11084 13097 ne
rect 11084 12960 11259 13097
tri 11259 12960 11396 13097 sw
tri 11497 12960 11634 13097 ne
rect 11634 12960 11809 13097
tri 11809 12960 11946 13097 sw
tri 12047 12960 12184 13097 ne
rect 12184 12960 12359 13097
tri 12359 12960 12496 13097 sw
tri 12597 12960 12734 13097 ne
rect 12734 12960 12909 13097
tri 12909 12960 13046 13097 sw
tri 13147 12960 13284 13097 ne
rect 13284 12960 13459 13097
tri 13459 12960 13596 13097 sw
rect -1025 12942 -310 12960
tri -448 12840 -346 12942 ne
rect -346 12840 -310 12942
rect -190 12840 -154 12960
rect -2525 12650 -447 12703
tri -447 12650 -394 12703 sw
tri -346 12650 -156 12840 ne
rect -156 12806 -154 12840
tri -154 12806 0 12960 sw
tri 84 12806 238 12960 ne
rect 238 12840 240 12960
rect 360 12840 396 12960
rect 238 12806 396 12840
tri 396 12806 550 12960 sw
tri 634 12806 788 12960 ne
rect 788 12840 790 12960
rect 910 12840 946 12960
rect 788 12806 946 12840
tri 946 12806 1100 12960 sw
tri 1184 12806 1338 12960 ne
rect 1338 12840 1340 12960
rect 1460 12840 1496 12960
rect 1338 12806 1496 12840
tri 1496 12806 1650 12960 sw
tri 1734 12806 1888 12960 ne
rect 1888 12840 1890 12960
rect 2010 12840 2046 12960
rect 1888 12806 2046 12840
tri 2046 12806 2200 12960 sw
tri 2284 12806 2438 12960 ne
rect 2438 12840 2440 12960
rect 2560 12840 2596 12960
rect 2438 12806 2596 12840
tri 2596 12806 2750 12960 sw
tri 2834 12806 2988 12960 ne
rect 2988 12840 2990 12960
rect 3110 12840 3146 12960
rect 2988 12806 3146 12840
tri 3146 12806 3300 12960 sw
tri 3384 12806 3538 12960 ne
rect 3538 12840 3540 12960
rect 3660 12840 3696 12960
rect 3538 12806 3696 12840
tri 3696 12806 3850 12960 sw
tri 3934 12806 4088 12960 ne
rect 4088 12840 4090 12960
rect 4210 12840 4246 12960
rect 4088 12806 4246 12840
tri 4246 12806 4400 12960 sw
tri 4484 12806 4638 12960 ne
rect 4638 12840 4640 12960
rect 4760 12840 4796 12960
rect 4638 12806 4796 12840
tri 4796 12806 4950 12960 sw
tri 5034 12806 5188 12960 ne
rect 5188 12840 5190 12960
rect 5310 12840 5346 12960
rect 5188 12806 5346 12840
tri 5346 12806 5500 12960 sw
tri 5584 12806 5738 12960 ne
rect 5738 12840 5740 12960
rect 5860 12840 5896 12960
rect 5738 12806 5896 12840
tri 5896 12806 6050 12960 sw
tri 6134 12806 6288 12960 ne
rect 6288 12840 6290 12960
rect 6410 12840 6446 12960
rect 6288 12806 6446 12840
tri 6446 12806 6600 12960 sw
tri 6684 12806 6838 12960 ne
rect 6838 12840 6840 12960
rect 6960 12840 6996 12960
rect 6838 12806 6996 12840
tri 6996 12806 7150 12960 sw
tri 7234 12806 7388 12960 ne
rect 7388 12840 7390 12960
rect 7510 12840 7546 12960
rect 7388 12806 7546 12840
tri 7546 12806 7700 12960 sw
tri 7784 12806 7938 12960 ne
rect 7938 12840 7940 12960
rect 8060 12840 8096 12960
rect 7938 12806 8096 12840
tri 8096 12806 8250 12960 sw
tri 8334 12806 8488 12960 ne
rect 8488 12840 8490 12960
rect 8610 12840 8646 12960
rect 8488 12806 8646 12840
tri 8646 12806 8800 12960 sw
tri 8884 12806 9038 12960 ne
rect 9038 12840 9040 12960
rect 9160 12840 9196 12960
rect 9038 12806 9196 12840
tri 9196 12806 9350 12960 sw
tri 9434 12806 9588 12960 ne
rect 9588 12840 9590 12960
rect 9710 12840 9746 12960
rect 9588 12806 9746 12840
tri 9746 12806 9900 12960 sw
tri 9984 12806 10138 12960 ne
rect 10138 12840 10140 12960
rect 10260 12840 10296 12960
rect 10138 12806 10296 12840
tri 10296 12806 10450 12960 sw
tri 10534 12806 10688 12960 ne
rect 10688 12840 10690 12960
rect 10810 12840 10846 12960
rect 10688 12806 10846 12840
tri 10846 12806 11000 12960 sw
tri 11084 12806 11238 12960 ne
rect 11238 12840 11240 12960
rect 11360 12840 11396 12960
rect 11238 12806 11396 12840
tri 11396 12806 11550 12960 sw
tri 11634 12806 11788 12960 ne
rect 11788 12840 11790 12960
rect 11910 12840 11946 12960
rect 11788 12806 11946 12840
tri 11946 12806 12100 12960 sw
tri 12184 12806 12338 12960 ne
rect 12338 12840 12340 12960
rect 12460 12840 12496 12960
rect 12338 12806 12496 12840
tri 12496 12806 12650 12960 sw
tri 12734 12806 12888 12960 ne
rect 12888 12840 12890 12960
rect 13010 12840 13046 12960
rect 12888 12806 13046 12840
tri 13046 12806 13200 12960 sw
tri 13284 12806 13438 12960 ne
rect 13438 12840 13440 12960
rect 13560 12858 13596 12960
tri 13596 12858 13698 12960 sw
rect 13560 12840 14275 12858
rect 13438 12806 14275 12840
rect -156 12650 0 12806
tri 0 12650 156 12806 sw
tri 238 12650 394 12806 ne
rect 394 12650 550 12806
tri 550 12650 706 12806 sw
tri 788 12650 944 12806 ne
rect 944 12650 1100 12806
tri 1100 12650 1256 12806 sw
tri 1338 12650 1494 12806 ne
rect 1494 12650 1650 12806
tri 1650 12650 1806 12806 sw
tri 1888 12650 2044 12806 ne
rect 2044 12650 2200 12806
tri 2200 12650 2356 12806 sw
tri 2438 12650 2594 12806 ne
rect 2594 12650 2750 12806
tri 2750 12650 2906 12806 sw
tri 2988 12650 3144 12806 ne
rect 3144 12650 3300 12806
tri 3300 12650 3456 12806 sw
tri 3538 12650 3694 12806 ne
rect 3694 12650 3850 12806
tri 3850 12650 4006 12806 sw
tri 4088 12650 4244 12806 ne
rect 4244 12650 4400 12806
tri 4400 12650 4556 12806 sw
tri 4638 12650 4794 12806 ne
rect 4794 12650 4950 12806
tri 4950 12650 5106 12806 sw
tri 5188 12650 5344 12806 ne
rect 5344 12650 5500 12806
tri 5500 12650 5656 12806 sw
tri 5738 12650 5894 12806 ne
rect 5894 12650 6050 12806
tri 6050 12650 6206 12806 sw
tri 6288 12650 6444 12806 ne
rect 6444 12650 6600 12806
tri 6600 12650 6756 12806 sw
tri 6838 12650 6994 12806 ne
rect 6994 12650 7150 12806
tri 7150 12650 7306 12806 sw
tri 7388 12650 7544 12806 ne
rect 7544 12650 7700 12806
tri 7700 12650 7856 12806 sw
tri 7938 12650 8094 12806 ne
rect 8094 12650 8250 12806
tri 8250 12650 8406 12806 sw
tri 8488 12650 8644 12806 ne
rect 8644 12650 8800 12806
tri 8800 12650 8956 12806 sw
tri 9038 12650 9194 12806 ne
rect 9194 12650 9350 12806
tri 9350 12650 9506 12806 sw
tri 9588 12650 9744 12806 ne
rect 9744 12650 9900 12806
tri 9900 12650 10056 12806 sw
tri 10138 12650 10294 12806 ne
rect 10294 12650 10450 12806
tri 10450 12650 10606 12806 sw
tri 10688 12650 10844 12806 ne
rect 10844 12650 11000 12806
tri 11000 12650 11156 12806 sw
tri 11238 12650 11394 12806 ne
rect 11394 12650 11550 12806
tri 11550 12650 11706 12806 sw
tri 11788 12650 11944 12806 ne
rect 11944 12650 12100 12806
tri 12100 12650 12256 12806 sw
tri 12338 12650 12494 12806 ne
rect 12494 12650 12650 12806
tri 12650 12650 12806 12806 sw
tri 12888 12650 13044 12806 ne
rect 13044 12650 13200 12806
tri 13200 12650 13356 12806 sw
tri 13438 12650 13594 12806 ne
rect 13594 12650 14275 12806
rect -2525 12547 -394 12650
tri -394 12547 -291 12650 sw
tri -156 12547 -53 12650 ne
rect -53 12547 156 12650
tri 156 12547 259 12650 sw
tri 394 12547 497 12650 ne
rect 497 12547 706 12650
tri 706 12547 809 12650 sw
tri 944 12547 1047 12650 ne
rect 1047 12547 1256 12650
tri 1256 12547 1359 12650 sw
tri 1494 12547 1597 12650 ne
rect 1597 12547 1806 12650
tri 1806 12547 1909 12650 sw
tri 2044 12547 2147 12650 ne
rect 2147 12547 2356 12650
tri 2356 12547 2459 12650 sw
tri 2594 12547 2697 12650 ne
rect 2697 12547 2906 12650
tri 2906 12547 3009 12650 sw
tri 3144 12547 3247 12650 ne
rect 3247 12547 3456 12650
tri 3456 12547 3559 12650 sw
tri 3694 12547 3797 12650 ne
rect 3797 12547 4006 12650
tri 4006 12547 4109 12650 sw
tri 4244 12547 4347 12650 ne
rect 4347 12547 4556 12650
tri 4556 12547 4659 12650 sw
tri 4794 12547 4897 12650 ne
rect 4897 12547 5106 12650
tri 5106 12547 5209 12650 sw
tri 5344 12547 5447 12650 ne
rect 5447 12547 5656 12650
tri 5656 12547 5759 12650 sw
tri 5894 12547 5997 12650 ne
rect 5997 12547 6206 12650
tri 6206 12547 6309 12650 sw
tri 6444 12547 6547 12650 ne
rect 6547 12547 6756 12650
tri 6756 12547 6859 12650 sw
tri 6994 12547 7097 12650 ne
rect 7097 12547 7306 12650
tri 7306 12547 7409 12650 sw
tri 7544 12547 7647 12650 ne
rect 7647 12547 7856 12650
tri 7856 12547 7959 12650 sw
tri 8094 12547 8197 12650 ne
rect 8197 12547 8406 12650
tri 8406 12547 8509 12650 sw
tri 8644 12547 8747 12650 ne
rect 8747 12547 8956 12650
tri 8956 12547 9059 12650 sw
tri 9194 12547 9297 12650 ne
rect 9297 12547 9506 12650
tri 9506 12547 9609 12650 sw
tri 9744 12547 9847 12650 ne
rect 9847 12547 10056 12650
tri 10056 12547 10159 12650 sw
tri 10294 12547 10397 12650 ne
rect 10397 12547 10606 12650
tri 10606 12547 10709 12650 sw
tri 10844 12547 10947 12650 ne
rect 10947 12547 11156 12650
tri 11156 12547 11259 12650 sw
tri 11394 12547 11497 12650 ne
rect 11497 12547 11706 12650
tri 11706 12547 11809 12650 sw
tri 11944 12547 12047 12650 ne
rect 12047 12547 12256 12650
tri 12256 12547 12359 12650 sw
tri 12494 12547 12597 12650 ne
rect 12597 12547 12806 12650
tri 12806 12547 12909 12650 sw
tri 13044 12547 13147 12650 ne
rect 13147 12547 13356 12650
tri 13356 12547 13459 12650 sw
tri 13594 12547 13697 12650 ne
rect 13697 12547 14275 12650
rect -2525 12410 -291 12547
tri -291 12410 -154 12547 sw
tri -53 12410 84 12547 ne
rect 84 12410 259 12547
tri 259 12410 396 12547 sw
tri 497 12410 634 12547 ne
rect 634 12410 809 12547
tri 809 12410 946 12547 sw
tri 1047 12410 1184 12547 ne
rect 1184 12410 1359 12547
tri 1359 12410 1496 12547 sw
tri 1597 12410 1734 12547 ne
rect 1734 12410 1909 12547
tri 1909 12410 2046 12547 sw
tri 2147 12410 2284 12547 ne
rect 2284 12410 2459 12547
tri 2459 12410 2596 12547 sw
tri 2697 12410 2834 12547 ne
rect 2834 12410 3009 12547
tri 3009 12410 3146 12547 sw
tri 3247 12410 3384 12547 ne
rect 3384 12410 3559 12547
tri 3559 12410 3696 12547 sw
tri 3797 12410 3934 12547 ne
rect 3934 12410 4109 12547
tri 4109 12410 4246 12547 sw
tri 4347 12410 4484 12547 ne
rect 4484 12410 4659 12547
tri 4659 12410 4796 12547 sw
tri 4897 12410 5034 12547 ne
rect 5034 12410 5209 12547
tri 5209 12410 5346 12547 sw
tri 5447 12410 5584 12547 ne
rect 5584 12410 5759 12547
tri 5759 12410 5896 12547 sw
tri 5997 12410 6134 12547 ne
rect 6134 12410 6309 12547
tri 6309 12410 6446 12547 sw
tri 6547 12410 6684 12547 ne
rect 6684 12410 6859 12547
tri 6859 12410 6996 12547 sw
tri 7097 12410 7234 12547 ne
rect 7234 12410 7409 12547
tri 7409 12410 7546 12547 sw
tri 7647 12410 7784 12547 ne
rect 7784 12410 7959 12547
tri 7959 12410 8096 12547 sw
tri 8197 12410 8334 12547 ne
rect 8334 12410 8509 12547
tri 8509 12410 8646 12547 sw
tri 8747 12410 8884 12547 ne
rect 8884 12410 9059 12547
tri 9059 12410 9196 12547 sw
tri 9297 12410 9434 12547 ne
rect 9434 12410 9609 12547
tri 9609 12410 9746 12547 sw
tri 9847 12410 9984 12547 ne
rect 9984 12410 10159 12547
tri 10159 12410 10296 12547 sw
tri 10397 12410 10534 12547 ne
rect 10534 12410 10709 12547
tri 10709 12410 10846 12547 sw
tri 10947 12410 11084 12547 ne
rect 11084 12410 11259 12547
tri 11259 12410 11396 12547 sw
tri 11497 12410 11634 12547 ne
rect 11634 12410 11809 12547
tri 11809 12410 11946 12547 sw
tri 12047 12410 12184 12547 ne
rect 12184 12410 12359 12547
tri 12359 12410 12496 12547 sw
tri 12597 12410 12734 12547 ne
rect 12734 12410 12909 12547
tri 12909 12410 13046 12547 sw
tri 13147 12410 13284 12547 ne
rect 13284 12410 13459 12547
tri 13459 12410 13596 12547 sw
rect -2525 12392 -310 12410
rect -2525 11603 -1525 12392
tri -448 12290 -346 12392 ne
rect -346 12290 -310 12392
rect -190 12290 -154 12410
rect -1025 12100 -447 12153
tri -447 12100 -394 12153 sw
tri -346 12100 -156 12290 ne
rect -156 12256 -154 12290
tri -154 12256 0 12410 sw
tri 84 12256 238 12410 ne
rect 238 12290 240 12410
rect 360 12290 396 12410
rect 238 12256 396 12290
tri 396 12256 550 12410 sw
tri 634 12256 788 12410 ne
rect 788 12290 790 12410
rect 910 12290 946 12410
rect 788 12256 946 12290
tri 946 12256 1100 12410 sw
tri 1184 12256 1338 12410 ne
rect 1338 12290 1340 12410
rect 1460 12290 1496 12410
rect 1338 12256 1496 12290
tri 1496 12256 1650 12410 sw
tri 1734 12256 1888 12410 ne
rect 1888 12290 1890 12410
rect 2010 12290 2046 12410
rect 1888 12256 2046 12290
tri 2046 12256 2200 12410 sw
tri 2284 12256 2438 12410 ne
rect 2438 12290 2440 12410
rect 2560 12290 2596 12410
rect 2438 12256 2596 12290
tri 2596 12256 2750 12410 sw
tri 2834 12256 2988 12410 ne
rect 2988 12290 2990 12410
rect 3110 12290 3146 12410
rect 2988 12256 3146 12290
tri 3146 12256 3300 12410 sw
tri 3384 12256 3538 12410 ne
rect 3538 12290 3540 12410
rect 3660 12290 3696 12410
rect 3538 12256 3696 12290
tri 3696 12256 3850 12410 sw
tri 3934 12256 4088 12410 ne
rect 4088 12290 4090 12410
rect 4210 12290 4246 12410
rect 4088 12256 4246 12290
tri 4246 12256 4400 12410 sw
tri 4484 12256 4638 12410 ne
rect 4638 12290 4640 12410
rect 4760 12290 4796 12410
rect 4638 12256 4796 12290
tri 4796 12256 4950 12410 sw
tri 5034 12256 5188 12410 ne
rect 5188 12290 5190 12410
rect 5310 12290 5346 12410
rect 5188 12256 5346 12290
tri 5346 12256 5500 12410 sw
tri 5584 12256 5738 12410 ne
rect 5738 12290 5740 12410
rect 5860 12290 5896 12410
rect 5738 12256 5896 12290
tri 5896 12256 6050 12410 sw
tri 6134 12256 6288 12410 ne
rect 6288 12290 6290 12410
rect 6410 12290 6446 12410
rect 6288 12256 6446 12290
tri 6446 12256 6600 12410 sw
tri 6684 12256 6838 12410 ne
rect 6838 12290 6840 12410
rect 6960 12290 6996 12410
rect 6838 12256 6996 12290
tri 6996 12256 7150 12410 sw
tri 7234 12256 7388 12410 ne
rect 7388 12290 7390 12410
rect 7510 12290 7546 12410
rect 7388 12256 7546 12290
tri 7546 12256 7700 12410 sw
tri 7784 12256 7938 12410 ne
rect 7938 12290 7940 12410
rect 8060 12290 8096 12410
rect 7938 12256 8096 12290
tri 8096 12256 8250 12410 sw
tri 8334 12256 8488 12410 ne
rect 8488 12290 8490 12410
rect 8610 12290 8646 12410
rect 8488 12256 8646 12290
tri 8646 12256 8800 12410 sw
tri 8884 12256 9038 12410 ne
rect 9038 12290 9040 12410
rect 9160 12290 9196 12410
rect 9038 12256 9196 12290
tri 9196 12256 9350 12410 sw
tri 9434 12256 9588 12410 ne
rect 9588 12290 9590 12410
rect 9710 12290 9746 12410
rect 9588 12256 9746 12290
tri 9746 12256 9900 12410 sw
tri 9984 12256 10138 12410 ne
rect 10138 12290 10140 12410
rect 10260 12290 10296 12410
rect 10138 12256 10296 12290
tri 10296 12256 10450 12410 sw
tri 10534 12256 10688 12410 ne
rect 10688 12290 10690 12410
rect 10810 12290 10846 12410
rect 10688 12256 10846 12290
tri 10846 12256 11000 12410 sw
tri 11084 12256 11238 12410 ne
rect 11238 12290 11240 12410
rect 11360 12290 11396 12410
rect 11238 12256 11396 12290
tri 11396 12256 11550 12410 sw
tri 11634 12256 11788 12410 ne
rect 11788 12290 11790 12410
rect 11910 12290 11946 12410
rect 11788 12256 11946 12290
tri 11946 12256 12100 12410 sw
tri 12184 12256 12338 12410 ne
rect 12338 12290 12340 12410
rect 12460 12290 12496 12410
rect 12338 12256 12496 12290
tri 12496 12256 12650 12410 sw
tri 12734 12256 12888 12410 ne
rect 12888 12290 12890 12410
rect 13010 12290 13046 12410
rect 12888 12256 13046 12290
tri 13046 12256 13200 12410 sw
tri 13284 12256 13438 12410 ne
rect 13438 12290 13440 12410
rect 13560 12308 13596 12410
tri 13596 12308 13698 12410 sw
rect 14775 12308 15775 13097
rect 13560 12290 15775 12308
rect 13438 12256 15775 12290
rect -156 12100 0 12256
tri 0 12100 156 12256 sw
tri 238 12100 394 12256 ne
rect 394 12100 550 12256
tri 550 12100 706 12256 sw
tri 788 12100 944 12256 ne
rect 944 12100 1100 12256
tri 1100 12100 1256 12256 sw
tri 1338 12100 1494 12256 ne
rect 1494 12100 1650 12256
tri 1650 12100 1806 12256 sw
tri 1888 12100 2044 12256 ne
rect 2044 12100 2200 12256
tri 2200 12100 2356 12256 sw
tri 2438 12100 2594 12256 ne
rect 2594 12100 2750 12256
tri 2750 12100 2906 12256 sw
tri 2988 12100 3144 12256 ne
rect 3144 12100 3300 12256
tri 3300 12100 3456 12256 sw
tri 3538 12100 3694 12256 ne
rect 3694 12100 3850 12256
tri 3850 12100 4006 12256 sw
tri 4088 12100 4244 12256 ne
rect 4244 12100 4400 12256
tri 4400 12100 4556 12256 sw
tri 4638 12100 4794 12256 ne
rect 4794 12100 4950 12256
tri 4950 12100 5106 12256 sw
tri 5188 12100 5344 12256 ne
rect 5344 12100 5500 12256
tri 5500 12100 5656 12256 sw
tri 5738 12100 5894 12256 ne
rect 5894 12100 6050 12256
tri 6050 12100 6206 12256 sw
tri 6288 12100 6444 12256 ne
rect 6444 12100 6600 12256
tri 6600 12100 6756 12256 sw
tri 6838 12100 6994 12256 ne
rect 6994 12100 7150 12256
tri 7150 12100 7306 12256 sw
tri 7388 12100 7544 12256 ne
rect 7544 12100 7700 12256
tri 7700 12100 7856 12256 sw
tri 7938 12100 8094 12256 ne
rect 8094 12100 8250 12256
tri 8250 12100 8406 12256 sw
tri 8488 12100 8644 12256 ne
rect 8644 12100 8800 12256
tri 8800 12100 8956 12256 sw
tri 9038 12100 9194 12256 ne
rect 9194 12100 9350 12256
tri 9350 12100 9506 12256 sw
tri 9588 12100 9744 12256 ne
rect 9744 12100 9900 12256
tri 9900 12100 10056 12256 sw
tri 10138 12100 10294 12256 ne
rect 10294 12100 10450 12256
tri 10450 12100 10606 12256 sw
tri 10688 12100 10844 12256 ne
rect 10844 12100 11000 12256
tri 11000 12100 11156 12256 sw
tri 11238 12100 11394 12256 ne
rect 11394 12100 11550 12256
tri 11550 12100 11706 12256 sw
tri 11788 12100 11944 12256 ne
rect 11944 12100 12100 12256
tri 12100 12100 12256 12256 sw
tri 12338 12100 12494 12256 ne
rect 12494 12100 12650 12256
tri 12650 12100 12806 12256 sw
tri 12888 12100 13044 12256 ne
rect 13044 12100 13200 12256
tri 13200 12100 13356 12256 sw
tri 13438 12100 13594 12256 ne
rect 13594 12100 15775 12256
rect -1025 11997 -394 12100
tri -394 11997 -291 12100 sw
tri -156 11997 -53 12100 ne
rect -53 11997 156 12100
tri 156 11997 259 12100 sw
tri 394 11997 497 12100 ne
rect 497 11997 706 12100
tri 706 11997 809 12100 sw
tri 944 11997 1047 12100 ne
rect 1047 11997 1256 12100
tri 1256 11997 1359 12100 sw
tri 1494 11997 1597 12100 ne
rect 1597 11997 1806 12100
tri 1806 11997 1909 12100 sw
tri 2044 11997 2147 12100 ne
rect 2147 11997 2356 12100
tri 2356 11997 2459 12100 sw
tri 2594 11997 2697 12100 ne
rect 2697 11997 2906 12100
tri 2906 11997 3009 12100 sw
tri 3144 11997 3247 12100 ne
rect 3247 11997 3456 12100
tri 3456 11997 3559 12100 sw
tri 3694 11997 3797 12100 ne
rect 3797 11997 4006 12100
tri 4006 11997 4109 12100 sw
tri 4244 11997 4347 12100 ne
rect 4347 11997 4556 12100
tri 4556 11997 4659 12100 sw
tri 4794 11997 4897 12100 ne
rect 4897 11997 5106 12100
tri 5106 11997 5209 12100 sw
tri 5344 11997 5447 12100 ne
rect 5447 11997 5656 12100
tri 5656 11997 5759 12100 sw
tri 5894 11997 5997 12100 ne
rect 5997 11997 6206 12100
tri 6206 11997 6309 12100 sw
tri 6444 11997 6547 12100 ne
rect 6547 11997 6756 12100
tri 6756 11997 6859 12100 sw
tri 6994 11997 7097 12100 ne
rect 7097 11997 7306 12100
tri 7306 11997 7409 12100 sw
tri 7544 11997 7647 12100 ne
rect 7647 11997 7856 12100
tri 7856 11997 7959 12100 sw
tri 8094 11997 8197 12100 ne
rect 8197 11997 8406 12100
tri 8406 11997 8509 12100 sw
tri 8644 11997 8747 12100 ne
rect 8747 11997 8956 12100
tri 8956 11997 9059 12100 sw
tri 9194 11997 9297 12100 ne
rect 9297 11997 9506 12100
tri 9506 11997 9609 12100 sw
tri 9744 11997 9847 12100 ne
rect 9847 11997 10056 12100
tri 10056 11997 10159 12100 sw
tri 10294 11997 10397 12100 ne
rect 10397 11997 10606 12100
tri 10606 11997 10709 12100 sw
tri 10844 11997 10947 12100 ne
rect 10947 11997 11156 12100
tri 11156 11997 11259 12100 sw
tri 11394 11997 11497 12100 ne
rect 11497 11997 11706 12100
tri 11706 11997 11809 12100 sw
tri 11944 11997 12047 12100 ne
rect 12047 11997 12256 12100
tri 12256 11997 12359 12100 sw
tri 12494 11997 12597 12100 ne
rect 12597 11997 12806 12100
tri 12806 11997 12909 12100 sw
tri 13044 11997 13147 12100 ne
rect 13147 11997 13356 12100
tri 13356 11997 13459 12100 sw
tri 13594 11997 13697 12100 ne
rect 13697 11997 15775 12100
rect -1025 11860 -291 11997
tri -291 11860 -154 11997 sw
tri -53 11860 84 11997 ne
rect 84 11860 259 11997
tri 259 11860 396 11997 sw
tri 497 11860 634 11997 ne
rect 634 11860 809 11997
tri 809 11860 946 11997 sw
tri 1047 11860 1184 11997 ne
rect 1184 11860 1359 11997
tri 1359 11860 1496 11997 sw
tri 1597 11860 1734 11997 ne
rect 1734 11860 1909 11997
tri 1909 11860 2046 11997 sw
tri 2147 11860 2284 11997 ne
rect 2284 11860 2459 11997
tri 2459 11860 2596 11997 sw
tri 2697 11860 2834 11997 ne
rect 2834 11860 3009 11997
tri 3009 11860 3146 11997 sw
tri 3247 11860 3384 11997 ne
rect 3384 11860 3559 11997
tri 3559 11860 3696 11997 sw
tri 3797 11860 3934 11997 ne
rect 3934 11860 4109 11997
tri 4109 11860 4246 11997 sw
tri 4347 11860 4484 11997 ne
rect 4484 11860 4659 11997
tri 4659 11860 4796 11997 sw
tri 4897 11860 5034 11997 ne
rect 5034 11860 5209 11997
tri 5209 11860 5346 11997 sw
tri 5447 11860 5584 11997 ne
rect 5584 11860 5759 11997
tri 5759 11860 5896 11997 sw
tri 5997 11860 6134 11997 ne
rect 6134 11860 6309 11997
tri 6309 11860 6446 11997 sw
tri 6547 11860 6684 11997 ne
rect 6684 11860 6859 11997
tri 6859 11860 6996 11997 sw
tri 7097 11860 7234 11997 ne
rect 7234 11860 7409 11997
tri 7409 11860 7546 11997 sw
tri 7647 11860 7784 11997 ne
rect 7784 11860 7959 11997
tri 7959 11860 8096 11997 sw
tri 8197 11860 8334 11997 ne
rect 8334 11860 8509 11997
tri 8509 11860 8646 11997 sw
tri 8747 11860 8884 11997 ne
rect 8884 11860 9059 11997
tri 9059 11860 9196 11997 sw
tri 9297 11860 9434 11997 ne
rect 9434 11860 9609 11997
tri 9609 11860 9746 11997 sw
tri 9847 11860 9984 11997 ne
rect 9984 11860 10159 11997
tri 10159 11860 10296 11997 sw
tri 10397 11860 10534 11997 ne
rect 10534 11860 10709 11997
tri 10709 11860 10846 11997 sw
tri 10947 11860 11084 11997 ne
rect 11084 11860 11259 11997
tri 11259 11860 11396 11997 sw
tri 11497 11860 11634 11997 ne
rect 11634 11860 11809 11997
tri 11809 11860 11946 11997 sw
tri 12047 11860 12184 11997 ne
rect 12184 11860 12359 11997
tri 12359 11860 12496 11997 sw
tri 12597 11860 12734 11997 ne
rect 12734 11860 12909 11997
tri 12909 11860 13046 11997 sw
tri 13147 11860 13284 11997 ne
rect 13284 11860 13459 11997
tri 13459 11860 13596 11997 sw
rect -1025 11842 -310 11860
tri -448 11740 -346 11842 ne
rect -346 11740 -310 11842
rect -190 11740 -154 11860
rect -2525 11550 -447 11603
tri -447 11550 -394 11603 sw
tri -346 11550 -156 11740 ne
rect -156 11706 -154 11740
tri -154 11706 0 11860 sw
tri 84 11706 238 11860 ne
rect 238 11740 240 11860
rect 360 11740 396 11860
rect 238 11706 396 11740
tri 396 11706 550 11860 sw
tri 634 11706 788 11860 ne
rect 788 11740 790 11860
rect 910 11740 946 11860
rect 788 11706 946 11740
tri 946 11706 1100 11860 sw
tri 1184 11706 1338 11860 ne
rect 1338 11740 1340 11860
rect 1460 11740 1496 11860
rect 1338 11706 1496 11740
tri 1496 11706 1650 11860 sw
tri 1734 11706 1888 11860 ne
rect 1888 11740 1890 11860
rect 2010 11740 2046 11860
rect 1888 11706 2046 11740
tri 2046 11706 2200 11860 sw
tri 2284 11706 2438 11860 ne
rect 2438 11740 2440 11860
rect 2560 11740 2596 11860
rect 2438 11706 2596 11740
tri 2596 11706 2750 11860 sw
tri 2834 11706 2988 11860 ne
rect 2988 11740 2990 11860
rect 3110 11740 3146 11860
rect 2988 11706 3146 11740
tri 3146 11706 3300 11860 sw
tri 3384 11706 3538 11860 ne
rect 3538 11740 3540 11860
rect 3660 11740 3696 11860
rect 3538 11706 3696 11740
tri 3696 11706 3850 11860 sw
tri 3934 11706 4088 11860 ne
rect 4088 11740 4090 11860
rect 4210 11740 4246 11860
rect 4088 11706 4246 11740
tri 4246 11706 4400 11860 sw
tri 4484 11706 4638 11860 ne
rect 4638 11740 4640 11860
rect 4760 11740 4796 11860
rect 4638 11706 4796 11740
tri 4796 11706 4950 11860 sw
tri 5034 11706 5188 11860 ne
rect 5188 11740 5190 11860
rect 5310 11740 5346 11860
rect 5188 11706 5346 11740
tri 5346 11706 5500 11860 sw
tri 5584 11706 5738 11860 ne
rect 5738 11740 5740 11860
rect 5860 11740 5896 11860
rect 5738 11706 5896 11740
tri 5896 11706 6050 11860 sw
tri 6134 11706 6288 11860 ne
rect 6288 11740 6290 11860
rect 6410 11740 6446 11860
rect 6288 11706 6446 11740
tri 6446 11706 6600 11860 sw
tri 6684 11706 6838 11860 ne
rect 6838 11740 6840 11860
rect 6960 11740 6996 11860
rect 6838 11706 6996 11740
tri 6996 11706 7150 11860 sw
tri 7234 11706 7388 11860 ne
rect 7388 11740 7390 11860
rect 7510 11740 7546 11860
rect 7388 11706 7546 11740
tri 7546 11706 7700 11860 sw
tri 7784 11706 7938 11860 ne
rect 7938 11740 7940 11860
rect 8060 11740 8096 11860
rect 7938 11706 8096 11740
tri 8096 11706 8250 11860 sw
tri 8334 11706 8488 11860 ne
rect 8488 11740 8490 11860
rect 8610 11740 8646 11860
rect 8488 11706 8646 11740
tri 8646 11706 8800 11860 sw
tri 8884 11706 9038 11860 ne
rect 9038 11740 9040 11860
rect 9160 11740 9196 11860
rect 9038 11706 9196 11740
tri 9196 11706 9350 11860 sw
tri 9434 11706 9588 11860 ne
rect 9588 11740 9590 11860
rect 9710 11740 9746 11860
rect 9588 11706 9746 11740
tri 9746 11706 9900 11860 sw
tri 9984 11706 10138 11860 ne
rect 10138 11740 10140 11860
rect 10260 11740 10296 11860
rect 10138 11706 10296 11740
tri 10296 11706 10450 11860 sw
tri 10534 11706 10688 11860 ne
rect 10688 11740 10690 11860
rect 10810 11740 10846 11860
rect 10688 11706 10846 11740
tri 10846 11706 11000 11860 sw
tri 11084 11706 11238 11860 ne
rect 11238 11740 11240 11860
rect 11360 11740 11396 11860
rect 11238 11706 11396 11740
tri 11396 11706 11550 11860 sw
tri 11634 11706 11788 11860 ne
rect 11788 11740 11790 11860
rect 11910 11740 11946 11860
rect 11788 11706 11946 11740
tri 11946 11706 12100 11860 sw
tri 12184 11706 12338 11860 ne
rect 12338 11740 12340 11860
rect 12460 11740 12496 11860
rect 12338 11706 12496 11740
tri 12496 11706 12650 11860 sw
tri 12734 11706 12888 11860 ne
rect 12888 11740 12890 11860
rect 13010 11740 13046 11860
rect 12888 11706 13046 11740
tri 13046 11706 13200 11860 sw
tri 13284 11706 13438 11860 ne
rect 13438 11740 13440 11860
rect 13560 11758 13596 11860
tri 13596 11758 13698 11860 sw
rect 13560 11740 14275 11758
rect 13438 11706 14275 11740
rect -156 11550 0 11706
tri 0 11550 156 11706 sw
tri 238 11550 394 11706 ne
rect 394 11550 550 11706
tri 550 11550 706 11706 sw
tri 788 11550 944 11706 ne
rect 944 11550 1100 11706
tri 1100 11550 1256 11706 sw
tri 1338 11550 1494 11706 ne
rect 1494 11550 1650 11706
tri 1650 11550 1806 11706 sw
tri 1888 11550 2044 11706 ne
rect 2044 11550 2200 11706
tri 2200 11550 2356 11706 sw
tri 2438 11550 2594 11706 ne
rect 2594 11550 2750 11706
tri 2750 11550 2906 11706 sw
tri 2988 11550 3144 11706 ne
rect 3144 11550 3300 11706
tri 3300 11550 3456 11706 sw
tri 3538 11550 3694 11706 ne
rect 3694 11550 3850 11706
tri 3850 11550 4006 11706 sw
tri 4088 11550 4244 11706 ne
rect 4244 11550 4400 11706
tri 4400 11550 4556 11706 sw
tri 4638 11550 4794 11706 ne
rect 4794 11550 4950 11706
tri 4950 11550 5106 11706 sw
tri 5188 11550 5344 11706 ne
rect 5344 11550 5500 11706
tri 5500 11550 5656 11706 sw
tri 5738 11550 5894 11706 ne
rect 5894 11550 6050 11706
tri 6050 11550 6206 11706 sw
tri 6288 11550 6444 11706 ne
rect 6444 11550 6600 11706
tri 6600 11550 6756 11706 sw
tri 6838 11550 6994 11706 ne
rect 6994 11550 7150 11706
tri 7150 11550 7306 11706 sw
tri 7388 11550 7544 11706 ne
rect 7544 11550 7700 11706
tri 7700 11550 7856 11706 sw
tri 7938 11550 8094 11706 ne
rect 8094 11550 8250 11706
tri 8250 11550 8406 11706 sw
tri 8488 11550 8644 11706 ne
rect 8644 11550 8800 11706
tri 8800 11550 8956 11706 sw
tri 9038 11550 9194 11706 ne
rect 9194 11550 9350 11706
tri 9350 11550 9506 11706 sw
tri 9588 11550 9744 11706 ne
rect 9744 11550 9900 11706
tri 9900 11550 10056 11706 sw
tri 10138 11550 10294 11706 ne
rect 10294 11550 10450 11706
tri 10450 11550 10606 11706 sw
tri 10688 11550 10844 11706 ne
rect 10844 11550 11000 11706
tri 11000 11550 11156 11706 sw
tri 11238 11550 11394 11706 ne
rect 11394 11550 11550 11706
tri 11550 11550 11706 11706 sw
tri 11788 11550 11944 11706 ne
rect 11944 11550 12100 11706
tri 12100 11550 12256 11706 sw
tri 12338 11550 12494 11706 ne
rect 12494 11550 12650 11706
tri 12650 11550 12806 11706 sw
tri 12888 11550 13044 11706 ne
rect 13044 11550 13200 11706
tri 13200 11550 13356 11706 sw
tri 13438 11550 13594 11706 ne
rect 13594 11550 14275 11706
rect -2525 11447 -394 11550
tri -394 11447 -291 11550 sw
tri -156 11447 -53 11550 ne
rect -53 11447 156 11550
tri 156 11447 259 11550 sw
tri 394 11447 497 11550 ne
rect 497 11447 706 11550
tri 706 11447 809 11550 sw
tri 944 11447 1047 11550 ne
rect 1047 11447 1256 11550
tri 1256 11447 1359 11550 sw
tri 1494 11447 1597 11550 ne
rect 1597 11447 1806 11550
tri 1806 11447 1909 11550 sw
tri 2044 11447 2147 11550 ne
rect 2147 11447 2356 11550
tri 2356 11447 2459 11550 sw
tri 2594 11447 2697 11550 ne
rect 2697 11447 2906 11550
tri 2906 11447 3009 11550 sw
tri 3144 11447 3247 11550 ne
rect 3247 11447 3456 11550
tri 3456 11447 3559 11550 sw
tri 3694 11447 3797 11550 ne
rect 3797 11447 4006 11550
tri 4006 11447 4109 11550 sw
tri 4244 11447 4347 11550 ne
rect 4347 11447 4556 11550
tri 4556 11447 4659 11550 sw
tri 4794 11447 4897 11550 ne
rect 4897 11447 5106 11550
tri 5106 11447 5209 11550 sw
tri 5344 11447 5447 11550 ne
rect 5447 11447 5656 11550
tri 5656 11447 5759 11550 sw
tri 5894 11447 5997 11550 ne
rect 5997 11447 6206 11550
tri 6206 11447 6309 11550 sw
tri 6444 11447 6547 11550 ne
rect 6547 11447 6756 11550
tri 6756 11447 6859 11550 sw
tri 6994 11447 7097 11550 ne
rect 7097 11447 7306 11550
tri 7306 11447 7409 11550 sw
tri 7544 11447 7647 11550 ne
rect 7647 11447 7856 11550
tri 7856 11447 7959 11550 sw
tri 8094 11447 8197 11550 ne
rect 8197 11447 8406 11550
tri 8406 11447 8509 11550 sw
tri 8644 11447 8747 11550 ne
rect 8747 11447 8956 11550
tri 8956 11447 9059 11550 sw
tri 9194 11447 9297 11550 ne
rect 9297 11447 9506 11550
tri 9506 11447 9609 11550 sw
tri 9744 11447 9847 11550 ne
rect 9847 11447 10056 11550
tri 10056 11447 10159 11550 sw
tri 10294 11447 10397 11550 ne
rect 10397 11447 10606 11550
tri 10606 11447 10709 11550 sw
tri 10844 11447 10947 11550 ne
rect 10947 11447 11156 11550
tri 11156 11447 11259 11550 sw
tri 11394 11447 11497 11550 ne
rect 11497 11447 11706 11550
tri 11706 11447 11809 11550 sw
tri 11944 11447 12047 11550 ne
rect 12047 11447 12256 11550
tri 12256 11447 12359 11550 sw
tri 12494 11447 12597 11550 ne
rect 12597 11447 12806 11550
tri 12806 11447 12909 11550 sw
tri 13044 11447 13147 11550 ne
rect 13147 11447 13356 11550
tri 13356 11447 13459 11550 sw
tri 13594 11447 13697 11550 ne
rect 13697 11447 14275 11550
rect -2525 11310 -291 11447
tri -291 11310 -154 11447 sw
tri -53 11310 84 11447 ne
rect 84 11310 259 11447
tri 259 11310 396 11447 sw
tri 497 11310 634 11447 ne
rect 634 11310 809 11447
tri 809 11310 946 11447 sw
tri 1047 11310 1184 11447 ne
rect 1184 11310 1359 11447
tri 1359 11310 1496 11447 sw
tri 1597 11310 1734 11447 ne
rect 1734 11310 1909 11447
tri 1909 11310 2046 11447 sw
tri 2147 11310 2284 11447 ne
rect 2284 11310 2459 11447
tri 2459 11310 2596 11447 sw
tri 2697 11310 2834 11447 ne
rect 2834 11310 3009 11447
tri 3009 11310 3146 11447 sw
tri 3247 11310 3384 11447 ne
rect 3384 11310 3559 11447
tri 3559 11310 3696 11447 sw
tri 3797 11310 3934 11447 ne
rect 3934 11310 4109 11447
tri 4109 11310 4246 11447 sw
tri 4347 11310 4484 11447 ne
rect 4484 11310 4659 11447
tri 4659 11310 4796 11447 sw
tri 4897 11310 5034 11447 ne
rect 5034 11310 5209 11447
tri 5209 11310 5346 11447 sw
tri 5447 11310 5584 11447 ne
rect 5584 11310 5759 11447
tri 5759 11310 5896 11447 sw
tri 5997 11310 6134 11447 ne
rect 6134 11310 6309 11447
tri 6309 11310 6446 11447 sw
tri 6547 11310 6684 11447 ne
rect 6684 11310 6859 11447
tri 6859 11310 6996 11447 sw
tri 7097 11310 7234 11447 ne
rect 7234 11310 7409 11447
tri 7409 11310 7546 11447 sw
tri 7647 11310 7784 11447 ne
rect 7784 11310 7959 11447
tri 7959 11310 8096 11447 sw
tri 8197 11310 8334 11447 ne
rect 8334 11310 8509 11447
tri 8509 11310 8646 11447 sw
tri 8747 11310 8884 11447 ne
rect 8884 11310 9059 11447
tri 9059 11310 9196 11447 sw
tri 9297 11310 9434 11447 ne
rect 9434 11310 9609 11447
tri 9609 11310 9746 11447 sw
tri 9847 11310 9984 11447 ne
rect 9984 11310 10159 11447
tri 10159 11310 10296 11447 sw
tri 10397 11310 10534 11447 ne
rect 10534 11310 10709 11447
tri 10709 11310 10846 11447 sw
tri 10947 11310 11084 11447 ne
rect 11084 11310 11259 11447
tri 11259 11310 11396 11447 sw
tri 11497 11310 11634 11447 ne
rect 11634 11310 11809 11447
tri 11809 11310 11946 11447 sw
tri 12047 11310 12184 11447 ne
rect 12184 11310 12359 11447
tri 12359 11310 12496 11447 sw
tri 12597 11310 12734 11447 ne
rect 12734 11310 12909 11447
tri 12909 11310 13046 11447 sw
tri 13147 11310 13284 11447 ne
rect 13284 11310 13459 11447
tri 13459 11310 13596 11447 sw
rect -2525 11292 -310 11310
rect -2525 10503 -1525 11292
tri -448 11190 -346 11292 ne
rect -346 11190 -310 11292
rect -190 11190 -154 11310
rect -1025 11000 -447 11053
tri -447 11000 -394 11053 sw
tri -346 11000 -156 11190 ne
rect -156 11156 -154 11190
tri -154 11156 0 11310 sw
tri 84 11156 238 11310 ne
rect 238 11190 240 11310
rect 360 11190 396 11310
rect 238 11156 396 11190
tri 396 11156 550 11310 sw
tri 634 11156 788 11310 ne
rect 788 11190 790 11310
rect 910 11190 946 11310
rect 788 11156 946 11190
tri 946 11156 1100 11310 sw
tri 1184 11156 1338 11310 ne
rect 1338 11190 1340 11310
rect 1460 11190 1496 11310
rect 1338 11156 1496 11190
tri 1496 11156 1650 11310 sw
tri 1734 11156 1888 11310 ne
rect 1888 11190 1890 11310
rect 2010 11190 2046 11310
rect 1888 11156 2046 11190
tri 2046 11156 2200 11310 sw
tri 2284 11156 2438 11310 ne
rect 2438 11190 2440 11310
rect 2560 11190 2596 11310
rect 2438 11156 2596 11190
tri 2596 11156 2750 11310 sw
tri 2834 11156 2988 11310 ne
rect 2988 11190 2990 11310
rect 3110 11190 3146 11310
rect 2988 11156 3146 11190
tri 3146 11156 3300 11310 sw
tri 3384 11156 3538 11310 ne
rect 3538 11190 3540 11310
rect 3660 11190 3696 11310
rect 3538 11156 3696 11190
tri 3696 11156 3850 11310 sw
tri 3934 11156 4088 11310 ne
rect 4088 11190 4090 11310
rect 4210 11190 4246 11310
rect 4088 11156 4246 11190
tri 4246 11156 4400 11310 sw
tri 4484 11156 4638 11310 ne
rect 4638 11190 4640 11310
rect 4760 11190 4796 11310
rect 4638 11156 4796 11190
tri 4796 11156 4950 11310 sw
tri 5034 11156 5188 11310 ne
rect 5188 11190 5190 11310
rect 5310 11190 5346 11310
rect 5188 11156 5346 11190
tri 5346 11156 5500 11310 sw
tri 5584 11156 5738 11310 ne
rect 5738 11190 5740 11310
rect 5860 11190 5896 11310
rect 5738 11156 5896 11190
tri 5896 11156 6050 11310 sw
tri 6134 11156 6288 11310 ne
rect 6288 11190 6290 11310
rect 6410 11190 6446 11310
rect 6288 11156 6446 11190
tri 6446 11156 6600 11310 sw
tri 6684 11156 6838 11310 ne
rect 6838 11190 6840 11310
rect 6960 11190 6996 11310
rect 6838 11156 6996 11190
tri 6996 11156 7150 11310 sw
tri 7234 11156 7388 11310 ne
rect 7388 11190 7390 11310
rect 7510 11190 7546 11310
rect 7388 11156 7546 11190
tri 7546 11156 7700 11310 sw
tri 7784 11156 7938 11310 ne
rect 7938 11190 7940 11310
rect 8060 11190 8096 11310
rect 7938 11156 8096 11190
tri 8096 11156 8250 11310 sw
tri 8334 11156 8488 11310 ne
rect 8488 11190 8490 11310
rect 8610 11190 8646 11310
rect 8488 11156 8646 11190
tri 8646 11156 8800 11310 sw
tri 8884 11156 9038 11310 ne
rect 9038 11190 9040 11310
rect 9160 11190 9196 11310
rect 9038 11156 9196 11190
tri 9196 11156 9350 11310 sw
tri 9434 11156 9588 11310 ne
rect 9588 11190 9590 11310
rect 9710 11190 9746 11310
rect 9588 11156 9746 11190
tri 9746 11156 9900 11310 sw
tri 9984 11156 10138 11310 ne
rect 10138 11190 10140 11310
rect 10260 11190 10296 11310
rect 10138 11156 10296 11190
tri 10296 11156 10450 11310 sw
tri 10534 11156 10688 11310 ne
rect 10688 11190 10690 11310
rect 10810 11190 10846 11310
rect 10688 11156 10846 11190
tri 10846 11156 11000 11310 sw
tri 11084 11156 11238 11310 ne
rect 11238 11190 11240 11310
rect 11360 11190 11396 11310
rect 11238 11156 11396 11190
tri 11396 11156 11550 11310 sw
tri 11634 11156 11788 11310 ne
rect 11788 11190 11790 11310
rect 11910 11190 11946 11310
rect 11788 11156 11946 11190
tri 11946 11156 12100 11310 sw
tri 12184 11156 12338 11310 ne
rect 12338 11190 12340 11310
rect 12460 11190 12496 11310
rect 12338 11156 12496 11190
tri 12496 11156 12650 11310 sw
tri 12734 11156 12888 11310 ne
rect 12888 11190 12890 11310
rect 13010 11190 13046 11310
rect 12888 11156 13046 11190
tri 13046 11156 13200 11310 sw
tri 13284 11156 13438 11310 ne
rect 13438 11190 13440 11310
rect 13560 11208 13596 11310
tri 13596 11208 13698 11310 sw
rect 14775 11208 15775 11997
rect 13560 11190 15775 11208
rect 13438 11156 15775 11190
rect -156 11000 0 11156
tri 0 11000 156 11156 sw
tri 238 11000 394 11156 ne
rect 394 11000 550 11156
tri 550 11000 706 11156 sw
tri 788 11000 944 11156 ne
rect 944 11000 1100 11156
tri 1100 11000 1256 11156 sw
tri 1338 11000 1494 11156 ne
rect 1494 11000 1650 11156
tri 1650 11000 1806 11156 sw
tri 1888 11000 2044 11156 ne
rect 2044 11000 2200 11156
tri 2200 11000 2356 11156 sw
tri 2438 11000 2594 11156 ne
rect 2594 11000 2750 11156
tri 2750 11000 2906 11156 sw
tri 2988 11000 3144 11156 ne
rect 3144 11000 3300 11156
tri 3300 11000 3456 11156 sw
tri 3538 11000 3694 11156 ne
rect 3694 11000 3850 11156
tri 3850 11000 4006 11156 sw
tri 4088 11000 4244 11156 ne
rect 4244 11000 4400 11156
tri 4400 11000 4556 11156 sw
tri 4638 11000 4794 11156 ne
rect 4794 11000 4950 11156
tri 4950 11000 5106 11156 sw
tri 5188 11000 5344 11156 ne
rect 5344 11000 5500 11156
tri 5500 11000 5656 11156 sw
tri 5738 11000 5894 11156 ne
rect 5894 11000 6050 11156
tri 6050 11000 6206 11156 sw
tri 6288 11000 6444 11156 ne
rect 6444 11000 6600 11156
tri 6600 11000 6756 11156 sw
tri 6838 11000 6994 11156 ne
rect 6994 11000 7150 11156
tri 7150 11000 7306 11156 sw
tri 7388 11000 7544 11156 ne
rect 7544 11000 7700 11156
tri 7700 11000 7856 11156 sw
tri 7938 11000 8094 11156 ne
rect 8094 11000 8250 11156
tri 8250 11000 8406 11156 sw
tri 8488 11000 8644 11156 ne
rect 8644 11000 8800 11156
tri 8800 11000 8956 11156 sw
tri 9038 11000 9194 11156 ne
rect 9194 11000 9350 11156
tri 9350 11000 9506 11156 sw
tri 9588 11000 9744 11156 ne
rect 9744 11000 9900 11156
tri 9900 11000 10056 11156 sw
tri 10138 11000 10294 11156 ne
rect 10294 11000 10450 11156
tri 10450 11000 10606 11156 sw
tri 10688 11000 10844 11156 ne
rect 10844 11000 11000 11156
tri 11000 11000 11156 11156 sw
tri 11238 11000 11394 11156 ne
rect 11394 11000 11550 11156
tri 11550 11000 11706 11156 sw
tri 11788 11000 11944 11156 ne
rect 11944 11000 12100 11156
tri 12100 11000 12256 11156 sw
tri 12338 11000 12494 11156 ne
rect 12494 11000 12650 11156
tri 12650 11000 12806 11156 sw
tri 12888 11000 13044 11156 ne
rect 13044 11000 13200 11156
tri 13200 11000 13356 11156 sw
tri 13438 11000 13594 11156 ne
rect 13594 11000 15775 11156
rect -1025 10897 -394 11000
tri -394 10897 -291 11000 sw
tri -156 10897 -53 11000 ne
rect -53 10897 156 11000
tri 156 10897 259 11000 sw
tri 394 10897 497 11000 ne
rect 497 10897 706 11000
tri 706 10897 809 11000 sw
tri 944 10897 1047 11000 ne
rect 1047 10897 1256 11000
tri 1256 10897 1359 11000 sw
tri 1494 10897 1597 11000 ne
rect 1597 10897 1806 11000
tri 1806 10897 1909 11000 sw
tri 2044 10897 2147 11000 ne
rect 2147 10897 2356 11000
tri 2356 10897 2459 11000 sw
tri 2594 10897 2697 11000 ne
rect 2697 10897 2906 11000
tri 2906 10897 3009 11000 sw
tri 3144 10897 3247 11000 ne
rect 3247 10897 3456 11000
tri 3456 10897 3559 11000 sw
tri 3694 10897 3797 11000 ne
rect 3797 10897 4006 11000
tri 4006 10897 4109 11000 sw
tri 4244 10897 4347 11000 ne
rect 4347 10897 4556 11000
tri 4556 10897 4659 11000 sw
tri 4794 10897 4897 11000 ne
rect 4897 10897 5106 11000
tri 5106 10897 5209 11000 sw
tri 5344 10897 5447 11000 ne
rect 5447 10897 5656 11000
tri 5656 10897 5759 11000 sw
tri 5894 10897 5997 11000 ne
rect 5997 10897 6206 11000
tri 6206 10897 6309 11000 sw
tri 6444 10897 6547 11000 ne
rect 6547 10897 6756 11000
tri 6756 10897 6859 11000 sw
tri 6994 10897 7097 11000 ne
rect 7097 10897 7306 11000
tri 7306 10897 7409 11000 sw
tri 7544 10897 7647 11000 ne
rect 7647 10897 7856 11000
tri 7856 10897 7959 11000 sw
tri 8094 10897 8197 11000 ne
rect 8197 10897 8406 11000
tri 8406 10897 8509 11000 sw
tri 8644 10897 8747 11000 ne
rect 8747 10897 8956 11000
tri 8956 10897 9059 11000 sw
tri 9194 10897 9297 11000 ne
rect 9297 10897 9506 11000
tri 9506 10897 9609 11000 sw
tri 9744 10897 9847 11000 ne
rect 9847 10897 10056 11000
tri 10056 10897 10159 11000 sw
tri 10294 10897 10397 11000 ne
rect 10397 10897 10606 11000
tri 10606 10897 10709 11000 sw
tri 10844 10897 10947 11000 ne
rect 10947 10897 11156 11000
tri 11156 10897 11259 11000 sw
tri 11394 10897 11497 11000 ne
rect 11497 10897 11706 11000
tri 11706 10897 11809 11000 sw
tri 11944 10897 12047 11000 ne
rect 12047 10897 12256 11000
tri 12256 10897 12359 11000 sw
tri 12494 10897 12597 11000 ne
rect 12597 10897 12806 11000
tri 12806 10897 12909 11000 sw
tri 13044 10897 13147 11000 ne
rect 13147 10897 13356 11000
tri 13356 10897 13459 11000 sw
tri 13594 10897 13697 11000 ne
rect 13697 10897 15775 11000
rect -1025 10760 -291 10897
tri -291 10760 -154 10897 sw
tri -53 10760 84 10897 ne
rect 84 10760 259 10897
tri 259 10760 396 10897 sw
tri 497 10760 634 10897 ne
rect 634 10760 809 10897
tri 809 10760 946 10897 sw
tri 1047 10760 1184 10897 ne
rect 1184 10760 1359 10897
tri 1359 10760 1496 10897 sw
tri 1597 10760 1734 10897 ne
rect 1734 10760 1909 10897
tri 1909 10760 2046 10897 sw
tri 2147 10760 2284 10897 ne
rect 2284 10760 2459 10897
tri 2459 10760 2596 10897 sw
tri 2697 10760 2834 10897 ne
rect 2834 10760 3009 10897
tri 3009 10760 3146 10897 sw
tri 3247 10760 3384 10897 ne
rect 3384 10760 3559 10897
tri 3559 10760 3696 10897 sw
tri 3797 10760 3934 10897 ne
rect 3934 10760 4109 10897
tri 4109 10760 4246 10897 sw
tri 4347 10760 4484 10897 ne
rect 4484 10760 4659 10897
tri 4659 10760 4796 10897 sw
tri 4897 10760 5034 10897 ne
rect 5034 10760 5209 10897
tri 5209 10760 5346 10897 sw
tri 5447 10760 5584 10897 ne
rect 5584 10760 5759 10897
tri 5759 10760 5896 10897 sw
tri 5997 10760 6134 10897 ne
rect 6134 10760 6309 10897
tri 6309 10760 6446 10897 sw
tri 6547 10760 6684 10897 ne
rect 6684 10760 6859 10897
tri 6859 10760 6996 10897 sw
tri 7097 10760 7234 10897 ne
rect 7234 10760 7409 10897
tri 7409 10760 7546 10897 sw
tri 7647 10760 7784 10897 ne
rect 7784 10760 7959 10897
tri 7959 10760 8096 10897 sw
tri 8197 10760 8334 10897 ne
rect 8334 10760 8509 10897
tri 8509 10760 8646 10897 sw
tri 8747 10760 8884 10897 ne
rect 8884 10760 9059 10897
tri 9059 10760 9196 10897 sw
tri 9297 10760 9434 10897 ne
rect 9434 10760 9609 10897
tri 9609 10760 9746 10897 sw
tri 9847 10760 9984 10897 ne
rect 9984 10760 10159 10897
tri 10159 10760 10296 10897 sw
tri 10397 10760 10534 10897 ne
rect 10534 10760 10709 10897
tri 10709 10760 10846 10897 sw
tri 10947 10760 11084 10897 ne
rect 11084 10760 11259 10897
tri 11259 10760 11396 10897 sw
tri 11497 10760 11634 10897 ne
rect 11634 10760 11809 10897
tri 11809 10760 11946 10897 sw
tri 12047 10760 12184 10897 ne
rect 12184 10760 12359 10897
tri 12359 10760 12496 10897 sw
tri 12597 10760 12734 10897 ne
rect 12734 10760 12909 10897
tri 12909 10760 13046 10897 sw
tri 13147 10760 13284 10897 ne
rect 13284 10760 13459 10897
tri 13459 10760 13596 10897 sw
rect -1025 10742 -310 10760
tri -448 10640 -346 10742 ne
rect -346 10640 -310 10742
rect -190 10640 -154 10760
rect -2525 10450 -447 10503
tri -447 10450 -394 10503 sw
tri -346 10450 -156 10640 ne
rect -156 10606 -154 10640
tri -154 10606 0 10760 sw
tri 84 10606 238 10760 ne
rect 238 10640 240 10760
rect 360 10640 396 10760
rect 238 10606 396 10640
tri 396 10606 550 10760 sw
tri 634 10606 788 10760 ne
rect 788 10640 790 10760
rect 910 10640 946 10760
rect 788 10606 946 10640
tri 946 10606 1100 10760 sw
tri 1184 10606 1338 10760 ne
rect 1338 10640 1340 10760
rect 1460 10640 1496 10760
rect 1338 10606 1496 10640
tri 1496 10606 1650 10760 sw
tri 1734 10606 1888 10760 ne
rect 1888 10640 1890 10760
rect 2010 10640 2046 10760
rect 1888 10606 2046 10640
tri 2046 10606 2200 10760 sw
tri 2284 10606 2438 10760 ne
rect 2438 10640 2440 10760
rect 2560 10640 2596 10760
rect 2438 10606 2596 10640
tri 2596 10606 2750 10760 sw
tri 2834 10606 2988 10760 ne
rect 2988 10640 2990 10760
rect 3110 10640 3146 10760
rect 2988 10606 3146 10640
tri 3146 10606 3300 10760 sw
tri 3384 10606 3538 10760 ne
rect 3538 10640 3540 10760
rect 3660 10640 3696 10760
rect 3538 10606 3696 10640
tri 3696 10606 3850 10760 sw
tri 3934 10606 4088 10760 ne
rect 4088 10640 4090 10760
rect 4210 10640 4246 10760
rect 4088 10606 4246 10640
tri 4246 10606 4400 10760 sw
tri 4484 10606 4638 10760 ne
rect 4638 10640 4640 10760
rect 4760 10640 4796 10760
rect 4638 10606 4796 10640
tri 4796 10606 4950 10760 sw
tri 5034 10606 5188 10760 ne
rect 5188 10640 5190 10760
rect 5310 10640 5346 10760
rect 5188 10606 5346 10640
tri 5346 10606 5500 10760 sw
tri 5584 10606 5738 10760 ne
rect 5738 10640 5740 10760
rect 5860 10640 5896 10760
rect 5738 10606 5896 10640
tri 5896 10606 6050 10760 sw
tri 6134 10606 6288 10760 ne
rect 6288 10640 6290 10760
rect 6410 10640 6446 10760
rect 6288 10606 6446 10640
tri 6446 10606 6600 10760 sw
tri 6684 10606 6838 10760 ne
rect 6838 10640 6840 10760
rect 6960 10640 6996 10760
rect 6838 10606 6996 10640
tri 6996 10606 7150 10760 sw
tri 7234 10606 7388 10760 ne
rect 7388 10640 7390 10760
rect 7510 10640 7546 10760
rect 7388 10606 7546 10640
tri 7546 10606 7700 10760 sw
tri 7784 10606 7938 10760 ne
rect 7938 10640 7940 10760
rect 8060 10640 8096 10760
rect 7938 10606 8096 10640
tri 8096 10606 8250 10760 sw
tri 8334 10606 8488 10760 ne
rect 8488 10640 8490 10760
rect 8610 10640 8646 10760
rect 8488 10606 8646 10640
tri 8646 10606 8800 10760 sw
tri 8884 10606 9038 10760 ne
rect 9038 10640 9040 10760
rect 9160 10640 9196 10760
rect 9038 10606 9196 10640
tri 9196 10606 9350 10760 sw
tri 9434 10606 9588 10760 ne
rect 9588 10640 9590 10760
rect 9710 10640 9746 10760
rect 9588 10606 9746 10640
tri 9746 10606 9900 10760 sw
tri 9984 10606 10138 10760 ne
rect 10138 10640 10140 10760
rect 10260 10640 10296 10760
rect 10138 10606 10296 10640
tri 10296 10606 10450 10760 sw
tri 10534 10606 10688 10760 ne
rect 10688 10640 10690 10760
rect 10810 10640 10846 10760
rect 10688 10606 10846 10640
tri 10846 10606 11000 10760 sw
tri 11084 10606 11238 10760 ne
rect 11238 10640 11240 10760
rect 11360 10640 11396 10760
rect 11238 10606 11396 10640
tri 11396 10606 11550 10760 sw
tri 11634 10606 11788 10760 ne
rect 11788 10640 11790 10760
rect 11910 10640 11946 10760
rect 11788 10606 11946 10640
tri 11946 10606 12100 10760 sw
tri 12184 10606 12338 10760 ne
rect 12338 10640 12340 10760
rect 12460 10640 12496 10760
rect 12338 10606 12496 10640
tri 12496 10606 12650 10760 sw
tri 12734 10606 12888 10760 ne
rect 12888 10640 12890 10760
rect 13010 10640 13046 10760
rect 12888 10606 13046 10640
tri 13046 10606 13200 10760 sw
tri 13284 10606 13438 10760 ne
rect 13438 10640 13440 10760
rect 13560 10658 13596 10760
tri 13596 10658 13698 10760 sw
rect 13560 10640 14275 10658
rect 13438 10606 14275 10640
rect -156 10450 0 10606
tri 0 10450 156 10606 sw
tri 238 10450 394 10606 ne
rect 394 10450 550 10606
tri 550 10450 706 10606 sw
tri 788 10450 944 10606 ne
rect 944 10450 1100 10606
tri 1100 10450 1256 10606 sw
tri 1338 10450 1494 10606 ne
rect 1494 10450 1650 10606
tri 1650 10450 1806 10606 sw
tri 1888 10450 2044 10606 ne
rect 2044 10450 2200 10606
tri 2200 10450 2356 10606 sw
tri 2438 10450 2594 10606 ne
rect 2594 10450 2750 10606
tri 2750 10450 2906 10606 sw
tri 2988 10450 3144 10606 ne
rect 3144 10450 3300 10606
tri 3300 10450 3456 10606 sw
tri 3538 10450 3694 10606 ne
rect 3694 10450 3850 10606
tri 3850 10450 4006 10606 sw
tri 4088 10450 4244 10606 ne
rect 4244 10450 4400 10606
tri 4400 10450 4556 10606 sw
tri 4638 10450 4794 10606 ne
rect 4794 10450 4950 10606
tri 4950 10450 5106 10606 sw
tri 5188 10450 5344 10606 ne
rect 5344 10450 5500 10606
tri 5500 10450 5656 10606 sw
tri 5738 10450 5894 10606 ne
rect 5894 10450 6050 10606
tri 6050 10450 6206 10606 sw
tri 6288 10450 6444 10606 ne
rect 6444 10450 6600 10606
tri 6600 10450 6756 10606 sw
tri 6838 10450 6994 10606 ne
rect 6994 10450 7150 10606
tri 7150 10450 7306 10606 sw
tri 7388 10450 7544 10606 ne
rect 7544 10450 7700 10606
tri 7700 10450 7856 10606 sw
tri 7938 10450 8094 10606 ne
rect 8094 10450 8250 10606
tri 8250 10450 8406 10606 sw
tri 8488 10450 8644 10606 ne
rect 8644 10450 8800 10606
tri 8800 10450 8956 10606 sw
tri 9038 10450 9194 10606 ne
rect 9194 10450 9350 10606
tri 9350 10450 9506 10606 sw
tri 9588 10450 9744 10606 ne
rect 9744 10450 9900 10606
tri 9900 10450 10056 10606 sw
tri 10138 10450 10294 10606 ne
rect 10294 10450 10450 10606
tri 10450 10450 10606 10606 sw
tri 10688 10450 10844 10606 ne
rect 10844 10450 11000 10606
tri 11000 10450 11156 10606 sw
tri 11238 10450 11394 10606 ne
rect 11394 10450 11550 10606
tri 11550 10450 11706 10606 sw
tri 11788 10450 11944 10606 ne
rect 11944 10450 12100 10606
tri 12100 10450 12256 10606 sw
tri 12338 10450 12494 10606 ne
rect 12494 10450 12650 10606
tri 12650 10450 12806 10606 sw
tri 12888 10450 13044 10606 ne
rect 13044 10450 13200 10606
tri 13200 10450 13356 10606 sw
tri 13438 10450 13594 10606 ne
rect 13594 10450 14275 10606
rect -2525 10347 -394 10450
tri -394 10347 -291 10450 sw
tri -156 10347 -53 10450 ne
rect -53 10347 156 10450
tri 156 10347 259 10450 sw
tri 394 10347 497 10450 ne
rect 497 10347 706 10450
tri 706 10347 809 10450 sw
tri 944 10347 1047 10450 ne
rect 1047 10347 1256 10450
tri 1256 10347 1359 10450 sw
tri 1494 10347 1597 10450 ne
rect 1597 10347 1806 10450
tri 1806 10347 1909 10450 sw
tri 2044 10347 2147 10450 ne
rect 2147 10347 2356 10450
tri 2356 10347 2459 10450 sw
tri 2594 10347 2697 10450 ne
rect 2697 10347 2906 10450
tri 2906 10347 3009 10450 sw
tri 3144 10347 3247 10450 ne
rect 3247 10347 3456 10450
tri 3456 10347 3559 10450 sw
tri 3694 10347 3797 10450 ne
rect 3797 10347 4006 10450
tri 4006 10347 4109 10450 sw
tri 4244 10347 4347 10450 ne
rect 4347 10347 4556 10450
tri 4556 10347 4659 10450 sw
tri 4794 10347 4897 10450 ne
rect 4897 10347 5106 10450
tri 5106 10347 5209 10450 sw
tri 5344 10347 5447 10450 ne
rect 5447 10347 5656 10450
tri 5656 10347 5759 10450 sw
tri 5894 10347 5997 10450 ne
rect 5997 10347 6206 10450
tri 6206 10347 6309 10450 sw
tri 6444 10347 6547 10450 ne
rect 6547 10347 6756 10450
tri 6756 10347 6859 10450 sw
tri 6994 10347 7097 10450 ne
rect 7097 10347 7306 10450
tri 7306 10347 7409 10450 sw
tri 7544 10347 7647 10450 ne
rect 7647 10347 7856 10450
tri 7856 10347 7959 10450 sw
tri 8094 10347 8197 10450 ne
rect 8197 10347 8406 10450
tri 8406 10347 8509 10450 sw
tri 8644 10347 8747 10450 ne
rect 8747 10347 8956 10450
tri 8956 10347 9059 10450 sw
tri 9194 10347 9297 10450 ne
rect 9297 10347 9506 10450
tri 9506 10347 9609 10450 sw
tri 9744 10347 9847 10450 ne
rect 9847 10347 10056 10450
tri 10056 10347 10159 10450 sw
tri 10294 10347 10397 10450 ne
rect 10397 10347 10606 10450
tri 10606 10347 10709 10450 sw
tri 10844 10347 10947 10450 ne
rect 10947 10347 11156 10450
tri 11156 10347 11259 10450 sw
tri 11394 10347 11497 10450 ne
rect 11497 10347 11706 10450
tri 11706 10347 11809 10450 sw
tri 11944 10347 12047 10450 ne
rect 12047 10347 12256 10450
tri 12256 10347 12359 10450 sw
tri 12494 10347 12597 10450 ne
rect 12597 10347 12806 10450
tri 12806 10347 12909 10450 sw
tri 13044 10347 13147 10450 ne
rect 13147 10347 13356 10450
tri 13356 10347 13459 10450 sw
tri 13594 10347 13697 10450 ne
rect 13697 10347 14275 10450
rect -2525 10210 -291 10347
tri -291 10210 -154 10347 sw
tri -53 10210 84 10347 ne
rect 84 10210 259 10347
tri 259 10210 396 10347 sw
tri 497 10210 634 10347 ne
rect 634 10210 809 10347
tri 809 10210 946 10347 sw
tri 1047 10210 1184 10347 ne
rect 1184 10210 1359 10347
tri 1359 10210 1496 10347 sw
tri 1597 10210 1734 10347 ne
rect 1734 10210 1909 10347
tri 1909 10210 2046 10347 sw
tri 2147 10210 2284 10347 ne
rect 2284 10210 2459 10347
tri 2459 10210 2596 10347 sw
tri 2697 10210 2834 10347 ne
rect 2834 10210 3009 10347
tri 3009 10210 3146 10347 sw
tri 3247 10210 3384 10347 ne
rect 3384 10210 3559 10347
tri 3559 10210 3696 10347 sw
tri 3797 10210 3934 10347 ne
rect 3934 10210 4109 10347
tri 4109 10210 4246 10347 sw
tri 4347 10210 4484 10347 ne
rect 4484 10210 4659 10347
tri 4659 10210 4796 10347 sw
tri 4897 10210 5034 10347 ne
rect 5034 10210 5209 10347
tri 5209 10210 5346 10347 sw
tri 5447 10210 5584 10347 ne
rect 5584 10210 5759 10347
tri 5759 10210 5896 10347 sw
tri 5997 10210 6134 10347 ne
rect 6134 10210 6309 10347
tri 6309 10210 6446 10347 sw
tri 6547 10210 6684 10347 ne
rect 6684 10210 6859 10347
tri 6859 10210 6996 10347 sw
tri 7097 10210 7234 10347 ne
rect 7234 10210 7409 10347
tri 7409 10210 7546 10347 sw
tri 7647 10210 7784 10347 ne
rect 7784 10210 7959 10347
tri 7959 10210 8096 10347 sw
tri 8197 10210 8334 10347 ne
rect 8334 10210 8509 10347
tri 8509 10210 8646 10347 sw
tri 8747 10210 8884 10347 ne
rect 8884 10210 9059 10347
tri 9059 10210 9196 10347 sw
tri 9297 10210 9434 10347 ne
rect 9434 10210 9609 10347
tri 9609 10210 9746 10347 sw
tri 9847 10210 9984 10347 ne
rect 9984 10210 10159 10347
tri 10159 10210 10296 10347 sw
tri 10397 10210 10534 10347 ne
rect 10534 10210 10709 10347
tri 10709 10210 10846 10347 sw
tri 10947 10210 11084 10347 ne
rect 11084 10210 11259 10347
tri 11259 10210 11396 10347 sw
tri 11497 10210 11634 10347 ne
rect 11634 10210 11809 10347
tri 11809 10210 11946 10347 sw
tri 12047 10210 12184 10347 ne
rect 12184 10210 12359 10347
tri 12359 10210 12496 10347 sw
tri 12597 10210 12734 10347 ne
rect 12734 10210 12909 10347
tri 12909 10210 13046 10347 sw
tri 13147 10210 13284 10347 ne
rect 13284 10210 13459 10347
tri 13459 10210 13596 10347 sw
rect -2525 10192 -310 10210
rect -2525 9403 -1525 10192
tri -448 10090 -346 10192 ne
rect -346 10090 -310 10192
rect -190 10090 -154 10210
rect -1025 9900 -447 9953
tri -447 9900 -394 9953 sw
tri -346 9900 -156 10090 ne
rect -156 10056 -154 10090
tri -154 10056 0 10210 sw
tri 84 10056 238 10210 ne
rect 238 10090 240 10210
rect 360 10090 396 10210
rect 238 10056 396 10090
tri 396 10056 550 10210 sw
tri 634 10056 788 10210 ne
rect 788 10090 790 10210
rect 910 10090 946 10210
rect 788 10056 946 10090
tri 946 10056 1100 10210 sw
tri 1184 10056 1338 10210 ne
rect 1338 10090 1340 10210
rect 1460 10090 1496 10210
rect 1338 10056 1496 10090
tri 1496 10056 1650 10210 sw
tri 1734 10056 1888 10210 ne
rect 1888 10090 1890 10210
rect 2010 10090 2046 10210
rect 1888 10056 2046 10090
tri 2046 10056 2200 10210 sw
tri 2284 10056 2438 10210 ne
rect 2438 10090 2440 10210
rect 2560 10090 2596 10210
rect 2438 10056 2596 10090
tri 2596 10056 2750 10210 sw
tri 2834 10056 2988 10210 ne
rect 2988 10090 2990 10210
rect 3110 10090 3146 10210
rect 2988 10056 3146 10090
tri 3146 10056 3300 10210 sw
tri 3384 10056 3538 10210 ne
rect 3538 10090 3540 10210
rect 3660 10090 3696 10210
rect 3538 10056 3696 10090
tri 3696 10056 3850 10210 sw
tri 3934 10056 4088 10210 ne
rect 4088 10090 4090 10210
rect 4210 10090 4246 10210
rect 4088 10056 4246 10090
tri 4246 10056 4400 10210 sw
tri 4484 10056 4638 10210 ne
rect 4638 10090 4640 10210
rect 4760 10090 4796 10210
rect 4638 10056 4796 10090
tri 4796 10056 4950 10210 sw
tri 5034 10056 5188 10210 ne
rect 5188 10090 5190 10210
rect 5310 10090 5346 10210
rect 5188 10056 5346 10090
tri 5346 10056 5500 10210 sw
tri 5584 10056 5738 10210 ne
rect 5738 10090 5740 10210
rect 5860 10090 5896 10210
rect 5738 10056 5896 10090
tri 5896 10056 6050 10210 sw
tri 6134 10056 6288 10210 ne
rect 6288 10090 6290 10210
rect 6410 10090 6446 10210
rect 6288 10056 6446 10090
tri 6446 10056 6600 10210 sw
tri 6684 10056 6838 10210 ne
rect 6838 10090 6840 10210
rect 6960 10090 6996 10210
rect 6838 10056 6996 10090
tri 6996 10056 7150 10210 sw
tri 7234 10056 7388 10210 ne
rect 7388 10090 7390 10210
rect 7510 10090 7546 10210
rect 7388 10056 7546 10090
tri 7546 10056 7700 10210 sw
tri 7784 10056 7938 10210 ne
rect 7938 10090 7940 10210
rect 8060 10090 8096 10210
rect 7938 10056 8096 10090
tri 8096 10056 8250 10210 sw
tri 8334 10056 8488 10210 ne
rect 8488 10090 8490 10210
rect 8610 10090 8646 10210
rect 8488 10056 8646 10090
tri 8646 10056 8800 10210 sw
tri 8884 10056 9038 10210 ne
rect 9038 10090 9040 10210
rect 9160 10090 9196 10210
rect 9038 10056 9196 10090
tri 9196 10056 9350 10210 sw
tri 9434 10056 9588 10210 ne
rect 9588 10090 9590 10210
rect 9710 10090 9746 10210
rect 9588 10056 9746 10090
tri 9746 10056 9900 10210 sw
tri 9984 10056 10138 10210 ne
rect 10138 10090 10140 10210
rect 10260 10090 10296 10210
rect 10138 10056 10296 10090
tri 10296 10056 10450 10210 sw
tri 10534 10056 10688 10210 ne
rect 10688 10090 10690 10210
rect 10810 10090 10846 10210
rect 10688 10056 10846 10090
tri 10846 10056 11000 10210 sw
tri 11084 10056 11238 10210 ne
rect 11238 10090 11240 10210
rect 11360 10090 11396 10210
rect 11238 10056 11396 10090
tri 11396 10056 11550 10210 sw
tri 11634 10056 11788 10210 ne
rect 11788 10090 11790 10210
rect 11910 10090 11946 10210
rect 11788 10056 11946 10090
tri 11946 10056 12100 10210 sw
tri 12184 10056 12338 10210 ne
rect 12338 10090 12340 10210
rect 12460 10090 12496 10210
rect 12338 10056 12496 10090
tri 12496 10056 12650 10210 sw
tri 12734 10056 12888 10210 ne
rect 12888 10090 12890 10210
rect 13010 10090 13046 10210
rect 12888 10056 13046 10090
tri 13046 10056 13200 10210 sw
tri 13284 10056 13438 10210 ne
rect 13438 10090 13440 10210
rect 13560 10108 13596 10210
tri 13596 10108 13698 10210 sw
rect 14775 10108 15775 10897
rect 13560 10090 15775 10108
rect 13438 10056 15775 10090
rect -156 9900 0 10056
tri 0 9900 156 10056 sw
tri 238 9900 394 10056 ne
rect 394 9900 550 10056
tri 550 9900 706 10056 sw
tri 788 9900 944 10056 ne
rect 944 9900 1100 10056
tri 1100 9900 1256 10056 sw
tri 1338 9900 1494 10056 ne
rect 1494 9900 1650 10056
tri 1650 9900 1806 10056 sw
tri 1888 9900 2044 10056 ne
rect 2044 9900 2200 10056
tri 2200 9900 2356 10056 sw
tri 2438 9900 2594 10056 ne
rect 2594 9900 2750 10056
tri 2750 9900 2906 10056 sw
tri 2988 9900 3144 10056 ne
rect 3144 9900 3300 10056
tri 3300 9900 3456 10056 sw
tri 3538 9900 3694 10056 ne
rect 3694 9900 3850 10056
tri 3850 9900 4006 10056 sw
tri 4088 9900 4244 10056 ne
rect 4244 9900 4400 10056
tri 4400 9900 4556 10056 sw
tri 4638 9900 4794 10056 ne
rect 4794 9900 4950 10056
tri 4950 9900 5106 10056 sw
tri 5188 9900 5344 10056 ne
rect 5344 9900 5500 10056
tri 5500 9900 5656 10056 sw
tri 5738 9900 5894 10056 ne
rect 5894 9900 6050 10056
tri 6050 9900 6206 10056 sw
tri 6288 9900 6444 10056 ne
rect 6444 9900 6600 10056
tri 6600 9900 6756 10056 sw
tri 6838 9900 6994 10056 ne
rect 6994 9900 7150 10056
tri 7150 9900 7306 10056 sw
tri 7388 9900 7544 10056 ne
rect 7544 9900 7700 10056
tri 7700 9900 7856 10056 sw
tri 7938 9900 8094 10056 ne
rect 8094 9900 8250 10056
tri 8250 9900 8406 10056 sw
tri 8488 9900 8644 10056 ne
rect 8644 9900 8800 10056
tri 8800 9900 8956 10056 sw
tri 9038 9900 9194 10056 ne
rect 9194 9900 9350 10056
tri 9350 9900 9506 10056 sw
tri 9588 9900 9744 10056 ne
rect 9744 9900 9900 10056
tri 9900 9900 10056 10056 sw
tri 10138 9900 10294 10056 ne
rect 10294 9900 10450 10056
tri 10450 9900 10606 10056 sw
tri 10688 9900 10844 10056 ne
rect 10844 9900 11000 10056
tri 11000 9900 11156 10056 sw
tri 11238 9900 11394 10056 ne
rect 11394 9900 11550 10056
tri 11550 9900 11706 10056 sw
tri 11788 9900 11944 10056 ne
rect 11944 9900 12100 10056
tri 12100 9900 12256 10056 sw
tri 12338 9900 12494 10056 ne
rect 12494 9900 12650 10056
tri 12650 9900 12806 10056 sw
tri 12888 9900 13044 10056 ne
rect 13044 9900 13200 10056
tri 13200 9900 13356 10056 sw
tri 13438 9900 13594 10056 ne
rect 13594 9900 15775 10056
rect -1025 9797 -394 9900
tri -394 9797 -291 9900 sw
tri -156 9797 -53 9900 ne
rect -53 9797 156 9900
tri 156 9797 259 9900 sw
tri 394 9797 497 9900 ne
rect 497 9797 706 9900
tri 706 9797 809 9900 sw
tri 944 9797 1047 9900 ne
rect 1047 9797 1256 9900
tri 1256 9797 1359 9900 sw
tri 1494 9797 1597 9900 ne
rect 1597 9797 1806 9900
tri 1806 9797 1909 9900 sw
tri 2044 9797 2147 9900 ne
rect 2147 9797 2356 9900
tri 2356 9797 2459 9900 sw
tri 2594 9797 2697 9900 ne
rect 2697 9797 2906 9900
tri 2906 9797 3009 9900 sw
tri 3144 9797 3247 9900 ne
rect 3247 9797 3456 9900
tri 3456 9797 3559 9900 sw
tri 3694 9797 3797 9900 ne
rect 3797 9797 4006 9900
tri 4006 9797 4109 9900 sw
tri 4244 9797 4347 9900 ne
rect 4347 9797 4556 9900
tri 4556 9797 4659 9900 sw
tri 4794 9797 4897 9900 ne
rect 4897 9797 5106 9900
tri 5106 9797 5209 9900 sw
tri 5344 9797 5447 9900 ne
rect 5447 9797 5656 9900
tri 5656 9797 5759 9900 sw
tri 5894 9797 5997 9900 ne
rect 5997 9797 6206 9900
tri 6206 9797 6309 9900 sw
tri 6444 9797 6547 9900 ne
rect 6547 9797 6756 9900
tri 6756 9797 6859 9900 sw
tri 6994 9797 7097 9900 ne
rect 7097 9797 7306 9900
tri 7306 9797 7409 9900 sw
tri 7544 9797 7647 9900 ne
rect 7647 9797 7856 9900
tri 7856 9797 7959 9900 sw
tri 8094 9797 8197 9900 ne
rect 8197 9797 8406 9900
tri 8406 9797 8509 9900 sw
tri 8644 9797 8747 9900 ne
rect 8747 9797 8956 9900
tri 8956 9797 9059 9900 sw
tri 9194 9797 9297 9900 ne
rect 9297 9797 9506 9900
tri 9506 9797 9609 9900 sw
tri 9744 9797 9847 9900 ne
rect 9847 9797 10056 9900
tri 10056 9797 10159 9900 sw
tri 10294 9797 10397 9900 ne
rect 10397 9797 10606 9900
tri 10606 9797 10709 9900 sw
tri 10844 9797 10947 9900 ne
rect 10947 9797 11156 9900
tri 11156 9797 11259 9900 sw
tri 11394 9797 11497 9900 ne
rect 11497 9797 11706 9900
tri 11706 9797 11809 9900 sw
tri 11944 9797 12047 9900 ne
rect 12047 9797 12256 9900
tri 12256 9797 12359 9900 sw
tri 12494 9797 12597 9900 ne
rect 12597 9797 12806 9900
tri 12806 9797 12909 9900 sw
tri 13044 9797 13147 9900 ne
rect 13147 9797 13356 9900
tri 13356 9797 13459 9900 sw
tri 13594 9797 13697 9900 ne
rect 13697 9797 15775 9900
rect -1025 9660 -291 9797
tri -291 9660 -154 9797 sw
tri -53 9660 84 9797 ne
rect 84 9660 259 9797
tri 259 9660 396 9797 sw
tri 497 9660 634 9797 ne
rect 634 9660 809 9797
tri 809 9660 946 9797 sw
tri 1047 9660 1184 9797 ne
rect 1184 9660 1359 9797
tri 1359 9660 1496 9797 sw
tri 1597 9660 1734 9797 ne
rect 1734 9660 1909 9797
tri 1909 9660 2046 9797 sw
tri 2147 9660 2284 9797 ne
rect 2284 9660 2459 9797
tri 2459 9660 2596 9797 sw
tri 2697 9660 2834 9797 ne
rect 2834 9660 3009 9797
tri 3009 9660 3146 9797 sw
tri 3247 9660 3384 9797 ne
rect 3384 9660 3559 9797
tri 3559 9660 3696 9797 sw
tri 3797 9660 3934 9797 ne
rect 3934 9660 4109 9797
tri 4109 9660 4246 9797 sw
tri 4347 9660 4484 9797 ne
rect 4484 9660 4659 9797
tri 4659 9660 4796 9797 sw
tri 4897 9660 5034 9797 ne
rect 5034 9660 5209 9797
tri 5209 9660 5346 9797 sw
tri 5447 9660 5584 9797 ne
rect 5584 9660 5759 9797
tri 5759 9660 5896 9797 sw
tri 5997 9660 6134 9797 ne
rect 6134 9660 6309 9797
tri 6309 9660 6446 9797 sw
tri 6547 9660 6684 9797 ne
rect 6684 9660 6859 9797
tri 6859 9660 6996 9797 sw
tri 7097 9660 7234 9797 ne
rect 7234 9660 7409 9797
tri 7409 9660 7546 9797 sw
tri 7647 9660 7784 9797 ne
rect 7784 9660 7959 9797
tri 7959 9660 8096 9797 sw
tri 8197 9660 8334 9797 ne
rect 8334 9660 8509 9797
tri 8509 9660 8646 9797 sw
tri 8747 9660 8884 9797 ne
rect 8884 9660 9059 9797
tri 9059 9660 9196 9797 sw
tri 9297 9660 9434 9797 ne
rect 9434 9660 9609 9797
tri 9609 9660 9746 9797 sw
tri 9847 9660 9984 9797 ne
rect 9984 9660 10159 9797
tri 10159 9660 10296 9797 sw
tri 10397 9660 10534 9797 ne
rect 10534 9660 10709 9797
tri 10709 9660 10846 9797 sw
tri 10947 9660 11084 9797 ne
rect 11084 9660 11259 9797
tri 11259 9660 11396 9797 sw
tri 11497 9660 11634 9797 ne
rect 11634 9660 11809 9797
tri 11809 9660 11946 9797 sw
tri 12047 9660 12184 9797 ne
rect 12184 9660 12359 9797
tri 12359 9660 12496 9797 sw
tri 12597 9660 12734 9797 ne
rect 12734 9660 12909 9797
tri 12909 9660 13046 9797 sw
tri 13147 9660 13284 9797 ne
rect 13284 9660 13459 9797
tri 13459 9660 13596 9797 sw
rect -1025 9642 -310 9660
tri -448 9540 -346 9642 ne
rect -346 9540 -310 9642
rect -190 9540 -154 9660
rect -2525 9350 -447 9403
tri -447 9350 -394 9403 sw
tri -346 9350 -156 9540 ne
rect -156 9506 -154 9540
tri -154 9506 0 9660 sw
tri 84 9506 238 9660 ne
rect 238 9540 240 9660
rect 360 9540 396 9660
rect 238 9506 396 9540
tri 396 9506 550 9660 sw
tri 634 9506 788 9660 ne
rect 788 9540 790 9660
rect 910 9540 946 9660
rect 788 9506 946 9540
tri 946 9506 1100 9660 sw
tri 1184 9506 1338 9660 ne
rect 1338 9540 1340 9660
rect 1460 9540 1496 9660
rect 1338 9506 1496 9540
tri 1496 9506 1650 9660 sw
tri 1734 9506 1888 9660 ne
rect 1888 9540 1890 9660
rect 2010 9540 2046 9660
rect 1888 9506 2046 9540
tri 2046 9506 2200 9660 sw
tri 2284 9506 2438 9660 ne
rect 2438 9540 2440 9660
rect 2560 9540 2596 9660
rect 2438 9506 2596 9540
tri 2596 9506 2750 9660 sw
tri 2834 9506 2988 9660 ne
rect 2988 9540 2990 9660
rect 3110 9540 3146 9660
rect 2988 9506 3146 9540
tri 3146 9506 3300 9660 sw
tri 3384 9506 3538 9660 ne
rect 3538 9540 3540 9660
rect 3660 9540 3696 9660
rect 3538 9506 3696 9540
tri 3696 9506 3850 9660 sw
tri 3934 9506 4088 9660 ne
rect 4088 9540 4090 9660
rect 4210 9540 4246 9660
rect 4088 9506 4246 9540
tri 4246 9506 4400 9660 sw
tri 4484 9506 4638 9660 ne
rect 4638 9540 4640 9660
rect 4760 9540 4796 9660
rect 4638 9506 4796 9540
tri 4796 9506 4950 9660 sw
tri 5034 9506 5188 9660 ne
rect 5188 9540 5190 9660
rect 5310 9540 5346 9660
rect 5188 9506 5346 9540
tri 5346 9506 5500 9660 sw
tri 5584 9506 5738 9660 ne
rect 5738 9540 5740 9660
rect 5860 9540 5896 9660
rect 5738 9506 5896 9540
tri 5896 9506 6050 9660 sw
tri 6134 9506 6288 9660 ne
rect 6288 9540 6290 9660
rect 6410 9540 6446 9660
rect 6288 9506 6446 9540
tri 6446 9506 6600 9660 sw
tri 6684 9506 6838 9660 ne
rect 6838 9540 6840 9660
rect 6960 9540 6996 9660
rect 6838 9506 6996 9540
tri 6996 9506 7150 9660 sw
tri 7234 9506 7388 9660 ne
rect 7388 9540 7390 9660
rect 7510 9540 7546 9660
rect 7388 9506 7546 9540
tri 7546 9506 7700 9660 sw
tri 7784 9506 7938 9660 ne
rect 7938 9540 7940 9660
rect 8060 9540 8096 9660
rect 7938 9506 8096 9540
tri 8096 9506 8250 9660 sw
tri 8334 9506 8488 9660 ne
rect 8488 9540 8490 9660
rect 8610 9540 8646 9660
rect 8488 9506 8646 9540
tri 8646 9506 8800 9660 sw
tri 8884 9506 9038 9660 ne
rect 9038 9540 9040 9660
rect 9160 9540 9196 9660
rect 9038 9506 9196 9540
tri 9196 9506 9350 9660 sw
tri 9434 9506 9588 9660 ne
rect 9588 9540 9590 9660
rect 9710 9540 9746 9660
rect 9588 9506 9746 9540
tri 9746 9506 9900 9660 sw
tri 9984 9506 10138 9660 ne
rect 10138 9540 10140 9660
rect 10260 9540 10296 9660
rect 10138 9506 10296 9540
tri 10296 9506 10450 9660 sw
tri 10534 9506 10688 9660 ne
rect 10688 9540 10690 9660
rect 10810 9540 10846 9660
rect 10688 9506 10846 9540
tri 10846 9506 11000 9660 sw
tri 11084 9506 11238 9660 ne
rect 11238 9540 11240 9660
rect 11360 9540 11396 9660
rect 11238 9506 11396 9540
tri 11396 9506 11550 9660 sw
tri 11634 9506 11788 9660 ne
rect 11788 9540 11790 9660
rect 11910 9540 11946 9660
rect 11788 9506 11946 9540
tri 11946 9506 12100 9660 sw
tri 12184 9506 12338 9660 ne
rect 12338 9540 12340 9660
rect 12460 9540 12496 9660
rect 12338 9506 12496 9540
tri 12496 9506 12650 9660 sw
tri 12734 9506 12888 9660 ne
rect 12888 9540 12890 9660
rect 13010 9540 13046 9660
rect 12888 9506 13046 9540
tri 13046 9506 13200 9660 sw
tri 13284 9506 13438 9660 ne
rect 13438 9540 13440 9660
rect 13560 9558 13596 9660
tri 13596 9558 13698 9660 sw
rect 13560 9540 14275 9558
rect 13438 9506 14275 9540
rect -156 9350 0 9506
tri 0 9350 156 9506 sw
tri 238 9350 394 9506 ne
rect 394 9350 550 9506
tri 550 9350 706 9506 sw
tri 788 9350 944 9506 ne
rect 944 9350 1100 9506
tri 1100 9350 1256 9506 sw
tri 1338 9350 1494 9506 ne
rect 1494 9350 1650 9506
tri 1650 9350 1806 9506 sw
tri 1888 9350 2044 9506 ne
rect 2044 9350 2200 9506
tri 2200 9350 2356 9506 sw
tri 2438 9350 2594 9506 ne
rect 2594 9350 2750 9506
tri 2750 9350 2906 9506 sw
tri 2988 9350 3144 9506 ne
rect 3144 9350 3300 9506
tri 3300 9350 3456 9506 sw
tri 3538 9350 3694 9506 ne
rect 3694 9350 3850 9506
tri 3850 9350 4006 9506 sw
tri 4088 9350 4244 9506 ne
rect 4244 9350 4400 9506
tri 4400 9350 4556 9506 sw
tri 4638 9350 4794 9506 ne
rect 4794 9350 4950 9506
tri 4950 9350 5106 9506 sw
tri 5188 9350 5344 9506 ne
rect 5344 9350 5500 9506
tri 5500 9350 5656 9506 sw
tri 5738 9350 5894 9506 ne
rect 5894 9350 6050 9506
tri 6050 9350 6206 9506 sw
tri 6288 9350 6444 9506 ne
rect 6444 9350 6600 9506
tri 6600 9350 6756 9506 sw
tri 6838 9350 6994 9506 ne
rect 6994 9350 7150 9506
tri 7150 9350 7306 9506 sw
tri 7388 9350 7544 9506 ne
rect 7544 9350 7700 9506
tri 7700 9350 7856 9506 sw
tri 7938 9350 8094 9506 ne
rect 8094 9350 8250 9506
tri 8250 9350 8406 9506 sw
tri 8488 9350 8644 9506 ne
rect 8644 9350 8800 9506
tri 8800 9350 8956 9506 sw
tri 9038 9350 9194 9506 ne
rect 9194 9350 9350 9506
tri 9350 9350 9506 9506 sw
tri 9588 9350 9744 9506 ne
rect 9744 9350 9900 9506
tri 9900 9350 10056 9506 sw
tri 10138 9350 10294 9506 ne
rect 10294 9350 10450 9506
tri 10450 9350 10606 9506 sw
tri 10688 9350 10844 9506 ne
rect 10844 9350 11000 9506
tri 11000 9350 11156 9506 sw
tri 11238 9350 11394 9506 ne
rect 11394 9350 11550 9506
tri 11550 9350 11706 9506 sw
tri 11788 9350 11944 9506 ne
rect 11944 9350 12100 9506
tri 12100 9350 12256 9506 sw
tri 12338 9350 12494 9506 ne
rect 12494 9350 12650 9506
tri 12650 9350 12806 9506 sw
tri 12888 9350 13044 9506 ne
rect 13044 9350 13200 9506
tri 13200 9350 13356 9506 sw
tri 13438 9350 13594 9506 ne
rect 13594 9350 14275 9506
rect -2525 9247 -394 9350
tri -394 9247 -291 9350 sw
tri -156 9247 -53 9350 ne
rect -53 9247 156 9350
tri 156 9247 259 9350 sw
tri 394 9247 497 9350 ne
rect 497 9247 706 9350
tri 706 9247 809 9350 sw
tri 944 9247 1047 9350 ne
rect 1047 9247 1256 9350
tri 1256 9247 1359 9350 sw
tri 1494 9247 1597 9350 ne
rect 1597 9247 1806 9350
tri 1806 9247 1909 9350 sw
tri 2044 9247 2147 9350 ne
rect 2147 9247 2356 9350
tri 2356 9247 2459 9350 sw
tri 2594 9247 2697 9350 ne
rect 2697 9247 2906 9350
tri 2906 9247 3009 9350 sw
tri 3144 9247 3247 9350 ne
rect 3247 9247 3456 9350
tri 3456 9247 3559 9350 sw
tri 3694 9247 3797 9350 ne
rect 3797 9247 4006 9350
tri 4006 9247 4109 9350 sw
tri 4244 9247 4347 9350 ne
rect 4347 9247 4556 9350
tri 4556 9247 4659 9350 sw
tri 4794 9247 4897 9350 ne
rect 4897 9247 5106 9350
tri 5106 9247 5209 9350 sw
tri 5344 9247 5447 9350 ne
rect 5447 9247 5656 9350
tri 5656 9247 5759 9350 sw
tri 5894 9247 5997 9350 ne
rect 5997 9247 6206 9350
tri 6206 9247 6309 9350 sw
tri 6444 9247 6547 9350 ne
rect 6547 9247 6756 9350
tri 6756 9247 6859 9350 sw
tri 6994 9247 7097 9350 ne
rect 7097 9247 7306 9350
tri 7306 9247 7409 9350 sw
tri 7544 9247 7647 9350 ne
rect 7647 9247 7856 9350
tri 7856 9247 7959 9350 sw
tri 8094 9247 8197 9350 ne
rect 8197 9247 8406 9350
tri 8406 9247 8509 9350 sw
tri 8644 9247 8747 9350 ne
rect 8747 9247 8956 9350
tri 8956 9247 9059 9350 sw
tri 9194 9247 9297 9350 ne
rect 9297 9247 9506 9350
tri 9506 9247 9609 9350 sw
tri 9744 9247 9847 9350 ne
rect 9847 9247 10056 9350
tri 10056 9247 10159 9350 sw
tri 10294 9247 10397 9350 ne
rect 10397 9247 10606 9350
tri 10606 9247 10709 9350 sw
tri 10844 9247 10947 9350 ne
rect 10947 9247 11156 9350
tri 11156 9247 11259 9350 sw
tri 11394 9247 11497 9350 ne
rect 11497 9247 11706 9350
tri 11706 9247 11809 9350 sw
tri 11944 9247 12047 9350 ne
rect 12047 9247 12256 9350
tri 12256 9247 12359 9350 sw
tri 12494 9247 12597 9350 ne
rect 12597 9247 12806 9350
tri 12806 9247 12909 9350 sw
tri 13044 9247 13147 9350 ne
rect 13147 9247 13356 9350
tri 13356 9247 13459 9350 sw
tri 13594 9247 13697 9350 ne
rect 13697 9247 14275 9350
rect -2525 9110 -291 9247
tri -291 9110 -154 9247 sw
tri -53 9110 84 9247 ne
rect 84 9110 259 9247
tri 259 9110 396 9247 sw
tri 497 9110 634 9247 ne
rect 634 9110 809 9247
tri 809 9110 946 9247 sw
tri 1047 9110 1184 9247 ne
rect 1184 9110 1359 9247
tri 1359 9110 1496 9247 sw
tri 1597 9110 1734 9247 ne
rect 1734 9110 1909 9247
tri 1909 9110 2046 9247 sw
tri 2147 9110 2284 9247 ne
rect 2284 9110 2459 9247
tri 2459 9110 2596 9247 sw
tri 2697 9110 2834 9247 ne
rect 2834 9110 3009 9247
tri 3009 9110 3146 9247 sw
tri 3247 9110 3384 9247 ne
rect 3384 9110 3559 9247
tri 3559 9110 3696 9247 sw
tri 3797 9110 3934 9247 ne
rect 3934 9110 4109 9247
tri 4109 9110 4246 9247 sw
tri 4347 9110 4484 9247 ne
rect 4484 9110 4659 9247
tri 4659 9110 4796 9247 sw
tri 4897 9110 5034 9247 ne
rect 5034 9110 5209 9247
tri 5209 9110 5346 9247 sw
tri 5447 9110 5584 9247 ne
rect 5584 9110 5759 9247
tri 5759 9110 5896 9247 sw
tri 5997 9110 6134 9247 ne
rect 6134 9110 6309 9247
tri 6309 9110 6446 9247 sw
tri 6547 9110 6684 9247 ne
rect 6684 9110 6859 9247
tri 6859 9110 6996 9247 sw
tri 7097 9110 7234 9247 ne
rect 7234 9110 7409 9247
tri 7409 9110 7546 9247 sw
tri 7647 9110 7784 9247 ne
rect 7784 9110 7959 9247
tri 7959 9110 8096 9247 sw
tri 8197 9110 8334 9247 ne
rect 8334 9110 8509 9247
tri 8509 9110 8646 9247 sw
tri 8747 9110 8884 9247 ne
rect 8884 9110 9059 9247
tri 9059 9110 9196 9247 sw
tri 9297 9110 9434 9247 ne
rect 9434 9110 9609 9247
tri 9609 9110 9746 9247 sw
tri 9847 9110 9984 9247 ne
rect 9984 9110 10159 9247
tri 10159 9110 10296 9247 sw
tri 10397 9110 10534 9247 ne
rect 10534 9110 10709 9247
tri 10709 9110 10846 9247 sw
tri 10947 9110 11084 9247 ne
rect 11084 9110 11259 9247
tri 11259 9110 11396 9247 sw
tri 11497 9110 11634 9247 ne
rect 11634 9110 11809 9247
tri 11809 9110 11946 9247 sw
tri 12047 9110 12184 9247 ne
rect 12184 9110 12359 9247
tri 12359 9110 12496 9247 sw
tri 12597 9110 12734 9247 ne
rect 12734 9110 12909 9247
tri 12909 9110 13046 9247 sw
tri 13147 9110 13284 9247 ne
rect 13284 9110 13459 9247
tri 13459 9110 13596 9247 sw
rect -2525 9092 -310 9110
rect -2525 8303 -1525 9092
tri -448 8990 -346 9092 ne
rect -346 8990 -310 9092
rect -190 8990 -154 9110
rect -1025 8800 -447 8853
tri -447 8800 -394 8853 sw
tri -346 8800 -156 8990 ne
rect -156 8956 -154 8990
tri -154 8956 0 9110 sw
tri 84 8956 238 9110 ne
rect 238 8990 240 9110
rect 360 8990 396 9110
rect 238 8956 396 8990
tri 396 8956 550 9110 sw
tri 634 8956 788 9110 ne
rect 788 8990 790 9110
rect 910 8990 946 9110
rect 788 8956 946 8990
tri 946 8956 1100 9110 sw
tri 1184 8956 1338 9110 ne
rect 1338 8990 1340 9110
rect 1460 8990 1496 9110
rect 1338 8956 1496 8990
tri 1496 8956 1650 9110 sw
tri 1734 8956 1888 9110 ne
rect 1888 8990 1890 9110
rect 2010 8990 2046 9110
rect 1888 8956 2046 8990
tri 2046 8956 2200 9110 sw
tri 2284 8956 2438 9110 ne
rect 2438 8990 2440 9110
rect 2560 8990 2596 9110
rect 2438 8956 2596 8990
tri 2596 8956 2750 9110 sw
tri 2834 8956 2988 9110 ne
rect 2988 8990 2990 9110
rect 3110 8990 3146 9110
rect 2988 8956 3146 8990
tri 3146 8956 3300 9110 sw
tri 3384 8956 3538 9110 ne
rect 3538 8990 3540 9110
rect 3660 8990 3696 9110
rect 3538 8956 3696 8990
tri 3696 8956 3850 9110 sw
tri 3934 8956 4088 9110 ne
rect 4088 8990 4090 9110
rect 4210 8990 4246 9110
rect 4088 8956 4246 8990
tri 4246 8956 4400 9110 sw
tri 4484 8956 4638 9110 ne
rect 4638 8990 4640 9110
rect 4760 8990 4796 9110
rect 4638 8956 4796 8990
tri 4796 8956 4950 9110 sw
tri 5034 8956 5188 9110 ne
rect 5188 8990 5190 9110
rect 5310 8990 5346 9110
rect 5188 8956 5346 8990
tri 5346 8956 5500 9110 sw
tri 5584 8956 5738 9110 ne
rect 5738 8990 5740 9110
rect 5860 8990 5896 9110
rect 5738 8956 5896 8990
tri 5896 8956 6050 9110 sw
tri 6134 8956 6288 9110 ne
rect 6288 8990 6290 9110
rect 6410 8990 6446 9110
rect 6288 8956 6446 8990
tri 6446 8956 6600 9110 sw
tri 6684 8956 6838 9110 ne
rect 6838 8990 6840 9110
rect 6960 8990 6996 9110
rect 6838 8956 6996 8990
tri 6996 8956 7150 9110 sw
tri 7234 8956 7388 9110 ne
rect 7388 8990 7390 9110
rect 7510 8990 7546 9110
rect 7388 8956 7546 8990
tri 7546 8956 7700 9110 sw
tri 7784 8956 7938 9110 ne
rect 7938 8990 7940 9110
rect 8060 8990 8096 9110
rect 7938 8956 8096 8990
tri 8096 8956 8250 9110 sw
tri 8334 8956 8488 9110 ne
rect 8488 8990 8490 9110
rect 8610 8990 8646 9110
rect 8488 8956 8646 8990
tri 8646 8956 8800 9110 sw
tri 8884 8956 9038 9110 ne
rect 9038 8990 9040 9110
rect 9160 8990 9196 9110
rect 9038 8956 9196 8990
tri 9196 8956 9350 9110 sw
tri 9434 8956 9588 9110 ne
rect 9588 8990 9590 9110
rect 9710 8990 9746 9110
rect 9588 8956 9746 8990
tri 9746 8956 9900 9110 sw
tri 9984 8956 10138 9110 ne
rect 10138 8990 10140 9110
rect 10260 8990 10296 9110
rect 10138 8956 10296 8990
tri 10296 8956 10450 9110 sw
tri 10534 8956 10688 9110 ne
rect 10688 8990 10690 9110
rect 10810 8990 10846 9110
rect 10688 8956 10846 8990
tri 10846 8956 11000 9110 sw
tri 11084 8956 11238 9110 ne
rect 11238 8990 11240 9110
rect 11360 8990 11396 9110
rect 11238 8956 11396 8990
tri 11396 8956 11550 9110 sw
tri 11634 8956 11788 9110 ne
rect 11788 8990 11790 9110
rect 11910 8990 11946 9110
rect 11788 8956 11946 8990
tri 11946 8956 12100 9110 sw
tri 12184 8956 12338 9110 ne
rect 12338 8990 12340 9110
rect 12460 8990 12496 9110
rect 12338 8956 12496 8990
tri 12496 8956 12650 9110 sw
tri 12734 8956 12888 9110 ne
rect 12888 8990 12890 9110
rect 13010 8990 13046 9110
rect 12888 8956 13046 8990
tri 13046 8956 13200 9110 sw
tri 13284 8956 13438 9110 ne
rect 13438 8990 13440 9110
rect 13560 9008 13596 9110
tri 13596 9008 13698 9110 sw
rect 14775 9008 15775 9797
rect 13560 8990 15775 9008
rect 13438 8956 15775 8990
rect -156 8800 0 8956
tri 0 8800 156 8956 sw
tri 238 8800 394 8956 ne
rect 394 8800 550 8956
tri 550 8800 706 8956 sw
tri 788 8800 944 8956 ne
rect 944 8800 1100 8956
tri 1100 8800 1256 8956 sw
tri 1338 8800 1494 8956 ne
rect 1494 8800 1650 8956
tri 1650 8800 1806 8956 sw
tri 1888 8800 2044 8956 ne
rect 2044 8800 2200 8956
tri 2200 8800 2356 8956 sw
tri 2438 8800 2594 8956 ne
rect 2594 8800 2750 8956
tri 2750 8800 2906 8956 sw
tri 2988 8800 3144 8956 ne
rect 3144 8800 3300 8956
tri 3300 8800 3456 8956 sw
tri 3538 8800 3694 8956 ne
rect 3694 8800 3850 8956
tri 3850 8800 4006 8956 sw
tri 4088 8800 4244 8956 ne
rect 4244 8800 4400 8956
tri 4400 8800 4556 8956 sw
tri 4638 8800 4794 8956 ne
rect 4794 8800 4950 8956
tri 4950 8800 5106 8956 sw
tri 5188 8800 5344 8956 ne
rect 5344 8800 5500 8956
tri 5500 8800 5656 8956 sw
tri 5738 8800 5894 8956 ne
rect 5894 8800 6050 8956
tri 6050 8800 6206 8956 sw
tri 6288 8800 6444 8956 ne
rect 6444 8800 6600 8956
tri 6600 8800 6756 8956 sw
tri 6838 8800 6994 8956 ne
rect 6994 8800 7150 8956
tri 7150 8800 7306 8956 sw
tri 7388 8800 7544 8956 ne
rect 7544 8800 7700 8956
tri 7700 8800 7856 8956 sw
tri 7938 8800 8094 8956 ne
rect 8094 8800 8250 8956
tri 8250 8800 8406 8956 sw
tri 8488 8800 8644 8956 ne
rect 8644 8800 8800 8956
tri 8800 8800 8956 8956 sw
tri 9038 8800 9194 8956 ne
rect 9194 8800 9350 8956
tri 9350 8800 9506 8956 sw
tri 9588 8800 9744 8956 ne
rect 9744 8800 9900 8956
tri 9900 8800 10056 8956 sw
tri 10138 8800 10294 8956 ne
rect 10294 8800 10450 8956
tri 10450 8800 10606 8956 sw
tri 10688 8800 10844 8956 ne
rect 10844 8800 11000 8956
tri 11000 8800 11156 8956 sw
tri 11238 8800 11394 8956 ne
rect 11394 8800 11550 8956
tri 11550 8800 11706 8956 sw
tri 11788 8800 11944 8956 ne
rect 11944 8800 12100 8956
tri 12100 8800 12256 8956 sw
tri 12338 8800 12494 8956 ne
rect 12494 8800 12650 8956
tri 12650 8800 12806 8956 sw
tri 12888 8800 13044 8956 ne
rect 13044 8800 13200 8956
tri 13200 8800 13356 8956 sw
tri 13438 8800 13594 8956 ne
rect 13594 8800 15775 8956
rect -1025 8697 -394 8800
tri -394 8697 -291 8800 sw
tri -156 8697 -53 8800 ne
rect -53 8697 156 8800
tri 156 8697 259 8800 sw
tri 394 8697 497 8800 ne
rect 497 8697 706 8800
tri 706 8697 809 8800 sw
tri 944 8697 1047 8800 ne
rect 1047 8697 1256 8800
tri 1256 8697 1359 8800 sw
tri 1494 8697 1597 8800 ne
rect 1597 8697 1806 8800
tri 1806 8697 1909 8800 sw
tri 2044 8697 2147 8800 ne
rect 2147 8697 2356 8800
tri 2356 8697 2459 8800 sw
tri 2594 8697 2697 8800 ne
rect 2697 8697 2906 8800
tri 2906 8697 3009 8800 sw
tri 3144 8697 3247 8800 ne
rect 3247 8697 3456 8800
tri 3456 8697 3559 8800 sw
tri 3694 8697 3797 8800 ne
rect 3797 8697 4006 8800
tri 4006 8697 4109 8800 sw
tri 4244 8697 4347 8800 ne
rect 4347 8697 4556 8800
tri 4556 8697 4659 8800 sw
tri 4794 8697 4897 8800 ne
rect 4897 8697 5106 8800
tri 5106 8697 5209 8800 sw
tri 5344 8697 5447 8800 ne
rect 5447 8697 5656 8800
tri 5656 8697 5759 8800 sw
tri 5894 8697 5997 8800 ne
rect 5997 8697 6206 8800
tri 6206 8697 6309 8800 sw
tri 6444 8697 6547 8800 ne
rect 6547 8697 6756 8800
tri 6756 8697 6859 8800 sw
tri 6994 8697 7097 8800 ne
rect 7097 8697 7306 8800
tri 7306 8697 7409 8800 sw
tri 7544 8697 7647 8800 ne
rect 7647 8697 7856 8800
tri 7856 8697 7959 8800 sw
tri 8094 8697 8197 8800 ne
rect 8197 8697 8406 8800
tri 8406 8697 8509 8800 sw
tri 8644 8697 8747 8800 ne
rect 8747 8697 8956 8800
tri 8956 8697 9059 8800 sw
tri 9194 8697 9297 8800 ne
rect 9297 8697 9506 8800
tri 9506 8697 9609 8800 sw
tri 9744 8697 9847 8800 ne
rect 9847 8697 10056 8800
tri 10056 8697 10159 8800 sw
tri 10294 8697 10397 8800 ne
rect 10397 8697 10606 8800
tri 10606 8697 10709 8800 sw
tri 10844 8697 10947 8800 ne
rect 10947 8697 11156 8800
tri 11156 8697 11259 8800 sw
tri 11394 8697 11497 8800 ne
rect 11497 8697 11706 8800
tri 11706 8697 11809 8800 sw
tri 11944 8697 12047 8800 ne
rect 12047 8697 12256 8800
tri 12256 8697 12359 8800 sw
tri 12494 8697 12597 8800 ne
rect 12597 8697 12806 8800
tri 12806 8697 12909 8800 sw
tri 13044 8697 13147 8800 ne
rect 13147 8697 13356 8800
tri 13356 8697 13459 8800 sw
tri 13594 8697 13697 8800 ne
rect 13697 8697 15775 8800
rect -1025 8560 -291 8697
tri -291 8560 -154 8697 sw
tri -53 8560 84 8697 ne
rect 84 8560 259 8697
tri 259 8560 396 8697 sw
tri 497 8560 634 8697 ne
rect 634 8560 809 8697
tri 809 8560 946 8697 sw
tri 1047 8560 1184 8697 ne
rect 1184 8560 1359 8697
tri 1359 8560 1496 8697 sw
tri 1597 8560 1734 8697 ne
rect 1734 8560 1909 8697
tri 1909 8560 2046 8697 sw
tri 2147 8560 2284 8697 ne
rect 2284 8560 2459 8697
tri 2459 8560 2596 8697 sw
tri 2697 8560 2834 8697 ne
rect 2834 8560 3009 8697
tri 3009 8560 3146 8697 sw
tri 3247 8560 3384 8697 ne
rect 3384 8560 3559 8697
tri 3559 8560 3696 8697 sw
tri 3797 8560 3934 8697 ne
rect 3934 8560 4109 8697
tri 4109 8560 4246 8697 sw
tri 4347 8560 4484 8697 ne
rect 4484 8560 4659 8697
tri 4659 8560 4796 8697 sw
tri 4897 8560 5034 8697 ne
rect 5034 8560 5209 8697
tri 5209 8560 5346 8697 sw
tri 5447 8560 5584 8697 ne
rect 5584 8560 5759 8697
tri 5759 8560 5896 8697 sw
tri 5997 8560 6134 8697 ne
rect 6134 8560 6309 8697
tri 6309 8560 6446 8697 sw
tri 6547 8560 6684 8697 ne
rect 6684 8560 6859 8697
tri 6859 8560 6996 8697 sw
tri 7097 8560 7234 8697 ne
rect 7234 8560 7409 8697
tri 7409 8560 7546 8697 sw
tri 7647 8560 7784 8697 ne
rect 7784 8560 7959 8697
tri 7959 8560 8096 8697 sw
tri 8197 8560 8334 8697 ne
rect 8334 8560 8509 8697
tri 8509 8560 8646 8697 sw
tri 8747 8560 8884 8697 ne
rect 8884 8560 9059 8697
tri 9059 8560 9196 8697 sw
tri 9297 8560 9434 8697 ne
rect 9434 8560 9609 8697
tri 9609 8560 9746 8697 sw
tri 9847 8560 9984 8697 ne
rect 9984 8560 10159 8697
tri 10159 8560 10296 8697 sw
tri 10397 8560 10534 8697 ne
rect 10534 8560 10709 8697
tri 10709 8560 10846 8697 sw
tri 10947 8560 11084 8697 ne
rect 11084 8560 11259 8697
tri 11259 8560 11396 8697 sw
tri 11497 8560 11634 8697 ne
rect 11634 8560 11809 8697
tri 11809 8560 11946 8697 sw
tri 12047 8560 12184 8697 ne
rect 12184 8560 12359 8697
tri 12359 8560 12496 8697 sw
tri 12597 8560 12734 8697 ne
rect 12734 8560 12909 8697
tri 12909 8560 13046 8697 sw
tri 13147 8560 13284 8697 ne
rect 13284 8560 13459 8697
tri 13459 8560 13596 8697 sw
rect -1025 8542 -310 8560
tri -448 8440 -346 8542 ne
rect -346 8440 -310 8542
rect -190 8440 -154 8560
rect -2525 8250 -447 8303
tri -447 8250 -394 8303 sw
tri -346 8250 -156 8440 ne
rect -156 8406 -154 8440
tri -154 8406 0 8560 sw
tri 84 8406 238 8560 ne
rect 238 8440 240 8560
rect 360 8440 396 8560
rect 238 8406 396 8440
tri 396 8406 550 8560 sw
tri 634 8406 788 8560 ne
rect 788 8440 790 8560
rect 910 8440 946 8560
rect 788 8406 946 8440
tri 946 8406 1100 8560 sw
tri 1184 8406 1338 8560 ne
rect 1338 8440 1340 8560
rect 1460 8440 1496 8560
rect 1338 8406 1496 8440
tri 1496 8406 1650 8560 sw
tri 1734 8406 1888 8560 ne
rect 1888 8440 1890 8560
rect 2010 8440 2046 8560
rect 1888 8406 2046 8440
tri 2046 8406 2200 8560 sw
tri 2284 8406 2438 8560 ne
rect 2438 8440 2440 8560
rect 2560 8440 2596 8560
rect 2438 8406 2596 8440
tri 2596 8406 2750 8560 sw
tri 2834 8406 2988 8560 ne
rect 2988 8440 2990 8560
rect 3110 8440 3146 8560
rect 2988 8406 3146 8440
tri 3146 8406 3300 8560 sw
tri 3384 8406 3538 8560 ne
rect 3538 8440 3540 8560
rect 3660 8440 3696 8560
rect 3538 8406 3696 8440
tri 3696 8406 3850 8560 sw
tri 3934 8406 4088 8560 ne
rect 4088 8440 4090 8560
rect 4210 8440 4246 8560
rect 4088 8406 4246 8440
tri 4246 8406 4400 8560 sw
tri 4484 8406 4638 8560 ne
rect 4638 8440 4640 8560
rect 4760 8440 4796 8560
rect 4638 8406 4796 8440
tri 4796 8406 4950 8560 sw
tri 5034 8406 5188 8560 ne
rect 5188 8440 5190 8560
rect 5310 8440 5346 8560
rect 5188 8406 5346 8440
tri 5346 8406 5500 8560 sw
tri 5584 8406 5738 8560 ne
rect 5738 8440 5740 8560
rect 5860 8440 5896 8560
rect 5738 8406 5896 8440
tri 5896 8406 6050 8560 sw
tri 6134 8406 6288 8560 ne
rect 6288 8440 6290 8560
rect 6410 8440 6446 8560
rect 6288 8406 6446 8440
tri 6446 8406 6600 8560 sw
tri 6684 8406 6838 8560 ne
rect 6838 8440 6840 8560
rect 6960 8440 6996 8560
rect 6838 8406 6996 8440
tri 6996 8406 7150 8560 sw
tri 7234 8406 7388 8560 ne
rect 7388 8440 7390 8560
rect 7510 8440 7546 8560
rect 7388 8406 7546 8440
tri 7546 8406 7700 8560 sw
tri 7784 8406 7938 8560 ne
rect 7938 8440 7940 8560
rect 8060 8440 8096 8560
rect 7938 8406 8096 8440
tri 8096 8406 8250 8560 sw
tri 8334 8406 8488 8560 ne
rect 8488 8440 8490 8560
rect 8610 8440 8646 8560
rect 8488 8406 8646 8440
tri 8646 8406 8800 8560 sw
tri 8884 8406 9038 8560 ne
rect 9038 8440 9040 8560
rect 9160 8440 9196 8560
rect 9038 8406 9196 8440
tri 9196 8406 9350 8560 sw
tri 9434 8406 9588 8560 ne
rect 9588 8440 9590 8560
rect 9710 8440 9746 8560
rect 9588 8406 9746 8440
tri 9746 8406 9900 8560 sw
tri 9984 8406 10138 8560 ne
rect 10138 8440 10140 8560
rect 10260 8440 10296 8560
rect 10138 8406 10296 8440
tri 10296 8406 10450 8560 sw
tri 10534 8406 10688 8560 ne
rect 10688 8440 10690 8560
rect 10810 8440 10846 8560
rect 10688 8406 10846 8440
tri 10846 8406 11000 8560 sw
tri 11084 8406 11238 8560 ne
rect 11238 8440 11240 8560
rect 11360 8440 11396 8560
rect 11238 8406 11396 8440
tri 11396 8406 11550 8560 sw
tri 11634 8406 11788 8560 ne
rect 11788 8440 11790 8560
rect 11910 8440 11946 8560
rect 11788 8406 11946 8440
tri 11946 8406 12100 8560 sw
tri 12184 8406 12338 8560 ne
rect 12338 8440 12340 8560
rect 12460 8440 12496 8560
rect 12338 8406 12496 8440
tri 12496 8406 12650 8560 sw
tri 12734 8406 12888 8560 ne
rect 12888 8440 12890 8560
rect 13010 8440 13046 8560
rect 12888 8406 13046 8440
tri 13046 8406 13200 8560 sw
tri 13284 8406 13438 8560 ne
rect 13438 8440 13440 8560
rect 13560 8458 13596 8560
tri 13596 8458 13698 8560 sw
rect 13560 8440 14275 8458
rect 13438 8406 14275 8440
rect -156 8250 0 8406
tri 0 8250 156 8406 sw
tri 238 8250 394 8406 ne
rect 394 8250 550 8406
tri 550 8250 706 8406 sw
tri 788 8250 944 8406 ne
rect 944 8250 1100 8406
tri 1100 8250 1256 8406 sw
tri 1338 8250 1494 8406 ne
rect 1494 8250 1650 8406
tri 1650 8250 1806 8406 sw
tri 1888 8250 2044 8406 ne
rect 2044 8250 2200 8406
tri 2200 8250 2356 8406 sw
tri 2438 8250 2594 8406 ne
rect 2594 8250 2750 8406
tri 2750 8250 2906 8406 sw
tri 2988 8250 3144 8406 ne
rect 3144 8250 3300 8406
tri 3300 8250 3456 8406 sw
tri 3538 8250 3694 8406 ne
rect 3694 8250 3850 8406
tri 3850 8250 4006 8406 sw
tri 4088 8250 4244 8406 ne
rect 4244 8250 4400 8406
tri 4400 8250 4556 8406 sw
tri 4638 8250 4794 8406 ne
rect 4794 8250 4950 8406
tri 4950 8250 5106 8406 sw
tri 5188 8250 5344 8406 ne
rect 5344 8250 5500 8406
tri 5500 8250 5656 8406 sw
tri 5738 8250 5894 8406 ne
rect 5894 8250 6050 8406
tri 6050 8250 6206 8406 sw
tri 6288 8250 6444 8406 ne
rect 6444 8250 6600 8406
tri 6600 8250 6756 8406 sw
tri 6838 8250 6994 8406 ne
rect 6994 8250 7150 8406
tri 7150 8250 7306 8406 sw
tri 7388 8250 7544 8406 ne
rect 7544 8250 7700 8406
tri 7700 8250 7856 8406 sw
tri 7938 8250 8094 8406 ne
rect 8094 8250 8250 8406
tri 8250 8250 8406 8406 sw
tri 8488 8250 8644 8406 ne
rect 8644 8250 8800 8406
tri 8800 8250 8956 8406 sw
tri 9038 8250 9194 8406 ne
rect 9194 8250 9350 8406
tri 9350 8250 9506 8406 sw
tri 9588 8250 9744 8406 ne
rect 9744 8250 9900 8406
tri 9900 8250 10056 8406 sw
tri 10138 8250 10294 8406 ne
rect 10294 8250 10450 8406
tri 10450 8250 10606 8406 sw
tri 10688 8250 10844 8406 ne
rect 10844 8250 11000 8406
tri 11000 8250 11156 8406 sw
tri 11238 8250 11394 8406 ne
rect 11394 8250 11550 8406
tri 11550 8250 11706 8406 sw
tri 11788 8250 11944 8406 ne
rect 11944 8250 12100 8406
tri 12100 8250 12256 8406 sw
tri 12338 8250 12494 8406 ne
rect 12494 8250 12650 8406
tri 12650 8250 12806 8406 sw
tri 12888 8250 13044 8406 ne
rect 13044 8250 13200 8406
tri 13200 8250 13356 8406 sw
tri 13438 8250 13594 8406 ne
rect 13594 8250 14275 8406
rect -2525 8147 -394 8250
tri -394 8147 -291 8250 sw
tri -156 8147 -53 8250 ne
rect -53 8147 156 8250
tri 156 8147 259 8250 sw
tri 394 8147 497 8250 ne
rect 497 8147 706 8250
tri 706 8147 809 8250 sw
tri 944 8147 1047 8250 ne
rect 1047 8147 1256 8250
tri 1256 8147 1359 8250 sw
tri 1494 8147 1597 8250 ne
rect 1597 8147 1806 8250
tri 1806 8147 1909 8250 sw
tri 2044 8147 2147 8250 ne
rect 2147 8147 2356 8250
tri 2356 8147 2459 8250 sw
tri 2594 8147 2697 8250 ne
rect 2697 8147 2906 8250
tri 2906 8147 3009 8250 sw
tri 3144 8147 3247 8250 ne
rect 3247 8147 3456 8250
tri 3456 8147 3559 8250 sw
tri 3694 8147 3797 8250 ne
rect 3797 8147 4006 8250
tri 4006 8147 4109 8250 sw
tri 4244 8147 4347 8250 ne
rect 4347 8147 4556 8250
tri 4556 8147 4659 8250 sw
tri 4794 8147 4897 8250 ne
rect 4897 8147 5106 8250
tri 5106 8147 5209 8250 sw
tri 5344 8147 5447 8250 ne
rect 5447 8147 5656 8250
tri 5656 8147 5759 8250 sw
tri 5894 8147 5997 8250 ne
rect 5997 8147 6206 8250
tri 6206 8147 6309 8250 sw
tri 6444 8147 6547 8250 ne
rect 6547 8147 6756 8250
tri 6756 8147 6859 8250 sw
tri 6994 8147 7097 8250 ne
rect 7097 8147 7306 8250
tri 7306 8147 7409 8250 sw
tri 7544 8147 7647 8250 ne
rect 7647 8147 7856 8250
tri 7856 8147 7959 8250 sw
tri 8094 8147 8197 8250 ne
rect 8197 8147 8406 8250
tri 8406 8147 8509 8250 sw
tri 8644 8147 8747 8250 ne
rect 8747 8147 8956 8250
tri 8956 8147 9059 8250 sw
tri 9194 8147 9297 8250 ne
rect 9297 8147 9506 8250
tri 9506 8147 9609 8250 sw
tri 9744 8147 9847 8250 ne
rect 9847 8147 10056 8250
tri 10056 8147 10159 8250 sw
tri 10294 8147 10397 8250 ne
rect 10397 8147 10606 8250
tri 10606 8147 10709 8250 sw
tri 10844 8147 10947 8250 ne
rect 10947 8147 11156 8250
tri 11156 8147 11259 8250 sw
tri 11394 8147 11497 8250 ne
rect 11497 8147 11706 8250
tri 11706 8147 11809 8250 sw
tri 11944 8147 12047 8250 ne
rect 12047 8147 12256 8250
tri 12256 8147 12359 8250 sw
tri 12494 8147 12597 8250 ne
rect 12597 8147 12806 8250
tri 12806 8147 12909 8250 sw
tri 13044 8147 13147 8250 ne
rect 13147 8147 13356 8250
tri 13356 8147 13459 8250 sw
tri 13594 8147 13697 8250 ne
rect 13697 8147 14275 8250
rect -2525 8010 -291 8147
tri -291 8010 -154 8147 sw
tri -53 8010 84 8147 ne
rect 84 8010 259 8147
tri 259 8010 396 8147 sw
tri 497 8010 634 8147 ne
rect 634 8010 809 8147
tri 809 8010 946 8147 sw
tri 1047 8010 1184 8147 ne
rect 1184 8010 1359 8147
tri 1359 8010 1496 8147 sw
tri 1597 8010 1734 8147 ne
rect 1734 8010 1909 8147
tri 1909 8010 2046 8147 sw
tri 2147 8010 2284 8147 ne
rect 2284 8010 2459 8147
tri 2459 8010 2596 8147 sw
tri 2697 8010 2834 8147 ne
rect 2834 8010 3009 8147
tri 3009 8010 3146 8147 sw
tri 3247 8010 3384 8147 ne
rect 3384 8010 3559 8147
tri 3559 8010 3696 8147 sw
tri 3797 8010 3934 8147 ne
rect 3934 8010 4109 8147
tri 4109 8010 4246 8147 sw
tri 4347 8010 4484 8147 ne
rect 4484 8010 4659 8147
tri 4659 8010 4796 8147 sw
tri 4897 8010 5034 8147 ne
rect 5034 8010 5209 8147
tri 5209 8010 5346 8147 sw
tri 5447 8010 5584 8147 ne
rect 5584 8010 5759 8147
tri 5759 8010 5896 8147 sw
tri 5997 8010 6134 8147 ne
rect 6134 8010 6309 8147
tri 6309 8010 6446 8147 sw
tri 6547 8010 6684 8147 ne
rect 6684 8010 6859 8147
tri 6859 8010 6996 8147 sw
tri 7097 8010 7234 8147 ne
rect 7234 8010 7409 8147
tri 7409 8010 7546 8147 sw
tri 7647 8010 7784 8147 ne
rect 7784 8010 7959 8147
tri 7959 8010 8096 8147 sw
tri 8197 8010 8334 8147 ne
rect 8334 8010 8509 8147
tri 8509 8010 8646 8147 sw
tri 8747 8010 8884 8147 ne
rect 8884 8010 9059 8147
tri 9059 8010 9196 8147 sw
tri 9297 8010 9434 8147 ne
rect 9434 8010 9609 8147
tri 9609 8010 9746 8147 sw
tri 9847 8010 9984 8147 ne
rect 9984 8010 10159 8147
tri 10159 8010 10296 8147 sw
tri 10397 8010 10534 8147 ne
rect 10534 8010 10709 8147
tri 10709 8010 10846 8147 sw
tri 10947 8010 11084 8147 ne
rect 11084 8010 11259 8147
tri 11259 8010 11396 8147 sw
tri 11497 8010 11634 8147 ne
rect 11634 8010 11809 8147
tri 11809 8010 11946 8147 sw
tri 12047 8010 12184 8147 ne
rect 12184 8010 12359 8147
tri 12359 8010 12496 8147 sw
tri 12597 8010 12734 8147 ne
rect 12734 8010 12909 8147
tri 12909 8010 13046 8147 sw
tri 13147 8010 13284 8147 ne
rect 13284 8010 13459 8147
tri 13459 8010 13596 8147 sw
rect -2525 7992 -310 8010
rect -2525 7203 -1525 7992
tri -448 7890 -346 7992 ne
rect -346 7890 -310 7992
rect -190 7890 -154 8010
rect -1025 7700 -447 7753
tri -447 7700 -394 7753 sw
tri -346 7700 -156 7890 ne
rect -156 7856 -154 7890
tri -154 7856 0 8010 sw
tri 84 7856 238 8010 ne
rect 238 7890 240 8010
rect 360 7890 396 8010
rect 238 7856 396 7890
tri 396 7856 550 8010 sw
tri 634 7856 788 8010 ne
rect 788 7890 790 8010
rect 910 7890 946 8010
rect 788 7856 946 7890
tri 946 7856 1100 8010 sw
tri 1184 7856 1338 8010 ne
rect 1338 7890 1340 8010
rect 1460 7890 1496 8010
rect 1338 7856 1496 7890
tri 1496 7856 1650 8010 sw
tri 1734 7856 1888 8010 ne
rect 1888 7890 1890 8010
rect 2010 7890 2046 8010
rect 1888 7856 2046 7890
tri 2046 7856 2200 8010 sw
tri 2284 7856 2438 8010 ne
rect 2438 7890 2440 8010
rect 2560 7890 2596 8010
rect 2438 7856 2596 7890
tri 2596 7856 2750 8010 sw
tri 2834 7856 2988 8010 ne
rect 2988 7890 2990 8010
rect 3110 7890 3146 8010
rect 2988 7856 3146 7890
tri 3146 7856 3300 8010 sw
tri 3384 7856 3538 8010 ne
rect 3538 7890 3540 8010
rect 3660 7890 3696 8010
rect 3538 7856 3696 7890
tri 3696 7856 3850 8010 sw
tri 3934 7856 4088 8010 ne
rect 4088 7890 4090 8010
rect 4210 7890 4246 8010
rect 4088 7856 4246 7890
tri 4246 7856 4400 8010 sw
tri 4484 7856 4638 8010 ne
rect 4638 7890 4640 8010
rect 4760 7890 4796 8010
rect 4638 7856 4796 7890
tri 4796 7856 4950 8010 sw
tri 5034 7856 5188 8010 ne
rect 5188 7890 5190 8010
rect 5310 7890 5346 8010
rect 5188 7856 5346 7890
tri 5346 7856 5500 8010 sw
tri 5584 7856 5738 8010 ne
rect 5738 7890 5740 8010
rect 5860 7890 5896 8010
rect 5738 7856 5896 7890
tri 5896 7856 6050 8010 sw
tri 6134 7856 6288 8010 ne
rect 6288 7890 6290 8010
rect 6410 7890 6446 8010
rect 6288 7856 6446 7890
tri 6446 7856 6600 8010 sw
tri 6684 7856 6838 8010 ne
rect 6838 7890 6840 8010
rect 6960 7890 6996 8010
rect 6838 7856 6996 7890
tri 6996 7856 7150 8010 sw
tri 7234 7856 7388 8010 ne
rect 7388 7890 7390 8010
rect 7510 7890 7546 8010
rect 7388 7856 7546 7890
tri 7546 7856 7700 8010 sw
tri 7784 7856 7938 8010 ne
rect 7938 7890 7940 8010
rect 8060 7890 8096 8010
rect 7938 7856 8096 7890
tri 8096 7856 8250 8010 sw
tri 8334 7856 8488 8010 ne
rect 8488 7890 8490 8010
rect 8610 7890 8646 8010
rect 8488 7856 8646 7890
tri 8646 7856 8800 8010 sw
tri 8884 7856 9038 8010 ne
rect 9038 7890 9040 8010
rect 9160 7890 9196 8010
rect 9038 7856 9196 7890
tri 9196 7856 9350 8010 sw
tri 9434 7856 9588 8010 ne
rect 9588 7890 9590 8010
rect 9710 7890 9746 8010
rect 9588 7856 9746 7890
tri 9746 7856 9900 8010 sw
tri 9984 7856 10138 8010 ne
rect 10138 7890 10140 8010
rect 10260 7890 10296 8010
rect 10138 7856 10296 7890
tri 10296 7856 10450 8010 sw
tri 10534 7856 10688 8010 ne
rect 10688 7890 10690 8010
rect 10810 7890 10846 8010
rect 10688 7856 10846 7890
tri 10846 7856 11000 8010 sw
tri 11084 7856 11238 8010 ne
rect 11238 7890 11240 8010
rect 11360 7890 11396 8010
rect 11238 7856 11396 7890
tri 11396 7856 11550 8010 sw
tri 11634 7856 11788 8010 ne
rect 11788 7890 11790 8010
rect 11910 7890 11946 8010
rect 11788 7856 11946 7890
tri 11946 7856 12100 8010 sw
tri 12184 7856 12338 8010 ne
rect 12338 7890 12340 8010
rect 12460 7890 12496 8010
rect 12338 7856 12496 7890
tri 12496 7856 12650 8010 sw
tri 12734 7856 12888 8010 ne
rect 12888 7890 12890 8010
rect 13010 7890 13046 8010
rect 12888 7856 13046 7890
tri 13046 7856 13200 8010 sw
tri 13284 7856 13438 8010 ne
rect 13438 7890 13440 8010
rect 13560 7908 13596 8010
tri 13596 7908 13698 8010 sw
rect 14775 7908 15775 8697
rect 13560 7890 15775 7908
rect 13438 7856 15775 7890
rect -156 7700 0 7856
tri 0 7700 156 7856 sw
tri 238 7700 394 7856 ne
rect 394 7700 550 7856
tri 550 7700 706 7856 sw
tri 788 7700 944 7856 ne
rect 944 7700 1100 7856
tri 1100 7700 1256 7856 sw
tri 1338 7700 1494 7856 ne
rect 1494 7700 1650 7856
tri 1650 7700 1806 7856 sw
tri 1888 7700 2044 7856 ne
rect 2044 7700 2200 7856
tri 2200 7700 2356 7856 sw
tri 2438 7700 2594 7856 ne
rect 2594 7700 2750 7856
tri 2750 7700 2906 7856 sw
tri 2988 7700 3144 7856 ne
rect 3144 7700 3300 7856
tri 3300 7700 3456 7856 sw
tri 3538 7700 3694 7856 ne
rect 3694 7700 3850 7856
tri 3850 7700 4006 7856 sw
tri 4088 7700 4244 7856 ne
rect 4244 7700 4400 7856
tri 4400 7700 4556 7856 sw
tri 4638 7700 4794 7856 ne
rect 4794 7700 4950 7856
tri 4950 7700 5106 7856 sw
tri 5188 7700 5344 7856 ne
rect 5344 7700 5500 7856
tri 5500 7700 5656 7856 sw
tri 5738 7700 5894 7856 ne
rect 5894 7700 6050 7856
tri 6050 7700 6206 7856 sw
tri 6288 7700 6444 7856 ne
rect 6444 7700 6600 7856
tri 6600 7700 6756 7856 sw
tri 6838 7700 6994 7856 ne
rect 6994 7700 7150 7856
tri 7150 7700 7306 7856 sw
tri 7388 7700 7544 7856 ne
rect 7544 7700 7700 7856
tri 7700 7700 7856 7856 sw
tri 7938 7700 8094 7856 ne
rect 8094 7700 8250 7856
tri 8250 7700 8406 7856 sw
tri 8488 7700 8644 7856 ne
rect 8644 7700 8800 7856
tri 8800 7700 8956 7856 sw
tri 9038 7700 9194 7856 ne
rect 9194 7700 9350 7856
tri 9350 7700 9506 7856 sw
tri 9588 7700 9744 7856 ne
rect 9744 7700 9900 7856
tri 9900 7700 10056 7856 sw
tri 10138 7700 10294 7856 ne
rect 10294 7700 10450 7856
tri 10450 7700 10606 7856 sw
tri 10688 7700 10844 7856 ne
rect 10844 7700 11000 7856
tri 11000 7700 11156 7856 sw
tri 11238 7700 11394 7856 ne
rect 11394 7700 11550 7856
tri 11550 7700 11706 7856 sw
tri 11788 7700 11944 7856 ne
rect 11944 7700 12100 7856
tri 12100 7700 12256 7856 sw
tri 12338 7700 12494 7856 ne
rect 12494 7700 12650 7856
tri 12650 7700 12806 7856 sw
tri 12888 7700 13044 7856 ne
rect 13044 7700 13200 7856
tri 13200 7700 13356 7856 sw
tri 13438 7700 13594 7856 ne
rect 13594 7700 15775 7856
rect -1025 7597 -394 7700
tri -394 7597 -291 7700 sw
tri -156 7597 -53 7700 ne
rect -53 7597 156 7700
tri 156 7597 259 7700 sw
tri 394 7597 497 7700 ne
rect 497 7597 706 7700
tri 706 7597 809 7700 sw
tri 944 7597 1047 7700 ne
rect 1047 7597 1256 7700
tri 1256 7597 1359 7700 sw
tri 1494 7597 1597 7700 ne
rect 1597 7597 1806 7700
tri 1806 7597 1909 7700 sw
tri 2044 7597 2147 7700 ne
rect 2147 7597 2356 7700
tri 2356 7597 2459 7700 sw
tri 2594 7597 2697 7700 ne
rect 2697 7597 2906 7700
tri 2906 7597 3009 7700 sw
tri 3144 7597 3247 7700 ne
rect 3247 7597 3456 7700
tri 3456 7597 3559 7700 sw
tri 3694 7597 3797 7700 ne
rect 3797 7597 4006 7700
tri 4006 7597 4109 7700 sw
tri 4244 7597 4347 7700 ne
rect 4347 7597 4556 7700
tri 4556 7597 4659 7700 sw
tri 4794 7597 4897 7700 ne
rect 4897 7597 5106 7700
tri 5106 7597 5209 7700 sw
tri 5344 7597 5447 7700 ne
rect 5447 7597 5656 7700
tri 5656 7597 5759 7700 sw
tri 5894 7597 5997 7700 ne
rect 5997 7597 6206 7700
tri 6206 7597 6309 7700 sw
tri 6444 7597 6547 7700 ne
rect 6547 7597 6756 7700
tri 6756 7597 6859 7700 sw
tri 6994 7597 7097 7700 ne
rect 7097 7597 7306 7700
tri 7306 7597 7409 7700 sw
tri 7544 7597 7647 7700 ne
rect 7647 7597 7856 7700
tri 7856 7597 7959 7700 sw
tri 8094 7597 8197 7700 ne
rect 8197 7597 8406 7700
tri 8406 7597 8509 7700 sw
tri 8644 7597 8747 7700 ne
rect 8747 7597 8956 7700
tri 8956 7597 9059 7700 sw
tri 9194 7597 9297 7700 ne
rect 9297 7597 9506 7700
tri 9506 7597 9609 7700 sw
tri 9744 7597 9847 7700 ne
rect 9847 7597 10056 7700
tri 10056 7597 10159 7700 sw
tri 10294 7597 10397 7700 ne
rect 10397 7597 10606 7700
tri 10606 7597 10709 7700 sw
tri 10844 7597 10947 7700 ne
rect 10947 7597 11156 7700
tri 11156 7597 11259 7700 sw
tri 11394 7597 11497 7700 ne
rect 11497 7597 11706 7700
tri 11706 7597 11809 7700 sw
tri 11944 7597 12047 7700 ne
rect 12047 7597 12256 7700
tri 12256 7597 12359 7700 sw
tri 12494 7597 12597 7700 ne
rect 12597 7597 12806 7700
tri 12806 7597 12909 7700 sw
tri 13044 7597 13147 7700 ne
rect 13147 7597 13356 7700
tri 13356 7597 13459 7700 sw
tri 13594 7597 13697 7700 ne
rect 13697 7597 15775 7700
rect -1025 7460 -291 7597
tri -291 7460 -154 7597 sw
tri -53 7460 84 7597 ne
rect 84 7460 259 7597
tri 259 7460 396 7597 sw
tri 497 7460 634 7597 ne
rect 634 7460 809 7597
tri 809 7460 946 7597 sw
tri 1047 7460 1184 7597 ne
rect 1184 7460 1359 7597
tri 1359 7460 1496 7597 sw
tri 1597 7460 1734 7597 ne
rect 1734 7460 1909 7597
tri 1909 7460 2046 7597 sw
tri 2147 7460 2284 7597 ne
rect 2284 7460 2459 7597
tri 2459 7460 2596 7597 sw
tri 2697 7460 2834 7597 ne
rect 2834 7460 3009 7597
tri 3009 7460 3146 7597 sw
tri 3247 7460 3384 7597 ne
rect 3384 7460 3559 7597
tri 3559 7460 3696 7597 sw
tri 3797 7460 3934 7597 ne
rect 3934 7460 4109 7597
tri 4109 7460 4246 7597 sw
tri 4347 7460 4484 7597 ne
rect 4484 7460 4659 7597
tri 4659 7460 4796 7597 sw
tri 4897 7460 5034 7597 ne
rect 5034 7460 5209 7597
tri 5209 7460 5346 7597 sw
tri 5447 7460 5584 7597 ne
rect 5584 7460 5759 7597
tri 5759 7460 5896 7597 sw
tri 5997 7460 6134 7597 ne
rect 6134 7460 6309 7597
tri 6309 7460 6446 7597 sw
tri 6547 7460 6684 7597 ne
rect 6684 7460 6859 7597
tri 6859 7460 6996 7597 sw
tri 7097 7460 7234 7597 ne
rect 7234 7460 7409 7597
tri 7409 7460 7546 7597 sw
tri 7647 7460 7784 7597 ne
rect 7784 7460 7959 7597
tri 7959 7460 8096 7597 sw
tri 8197 7460 8334 7597 ne
rect 8334 7460 8509 7597
tri 8509 7460 8646 7597 sw
tri 8747 7460 8884 7597 ne
rect 8884 7460 9059 7597
tri 9059 7460 9196 7597 sw
tri 9297 7460 9434 7597 ne
rect 9434 7460 9609 7597
tri 9609 7460 9746 7597 sw
tri 9847 7460 9984 7597 ne
rect 9984 7460 10159 7597
tri 10159 7460 10296 7597 sw
tri 10397 7460 10534 7597 ne
rect 10534 7460 10709 7597
tri 10709 7460 10846 7597 sw
tri 10947 7460 11084 7597 ne
rect 11084 7460 11259 7597
tri 11259 7460 11396 7597 sw
tri 11497 7460 11634 7597 ne
rect 11634 7460 11809 7597
tri 11809 7460 11946 7597 sw
tri 12047 7460 12184 7597 ne
rect 12184 7460 12359 7597
tri 12359 7460 12496 7597 sw
tri 12597 7460 12734 7597 ne
rect 12734 7460 12909 7597
tri 12909 7460 13046 7597 sw
tri 13147 7460 13284 7597 ne
rect 13284 7460 13459 7597
tri 13459 7460 13596 7597 sw
rect -1025 7442 -310 7460
tri -448 7340 -346 7442 ne
rect -346 7340 -310 7442
rect -190 7340 -154 7460
rect -2525 7150 -447 7203
tri -447 7150 -394 7203 sw
tri -346 7150 -156 7340 ne
rect -156 7306 -154 7340
tri -154 7306 0 7460 sw
tri 84 7306 238 7460 ne
rect 238 7340 240 7460
rect 360 7340 396 7460
rect 238 7306 396 7340
tri 396 7306 550 7460 sw
tri 634 7306 788 7460 ne
rect 788 7340 790 7460
rect 910 7340 946 7460
rect 788 7306 946 7340
tri 946 7306 1100 7460 sw
tri 1184 7306 1338 7460 ne
rect 1338 7340 1340 7460
rect 1460 7340 1496 7460
rect 1338 7306 1496 7340
tri 1496 7306 1650 7460 sw
tri 1734 7306 1888 7460 ne
rect 1888 7340 1890 7460
rect 2010 7340 2046 7460
rect 1888 7306 2046 7340
tri 2046 7306 2200 7460 sw
tri 2284 7306 2438 7460 ne
rect 2438 7340 2440 7460
rect 2560 7340 2596 7460
rect 2438 7306 2596 7340
tri 2596 7306 2750 7460 sw
tri 2834 7306 2988 7460 ne
rect 2988 7340 2990 7460
rect 3110 7340 3146 7460
rect 2988 7306 3146 7340
tri 3146 7306 3300 7460 sw
tri 3384 7306 3538 7460 ne
rect 3538 7340 3540 7460
rect 3660 7340 3696 7460
rect 3538 7306 3696 7340
tri 3696 7306 3850 7460 sw
tri 3934 7306 4088 7460 ne
rect 4088 7340 4090 7460
rect 4210 7340 4246 7460
rect 4088 7306 4246 7340
tri 4246 7306 4400 7460 sw
tri 4484 7306 4638 7460 ne
rect 4638 7340 4640 7460
rect 4760 7340 4796 7460
rect 4638 7306 4796 7340
tri 4796 7306 4950 7460 sw
tri 5034 7306 5188 7460 ne
rect 5188 7340 5190 7460
rect 5310 7340 5346 7460
rect 5188 7306 5346 7340
tri 5346 7306 5500 7460 sw
tri 5584 7306 5738 7460 ne
rect 5738 7340 5740 7460
rect 5860 7340 5896 7460
rect 5738 7306 5896 7340
tri 5896 7306 6050 7460 sw
tri 6134 7306 6288 7460 ne
rect 6288 7340 6290 7460
rect 6410 7340 6446 7460
rect 6288 7306 6446 7340
tri 6446 7306 6600 7460 sw
tri 6684 7306 6838 7460 ne
rect 6838 7340 6840 7460
rect 6960 7340 6996 7460
rect 6838 7306 6996 7340
tri 6996 7306 7150 7460 sw
tri 7234 7306 7388 7460 ne
rect 7388 7340 7390 7460
rect 7510 7340 7546 7460
rect 7388 7306 7546 7340
tri 7546 7306 7700 7460 sw
tri 7784 7306 7938 7460 ne
rect 7938 7340 7940 7460
rect 8060 7340 8096 7460
rect 7938 7306 8096 7340
tri 8096 7306 8250 7460 sw
tri 8334 7306 8488 7460 ne
rect 8488 7340 8490 7460
rect 8610 7340 8646 7460
rect 8488 7306 8646 7340
tri 8646 7306 8800 7460 sw
tri 8884 7306 9038 7460 ne
rect 9038 7340 9040 7460
rect 9160 7340 9196 7460
rect 9038 7306 9196 7340
tri 9196 7306 9350 7460 sw
tri 9434 7306 9588 7460 ne
rect 9588 7340 9590 7460
rect 9710 7340 9746 7460
rect 9588 7306 9746 7340
tri 9746 7306 9900 7460 sw
tri 9984 7306 10138 7460 ne
rect 10138 7340 10140 7460
rect 10260 7340 10296 7460
rect 10138 7306 10296 7340
tri 10296 7306 10450 7460 sw
tri 10534 7306 10688 7460 ne
rect 10688 7340 10690 7460
rect 10810 7340 10846 7460
rect 10688 7306 10846 7340
tri 10846 7306 11000 7460 sw
tri 11084 7306 11238 7460 ne
rect 11238 7340 11240 7460
rect 11360 7340 11396 7460
rect 11238 7306 11396 7340
tri 11396 7306 11550 7460 sw
tri 11634 7306 11788 7460 ne
rect 11788 7340 11790 7460
rect 11910 7340 11946 7460
rect 11788 7306 11946 7340
tri 11946 7306 12100 7460 sw
tri 12184 7306 12338 7460 ne
rect 12338 7340 12340 7460
rect 12460 7340 12496 7460
rect 12338 7306 12496 7340
tri 12496 7306 12650 7460 sw
tri 12734 7306 12888 7460 ne
rect 12888 7340 12890 7460
rect 13010 7340 13046 7460
rect 12888 7306 13046 7340
tri 13046 7306 13200 7460 sw
tri 13284 7306 13438 7460 ne
rect 13438 7340 13440 7460
rect 13560 7358 13596 7460
tri 13596 7358 13698 7460 sw
rect 13560 7340 14275 7358
rect 13438 7306 14275 7340
rect -156 7150 0 7306
tri 0 7150 156 7306 sw
tri 238 7150 394 7306 ne
rect 394 7150 550 7306
tri 550 7150 706 7306 sw
tri 788 7150 944 7306 ne
rect 944 7150 1100 7306
tri 1100 7150 1256 7306 sw
tri 1338 7150 1494 7306 ne
rect 1494 7150 1650 7306
tri 1650 7150 1806 7306 sw
tri 1888 7150 2044 7306 ne
rect 2044 7150 2200 7306
tri 2200 7150 2356 7306 sw
tri 2438 7150 2594 7306 ne
rect 2594 7150 2750 7306
tri 2750 7150 2906 7306 sw
tri 2988 7150 3144 7306 ne
rect 3144 7150 3300 7306
tri 3300 7150 3456 7306 sw
tri 3538 7150 3694 7306 ne
rect 3694 7150 3850 7306
tri 3850 7150 4006 7306 sw
tri 4088 7150 4244 7306 ne
rect 4244 7150 4400 7306
tri 4400 7150 4556 7306 sw
tri 4638 7150 4794 7306 ne
rect 4794 7150 4950 7306
tri 4950 7150 5106 7306 sw
tri 5188 7150 5344 7306 ne
rect 5344 7150 5500 7306
tri 5500 7150 5656 7306 sw
tri 5738 7150 5894 7306 ne
rect 5894 7150 6050 7306
tri 6050 7150 6206 7306 sw
tri 6288 7150 6444 7306 ne
rect 6444 7150 6600 7306
tri 6600 7150 6756 7306 sw
tri 6838 7150 6994 7306 ne
rect 6994 7150 7150 7306
tri 7150 7150 7306 7306 sw
tri 7388 7150 7544 7306 ne
rect 7544 7150 7700 7306
tri 7700 7150 7856 7306 sw
tri 7938 7150 8094 7306 ne
rect 8094 7150 8250 7306
tri 8250 7150 8406 7306 sw
tri 8488 7150 8644 7306 ne
rect 8644 7150 8800 7306
tri 8800 7150 8956 7306 sw
tri 9038 7150 9194 7306 ne
rect 9194 7150 9350 7306
tri 9350 7150 9506 7306 sw
tri 9588 7150 9744 7306 ne
rect 9744 7150 9900 7306
tri 9900 7150 10056 7306 sw
tri 10138 7150 10294 7306 ne
rect 10294 7150 10450 7306
tri 10450 7150 10606 7306 sw
tri 10688 7150 10844 7306 ne
rect 10844 7150 11000 7306
tri 11000 7150 11156 7306 sw
tri 11238 7150 11394 7306 ne
rect 11394 7150 11550 7306
tri 11550 7150 11706 7306 sw
tri 11788 7150 11944 7306 ne
rect 11944 7150 12100 7306
tri 12100 7150 12256 7306 sw
tri 12338 7150 12494 7306 ne
rect 12494 7150 12650 7306
tri 12650 7150 12806 7306 sw
tri 12888 7150 13044 7306 ne
rect 13044 7150 13200 7306
tri 13200 7150 13356 7306 sw
tri 13438 7150 13594 7306 ne
rect 13594 7150 14275 7306
rect -2525 7047 -394 7150
tri -394 7047 -291 7150 sw
tri -156 7047 -53 7150 ne
rect -53 7047 156 7150
tri 156 7047 259 7150 sw
tri 394 7047 497 7150 ne
rect 497 7047 706 7150
tri 706 7047 809 7150 sw
tri 944 7047 1047 7150 ne
rect 1047 7047 1256 7150
tri 1256 7047 1359 7150 sw
tri 1494 7047 1597 7150 ne
rect 1597 7047 1806 7150
tri 1806 7047 1909 7150 sw
tri 2044 7047 2147 7150 ne
rect 2147 7047 2356 7150
tri 2356 7047 2459 7150 sw
tri 2594 7047 2697 7150 ne
rect 2697 7047 2906 7150
tri 2906 7047 3009 7150 sw
tri 3144 7047 3247 7150 ne
rect 3247 7047 3456 7150
tri 3456 7047 3559 7150 sw
tri 3694 7047 3797 7150 ne
rect 3797 7047 4006 7150
tri 4006 7047 4109 7150 sw
tri 4244 7047 4347 7150 ne
rect 4347 7047 4556 7150
tri 4556 7047 4659 7150 sw
tri 4794 7047 4897 7150 ne
rect 4897 7047 5106 7150
tri 5106 7047 5209 7150 sw
tri 5344 7047 5447 7150 ne
rect 5447 7047 5656 7150
tri 5656 7047 5759 7150 sw
tri 5894 7047 5997 7150 ne
rect 5997 7047 6206 7150
tri 6206 7047 6309 7150 sw
tri 6444 7047 6547 7150 ne
rect 6547 7047 6756 7150
tri 6756 7047 6859 7150 sw
tri 6994 7047 7097 7150 ne
rect 7097 7047 7306 7150
tri 7306 7047 7409 7150 sw
tri 7544 7047 7647 7150 ne
rect 7647 7047 7856 7150
tri 7856 7047 7959 7150 sw
tri 8094 7047 8197 7150 ne
rect 8197 7047 8406 7150
tri 8406 7047 8509 7150 sw
tri 8644 7047 8747 7150 ne
rect 8747 7047 8956 7150
tri 8956 7047 9059 7150 sw
tri 9194 7047 9297 7150 ne
rect 9297 7047 9506 7150
tri 9506 7047 9609 7150 sw
tri 9744 7047 9847 7150 ne
rect 9847 7047 10056 7150
tri 10056 7047 10159 7150 sw
tri 10294 7047 10397 7150 ne
rect 10397 7047 10606 7150
tri 10606 7047 10709 7150 sw
tri 10844 7047 10947 7150 ne
rect 10947 7047 11156 7150
tri 11156 7047 11259 7150 sw
tri 11394 7047 11497 7150 ne
rect 11497 7047 11706 7150
tri 11706 7047 11809 7150 sw
tri 11944 7047 12047 7150 ne
rect 12047 7047 12256 7150
tri 12256 7047 12359 7150 sw
tri 12494 7047 12597 7150 ne
rect 12597 7047 12806 7150
tri 12806 7047 12909 7150 sw
tri 13044 7047 13147 7150 ne
rect 13147 7047 13356 7150
tri 13356 7047 13459 7150 sw
tri 13594 7047 13697 7150 ne
rect 13697 7047 14275 7150
rect -2525 6910 -291 7047
tri -291 6910 -154 7047 sw
tri -53 6910 84 7047 ne
rect 84 6910 259 7047
tri 259 6910 396 7047 sw
tri 497 6910 634 7047 ne
rect 634 6910 809 7047
tri 809 6910 946 7047 sw
tri 1047 6910 1184 7047 ne
rect 1184 6910 1359 7047
tri 1359 6910 1496 7047 sw
tri 1597 6910 1734 7047 ne
rect 1734 6910 1909 7047
tri 1909 6910 2046 7047 sw
tri 2147 6910 2284 7047 ne
rect 2284 6910 2459 7047
tri 2459 6910 2596 7047 sw
tri 2697 6910 2834 7047 ne
rect 2834 6910 3009 7047
tri 3009 6910 3146 7047 sw
tri 3247 6910 3384 7047 ne
rect 3384 6910 3559 7047
tri 3559 6910 3696 7047 sw
tri 3797 6910 3934 7047 ne
rect 3934 6910 4109 7047
tri 4109 6910 4246 7047 sw
tri 4347 6910 4484 7047 ne
rect 4484 6910 4659 7047
tri 4659 6910 4796 7047 sw
tri 4897 6910 5034 7047 ne
rect 5034 6910 5209 7047
tri 5209 6910 5346 7047 sw
tri 5447 6910 5584 7047 ne
rect 5584 6910 5759 7047
tri 5759 6910 5896 7047 sw
tri 5997 6910 6134 7047 ne
rect 6134 6910 6309 7047
tri 6309 6910 6446 7047 sw
tri 6547 6910 6684 7047 ne
rect 6684 6910 6859 7047
tri 6859 6910 6996 7047 sw
tri 7097 6910 7234 7047 ne
rect 7234 6910 7409 7047
tri 7409 6910 7546 7047 sw
tri 7647 6910 7784 7047 ne
rect 7784 6910 7959 7047
tri 7959 6910 8096 7047 sw
tri 8197 6910 8334 7047 ne
rect 8334 6910 8509 7047
tri 8509 6910 8646 7047 sw
tri 8747 6910 8884 7047 ne
rect 8884 6910 9059 7047
tri 9059 6910 9196 7047 sw
tri 9297 6910 9434 7047 ne
rect 9434 6910 9609 7047
tri 9609 6910 9746 7047 sw
tri 9847 6910 9984 7047 ne
rect 9984 6910 10159 7047
tri 10159 6910 10296 7047 sw
tri 10397 6910 10534 7047 ne
rect 10534 6910 10709 7047
tri 10709 6910 10846 7047 sw
tri 10947 6910 11084 7047 ne
rect 11084 6910 11259 7047
tri 11259 6910 11396 7047 sw
tri 11497 6910 11634 7047 ne
rect 11634 6910 11809 7047
tri 11809 6910 11946 7047 sw
tri 12047 6910 12184 7047 ne
rect 12184 6910 12359 7047
tri 12359 6910 12496 7047 sw
tri 12597 6910 12734 7047 ne
rect 12734 6910 12909 7047
tri 12909 6910 13046 7047 sw
tri 13147 6910 13284 7047 ne
rect 13284 6910 13459 7047
tri 13459 6910 13596 7047 sw
rect -2525 6892 -310 6910
rect -2525 6103 -1525 6892
tri -448 6790 -346 6892 ne
rect -346 6790 -310 6892
rect -190 6790 -154 6910
rect -1025 6600 -447 6653
tri -447 6600 -394 6653 sw
tri -346 6600 -156 6790 ne
rect -156 6756 -154 6790
tri -154 6756 0 6910 sw
tri 84 6756 238 6910 ne
rect 238 6790 240 6910
rect 360 6790 396 6910
rect 238 6756 396 6790
tri 396 6756 550 6910 sw
tri 634 6756 788 6910 ne
rect 788 6790 790 6910
rect 910 6790 946 6910
rect 788 6756 946 6790
tri 946 6756 1100 6910 sw
tri 1184 6756 1338 6910 ne
rect 1338 6790 1340 6910
rect 1460 6790 1496 6910
rect 1338 6756 1496 6790
tri 1496 6756 1650 6910 sw
tri 1734 6756 1888 6910 ne
rect 1888 6790 1890 6910
rect 2010 6790 2046 6910
rect 1888 6756 2046 6790
tri 2046 6756 2200 6910 sw
tri 2284 6756 2438 6910 ne
rect 2438 6790 2440 6910
rect 2560 6790 2596 6910
rect 2438 6756 2596 6790
tri 2596 6756 2750 6910 sw
tri 2834 6756 2988 6910 ne
rect 2988 6790 2990 6910
rect 3110 6790 3146 6910
rect 2988 6756 3146 6790
tri 3146 6756 3300 6910 sw
tri 3384 6756 3538 6910 ne
rect 3538 6790 3540 6910
rect 3660 6790 3696 6910
rect 3538 6756 3696 6790
tri 3696 6756 3850 6910 sw
tri 3934 6756 4088 6910 ne
rect 4088 6790 4090 6910
rect 4210 6790 4246 6910
rect 4088 6756 4246 6790
tri 4246 6756 4400 6910 sw
tri 4484 6756 4638 6910 ne
rect 4638 6790 4640 6910
rect 4760 6790 4796 6910
rect 4638 6756 4796 6790
tri 4796 6756 4950 6910 sw
tri 5034 6756 5188 6910 ne
rect 5188 6790 5190 6910
rect 5310 6790 5346 6910
rect 5188 6756 5346 6790
tri 5346 6756 5500 6910 sw
tri 5584 6756 5738 6910 ne
rect 5738 6790 5740 6910
rect 5860 6790 5896 6910
rect 5738 6756 5896 6790
tri 5896 6756 6050 6910 sw
tri 6134 6756 6288 6910 ne
rect 6288 6790 6290 6910
rect 6410 6790 6446 6910
rect 6288 6756 6446 6790
tri 6446 6756 6600 6910 sw
tri 6684 6756 6838 6910 ne
rect 6838 6790 6840 6910
rect 6960 6790 6996 6910
rect 6838 6756 6996 6790
tri 6996 6756 7150 6910 sw
tri 7234 6756 7388 6910 ne
rect 7388 6790 7390 6910
rect 7510 6790 7546 6910
rect 7388 6756 7546 6790
tri 7546 6756 7700 6910 sw
tri 7784 6756 7938 6910 ne
rect 7938 6790 7940 6910
rect 8060 6790 8096 6910
rect 7938 6756 8096 6790
tri 8096 6756 8250 6910 sw
tri 8334 6756 8488 6910 ne
rect 8488 6790 8490 6910
rect 8610 6790 8646 6910
rect 8488 6756 8646 6790
tri 8646 6756 8800 6910 sw
tri 8884 6756 9038 6910 ne
rect 9038 6790 9040 6910
rect 9160 6790 9196 6910
rect 9038 6756 9196 6790
tri 9196 6756 9350 6910 sw
tri 9434 6756 9588 6910 ne
rect 9588 6790 9590 6910
rect 9710 6790 9746 6910
rect 9588 6756 9746 6790
tri 9746 6756 9900 6910 sw
tri 9984 6756 10138 6910 ne
rect 10138 6790 10140 6910
rect 10260 6790 10296 6910
rect 10138 6756 10296 6790
tri 10296 6756 10450 6910 sw
tri 10534 6756 10688 6910 ne
rect 10688 6790 10690 6910
rect 10810 6790 10846 6910
rect 10688 6756 10846 6790
tri 10846 6756 11000 6910 sw
tri 11084 6756 11238 6910 ne
rect 11238 6790 11240 6910
rect 11360 6790 11396 6910
rect 11238 6756 11396 6790
tri 11396 6756 11550 6910 sw
tri 11634 6756 11788 6910 ne
rect 11788 6790 11790 6910
rect 11910 6790 11946 6910
rect 11788 6756 11946 6790
tri 11946 6756 12100 6910 sw
tri 12184 6756 12338 6910 ne
rect 12338 6790 12340 6910
rect 12460 6790 12496 6910
rect 12338 6756 12496 6790
tri 12496 6756 12650 6910 sw
tri 12734 6756 12888 6910 ne
rect 12888 6790 12890 6910
rect 13010 6790 13046 6910
rect 12888 6756 13046 6790
tri 13046 6756 13200 6910 sw
tri 13284 6756 13438 6910 ne
rect 13438 6790 13440 6910
rect 13560 6808 13596 6910
tri 13596 6808 13698 6910 sw
rect 14775 6808 15775 7597
rect 13560 6790 15775 6808
rect 13438 6756 15775 6790
rect -156 6600 0 6756
tri 0 6600 156 6756 sw
tri 238 6600 394 6756 ne
rect 394 6600 550 6756
tri 550 6600 706 6756 sw
tri 788 6600 944 6756 ne
rect 944 6600 1100 6756
tri 1100 6600 1256 6756 sw
tri 1338 6600 1494 6756 ne
rect 1494 6600 1650 6756
tri 1650 6600 1806 6756 sw
tri 1888 6600 2044 6756 ne
rect 2044 6600 2200 6756
tri 2200 6600 2356 6756 sw
tri 2438 6600 2594 6756 ne
rect 2594 6600 2750 6756
tri 2750 6600 2906 6756 sw
tri 2988 6600 3144 6756 ne
rect 3144 6600 3300 6756
tri 3300 6600 3456 6756 sw
tri 3538 6600 3694 6756 ne
rect 3694 6600 3850 6756
tri 3850 6600 4006 6756 sw
tri 4088 6600 4244 6756 ne
rect 4244 6600 4400 6756
tri 4400 6600 4556 6756 sw
tri 4638 6600 4794 6756 ne
rect 4794 6600 4950 6756
tri 4950 6600 5106 6756 sw
tri 5188 6600 5344 6756 ne
rect 5344 6600 5500 6756
tri 5500 6600 5656 6756 sw
tri 5738 6600 5894 6756 ne
rect 5894 6600 6050 6756
tri 6050 6600 6206 6756 sw
tri 6288 6600 6444 6756 ne
rect 6444 6600 6600 6756
tri 6600 6600 6756 6756 sw
tri 6838 6600 6994 6756 ne
rect 6994 6600 7150 6756
tri 7150 6600 7306 6756 sw
tri 7388 6600 7544 6756 ne
rect 7544 6600 7700 6756
tri 7700 6600 7856 6756 sw
tri 7938 6600 8094 6756 ne
rect 8094 6600 8250 6756
tri 8250 6600 8406 6756 sw
tri 8488 6600 8644 6756 ne
rect 8644 6600 8800 6756
tri 8800 6600 8956 6756 sw
tri 9038 6600 9194 6756 ne
rect 9194 6600 9350 6756
tri 9350 6600 9506 6756 sw
tri 9588 6600 9744 6756 ne
rect 9744 6600 9900 6756
tri 9900 6600 10056 6756 sw
tri 10138 6600 10294 6756 ne
rect 10294 6600 10450 6756
tri 10450 6600 10606 6756 sw
tri 10688 6600 10844 6756 ne
rect 10844 6600 11000 6756
tri 11000 6600 11156 6756 sw
tri 11238 6600 11394 6756 ne
rect 11394 6600 11550 6756
tri 11550 6600 11706 6756 sw
tri 11788 6600 11944 6756 ne
rect 11944 6600 12100 6756
tri 12100 6600 12256 6756 sw
tri 12338 6600 12494 6756 ne
rect 12494 6600 12650 6756
tri 12650 6600 12806 6756 sw
tri 12888 6600 13044 6756 ne
rect 13044 6600 13200 6756
tri 13200 6600 13356 6756 sw
tri 13438 6600 13594 6756 ne
rect 13594 6600 15775 6756
rect -1025 6497 -394 6600
tri -394 6497 -291 6600 sw
tri -156 6497 -53 6600 ne
rect -53 6497 156 6600
tri 156 6497 259 6600 sw
tri 394 6497 497 6600 ne
rect 497 6497 706 6600
tri 706 6497 809 6600 sw
tri 944 6497 1047 6600 ne
rect 1047 6497 1256 6600
tri 1256 6497 1359 6600 sw
tri 1494 6497 1597 6600 ne
rect 1597 6497 1806 6600
tri 1806 6497 1909 6600 sw
tri 2044 6497 2147 6600 ne
rect 2147 6497 2356 6600
tri 2356 6497 2459 6600 sw
tri 2594 6497 2697 6600 ne
rect 2697 6497 2906 6600
tri 2906 6497 3009 6600 sw
tri 3144 6497 3247 6600 ne
rect 3247 6497 3456 6600
tri 3456 6497 3559 6600 sw
tri 3694 6497 3797 6600 ne
rect 3797 6497 4006 6600
tri 4006 6497 4109 6600 sw
tri 4244 6497 4347 6600 ne
rect 4347 6497 4556 6600
tri 4556 6497 4659 6600 sw
tri 4794 6497 4897 6600 ne
rect 4897 6497 5106 6600
tri 5106 6497 5209 6600 sw
tri 5344 6497 5447 6600 ne
rect 5447 6497 5656 6600
tri 5656 6497 5759 6600 sw
tri 5894 6497 5997 6600 ne
rect 5997 6497 6206 6600
tri 6206 6497 6309 6600 sw
tri 6444 6497 6547 6600 ne
rect 6547 6497 6756 6600
tri 6756 6497 6859 6600 sw
tri 6994 6497 7097 6600 ne
rect 7097 6497 7306 6600
tri 7306 6497 7409 6600 sw
tri 7544 6497 7647 6600 ne
rect 7647 6497 7856 6600
tri 7856 6497 7959 6600 sw
tri 8094 6497 8197 6600 ne
rect 8197 6497 8406 6600
tri 8406 6497 8509 6600 sw
tri 8644 6497 8747 6600 ne
rect 8747 6497 8956 6600
tri 8956 6497 9059 6600 sw
tri 9194 6497 9297 6600 ne
rect 9297 6497 9506 6600
tri 9506 6497 9609 6600 sw
tri 9744 6497 9847 6600 ne
rect 9847 6497 10056 6600
tri 10056 6497 10159 6600 sw
tri 10294 6497 10397 6600 ne
rect 10397 6497 10606 6600
tri 10606 6497 10709 6600 sw
tri 10844 6497 10947 6600 ne
rect 10947 6497 11156 6600
tri 11156 6497 11259 6600 sw
tri 11394 6497 11497 6600 ne
rect 11497 6497 11706 6600
tri 11706 6497 11809 6600 sw
tri 11944 6497 12047 6600 ne
rect 12047 6497 12256 6600
tri 12256 6497 12359 6600 sw
tri 12494 6497 12597 6600 ne
rect 12597 6497 12806 6600
tri 12806 6497 12909 6600 sw
tri 13044 6497 13147 6600 ne
rect 13147 6497 13356 6600
tri 13356 6497 13459 6600 sw
tri 13594 6497 13697 6600 ne
rect 13697 6497 15775 6600
rect -1025 6360 -291 6497
tri -291 6360 -154 6497 sw
tri -53 6360 84 6497 ne
rect 84 6360 259 6497
tri 259 6360 396 6497 sw
tri 497 6360 634 6497 ne
rect 634 6360 809 6497
tri 809 6360 946 6497 sw
tri 1047 6360 1184 6497 ne
rect 1184 6360 1359 6497
tri 1359 6360 1496 6497 sw
tri 1597 6360 1734 6497 ne
rect 1734 6360 1909 6497
tri 1909 6360 2046 6497 sw
tri 2147 6360 2284 6497 ne
rect 2284 6360 2459 6497
tri 2459 6360 2596 6497 sw
tri 2697 6360 2834 6497 ne
rect 2834 6360 3009 6497
tri 3009 6360 3146 6497 sw
tri 3247 6360 3384 6497 ne
rect 3384 6360 3559 6497
tri 3559 6360 3696 6497 sw
tri 3797 6360 3934 6497 ne
rect 3934 6360 4109 6497
tri 4109 6360 4246 6497 sw
tri 4347 6360 4484 6497 ne
rect 4484 6360 4659 6497
tri 4659 6360 4796 6497 sw
tri 4897 6360 5034 6497 ne
rect 5034 6360 5209 6497
tri 5209 6360 5346 6497 sw
tri 5447 6360 5584 6497 ne
rect 5584 6360 5759 6497
tri 5759 6360 5896 6497 sw
tri 5997 6360 6134 6497 ne
rect 6134 6360 6309 6497
tri 6309 6360 6446 6497 sw
tri 6547 6360 6684 6497 ne
rect 6684 6360 6859 6497
tri 6859 6360 6996 6497 sw
tri 7097 6360 7234 6497 ne
rect 7234 6360 7409 6497
tri 7409 6360 7546 6497 sw
tri 7647 6360 7784 6497 ne
rect 7784 6360 7959 6497
tri 7959 6360 8096 6497 sw
tri 8197 6360 8334 6497 ne
rect 8334 6360 8509 6497
tri 8509 6360 8646 6497 sw
tri 8747 6360 8884 6497 ne
rect 8884 6360 9059 6497
tri 9059 6360 9196 6497 sw
tri 9297 6360 9434 6497 ne
rect 9434 6360 9609 6497
tri 9609 6360 9746 6497 sw
tri 9847 6360 9984 6497 ne
rect 9984 6360 10159 6497
tri 10159 6360 10296 6497 sw
tri 10397 6360 10534 6497 ne
rect 10534 6360 10709 6497
tri 10709 6360 10846 6497 sw
tri 10947 6360 11084 6497 ne
rect 11084 6360 11259 6497
tri 11259 6360 11396 6497 sw
tri 11497 6360 11634 6497 ne
rect 11634 6360 11809 6497
tri 11809 6360 11946 6497 sw
tri 12047 6360 12184 6497 ne
rect 12184 6360 12359 6497
tri 12359 6360 12496 6497 sw
tri 12597 6360 12734 6497 ne
rect 12734 6360 12909 6497
tri 12909 6360 13046 6497 sw
tri 13147 6360 13284 6497 ne
rect 13284 6360 13459 6497
tri 13459 6360 13596 6497 sw
rect -1025 6342 -310 6360
tri -448 6240 -346 6342 ne
rect -346 6240 -310 6342
rect -190 6240 -154 6360
rect -2525 6050 -447 6103
tri -447 6050 -394 6103 sw
tri -346 6050 -156 6240 ne
rect -156 6206 -154 6240
tri -154 6206 0 6360 sw
tri 84 6206 238 6360 ne
rect 238 6240 240 6360
rect 360 6240 396 6360
rect 238 6206 396 6240
tri 396 6206 550 6360 sw
tri 634 6206 788 6360 ne
rect 788 6240 790 6360
rect 910 6240 946 6360
rect 788 6206 946 6240
tri 946 6206 1100 6360 sw
tri 1184 6206 1338 6360 ne
rect 1338 6240 1340 6360
rect 1460 6240 1496 6360
rect 1338 6206 1496 6240
tri 1496 6206 1650 6360 sw
tri 1734 6206 1888 6360 ne
rect 1888 6240 1890 6360
rect 2010 6240 2046 6360
rect 1888 6206 2046 6240
tri 2046 6206 2200 6360 sw
tri 2284 6206 2438 6360 ne
rect 2438 6240 2440 6360
rect 2560 6240 2596 6360
rect 2438 6206 2596 6240
tri 2596 6206 2750 6360 sw
tri 2834 6206 2988 6360 ne
rect 2988 6240 2990 6360
rect 3110 6240 3146 6360
rect 2988 6206 3146 6240
tri 3146 6206 3300 6360 sw
tri 3384 6206 3538 6360 ne
rect 3538 6240 3540 6360
rect 3660 6240 3696 6360
rect 3538 6206 3696 6240
tri 3696 6206 3850 6360 sw
tri 3934 6206 4088 6360 ne
rect 4088 6240 4090 6360
rect 4210 6240 4246 6360
rect 4088 6206 4246 6240
tri 4246 6206 4400 6360 sw
tri 4484 6206 4638 6360 ne
rect 4638 6240 4640 6360
rect 4760 6240 4796 6360
rect 4638 6206 4796 6240
tri 4796 6206 4950 6360 sw
tri 5034 6206 5188 6360 ne
rect 5188 6240 5190 6360
rect 5310 6240 5346 6360
rect 5188 6206 5346 6240
tri 5346 6206 5500 6360 sw
tri 5584 6206 5738 6360 ne
rect 5738 6240 5740 6360
rect 5860 6240 5896 6360
rect 5738 6206 5896 6240
tri 5896 6206 6050 6360 sw
tri 6134 6206 6288 6360 ne
rect 6288 6240 6290 6360
rect 6410 6240 6446 6360
rect 6288 6206 6446 6240
tri 6446 6206 6600 6360 sw
tri 6684 6206 6838 6360 ne
rect 6838 6240 6840 6360
rect 6960 6240 6996 6360
rect 6838 6206 6996 6240
tri 6996 6206 7150 6360 sw
tri 7234 6206 7388 6360 ne
rect 7388 6240 7390 6360
rect 7510 6240 7546 6360
rect 7388 6206 7546 6240
tri 7546 6206 7700 6360 sw
tri 7784 6206 7938 6360 ne
rect 7938 6240 7940 6360
rect 8060 6240 8096 6360
rect 7938 6206 8096 6240
tri 8096 6206 8250 6360 sw
tri 8334 6206 8488 6360 ne
rect 8488 6240 8490 6360
rect 8610 6240 8646 6360
rect 8488 6206 8646 6240
tri 8646 6206 8800 6360 sw
tri 8884 6206 9038 6360 ne
rect 9038 6240 9040 6360
rect 9160 6240 9196 6360
rect 9038 6206 9196 6240
tri 9196 6206 9350 6360 sw
tri 9434 6206 9588 6360 ne
rect 9588 6240 9590 6360
rect 9710 6240 9746 6360
rect 9588 6206 9746 6240
tri 9746 6206 9900 6360 sw
tri 9984 6206 10138 6360 ne
rect 10138 6240 10140 6360
rect 10260 6240 10296 6360
rect 10138 6206 10296 6240
tri 10296 6206 10450 6360 sw
tri 10534 6206 10688 6360 ne
rect 10688 6240 10690 6360
rect 10810 6240 10846 6360
rect 10688 6206 10846 6240
tri 10846 6206 11000 6360 sw
tri 11084 6206 11238 6360 ne
rect 11238 6240 11240 6360
rect 11360 6240 11396 6360
rect 11238 6206 11396 6240
tri 11396 6206 11550 6360 sw
tri 11634 6206 11788 6360 ne
rect 11788 6240 11790 6360
rect 11910 6240 11946 6360
rect 11788 6206 11946 6240
tri 11946 6206 12100 6360 sw
tri 12184 6206 12338 6360 ne
rect 12338 6240 12340 6360
rect 12460 6240 12496 6360
rect 12338 6206 12496 6240
tri 12496 6206 12650 6360 sw
tri 12734 6206 12888 6360 ne
rect 12888 6240 12890 6360
rect 13010 6240 13046 6360
rect 12888 6206 13046 6240
tri 13046 6206 13200 6360 sw
tri 13284 6206 13438 6360 ne
rect 13438 6240 13440 6360
rect 13560 6258 13596 6360
tri 13596 6258 13698 6360 sw
rect 13560 6240 14275 6258
rect 13438 6206 14275 6240
rect -156 6050 0 6206
tri 0 6050 156 6206 sw
tri 238 6050 394 6206 ne
rect 394 6050 550 6206
tri 550 6050 706 6206 sw
tri 788 6050 944 6206 ne
rect 944 6050 1100 6206
tri 1100 6050 1256 6206 sw
tri 1338 6050 1494 6206 ne
rect 1494 6050 1650 6206
tri 1650 6050 1806 6206 sw
tri 1888 6050 2044 6206 ne
rect 2044 6050 2200 6206
tri 2200 6050 2356 6206 sw
tri 2438 6050 2594 6206 ne
rect 2594 6050 2750 6206
tri 2750 6050 2906 6206 sw
tri 2988 6050 3144 6206 ne
rect 3144 6050 3300 6206
tri 3300 6050 3456 6206 sw
tri 3538 6050 3694 6206 ne
rect 3694 6050 3850 6206
tri 3850 6050 4006 6206 sw
tri 4088 6050 4244 6206 ne
rect 4244 6050 4400 6206
tri 4400 6050 4556 6206 sw
tri 4638 6050 4794 6206 ne
rect 4794 6050 4950 6206
tri 4950 6050 5106 6206 sw
tri 5188 6050 5344 6206 ne
rect 5344 6050 5500 6206
tri 5500 6050 5656 6206 sw
tri 5738 6050 5894 6206 ne
rect 5894 6050 6050 6206
tri 6050 6050 6206 6206 sw
tri 6288 6050 6444 6206 ne
rect 6444 6050 6600 6206
tri 6600 6050 6756 6206 sw
tri 6838 6050 6994 6206 ne
rect 6994 6050 7150 6206
tri 7150 6050 7306 6206 sw
tri 7388 6050 7544 6206 ne
rect 7544 6050 7700 6206
tri 7700 6050 7856 6206 sw
tri 7938 6050 8094 6206 ne
rect 8094 6050 8250 6206
tri 8250 6050 8406 6206 sw
tri 8488 6050 8644 6206 ne
rect 8644 6050 8800 6206
tri 8800 6050 8956 6206 sw
tri 9038 6050 9194 6206 ne
rect 9194 6050 9350 6206
tri 9350 6050 9506 6206 sw
tri 9588 6050 9744 6206 ne
rect 9744 6050 9900 6206
tri 9900 6050 10056 6206 sw
tri 10138 6050 10294 6206 ne
rect 10294 6050 10450 6206
tri 10450 6050 10606 6206 sw
tri 10688 6050 10844 6206 ne
rect 10844 6050 11000 6206
tri 11000 6050 11156 6206 sw
tri 11238 6050 11394 6206 ne
rect 11394 6050 11550 6206
tri 11550 6050 11706 6206 sw
tri 11788 6050 11944 6206 ne
rect 11944 6050 12100 6206
tri 12100 6050 12256 6206 sw
tri 12338 6050 12494 6206 ne
rect 12494 6050 12650 6206
tri 12650 6050 12806 6206 sw
tri 12888 6050 13044 6206 ne
rect 13044 6050 13200 6206
tri 13200 6050 13356 6206 sw
tri 13438 6050 13594 6206 ne
rect 13594 6050 14275 6206
rect -2525 5947 -394 6050
tri -394 5947 -291 6050 sw
tri -156 5947 -53 6050 ne
rect -53 5947 156 6050
tri 156 5947 259 6050 sw
tri 394 5947 497 6050 ne
rect 497 5947 706 6050
tri 706 5947 809 6050 sw
tri 944 5947 1047 6050 ne
rect 1047 5947 1256 6050
tri 1256 5947 1359 6050 sw
tri 1494 5947 1597 6050 ne
rect 1597 5947 1806 6050
tri 1806 5947 1909 6050 sw
tri 2044 5947 2147 6050 ne
rect 2147 5947 2356 6050
tri 2356 5947 2459 6050 sw
tri 2594 5947 2697 6050 ne
rect 2697 5947 2906 6050
tri 2906 5947 3009 6050 sw
tri 3144 5947 3247 6050 ne
rect 3247 5947 3456 6050
tri 3456 5947 3559 6050 sw
tri 3694 5947 3797 6050 ne
rect 3797 5947 4006 6050
tri 4006 5947 4109 6050 sw
tri 4244 5947 4347 6050 ne
rect 4347 5947 4556 6050
tri 4556 5947 4659 6050 sw
tri 4794 5947 4897 6050 ne
rect 4897 5947 5106 6050
tri 5106 5947 5209 6050 sw
tri 5344 5947 5447 6050 ne
rect 5447 5947 5656 6050
tri 5656 5947 5759 6050 sw
tri 5894 5947 5997 6050 ne
rect 5997 5947 6206 6050
tri 6206 5947 6309 6050 sw
tri 6444 5947 6547 6050 ne
rect 6547 5947 6756 6050
tri 6756 5947 6859 6050 sw
tri 6994 5947 7097 6050 ne
rect 7097 5947 7306 6050
tri 7306 5947 7409 6050 sw
tri 7544 5947 7647 6050 ne
rect 7647 5947 7856 6050
tri 7856 5947 7959 6050 sw
tri 8094 5947 8197 6050 ne
rect 8197 5947 8406 6050
tri 8406 5947 8509 6050 sw
tri 8644 5947 8747 6050 ne
rect 8747 5947 8956 6050
tri 8956 5947 9059 6050 sw
tri 9194 5947 9297 6050 ne
rect 9297 5947 9506 6050
tri 9506 5947 9609 6050 sw
tri 9744 5947 9847 6050 ne
rect 9847 5947 10056 6050
tri 10056 5947 10159 6050 sw
tri 10294 5947 10397 6050 ne
rect 10397 5947 10606 6050
tri 10606 5947 10709 6050 sw
tri 10844 5947 10947 6050 ne
rect 10947 5947 11156 6050
tri 11156 5947 11259 6050 sw
tri 11394 5947 11497 6050 ne
rect 11497 5947 11706 6050
tri 11706 5947 11809 6050 sw
tri 11944 5947 12047 6050 ne
rect 12047 5947 12256 6050
tri 12256 5947 12359 6050 sw
tri 12494 5947 12597 6050 ne
rect 12597 5947 12806 6050
tri 12806 5947 12909 6050 sw
tri 13044 5947 13147 6050 ne
rect 13147 5947 13356 6050
tri 13356 5947 13459 6050 sw
tri 13594 5947 13697 6050 ne
rect 13697 5947 14275 6050
rect -2525 5810 -291 5947
tri -291 5810 -154 5947 sw
tri -53 5810 84 5947 ne
rect 84 5810 259 5947
tri 259 5810 396 5947 sw
tri 497 5810 634 5947 ne
rect 634 5810 809 5947
tri 809 5810 946 5947 sw
tri 1047 5810 1184 5947 ne
rect 1184 5810 1359 5947
tri 1359 5810 1496 5947 sw
tri 1597 5810 1734 5947 ne
rect 1734 5810 1909 5947
tri 1909 5810 2046 5947 sw
tri 2147 5810 2284 5947 ne
rect 2284 5810 2459 5947
tri 2459 5810 2596 5947 sw
tri 2697 5810 2834 5947 ne
rect 2834 5810 3009 5947
tri 3009 5810 3146 5947 sw
tri 3247 5810 3384 5947 ne
rect 3384 5810 3559 5947
tri 3559 5810 3696 5947 sw
tri 3797 5810 3934 5947 ne
rect 3934 5810 4109 5947
tri 4109 5810 4246 5947 sw
tri 4347 5810 4484 5947 ne
rect 4484 5810 4659 5947
tri 4659 5810 4796 5947 sw
tri 4897 5810 5034 5947 ne
rect 5034 5810 5209 5947
tri 5209 5810 5346 5947 sw
tri 5447 5810 5584 5947 ne
rect 5584 5810 5759 5947
tri 5759 5810 5896 5947 sw
tri 5997 5810 6134 5947 ne
rect 6134 5810 6309 5947
tri 6309 5810 6446 5947 sw
tri 6547 5810 6684 5947 ne
rect 6684 5810 6859 5947
tri 6859 5810 6996 5947 sw
tri 7097 5810 7234 5947 ne
rect 7234 5810 7409 5947
tri 7409 5810 7546 5947 sw
tri 7647 5810 7784 5947 ne
rect 7784 5810 7959 5947
tri 7959 5810 8096 5947 sw
tri 8197 5810 8334 5947 ne
rect 8334 5810 8509 5947
tri 8509 5810 8646 5947 sw
tri 8747 5810 8884 5947 ne
rect 8884 5810 9059 5947
tri 9059 5810 9196 5947 sw
tri 9297 5810 9434 5947 ne
rect 9434 5810 9609 5947
tri 9609 5810 9746 5947 sw
tri 9847 5810 9984 5947 ne
rect 9984 5810 10159 5947
tri 10159 5810 10296 5947 sw
tri 10397 5810 10534 5947 ne
rect 10534 5810 10709 5947
tri 10709 5810 10846 5947 sw
tri 10947 5810 11084 5947 ne
rect 11084 5810 11259 5947
tri 11259 5810 11396 5947 sw
tri 11497 5810 11634 5947 ne
rect 11634 5810 11809 5947
tri 11809 5810 11946 5947 sw
tri 12047 5810 12184 5947 ne
rect 12184 5810 12359 5947
tri 12359 5810 12496 5947 sw
tri 12597 5810 12734 5947 ne
rect 12734 5810 12909 5947
tri 12909 5810 13046 5947 sw
tri 13147 5810 13284 5947 ne
rect 13284 5810 13459 5947
tri 13459 5810 13596 5947 sw
rect -2525 5792 -310 5810
rect -2525 5003 -1525 5792
tri -448 5690 -346 5792 ne
rect -346 5690 -310 5792
rect -190 5690 -154 5810
rect -1025 5500 -447 5553
tri -447 5500 -394 5553 sw
tri -346 5500 -156 5690 ne
rect -156 5656 -154 5690
tri -154 5656 0 5810 sw
tri 84 5656 238 5810 ne
rect 238 5690 240 5810
rect 360 5690 396 5810
rect 238 5656 396 5690
tri 396 5656 550 5810 sw
tri 634 5656 788 5810 ne
rect 788 5690 790 5810
rect 910 5690 946 5810
rect 788 5656 946 5690
tri 946 5656 1100 5810 sw
tri 1184 5656 1338 5810 ne
rect 1338 5690 1340 5810
rect 1460 5690 1496 5810
rect 1338 5656 1496 5690
tri 1496 5656 1650 5810 sw
tri 1734 5656 1888 5810 ne
rect 1888 5690 1890 5810
rect 2010 5690 2046 5810
rect 1888 5656 2046 5690
tri 2046 5656 2200 5810 sw
tri 2284 5656 2438 5810 ne
rect 2438 5690 2440 5810
rect 2560 5690 2596 5810
rect 2438 5656 2596 5690
tri 2596 5656 2750 5810 sw
tri 2834 5656 2988 5810 ne
rect 2988 5690 2990 5810
rect 3110 5690 3146 5810
rect 2988 5656 3146 5690
tri 3146 5656 3300 5810 sw
tri 3384 5656 3538 5810 ne
rect 3538 5690 3540 5810
rect 3660 5690 3696 5810
rect 3538 5656 3696 5690
tri 3696 5656 3850 5810 sw
tri 3934 5656 4088 5810 ne
rect 4088 5690 4090 5810
rect 4210 5690 4246 5810
rect 4088 5656 4246 5690
tri 4246 5656 4400 5810 sw
tri 4484 5656 4638 5810 ne
rect 4638 5690 4640 5810
rect 4760 5690 4796 5810
rect 4638 5656 4796 5690
tri 4796 5656 4950 5810 sw
tri 5034 5656 5188 5810 ne
rect 5188 5690 5190 5810
rect 5310 5690 5346 5810
rect 5188 5656 5346 5690
tri 5346 5656 5500 5810 sw
tri 5584 5656 5738 5810 ne
rect 5738 5690 5740 5810
rect 5860 5690 5896 5810
rect 5738 5656 5896 5690
tri 5896 5656 6050 5810 sw
tri 6134 5656 6288 5810 ne
rect 6288 5690 6290 5810
rect 6410 5690 6446 5810
rect 6288 5656 6446 5690
tri 6446 5656 6600 5810 sw
tri 6684 5656 6838 5810 ne
rect 6838 5690 6840 5810
rect 6960 5690 6996 5810
rect 6838 5656 6996 5690
tri 6996 5656 7150 5810 sw
tri 7234 5656 7388 5810 ne
rect 7388 5690 7390 5810
rect 7510 5690 7546 5810
rect 7388 5656 7546 5690
tri 7546 5656 7700 5810 sw
tri 7784 5656 7938 5810 ne
rect 7938 5690 7940 5810
rect 8060 5690 8096 5810
rect 7938 5656 8096 5690
tri 8096 5656 8250 5810 sw
tri 8334 5656 8488 5810 ne
rect 8488 5690 8490 5810
rect 8610 5690 8646 5810
rect 8488 5656 8646 5690
tri 8646 5656 8800 5810 sw
tri 8884 5656 9038 5810 ne
rect 9038 5690 9040 5810
rect 9160 5690 9196 5810
rect 9038 5656 9196 5690
tri 9196 5656 9350 5810 sw
tri 9434 5656 9588 5810 ne
rect 9588 5690 9590 5810
rect 9710 5690 9746 5810
rect 9588 5656 9746 5690
tri 9746 5656 9900 5810 sw
tri 9984 5656 10138 5810 ne
rect 10138 5690 10140 5810
rect 10260 5690 10296 5810
rect 10138 5656 10296 5690
tri 10296 5656 10450 5810 sw
tri 10534 5656 10688 5810 ne
rect 10688 5690 10690 5810
rect 10810 5690 10846 5810
rect 10688 5656 10846 5690
tri 10846 5656 11000 5810 sw
tri 11084 5656 11238 5810 ne
rect 11238 5690 11240 5810
rect 11360 5690 11396 5810
rect 11238 5656 11396 5690
tri 11396 5656 11550 5810 sw
tri 11634 5656 11788 5810 ne
rect 11788 5690 11790 5810
rect 11910 5690 11946 5810
rect 11788 5656 11946 5690
tri 11946 5656 12100 5810 sw
tri 12184 5656 12338 5810 ne
rect 12338 5690 12340 5810
rect 12460 5690 12496 5810
rect 12338 5656 12496 5690
tri 12496 5656 12650 5810 sw
tri 12734 5656 12888 5810 ne
rect 12888 5690 12890 5810
rect 13010 5690 13046 5810
rect 12888 5656 13046 5690
tri 13046 5656 13200 5810 sw
tri 13284 5656 13438 5810 ne
rect 13438 5690 13440 5810
rect 13560 5708 13596 5810
tri 13596 5708 13698 5810 sw
rect 14775 5708 15775 6497
rect 13560 5690 15775 5708
rect 13438 5656 15775 5690
rect -156 5500 0 5656
tri 0 5500 156 5656 sw
tri 238 5500 394 5656 ne
rect 394 5500 550 5656
tri 550 5500 706 5656 sw
tri 788 5500 944 5656 ne
rect 944 5500 1100 5656
tri 1100 5500 1256 5656 sw
tri 1338 5500 1494 5656 ne
rect 1494 5500 1650 5656
tri 1650 5500 1806 5656 sw
tri 1888 5500 2044 5656 ne
rect 2044 5500 2200 5656
tri 2200 5500 2356 5656 sw
tri 2438 5500 2594 5656 ne
rect 2594 5500 2750 5656
tri 2750 5500 2906 5656 sw
tri 2988 5500 3144 5656 ne
rect 3144 5500 3300 5656
tri 3300 5500 3456 5656 sw
tri 3538 5500 3694 5656 ne
rect 3694 5500 3850 5656
tri 3850 5500 4006 5656 sw
tri 4088 5500 4244 5656 ne
rect 4244 5500 4400 5656
tri 4400 5500 4556 5656 sw
tri 4638 5500 4794 5656 ne
rect 4794 5500 4950 5656
tri 4950 5500 5106 5656 sw
tri 5188 5500 5344 5656 ne
rect 5344 5500 5500 5656
tri 5500 5500 5656 5656 sw
tri 5738 5500 5894 5656 ne
rect 5894 5500 6050 5656
tri 6050 5500 6206 5656 sw
tri 6288 5500 6444 5656 ne
rect 6444 5500 6600 5656
tri 6600 5500 6756 5656 sw
tri 6838 5500 6994 5656 ne
rect 6994 5500 7150 5656
tri 7150 5500 7306 5656 sw
tri 7388 5500 7544 5656 ne
rect 7544 5500 7700 5656
tri 7700 5500 7856 5656 sw
tri 7938 5500 8094 5656 ne
rect 8094 5500 8250 5656
tri 8250 5500 8406 5656 sw
tri 8488 5500 8644 5656 ne
rect 8644 5500 8800 5656
tri 8800 5500 8956 5656 sw
tri 9038 5500 9194 5656 ne
rect 9194 5500 9350 5656
tri 9350 5500 9506 5656 sw
tri 9588 5500 9744 5656 ne
rect 9744 5500 9900 5656
tri 9900 5500 10056 5656 sw
tri 10138 5500 10294 5656 ne
rect 10294 5500 10450 5656
tri 10450 5500 10606 5656 sw
tri 10688 5500 10844 5656 ne
rect 10844 5500 11000 5656
tri 11000 5500 11156 5656 sw
tri 11238 5500 11394 5656 ne
rect 11394 5500 11550 5656
tri 11550 5500 11706 5656 sw
tri 11788 5500 11944 5656 ne
rect 11944 5500 12100 5656
tri 12100 5500 12256 5656 sw
tri 12338 5500 12494 5656 ne
rect 12494 5500 12650 5656
tri 12650 5500 12806 5656 sw
tri 12888 5500 13044 5656 ne
rect 13044 5500 13200 5656
tri 13200 5500 13356 5656 sw
tri 13438 5500 13594 5656 ne
rect 13594 5500 15775 5656
rect -1025 5397 -394 5500
tri -394 5397 -291 5500 sw
tri -156 5397 -53 5500 ne
rect -53 5397 156 5500
tri 156 5397 259 5500 sw
tri 394 5397 497 5500 ne
rect 497 5397 706 5500
tri 706 5397 809 5500 sw
tri 944 5397 1047 5500 ne
rect 1047 5397 1256 5500
tri 1256 5397 1359 5500 sw
tri 1494 5397 1597 5500 ne
rect 1597 5397 1806 5500
tri 1806 5397 1909 5500 sw
tri 2044 5397 2147 5500 ne
rect 2147 5397 2356 5500
tri 2356 5397 2459 5500 sw
tri 2594 5397 2697 5500 ne
rect 2697 5397 2906 5500
tri 2906 5397 3009 5500 sw
tri 3144 5397 3247 5500 ne
rect 3247 5397 3456 5500
tri 3456 5397 3559 5500 sw
tri 3694 5397 3797 5500 ne
rect 3797 5397 4006 5500
tri 4006 5397 4109 5500 sw
tri 4244 5397 4347 5500 ne
rect 4347 5397 4556 5500
tri 4556 5397 4659 5500 sw
tri 4794 5397 4897 5500 ne
rect 4897 5397 5106 5500
tri 5106 5397 5209 5500 sw
tri 5344 5397 5447 5500 ne
rect 5447 5397 5656 5500
tri 5656 5397 5759 5500 sw
tri 5894 5397 5997 5500 ne
rect 5997 5397 6206 5500
tri 6206 5397 6309 5500 sw
tri 6444 5397 6547 5500 ne
rect 6547 5397 6756 5500
tri 6756 5397 6859 5500 sw
tri 6994 5397 7097 5500 ne
rect 7097 5397 7306 5500
tri 7306 5397 7409 5500 sw
tri 7544 5397 7647 5500 ne
rect 7647 5397 7856 5500
tri 7856 5397 7959 5500 sw
tri 8094 5397 8197 5500 ne
rect 8197 5397 8406 5500
tri 8406 5397 8509 5500 sw
tri 8644 5397 8747 5500 ne
rect 8747 5397 8956 5500
tri 8956 5397 9059 5500 sw
tri 9194 5397 9297 5500 ne
rect 9297 5397 9506 5500
tri 9506 5397 9609 5500 sw
tri 9744 5397 9847 5500 ne
rect 9847 5397 10056 5500
tri 10056 5397 10159 5500 sw
tri 10294 5397 10397 5500 ne
rect 10397 5397 10606 5500
tri 10606 5397 10709 5500 sw
tri 10844 5397 10947 5500 ne
rect 10947 5397 11156 5500
tri 11156 5397 11259 5500 sw
tri 11394 5397 11497 5500 ne
rect 11497 5397 11706 5500
tri 11706 5397 11809 5500 sw
tri 11944 5397 12047 5500 ne
rect 12047 5397 12256 5500
tri 12256 5397 12359 5500 sw
tri 12494 5397 12597 5500 ne
rect 12597 5397 12806 5500
tri 12806 5397 12909 5500 sw
tri 13044 5397 13147 5500 ne
rect 13147 5397 13356 5500
tri 13356 5397 13459 5500 sw
tri 13594 5397 13697 5500 ne
rect 13697 5397 15775 5500
rect -1025 5260 -291 5397
tri -291 5260 -154 5397 sw
tri -53 5260 84 5397 ne
rect 84 5260 259 5397
tri 259 5260 396 5397 sw
tri 497 5260 634 5397 ne
rect 634 5260 809 5397
tri 809 5260 946 5397 sw
tri 1047 5260 1184 5397 ne
rect 1184 5260 1359 5397
tri 1359 5260 1496 5397 sw
tri 1597 5260 1734 5397 ne
rect 1734 5260 1909 5397
tri 1909 5260 2046 5397 sw
tri 2147 5260 2284 5397 ne
rect 2284 5260 2459 5397
tri 2459 5260 2596 5397 sw
tri 2697 5260 2834 5397 ne
rect 2834 5260 3009 5397
tri 3009 5260 3146 5397 sw
tri 3247 5260 3384 5397 ne
rect 3384 5260 3559 5397
tri 3559 5260 3696 5397 sw
tri 3797 5260 3934 5397 ne
rect 3934 5260 4109 5397
tri 4109 5260 4246 5397 sw
tri 4347 5260 4484 5397 ne
rect 4484 5260 4659 5397
tri 4659 5260 4796 5397 sw
tri 4897 5260 5034 5397 ne
rect 5034 5260 5209 5397
tri 5209 5260 5346 5397 sw
tri 5447 5260 5584 5397 ne
rect 5584 5260 5759 5397
tri 5759 5260 5896 5397 sw
tri 5997 5260 6134 5397 ne
rect 6134 5260 6309 5397
tri 6309 5260 6446 5397 sw
tri 6547 5260 6684 5397 ne
rect 6684 5260 6859 5397
tri 6859 5260 6996 5397 sw
tri 7097 5260 7234 5397 ne
rect 7234 5260 7409 5397
tri 7409 5260 7546 5397 sw
tri 7647 5260 7784 5397 ne
rect 7784 5260 7959 5397
tri 7959 5260 8096 5397 sw
tri 8197 5260 8334 5397 ne
rect 8334 5260 8509 5397
tri 8509 5260 8646 5397 sw
tri 8747 5260 8884 5397 ne
rect 8884 5260 9059 5397
tri 9059 5260 9196 5397 sw
tri 9297 5260 9434 5397 ne
rect 9434 5260 9609 5397
tri 9609 5260 9746 5397 sw
tri 9847 5260 9984 5397 ne
rect 9984 5260 10159 5397
tri 10159 5260 10296 5397 sw
tri 10397 5260 10534 5397 ne
rect 10534 5260 10709 5397
tri 10709 5260 10846 5397 sw
tri 10947 5260 11084 5397 ne
rect 11084 5260 11259 5397
tri 11259 5260 11396 5397 sw
tri 11497 5260 11634 5397 ne
rect 11634 5260 11809 5397
tri 11809 5260 11946 5397 sw
tri 12047 5260 12184 5397 ne
rect 12184 5260 12359 5397
tri 12359 5260 12496 5397 sw
tri 12597 5260 12734 5397 ne
rect 12734 5260 12909 5397
tri 12909 5260 13046 5397 sw
tri 13147 5260 13284 5397 ne
rect 13284 5260 13459 5397
tri 13459 5260 13596 5397 sw
rect -1025 5242 -310 5260
tri -448 5140 -346 5242 ne
rect -346 5140 -310 5242
rect -190 5140 -154 5260
rect -2525 4950 -447 5003
tri -447 4950 -394 5003 sw
tri -346 4950 -156 5140 ne
rect -156 5106 -154 5140
tri -154 5106 0 5260 sw
tri 84 5106 238 5260 ne
rect 238 5140 240 5260
rect 360 5140 396 5260
rect 238 5106 396 5140
tri 396 5106 550 5260 sw
tri 634 5106 788 5260 ne
rect 788 5140 790 5260
rect 910 5140 946 5260
rect 788 5106 946 5140
tri 946 5106 1100 5260 sw
tri 1184 5106 1338 5260 ne
rect 1338 5140 1340 5260
rect 1460 5140 1496 5260
rect 1338 5106 1496 5140
tri 1496 5106 1650 5260 sw
tri 1734 5106 1888 5260 ne
rect 1888 5140 1890 5260
rect 2010 5140 2046 5260
rect 1888 5106 2046 5140
tri 2046 5106 2200 5260 sw
tri 2284 5106 2438 5260 ne
rect 2438 5140 2440 5260
rect 2560 5140 2596 5260
rect 2438 5106 2596 5140
tri 2596 5106 2750 5260 sw
tri 2834 5106 2988 5260 ne
rect 2988 5140 2990 5260
rect 3110 5140 3146 5260
rect 2988 5106 3146 5140
tri 3146 5106 3300 5260 sw
tri 3384 5106 3538 5260 ne
rect 3538 5140 3540 5260
rect 3660 5140 3696 5260
rect 3538 5106 3696 5140
tri 3696 5106 3850 5260 sw
tri 3934 5106 4088 5260 ne
rect 4088 5140 4090 5260
rect 4210 5140 4246 5260
rect 4088 5106 4246 5140
tri 4246 5106 4400 5260 sw
tri 4484 5106 4638 5260 ne
rect 4638 5140 4640 5260
rect 4760 5140 4796 5260
rect 4638 5106 4796 5140
tri 4796 5106 4950 5260 sw
tri 5034 5106 5188 5260 ne
rect 5188 5140 5190 5260
rect 5310 5140 5346 5260
rect 5188 5106 5346 5140
tri 5346 5106 5500 5260 sw
tri 5584 5106 5738 5260 ne
rect 5738 5140 5740 5260
rect 5860 5140 5896 5260
rect 5738 5106 5896 5140
tri 5896 5106 6050 5260 sw
tri 6134 5106 6288 5260 ne
rect 6288 5140 6290 5260
rect 6410 5140 6446 5260
rect 6288 5106 6446 5140
tri 6446 5106 6600 5260 sw
tri 6684 5106 6838 5260 ne
rect 6838 5140 6840 5260
rect 6960 5140 6996 5260
rect 6838 5106 6996 5140
tri 6996 5106 7150 5260 sw
tri 7234 5106 7388 5260 ne
rect 7388 5140 7390 5260
rect 7510 5140 7546 5260
rect 7388 5106 7546 5140
tri 7546 5106 7700 5260 sw
tri 7784 5106 7938 5260 ne
rect 7938 5140 7940 5260
rect 8060 5140 8096 5260
rect 7938 5106 8096 5140
tri 8096 5106 8250 5260 sw
tri 8334 5106 8488 5260 ne
rect 8488 5140 8490 5260
rect 8610 5140 8646 5260
rect 8488 5106 8646 5140
tri 8646 5106 8800 5260 sw
tri 8884 5106 9038 5260 ne
rect 9038 5140 9040 5260
rect 9160 5140 9196 5260
rect 9038 5106 9196 5140
tri 9196 5106 9350 5260 sw
tri 9434 5106 9588 5260 ne
rect 9588 5140 9590 5260
rect 9710 5140 9746 5260
rect 9588 5106 9746 5140
tri 9746 5106 9900 5260 sw
tri 9984 5106 10138 5260 ne
rect 10138 5140 10140 5260
rect 10260 5140 10296 5260
rect 10138 5106 10296 5140
tri 10296 5106 10450 5260 sw
tri 10534 5106 10688 5260 ne
rect 10688 5140 10690 5260
rect 10810 5140 10846 5260
rect 10688 5106 10846 5140
tri 10846 5106 11000 5260 sw
tri 11084 5106 11238 5260 ne
rect 11238 5140 11240 5260
rect 11360 5140 11396 5260
rect 11238 5106 11396 5140
tri 11396 5106 11550 5260 sw
tri 11634 5106 11788 5260 ne
rect 11788 5140 11790 5260
rect 11910 5140 11946 5260
rect 11788 5106 11946 5140
tri 11946 5106 12100 5260 sw
tri 12184 5106 12338 5260 ne
rect 12338 5140 12340 5260
rect 12460 5140 12496 5260
rect 12338 5106 12496 5140
tri 12496 5106 12650 5260 sw
tri 12734 5106 12888 5260 ne
rect 12888 5140 12890 5260
rect 13010 5140 13046 5260
rect 12888 5106 13046 5140
tri 13046 5106 13200 5260 sw
tri 13284 5106 13438 5260 ne
rect 13438 5140 13440 5260
rect 13560 5158 13596 5260
tri 13596 5158 13698 5260 sw
rect 13560 5140 14275 5158
rect 13438 5106 14275 5140
rect -156 4950 0 5106
tri 0 4950 156 5106 sw
tri 238 4950 394 5106 ne
rect 394 4950 550 5106
tri 550 4950 706 5106 sw
tri 788 4950 944 5106 ne
rect 944 4950 1100 5106
tri 1100 4950 1256 5106 sw
tri 1338 4950 1494 5106 ne
rect 1494 4950 1650 5106
tri 1650 4950 1806 5106 sw
tri 1888 4950 2044 5106 ne
rect 2044 4950 2200 5106
tri 2200 4950 2356 5106 sw
tri 2438 4950 2594 5106 ne
rect 2594 4950 2750 5106
tri 2750 4950 2906 5106 sw
tri 2988 4950 3144 5106 ne
rect 3144 4950 3300 5106
tri 3300 4950 3456 5106 sw
tri 3538 4950 3694 5106 ne
rect 3694 4950 3850 5106
tri 3850 4950 4006 5106 sw
tri 4088 4950 4244 5106 ne
rect 4244 4950 4400 5106
tri 4400 4950 4556 5106 sw
tri 4638 4950 4794 5106 ne
rect 4794 4950 4950 5106
tri 4950 4950 5106 5106 sw
tri 5188 4950 5344 5106 ne
rect 5344 4950 5500 5106
tri 5500 4950 5656 5106 sw
tri 5738 4950 5894 5106 ne
rect 5894 4950 6050 5106
tri 6050 4950 6206 5106 sw
tri 6288 4950 6444 5106 ne
rect 6444 4950 6600 5106
tri 6600 4950 6756 5106 sw
tri 6838 4950 6994 5106 ne
rect 6994 4950 7150 5106
tri 7150 4950 7306 5106 sw
tri 7388 4950 7544 5106 ne
rect 7544 4950 7700 5106
tri 7700 4950 7856 5106 sw
tri 7938 4950 8094 5106 ne
rect 8094 4950 8250 5106
tri 8250 4950 8406 5106 sw
tri 8488 4950 8644 5106 ne
rect 8644 4950 8800 5106
tri 8800 4950 8956 5106 sw
tri 9038 4950 9194 5106 ne
rect 9194 4950 9350 5106
tri 9350 4950 9506 5106 sw
tri 9588 4950 9744 5106 ne
rect 9744 4950 9900 5106
tri 9900 4950 10056 5106 sw
tri 10138 4950 10294 5106 ne
rect 10294 4950 10450 5106
tri 10450 4950 10606 5106 sw
tri 10688 4950 10844 5106 ne
rect 10844 4950 11000 5106
tri 11000 4950 11156 5106 sw
tri 11238 4950 11394 5106 ne
rect 11394 4950 11550 5106
tri 11550 4950 11706 5106 sw
tri 11788 4950 11944 5106 ne
rect 11944 4950 12100 5106
tri 12100 4950 12256 5106 sw
tri 12338 4950 12494 5106 ne
rect 12494 4950 12650 5106
tri 12650 4950 12806 5106 sw
tri 12888 4950 13044 5106 ne
rect 13044 4950 13200 5106
tri 13200 4950 13356 5106 sw
tri 13438 4950 13594 5106 ne
rect 13594 4950 14275 5106
rect -2525 4847 -394 4950
tri -394 4847 -291 4950 sw
tri -156 4847 -53 4950 ne
rect -53 4847 156 4950
tri 156 4847 259 4950 sw
tri 394 4847 497 4950 ne
rect 497 4847 706 4950
tri 706 4847 809 4950 sw
tri 944 4847 1047 4950 ne
rect 1047 4847 1256 4950
tri 1256 4847 1359 4950 sw
tri 1494 4847 1597 4950 ne
rect 1597 4847 1806 4950
tri 1806 4847 1909 4950 sw
tri 2044 4847 2147 4950 ne
rect 2147 4847 2356 4950
tri 2356 4847 2459 4950 sw
tri 2594 4847 2697 4950 ne
rect 2697 4847 2906 4950
tri 2906 4847 3009 4950 sw
tri 3144 4847 3247 4950 ne
rect 3247 4847 3456 4950
tri 3456 4847 3559 4950 sw
tri 3694 4847 3797 4950 ne
rect 3797 4847 4006 4950
tri 4006 4847 4109 4950 sw
tri 4244 4847 4347 4950 ne
rect 4347 4847 4556 4950
tri 4556 4847 4659 4950 sw
tri 4794 4847 4897 4950 ne
rect 4897 4847 5106 4950
tri 5106 4847 5209 4950 sw
tri 5344 4847 5447 4950 ne
rect 5447 4847 5656 4950
tri 5656 4847 5759 4950 sw
tri 5894 4847 5997 4950 ne
rect 5997 4847 6206 4950
tri 6206 4847 6309 4950 sw
tri 6444 4847 6547 4950 ne
rect 6547 4847 6756 4950
tri 6756 4847 6859 4950 sw
tri 6994 4847 7097 4950 ne
rect 7097 4847 7306 4950
tri 7306 4847 7409 4950 sw
tri 7544 4847 7647 4950 ne
rect 7647 4847 7856 4950
tri 7856 4847 7959 4950 sw
tri 8094 4847 8197 4950 ne
rect 8197 4847 8406 4950
tri 8406 4847 8509 4950 sw
tri 8644 4847 8747 4950 ne
rect 8747 4847 8956 4950
tri 8956 4847 9059 4950 sw
tri 9194 4847 9297 4950 ne
rect 9297 4847 9506 4950
tri 9506 4847 9609 4950 sw
tri 9744 4847 9847 4950 ne
rect 9847 4847 10056 4950
tri 10056 4847 10159 4950 sw
tri 10294 4847 10397 4950 ne
rect 10397 4847 10606 4950
tri 10606 4847 10709 4950 sw
tri 10844 4847 10947 4950 ne
rect 10947 4847 11156 4950
tri 11156 4847 11259 4950 sw
tri 11394 4847 11497 4950 ne
rect 11497 4847 11706 4950
tri 11706 4847 11809 4950 sw
tri 11944 4847 12047 4950 ne
rect 12047 4847 12256 4950
tri 12256 4847 12359 4950 sw
tri 12494 4847 12597 4950 ne
rect 12597 4847 12806 4950
tri 12806 4847 12909 4950 sw
tri 13044 4847 13147 4950 ne
rect 13147 4847 13356 4950
tri 13356 4847 13459 4950 sw
tri 13594 4847 13697 4950 ne
rect 13697 4847 14275 4950
rect -2525 4710 -291 4847
tri -291 4710 -154 4847 sw
tri -53 4710 84 4847 ne
rect 84 4710 259 4847
tri 259 4710 396 4847 sw
tri 497 4710 634 4847 ne
rect 634 4710 809 4847
tri 809 4710 946 4847 sw
tri 1047 4710 1184 4847 ne
rect 1184 4710 1359 4847
tri 1359 4710 1496 4847 sw
tri 1597 4710 1734 4847 ne
rect 1734 4710 1909 4847
tri 1909 4710 2046 4847 sw
tri 2147 4710 2284 4847 ne
rect 2284 4710 2459 4847
tri 2459 4710 2596 4847 sw
tri 2697 4710 2834 4847 ne
rect 2834 4710 3009 4847
tri 3009 4710 3146 4847 sw
tri 3247 4710 3384 4847 ne
rect 3384 4710 3559 4847
tri 3559 4710 3696 4847 sw
tri 3797 4710 3934 4847 ne
rect 3934 4710 4109 4847
tri 4109 4710 4246 4847 sw
tri 4347 4710 4484 4847 ne
rect 4484 4710 4659 4847
tri 4659 4710 4796 4847 sw
tri 4897 4710 5034 4847 ne
rect 5034 4710 5209 4847
tri 5209 4710 5346 4847 sw
tri 5447 4710 5584 4847 ne
rect 5584 4710 5759 4847
tri 5759 4710 5896 4847 sw
tri 5997 4710 6134 4847 ne
rect 6134 4710 6309 4847
tri 6309 4710 6446 4847 sw
tri 6547 4710 6684 4847 ne
rect 6684 4710 6859 4847
tri 6859 4710 6996 4847 sw
tri 7097 4710 7234 4847 ne
rect 7234 4710 7409 4847
tri 7409 4710 7546 4847 sw
tri 7647 4710 7784 4847 ne
rect 7784 4710 7959 4847
tri 7959 4710 8096 4847 sw
tri 8197 4710 8334 4847 ne
rect 8334 4710 8509 4847
tri 8509 4710 8646 4847 sw
tri 8747 4710 8884 4847 ne
rect 8884 4710 9059 4847
tri 9059 4710 9196 4847 sw
tri 9297 4710 9434 4847 ne
rect 9434 4710 9609 4847
tri 9609 4710 9746 4847 sw
tri 9847 4710 9984 4847 ne
rect 9984 4710 10159 4847
tri 10159 4710 10296 4847 sw
tri 10397 4710 10534 4847 ne
rect 10534 4710 10709 4847
tri 10709 4710 10846 4847 sw
tri 10947 4710 11084 4847 ne
rect 11084 4710 11259 4847
tri 11259 4710 11396 4847 sw
tri 11497 4710 11634 4847 ne
rect 11634 4710 11809 4847
tri 11809 4710 11946 4847 sw
tri 12047 4710 12184 4847 ne
rect 12184 4710 12359 4847
tri 12359 4710 12496 4847 sw
tri 12597 4710 12734 4847 ne
rect 12734 4710 12909 4847
tri 12909 4710 13046 4847 sw
tri 13147 4710 13284 4847 ne
rect 13284 4710 13459 4847
tri 13459 4710 13596 4847 sw
rect -2525 4692 -310 4710
rect -2525 3903 -1525 4692
tri -448 4590 -346 4692 ne
rect -346 4590 -310 4692
rect -190 4590 -154 4710
rect -1025 4400 -447 4453
tri -447 4400 -394 4453 sw
tri -346 4400 -156 4590 ne
rect -156 4556 -154 4590
tri -154 4556 0 4710 sw
tri 84 4556 238 4710 ne
rect 238 4590 240 4710
rect 360 4590 396 4710
rect 238 4556 396 4590
tri 396 4556 550 4710 sw
tri 634 4556 788 4710 ne
rect 788 4590 790 4710
rect 910 4590 946 4710
rect 788 4556 946 4590
tri 946 4556 1100 4710 sw
tri 1184 4556 1338 4710 ne
rect 1338 4590 1340 4710
rect 1460 4590 1496 4710
rect 1338 4556 1496 4590
tri 1496 4556 1650 4710 sw
tri 1734 4556 1888 4710 ne
rect 1888 4590 1890 4710
rect 2010 4590 2046 4710
rect 1888 4556 2046 4590
tri 2046 4556 2200 4710 sw
tri 2284 4556 2438 4710 ne
rect 2438 4590 2440 4710
rect 2560 4590 2596 4710
rect 2438 4556 2596 4590
tri 2596 4556 2750 4710 sw
tri 2834 4556 2988 4710 ne
rect 2988 4590 2990 4710
rect 3110 4590 3146 4710
rect 2988 4556 3146 4590
tri 3146 4556 3300 4710 sw
tri 3384 4556 3538 4710 ne
rect 3538 4590 3540 4710
rect 3660 4590 3696 4710
rect 3538 4556 3696 4590
tri 3696 4556 3850 4710 sw
tri 3934 4556 4088 4710 ne
rect 4088 4590 4090 4710
rect 4210 4590 4246 4710
rect 4088 4556 4246 4590
tri 4246 4556 4400 4710 sw
tri 4484 4556 4638 4710 ne
rect 4638 4590 4640 4710
rect 4760 4590 4796 4710
rect 4638 4556 4796 4590
tri 4796 4556 4950 4710 sw
tri 5034 4556 5188 4710 ne
rect 5188 4590 5190 4710
rect 5310 4590 5346 4710
rect 5188 4556 5346 4590
tri 5346 4556 5500 4710 sw
tri 5584 4556 5738 4710 ne
rect 5738 4590 5740 4710
rect 5860 4590 5896 4710
rect 5738 4556 5896 4590
tri 5896 4556 6050 4710 sw
tri 6134 4556 6288 4710 ne
rect 6288 4590 6290 4710
rect 6410 4590 6446 4710
rect 6288 4556 6446 4590
tri 6446 4556 6600 4710 sw
tri 6684 4556 6838 4710 ne
rect 6838 4590 6840 4710
rect 6960 4590 6996 4710
rect 6838 4556 6996 4590
tri 6996 4556 7150 4710 sw
tri 7234 4556 7388 4710 ne
rect 7388 4590 7390 4710
rect 7510 4590 7546 4710
rect 7388 4556 7546 4590
tri 7546 4556 7700 4710 sw
tri 7784 4556 7938 4710 ne
rect 7938 4590 7940 4710
rect 8060 4590 8096 4710
rect 7938 4556 8096 4590
tri 8096 4556 8250 4710 sw
tri 8334 4556 8488 4710 ne
rect 8488 4590 8490 4710
rect 8610 4590 8646 4710
rect 8488 4556 8646 4590
tri 8646 4556 8800 4710 sw
tri 8884 4556 9038 4710 ne
rect 9038 4590 9040 4710
rect 9160 4590 9196 4710
rect 9038 4556 9196 4590
tri 9196 4556 9350 4710 sw
tri 9434 4556 9588 4710 ne
rect 9588 4590 9590 4710
rect 9710 4590 9746 4710
rect 9588 4556 9746 4590
tri 9746 4556 9900 4710 sw
tri 9984 4556 10138 4710 ne
rect 10138 4590 10140 4710
rect 10260 4590 10296 4710
rect 10138 4556 10296 4590
tri 10296 4556 10450 4710 sw
tri 10534 4556 10688 4710 ne
rect 10688 4590 10690 4710
rect 10810 4590 10846 4710
rect 10688 4556 10846 4590
tri 10846 4556 11000 4710 sw
tri 11084 4556 11238 4710 ne
rect 11238 4590 11240 4710
rect 11360 4590 11396 4710
rect 11238 4556 11396 4590
tri 11396 4556 11550 4710 sw
tri 11634 4556 11788 4710 ne
rect 11788 4590 11790 4710
rect 11910 4590 11946 4710
rect 11788 4556 11946 4590
tri 11946 4556 12100 4710 sw
tri 12184 4556 12338 4710 ne
rect 12338 4590 12340 4710
rect 12460 4590 12496 4710
rect 12338 4556 12496 4590
tri 12496 4556 12650 4710 sw
tri 12734 4556 12888 4710 ne
rect 12888 4590 12890 4710
rect 13010 4590 13046 4710
rect 12888 4556 13046 4590
tri 13046 4556 13200 4710 sw
tri 13284 4556 13438 4710 ne
rect 13438 4590 13440 4710
rect 13560 4608 13596 4710
tri 13596 4608 13698 4710 sw
rect 14775 4608 15775 5397
rect 13560 4590 15775 4608
rect 13438 4556 15775 4590
rect -156 4400 0 4556
tri 0 4400 156 4556 sw
tri 238 4400 394 4556 ne
rect 394 4400 550 4556
tri 550 4400 706 4556 sw
tri 788 4400 944 4556 ne
rect 944 4400 1100 4556
tri 1100 4400 1256 4556 sw
tri 1338 4400 1494 4556 ne
rect 1494 4400 1650 4556
tri 1650 4400 1806 4556 sw
tri 1888 4400 2044 4556 ne
rect 2044 4400 2200 4556
tri 2200 4400 2356 4556 sw
tri 2438 4400 2594 4556 ne
rect 2594 4400 2750 4556
tri 2750 4400 2906 4556 sw
tri 2988 4400 3144 4556 ne
rect 3144 4400 3300 4556
tri 3300 4400 3456 4556 sw
tri 3538 4400 3694 4556 ne
rect 3694 4400 3850 4556
tri 3850 4400 4006 4556 sw
tri 4088 4400 4244 4556 ne
rect 4244 4400 4400 4556
tri 4400 4400 4556 4556 sw
tri 4638 4400 4794 4556 ne
rect 4794 4400 4950 4556
tri 4950 4400 5106 4556 sw
tri 5188 4400 5344 4556 ne
rect 5344 4400 5500 4556
tri 5500 4400 5656 4556 sw
tri 5738 4400 5894 4556 ne
rect 5894 4400 6050 4556
tri 6050 4400 6206 4556 sw
tri 6288 4400 6444 4556 ne
rect 6444 4400 6600 4556
tri 6600 4400 6756 4556 sw
tri 6838 4400 6994 4556 ne
rect 6994 4400 7150 4556
tri 7150 4400 7306 4556 sw
tri 7388 4400 7544 4556 ne
rect 7544 4400 7700 4556
tri 7700 4400 7856 4556 sw
tri 7938 4400 8094 4556 ne
rect 8094 4400 8250 4556
tri 8250 4400 8406 4556 sw
tri 8488 4400 8644 4556 ne
rect 8644 4400 8800 4556
tri 8800 4400 8956 4556 sw
tri 9038 4400 9194 4556 ne
rect 9194 4400 9350 4556
tri 9350 4400 9506 4556 sw
tri 9588 4400 9744 4556 ne
rect 9744 4400 9900 4556
tri 9900 4400 10056 4556 sw
tri 10138 4400 10294 4556 ne
rect 10294 4400 10450 4556
tri 10450 4400 10606 4556 sw
tri 10688 4400 10844 4556 ne
rect 10844 4400 11000 4556
tri 11000 4400 11156 4556 sw
tri 11238 4400 11394 4556 ne
rect 11394 4400 11550 4556
tri 11550 4400 11706 4556 sw
tri 11788 4400 11944 4556 ne
rect 11944 4400 12100 4556
tri 12100 4400 12256 4556 sw
tri 12338 4400 12494 4556 ne
rect 12494 4400 12650 4556
tri 12650 4400 12806 4556 sw
tri 12888 4400 13044 4556 ne
rect 13044 4400 13200 4556
tri 13200 4400 13356 4556 sw
tri 13438 4400 13594 4556 ne
rect 13594 4400 15775 4556
rect -1025 4297 -394 4400
tri -394 4297 -291 4400 sw
tri -156 4297 -53 4400 ne
rect -53 4297 156 4400
tri 156 4297 259 4400 sw
tri 394 4297 497 4400 ne
rect 497 4297 706 4400
tri 706 4297 809 4400 sw
tri 944 4297 1047 4400 ne
rect 1047 4297 1256 4400
tri 1256 4297 1359 4400 sw
tri 1494 4297 1597 4400 ne
rect 1597 4297 1806 4400
tri 1806 4297 1909 4400 sw
tri 2044 4297 2147 4400 ne
rect 2147 4297 2356 4400
tri 2356 4297 2459 4400 sw
tri 2594 4297 2697 4400 ne
rect 2697 4297 2906 4400
tri 2906 4297 3009 4400 sw
tri 3144 4297 3247 4400 ne
rect 3247 4297 3456 4400
tri 3456 4297 3559 4400 sw
tri 3694 4297 3797 4400 ne
rect 3797 4297 4006 4400
tri 4006 4297 4109 4400 sw
tri 4244 4297 4347 4400 ne
rect 4347 4297 4556 4400
tri 4556 4297 4659 4400 sw
tri 4794 4297 4897 4400 ne
rect 4897 4297 5106 4400
tri 5106 4297 5209 4400 sw
tri 5344 4297 5447 4400 ne
rect 5447 4297 5656 4400
tri 5656 4297 5759 4400 sw
tri 5894 4297 5997 4400 ne
rect 5997 4297 6206 4400
tri 6206 4297 6309 4400 sw
tri 6444 4297 6547 4400 ne
rect 6547 4297 6756 4400
tri 6756 4297 6859 4400 sw
tri 6994 4297 7097 4400 ne
rect 7097 4297 7306 4400
tri 7306 4297 7409 4400 sw
tri 7544 4297 7647 4400 ne
rect 7647 4297 7856 4400
tri 7856 4297 7959 4400 sw
tri 8094 4297 8197 4400 ne
rect 8197 4297 8406 4400
tri 8406 4297 8509 4400 sw
tri 8644 4297 8747 4400 ne
rect 8747 4297 8956 4400
tri 8956 4297 9059 4400 sw
tri 9194 4297 9297 4400 ne
rect 9297 4297 9506 4400
tri 9506 4297 9609 4400 sw
tri 9744 4297 9847 4400 ne
rect 9847 4297 10056 4400
tri 10056 4297 10159 4400 sw
tri 10294 4297 10397 4400 ne
rect 10397 4297 10606 4400
tri 10606 4297 10709 4400 sw
tri 10844 4297 10947 4400 ne
rect 10947 4297 11156 4400
tri 11156 4297 11259 4400 sw
tri 11394 4297 11497 4400 ne
rect 11497 4297 11706 4400
tri 11706 4297 11809 4400 sw
tri 11944 4297 12047 4400 ne
rect 12047 4297 12256 4400
tri 12256 4297 12359 4400 sw
tri 12494 4297 12597 4400 ne
rect 12597 4297 12806 4400
tri 12806 4297 12909 4400 sw
tri 13044 4297 13147 4400 ne
rect 13147 4297 13356 4400
tri 13356 4297 13459 4400 sw
tri 13594 4297 13697 4400 ne
rect 13697 4297 15775 4400
rect -1025 4160 -291 4297
tri -291 4160 -154 4297 sw
tri -53 4160 84 4297 ne
rect 84 4160 259 4297
tri 259 4160 396 4297 sw
tri 497 4160 634 4297 ne
rect 634 4160 809 4297
tri 809 4160 946 4297 sw
tri 1047 4160 1184 4297 ne
rect 1184 4160 1359 4297
tri 1359 4160 1496 4297 sw
tri 1597 4160 1734 4297 ne
rect 1734 4160 1909 4297
tri 1909 4160 2046 4297 sw
tri 2147 4160 2284 4297 ne
rect 2284 4160 2459 4297
tri 2459 4160 2596 4297 sw
tri 2697 4160 2834 4297 ne
rect 2834 4160 3009 4297
tri 3009 4160 3146 4297 sw
tri 3247 4160 3384 4297 ne
rect 3384 4160 3559 4297
tri 3559 4160 3696 4297 sw
tri 3797 4160 3934 4297 ne
rect 3934 4160 4109 4297
tri 4109 4160 4246 4297 sw
tri 4347 4160 4484 4297 ne
rect 4484 4160 4659 4297
tri 4659 4160 4796 4297 sw
tri 4897 4160 5034 4297 ne
rect 5034 4160 5209 4297
tri 5209 4160 5346 4297 sw
tri 5447 4160 5584 4297 ne
rect 5584 4160 5759 4297
tri 5759 4160 5896 4297 sw
tri 5997 4160 6134 4297 ne
rect 6134 4160 6309 4297
tri 6309 4160 6446 4297 sw
tri 6547 4160 6684 4297 ne
rect 6684 4160 6859 4297
tri 6859 4160 6996 4297 sw
tri 7097 4160 7234 4297 ne
rect 7234 4160 7409 4297
tri 7409 4160 7546 4297 sw
tri 7647 4160 7784 4297 ne
rect 7784 4160 7959 4297
tri 7959 4160 8096 4297 sw
tri 8197 4160 8334 4297 ne
rect 8334 4160 8509 4297
tri 8509 4160 8646 4297 sw
tri 8747 4160 8884 4297 ne
rect 8884 4160 9059 4297
tri 9059 4160 9196 4297 sw
tri 9297 4160 9434 4297 ne
rect 9434 4160 9609 4297
tri 9609 4160 9746 4297 sw
tri 9847 4160 9984 4297 ne
rect 9984 4160 10159 4297
tri 10159 4160 10296 4297 sw
tri 10397 4160 10534 4297 ne
rect 10534 4160 10709 4297
tri 10709 4160 10846 4297 sw
tri 10947 4160 11084 4297 ne
rect 11084 4160 11259 4297
tri 11259 4160 11396 4297 sw
tri 11497 4160 11634 4297 ne
rect 11634 4160 11809 4297
tri 11809 4160 11946 4297 sw
tri 12047 4160 12184 4297 ne
rect 12184 4160 12359 4297
tri 12359 4160 12496 4297 sw
tri 12597 4160 12734 4297 ne
rect 12734 4160 12909 4297
tri 12909 4160 13046 4297 sw
tri 13147 4160 13284 4297 ne
rect 13284 4160 13459 4297
tri 13459 4160 13596 4297 sw
rect -1025 4142 -310 4160
tri -448 4040 -346 4142 ne
rect -346 4040 -310 4142
rect -190 4040 -154 4160
rect -2525 3850 -447 3903
tri -447 3850 -394 3903 sw
tri -346 3850 -156 4040 ne
rect -156 4006 -154 4040
tri -154 4006 0 4160 sw
tri 84 4006 238 4160 ne
rect 238 4040 240 4160
rect 360 4040 396 4160
rect 238 4006 396 4040
tri 396 4006 550 4160 sw
tri 634 4006 788 4160 ne
rect 788 4040 790 4160
rect 910 4040 946 4160
rect 788 4006 946 4040
tri 946 4006 1100 4160 sw
tri 1184 4006 1338 4160 ne
rect 1338 4040 1340 4160
rect 1460 4040 1496 4160
rect 1338 4006 1496 4040
tri 1496 4006 1650 4160 sw
tri 1734 4006 1888 4160 ne
rect 1888 4040 1890 4160
rect 2010 4040 2046 4160
rect 1888 4006 2046 4040
tri 2046 4006 2200 4160 sw
tri 2284 4006 2438 4160 ne
rect 2438 4040 2440 4160
rect 2560 4040 2596 4160
rect 2438 4006 2596 4040
tri 2596 4006 2750 4160 sw
tri 2834 4006 2988 4160 ne
rect 2988 4040 2990 4160
rect 3110 4040 3146 4160
rect 2988 4006 3146 4040
tri 3146 4006 3300 4160 sw
tri 3384 4006 3538 4160 ne
rect 3538 4040 3540 4160
rect 3660 4040 3696 4160
rect 3538 4006 3696 4040
tri 3696 4006 3850 4160 sw
tri 3934 4006 4088 4160 ne
rect 4088 4040 4090 4160
rect 4210 4040 4246 4160
rect 4088 4006 4246 4040
tri 4246 4006 4400 4160 sw
tri 4484 4006 4638 4160 ne
rect 4638 4040 4640 4160
rect 4760 4040 4796 4160
rect 4638 4006 4796 4040
tri 4796 4006 4950 4160 sw
tri 5034 4006 5188 4160 ne
rect 5188 4040 5190 4160
rect 5310 4040 5346 4160
rect 5188 4006 5346 4040
tri 5346 4006 5500 4160 sw
tri 5584 4006 5738 4160 ne
rect 5738 4040 5740 4160
rect 5860 4040 5896 4160
rect 5738 4006 5896 4040
tri 5896 4006 6050 4160 sw
tri 6134 4006 6288 4160 ne
rect 6288 4040 6290 4160
rect 6410 4040 6446 4160
rect 6288 4006 6446 4040
tri 6446 4006 6600 4160 sw
tri 6684 4006 6838 4160 ne
rect 6838 4040 6840 4160
rect 6960 4040 6996 4160
rect 6838 4006 6996 4040
tri 6996 4006 7150 4160 sw
tri 7234 4006 7388 4160 ne
rect 7388 4040 7390 4160
rect 7510 4040 7546 4160
rect 7388 4006 7546 4040
tri 7546 4006 7700 4160 sw
tri 7784 4006 7938 4160 ne
rect 7938 4040 7940 4160
rect 8060 4040 8096 4160
rect 7938 4006 8096 4040
tri 8096 4006 8250 4160 sw
tri 8334 4006 8488 4160 ne
rect 8488 4040 8490 4160
rect 8610 4040 8646 4160
rect 8488 4006 8646 4040
tri 8646 4006 8800 4160 sw
tri 8884 4006 9038 4160 ne
rect 9038 4040 9040 4160
rect 9160 4040 9196 4160
rect 9038 4006 9196 4040
tri 9196 4006 9350 4160 sw
tri 9434 4006 9588 4160 ne
rect 9588 4040 9590 4160
rect 9710 4040 9746 4160
rect 9588 4006 9746 4040
tri 9746 4006 9900 4160 sw
tri 9984 4006 10138 4160 ne
rect 10138 4040 10140 4160
rect 10260 4040 10296 4160
rect 10138 4006 10296 4040
tri 10296 4006 10450 4160 sw
tri 10534 4006 10688 4160 ne
rect 10688 4040 10690 4160
rect 10810 4040 10846 4160
rect 10688 4006 10846 4040
tri 10846 4006 11000 4160 sw
tri 11084 4006 11238 4160 ne
rect 11238 4040 11240 4160
rect 11360 4040 11396 4160
rect 11238 4006 11396 4040
tri 11396 4006 11550 4160 sw
tri 11634 4006 11788 4160 ne
rect 11788 4040 11790 4160
rect 11910 4040 11946 4160
rect 11788 4006 11946 4040
tri 11946 4006 12100 4160 sw
tri 12184 4006 12338 4160 ne
rect 12338 4040 12340 4160
rect 12460 4040 12496 4160
rect 12338 4006 12496 4040
tri 12496 4006 12650 4160 sw
tri 12734 4006 12888 4160 ne
rect 12888 4040 12890 4160
rect 13010 4040 13046 4160
rect 12888 4006 13046 4040
tri 13046 4006 13200 4160 sw
tri 13284 4006 13438 4160 ne
rect 13438 4040 13440 4160
rect 13560 4058 13596 4160
tri 13596 4058 13698 4160 sw
rect 13560 4040 14275 4058
rect 13438 4006 14275 4040
rect -156 3850 0 4006
tri 0 3850 156 4006 sw
tri 238 3850 394 4006 ne
rect 394 3850 550 4006
tri 550 3850 706 4006 sw
tri 788 3850 944 4006 ne
rect 944 3850 1100 4006
tri 1100 3850 1256 4006 sw
tri 1338 3850 1494 4006 ne
rect 1494 3850 1650 4006
tri 1650 3850 1806 4006 sw
tri 1888 3850 2044 4006 ne
rect 2044 3850 2200 4006
tri 2200 3850 2356 4006 sw
tri 2438 3850 2594 4006 ne
rect 2594 3850 2750 4006
tri 2750 3850 2906 4006 sw
tri 2988 3850 3144 4006 ne
rect 3144 3850 3300 4006
tri 3300 3850 3456 4006 sw
tri 3538 3850 3694 4006 ne
rect 3694 3850 3850 4006
tri 3850 3850 4006 4006 sw
tri 4088 3850 4244 4006 ne
rect 4244 3850 4400 4006
tri 4400 3850 4556 4006 sw
tri 4638 3850 4794 4006 ne
rect 4794 3850 4950 4006
tri 4950 3850 5106 4006 sw
tri 5188 3850 5344 4006 ne
rect 5344 3850 5500 4006
tri 5500 3850 5656 4006 sw
tri 5738 3850 5894 4006 ne
rect 5894 3850 6050 4006
tri 6050 3850 6206 4006 sw
tri 6288 3850 6444 4006 ne
rect 6444 3850 6600 4006
tri 6600 3850 6756 4006 sw
tri 6838 3850 6994 4006 ne
rect 6994 3850 7150 4006
tri 7150 3850 7306 4006 sw
tri 7388 3850 7544 4006 ne
rect 7544 3850 7700 4006
tri 7700 3850 7856 4006 sw
tri 7938 3850 8094 4006 ne
rect 8094 3850 8250 4006
tri 8250 3850 8406 4006 sw
tri 8488 3850 8644 4006 ne
rect 8644 3850 8800 4006
tri 8800 3850 8956 4006 sw
tri 9038 3850 9194 4006 ne
rect 9194 3850 9350 4006
tri 9350 3850 9506 4006 sw
tri 9588 3850 9744 4006 ne
rect 9744 3850 9900 4006
tri 9900 3850 10056 4006 sw
tri 10138 3850 10294 4006 ne
rect 10294 3850 10450 4006
tri 10450 3850 10606 4006 sw
tri 10688 3850 10844 4006 ne
rect 10844 3850 11000 4006
tri 11000 3850 11156 4006 sw
tri 11238 3850 11394 4006 ne
rect 11394 3850 11550 4006
tri 11550 3850 11706 4006 sw
tri 11788 3850 11944 4006 ne
rect 11944 3850 12100 4006
tri 12100 3850 12256 4006 sw
tri 12338 3850 12494 4006 ne
rect 12494 3850 12650 4006
tri 12650 3850 12806 4006 sw
tri 12888 3850 13044 4006 ne
rect 13044 3850 13200 4006
tri 13200 3850 13356 4006 sw
tri 13438 3850 13594 4006 ne
rect 13594 3850 14275 4006
rect -2525 3747 -394 3850
tri -394 3747 -291 3850 sw
tri -156 3747 -53 3850 ne
rect -53 3747 156 3850
tri 156 3747 259 3850 sw
tri 394 3747 497 3850 ne
rect 497 3747 706 3850
tri 706 3747 809 3850 sw
tri 944 3747 1047 3850 ne
rect 1047 3747 1256 3850
tri 1256 3747 1359 3850 sw
tri 1494 3747 1597 3850 ne
rect 1597 3747 1806 3850
tri 1806 3747 1909 3850 sw
tri 2044 3747 2147 3850 ne
rect 2147 3747 2356 3850
tri 2356 3747 2459 3850 sw
tri 2594 3747 2697 3850 ne
rect 2697 3747 2906 3850
tri 2906 3747 3009 3850 sw
tri 3144 3747 3247 3850 ne
rect 3247 3747 3456 3850
tri 3456 3747 3559 3850 sw
tri 3694 3747 3797 3850 ne
rect 3797 3747 4006 3850
tri 4006 3747 4109 3850 sw
tri 4244 3747 4347 3850 ne
rect 4347 3747 4556 3850
tri 4556 3747 4659 3850 sw
tri 4794 3747 4897 3850 ne
rect 4897 3747 5106 3850
tri 5106 3747 5209 3850 sw
tri 5344 3747 5447 3850 ne
rect 5447 3747 5656 3850
tri 5656 3747 5759 3850 sw
tri 5894 3747 5997 3850 ne
rect 5997 3747 6206 3850
tri 6206 3747 6309 3850 sw
tri 6444 3747 6547 3850 ne
rect 6547 3747 6756 3850
tri 6756 3747 6859 3850 sw
tri 6994 3747 7097 3850 ne
rect 7097 3747 7306 3850
tri 7306 3747 7409 3850 sw
tri 7544 3747 7647 3850 ne
rect 7647 3747 7856 3850
tri 7856 3747 7959 3850 sw
tri 8094 3747 8197 3850 ne
rect 8197 3747 8406 3850
tri 8406 3747 8509 3850 sw
tri 8644 3747 8747 3850 ne
rect 8747 3747 8956 3850
tri 8956 3747 9059 3850 sw
tri 9194 3747 9297 3850 ne
rect 9297 3747 9506 3850
tri 9506 3747 9609 3850 sw
tri 9744 3747 9847 3850 ne
rect 9847 3747 10056 3850
tri 10056 3747 10159 3850 sw
tri 10294 3747 10397 3850 ne
rect 10397 3747 10606 3850
tri 10606 3747 10709 3850 sw
tri 10844 3747 10947 3850 ne
rect 10947 3747 11156 3850
tri 11156 3747 11259 3850 sw
tri 11394 3747 11497 3850 ne
rect 11497 3747 11706 3850
tri 11706 3747 11809 3850 sw
tri 11944 3747 12047 3850 ne
rect 12047 3747 12256 3850
tri 12256 3747 12359 3850 sw
tri 12494 3747 12597 3850 ne
rect 12597 3747 12806 3850
tri 12806 3747 12909 3850 sw
tri 13044 3747 13147 3850 ne
rect 13147 3747 13356 3850
tri 13356 3747 13459 3850 sw
tri 13594 3747 13697 3850 ne
rect 13697 3747 14275 3850
rect -2525 3610 -291 3747
tri -291 3610 -154 3747 sw
tri -53 3610 84 3747 ne
rect 84 3610 259 3747
tri 259 3610 396 3747 sw
tri 497 3610 634 3747 ne
rect 634 3610 809 3747
tri 809 3610 946 3747 sw
tri 1047 3610 1184 3747 ne
rect 1184 3610 1359 3747
tri 1359 3610 1496 3747 sw
tri 1597 3610 1734 3747 ne
rect 1734 3610 1909 3747
tri 1909 3610 2046 3747 sw
tri 2147 3610 2284 3747 ne
rect 2284 3610 2459 3747
tri 2459 3610 2596 3747 sw
tri 2697 3610 2834 3747 ne
rect 2834 3610 3009 3747
tri 3009 3610 3146 3747 sw
tri 3247 3610 3384 3747 ne
rect 3384 3610 3559 3747
tri 3559 3610 3696 3747 sw
tri 3797 3610 3934 3747 ne
rect 3934 3610 4109 3747
tri 4109 3610 4246 3747 sw
tri 4347 3610 4484 3747 ne
rect 4484 3610 4659 3747
tri 4659 3610 4796 3747 sw
tri 4897 3610 5034 3747 ne
rect 5034 3610 5209 3747
tri 5209 3610 5346 3747 sw
tri 5447 3610 5584 3747 ne
rect 5584 3610 5759 3747
tri 5759 3610 5896 3747 sw
tri 5997 3610 6134 3747 ne
rect 6134 3610 6309 3747
tri 6309 3610 6446 3747 sw
tri 6547 3610 6684 3747 ne
rect 6684 3610 6859 3747
tri 6859 3610 6996 3747 sw
tri 7097 3610 7234 3747 ne
rect 7234 3610 7409 3747
tri 7409 3610 7546 3747 sw
tri 7647 3610 7784 3747 ne
rect 7784 3610 7959 3747
tri 7959 3610 8096 3747 sw
tri 8197 3610 8334 3747 ne
rect 8334 3610 8509 3747
tri 8509 3610 8646 3747 sw
tri 8747 3610 8884 3747 ne
rect 8884 3610 9059 3747
tri 9059 3610 9196 3747 sw
tri 9297 3610 9434 3747 ne
rect 9434 3610 9609 3747
tri 9609 3610 9746 3747 sw
tri 9847 3610 9984 3747 ne
rect 9984 3610 10159 3747
tri 10159 3610 10296 3747 sw
tri 10397 3610 10534 3747 ne
rect 10534 3610 10709 3747
tri 10709 3610 10846 3747 sw
tri 10947 3610 11084 3747 ne
rect 11084 3610 11259 3747
tri 11259 3610 11396 3747 sw
tri 11497 3610 11634 3747 ne
rect 11634 3610 11809 3747
tri 11809 3610 11946 3747 sw
tri 12047 3610 12184 3747 ne
rect 12184 3610 12359 3747
tri 12359 3610 12496 3747 sw
tri 12597 3610 12734 3747 ne
rect 12734 3610 12909 3747
tri 12909 3610 13046 3747 sw
tri 13147 3610 13284 3747 ne
rect 13284 3610 13459 3747
tri 13459 3610 13596 3747 sw
rect -2525 3592 -310 3610
rect -2525 2803 -1525 3592
tri -448 3490 -346 3592 ne
rect -346 3490 -310 3592
rect -190 3490 -154 3610
rect -1025 3300 -447 3353
tri -447 3300 -394 3353 sw
tri -346 3300 -156 3490 ne
rect -156 3456 -154 3490
tri -154 3456 0 3610 sw
tri 84 3456 238 3610 ne
rect 238 3490 240 3610
rect 360 3490 396 3610
rect 238 3456 396 3490
tri 396 3456 550 3610 sw
tri 634 3456 788 3610 ne
rect 788 3490 790 3610
rect 910 3490 946 3610
rect 788 3456 946 3490
tri 946 3456 1100 3610 sw
tri 1184 3456 1338 3610 ne
rect 1338 3490 1340 3610
rect 1460 3490 1496 3610
rect 1338 3456 1496 3490
tri 1496 3456 1650 3610 sw
tri 1734 3456 1888 3610 ne
rect 1888 3490 1890 3610
rect 2010 3490 2046 3610
rect 1888 3456 2046 3490
tri 2046 3456 2200 3610 sw
tri 2284 3456 2438 3610 ne
rect 2438 3490 2440 3610
rect 2560 3490 2596 3610
rect 2438 3456 2596 3490
tri 2596 3456 2750 3610 sw
tri 2834 3456 2988 3610 ne
rect 2988 3490 2990 3610
rect 3110 3490 3146 3610
rect 2988 3456 3146 3490
tri 3146 3456 3300 3610 sw
tri 3384 3456 3538 3610 ne
rect 3538 3490 3540 3610
rect 3660 3490 3696 3610
rect 3538 3456 3696 3490
tri 3696 3456 3850 3610 sw
tri 3934 3456 4088 3610 ne
rect 4088 3490 4090 3610
rect 4210 3490 4246 3610
rect 4088 3456 4246 3490
tri 4246 3456 4400 3610 sw
tri 4484 3456 4638 3610 ne
rect 4638 3490 4640 3610
rect 4760 3490 4796 3610
rect 4638 3456 4796 3490
tri 4796 3456 4950 3610 sw
tri 5034 3456 5188 3610 ne
rect 5188 3490 5190 3610
rect 5310 3490 5346 3610
rect 5188 3456 5346 3490
tri 5346 3456 5500 3610 sw
tri 5584 3456 5738 3610 ne
rect 5738 3490 5740 3610
rect 5860 3490 5896 3610
rect 5738 3456 5896 3490
tri 5896 3456 6050 3610 sw
tri 6134 3456 6288 3610 ne
rect 6288 3490 6290 3610
rect 6410 3490 6446 3610
rect 6288 3456 6446 3490
tri 6446 3456 6600 3610 sw
tri 6684 3456 6838 3610 ne
rect 6838 3490 6840 3610
rect 6960 3490 6996 3610
rect 6838 3456 6996 3490
tri 6996 3456 7150 3610 sw
tri 7234 3456 7388 3610 ne
rect 7388 3490 7390 3610
rect 7510 3490 7546 3610
rect 7388 3456 7546 3490
tri 7546 3456 7700 3610 sw
tri 7784 3456 7938 3610 ne
rect 7938 3490 7940 3610
rect 8060 3490 8096 3610
rect 7938 3456 8096 3490
tri 8096 3456 8250 3610 sw
tri 8334 3456 8488 3610 ne
rect 8488 3490 8490 3610
rect 8610 3490 8646 3610
rect 8488 3456 8646 3490
tri 8646 3456 8800 3610 sw
tri 8884 3456 9038 3610 ne
rect 9038 3490 9040 3610
rect 9160 3490 9196 3610
rect 9038 3456 9196 3490
tri 9196 3456 9350 3610 sw
tri 9434 3456 9588 3610 ne
rect 9588 3490 9590 3610
rect 9710 3490 9746 3610
rect 9588 3456 9746 3490
tri 9746 3456 9900 3610 sw
tri 9984 3456 10138 3610 ne
rect 10138 3490 10140 3610
rect 10260 3490 10296 3610
rect 10138 3456 10296 3490
tri 10296 3456 10450 3610 sw
tri 10534 3456 10688 3610 ne
rect 10688 3490 10690 3610
rect 10810 3490 10846 3610
rect 10688 3456 10846 3490
tri 10846 3456 11000 3610 sw
tri 11084 3456 11238 3610 ne
rect 11238 3490 11240 3610
rect 11360 3490 11396 3610
rect 11238 3456 11396 3490
tri 11396 3456 11550 3610 sw
tri 11634 3456 11788 3610 ne
rect 11788 3490 11790 3610
rect 11910 3490 11946 3610
rect 11788 3456 11946 3490
tri 11946 3456 12100 3610 sw
tri 12184 3456 12338 3610 ne
rect 12338 3490 12340 3610
rect 12460 3490 12496 3610
rect 12338 3456 12496 3490
tri 12496 3456 12650 3610 sw
tri 12734 3456 12888 3610 ne
rect 12888 3490 12890 3610
rect 13010 3490 13046 3610
rect 12888 3456 13046 3490
tri 13046 3456 13200 3610 sw
tri 13284 3456 13438 3610 ne
rect 13438 3490 13440 3610
rect 13560 3508 13596 3610
tri 13596 3508 13698 3610 sw
rect 14775 3508 15775 4297
rect 13560 3490 15775 3508
rect 13438 3456 15775 3490
rect -156 3300 0 3456
tri 0 3300 156 3456 sw
tri 238 3300 394 3456 ne
rect 394 3300 550 3456
tri 550 3300 706 3456 sw
tri 788 3300 944 3456 ne
rect 944 3300 1100 3456
tri 1100 3300 1256 3456 sw
tri 1338 3300 1494 3456 ne
rect 1494 3300 1650 3456
tri 1650 3300 1806 3456 sw
tri 1888 3300 2044 3456 ne
rect 2044 3300 2200 3456
tri 2200 3300 2356 3456 sw
tri 2438 3300 2594 3456 ne
rect 2594 3300 2750 3456
tri 2750 3300 2906 3456 sw
tri 2988 3300 3144 3456 ne
rect 3144 3300 3300 3456
tri 3300 3300 3456 3456 sw
tri 3538 3300 3694 3456 ne
rect 3694 3300 3850 3456
tri 3850 3300 4006 3456 sw
tri 4088 3300 4244 3456 ne
rect 4244 3300 4400 3456
tri 4400 3300 4556 3456 sw
tri 4638 3300 4794 3456 ne
rect 4794 3300 4950 3456
tri 4950 3300 5106 3456 sw
tri 5188 3300 5344 3456 ne
rect 5344 3300 5500 3456
tri 5500 3300 5656 3456 sw
tri 5738 3300 5894 3456 ne
rect 5894 3300 6050 3456
tri 6050 3300 6206 3456 sw
tri 6288 3300 6444 3456 ne
rect 6444 3300 6600 3456
tri 6600 3300 6756 3456 sw
tri 6838 3300 6994 3456 ne
rect 6994 3300 7150 3456
tri 7150 3300 7306 3456 sw
tri 7388 3300 7544 3456 ne
rect 7544 3300 7700 3456
tri 7700 3300 7856 3456 sw
tri 7938 3300 8094 3456 ne
rect 8094 3300 8250 3456
tri 8250 3300 8406 3456 sw
tri 8488 3300 8644 3456 ne
rect 8644 3300 8800 3456
tri 8800 3300 8956 3456 sw
tri 9038 3300 9194 3456 ne
rect 9194 3300 9350 3456
tri 9350 3300 9506 3456 sw
tri 9588 3300 9744 3456 ne
rect 9744 3300 9900 3456
tri 9900 3300 10056 3456 sw
tri 10138 3300 10294 3456 ne
rect 10294 3300 10450 3456
tri 10450 3300 10606 3456 sw
tri 10688 3300 10844 3456 ne
rect 10844 3300 11000 3456
tri 11000 3300 11156 3456 sw
tri 11238 3300 11394 3456 ne
rect 11394 3300 11550 3456
tri 11550 3300 11706 3456 sw
tri 11788 3300 11944 3456 ne
rect 11944 3300 12100 3456
tri 12100 3300 12256 3456 sw
tri 12338 3300 12494 3456 ne
rect 12494 3300 12650 3456
tri 12650 3300 12806 3456 sw
tri 12888 3300 13044 3456 ne
rect 13044 3300 13200 3456
tri 13200 3300 13356 3456 sw
tri 13438 3300 13594 3456 ne
rect 13594 3300 15775 3456
rect -1025 3197 -394 3300
tri -394 3197 -291 3300 sw
tri -156 3197 -53 3300 ne
rect -53 3197 156 3300
tri 156 3197 259 3300 sw
tri 394 3197 497 3300 ne
rect 497 3197 706 3300
tri 706 3197 809 3300 sw
tri 944 3197 1047 3300 ne
rect 1047 3197 1256 3300
tri 1256 3197 1359 3300 sw
tri 1494 3197 1597 3300 ne
rect 1597 3197 1806 3300
tri 1806 3197 1909 3300 sw
tri 2044 3197 2147 3300 ne
rect 2147 3197 2356 3300
tri 2356 3197 2459 3300 sw
tri 2594 3197 2697 3300 ne
rect 2697 3197 2906 3300
tri 2906 3197 3009 3300 sw
tri 3144 3197 3247 3300 ne
rect 3247 3197 3456 3300
tri 3456 3197 3559 3300 sw
tri 3694 3197 3797 3300 ne
rect 3797 3197 4006 3300
tri 4006 3197 4109 3300 sw
tri 4244 3197 4347 3300 ne
rect 4347 3197 4556 3300
tri 4556 3197 4659 3300 sw
tri 4794 3197 4897 3300 ne
rect 4897 3197 5106 3300
tri 5106 3197 5209 3300 sw
tri 5344 3197 5447 3300 ne
rect 5447 3197 5656 3300
tri 5656 3197 5759 3300 sw
tri 5894 3197 5997 3300 ne
rect 5997 3197 6206 3300
tri 6206 3197 6309 3300 sw
tri 6444 3197 6547 3300 ne
rect 6547 3197 6756 3300
tri 6756 3197 6859 3300 sw
tri 6994 3197 7097 3300 ne
rect 7097 3197 7306 3300
tri 7306 3197 7409 3300 sw
tri 7544 3197 7647 3300 ne
rect 7647 3197 7856 3300
tri 7856 3197 7959 3300 sw
tri 8094 3197 8197 3300 ne
rect 8197 3197 8406 3300
tri 8406 3197 8509 3300 sw
tri 8644 3197 8747 3300 ne
rect 8747 3197 8956 3300
tri 8956 3197 9059 3300 sw
tri 9194 3197 9297 3300 ne
rect 9297 3197 9506 3300
tri 9506 3197 9609 3300 sw
tri 9744 3197 9847 3300 ne
rect 9847 3197 10056 3300
tri 10056 3197 10159 3300 sw
tri 10294 3197 10397 3300 ne
rect 10397 3197 10606 3300
tri 10606 3197 10709 3300 sw
tri 10844 3197 10947 3300 ne
rect 10947 3197 11156 3300
tri 11156 3197 11259 3300 sw
tri 11394 3197 11497 3300 ne
rect 11497 3197 11706 3300
tri 11706 3197 11809 3300 sw
tri 11944 3197 12047 3300 ne
rect 12047 3197 12256 3300
tri 12256 3197 12359 3300 sw
tri 12494 3197 12597 3300 ne
rect 12597 3197 12806 3300
tri 12806 3197 12909 3300 sw
tri 13044 3197 13147 3300 ne
rect 13147 3197 13356 3300
tri 13356 3197 13459 3300 sw
tri 13594 3197 13697 3300 ne
rect 13697 3197 15775 3300
rect -1025 3060 -291 3197
tri -291 3060 -154 3197 sw
tri -53 3060 84 3197 ne
rect 84 3060 259 3197
tri 259 3060 396 3197 sw
tri 497 3060 634 3197 ne
rect 634 3060 809 3197
tri 809 3060 946 3197 sw
tri 1047 3060 1184 3197 ne
rect 1184 3060 1359 3197
tri 1359 3060 1496 3197 sw
tri 1597 3060 1734 3197 ne
rect 1734 3060 1909 3197
tri 1909 3060 2046 3197 sw
tri 2147 3060 2284 3197 ne
rect 2284 3060 2459 3197
tri 2459 3060 2596 3197 sw
tri 2697 3060 2834 3197 ne
rect 2834 3060 3009 3197
tri 3009 3060 3146 3197 sw
tri 3247 3060 3384 3197 ne
rect 3384 3060 3559 3197
tri 3559 3060 3696 3197 sw
tri 3797 3060 3934 3197 ne
rect 3934 3060 4109 3197
tri 4109 3060 4246 3197 sw
tri 4347 3060 4484 3197 ne
rect 4484 3060 4659 3197
tri 4659 3060 4796 3197 sw
tri 4897 3060 5034 3197 ne
rect 5034 3060 5209 3197
tri 5209 3060 5346 3197 sw
tri 5447 3060 5584 3197 ne
rect 5584 3060 5759 3197
tri 5759 3060 5896 3197 sw
tri 5997 3060 6134 3197 ne
rect 6134 3060 6309 3197
tri 6309 3060 6446 3197 sw
tri 6547 3060 6684 3197 ne
rect 6684 3060 6859 3197
tri 6859 3060 6996 3197 sw
tri 7097 3060 7234 3197 ne
rect 7234 3060 7409 3197
tri 7409 3060 7546 3197 sw
tri 7647 3060 7784 3197 ne
rect 7784 3060 7959 3197
tri 7959 3060 8096 3197 sw
tri 8197 3060 8334 3197 ne
rect 8334 3060 8509 3197
tri 8509 3060 8646 3197 sw
tri 8747 3060 8884 3197 ne
rect 8884 3060 9059 3197
tri 9059 3060 9196 3197 sw
tri 9297 3060 9434 3197 ne
rect 9434 3060 9609 3197
tri 9609 3060 9746 3197 sw
tri 9847 3060 9984 3197 ne
rect 9984 3060 10159 3197
tri 10159 3060 10296 3197 sw
tri 10397 3060 10534 3197 ne
rect 10534 3060 10709 3197
tri 10709 3060 10846 3197 sw
tri 10947 3060 11084 3197 ne
rect 11084 3060 11259 3197
tri 11259 3060 11396 3197 sw
tri 11497 3060 11634 3197 ne
rect 11634 3060 11809 3197
tri 11809 3060 11946 3197 sw
tri 12047 3060 12184 3197 ne
rect 12184 3060 12359 3197
tri 12359 3060 12496 3197 sw
tri 12597 3060 12734 3197 ne
rect 12734 3060 12909 3197
tri 12909 3060 13046 3197 sw
tri 13147 3060 13284 3197 ne
rect 13284 3060 13459 3197
tri 13459 3060 13596 3197 sw
rect -1025 3042 -310 3060
tri -448 2940 -346 3042 ne
rect -346 2940 -310 3042
rect -190 2940 -154 3060
rect -2525 2750 -447 2803
tri -447 2750 -394 2803 sw
tri -346 2750 -156 2940 ne
rect -156 2906 -154 2940
tri -154 2906 0 3060 sw
tri 84 2906 238 3060 ne
rect 238 2940 240 3060
rect 360 2940 396 3060
rect 238 2906 396 2940
tri 396 2906 550 3060 sw
tri 634 2906 788 3060 ne
rect 788 2940 790 3060
rect 910 2940 946 3060
rect 788 2906 946 2940
tri 946 2906 1100 3060 sw
tri 1184 2906 1338 3060 ne
rect 1338 2940 1340 3060
rect 1460 2940 1496 3060
rect 1338 2906 1496 2940
tri 1496 2906 1650 3060 sw
tri 1734 2906 1888 3060 ne
rect 1888 2940 1890 3060
rect 2010 2940 2046 3060
rect 1888 2906 2046 2940
tri 2046 2906 2200 3060 sw
tri 2284 2906 2438 3060 ne
rect 2438 2940 2440 3060
rect 2560 2940 2596 3060
rect 2438 2906 2596 2940
tri 2596 2906 2750 3060 sw
tri 2834 2906 2988 3060 ne
rect 2988 2940 2990 3060
rect 3110 2940 3146 3060
rect 2988 2906 3146 2940
tri 3146 2906 3300 3060 sw
tri 3384 2906 3538 3060 ne
rect 3538 2940 3540 3060
rect 3660 2940 3696 3060
rect 3538 2906 3696 2940
tri 3696 2906 3850 3060 sw
tri 3934 2906 4088 3060 ne
rect 4088 2940 4090 3060
rect 4210 2940 4246 3060
rect 4088 2906 4246 2940
tri 4246 2906 4400 3060 sw
tri 4484 2906 4638 3060 ne
rect 4638 2940 4640 3060
rect 4760 2940 4796 3060
rect 4638 2906 4796 2940
tri 4796 2906 4950 3060 sw
tri 5034 2906 5188 3060 ne
rect 5188 2940 5190 3060
rect 5310 2940 5346 3060
rect 5188 2906 5346 2940
tri 5346 2906 5500 3060 sw
tri 5584 2906 5738 3060 ne
rect 5738 2940 5740 3060
rect 5860 2940 5896 3060
rect 5738 2906 5896 2940
tri 5896 2906 6050 3060 sw
tri 6134 2906 6288 3060 ne
rect 6288 2940 6290 3060
rect 6410 2940 6446 3060
rect 6288 2906 6446 2940
tri 6446 2906 6600 3060 sw
tri 6684 2906 6838 3060 ne
rect 6838 2940 6840 3060
rect 6960 2940 6996 3060
rect 6838 2906 6996 2940
tri 6996 2906 7150 3060 sw
tri 7234 2906 7388 3060 ne
rect 7388 2940 7390 3060
rect 7510 2940 7546 3060
rect 7388 2906 7546 2940
tri 7546 2906 7700 3060 sw
tri 7784 2906 7938 3060 ne
rect 7938 2940 7940 3060
rect 8060 2940 8096 3060
rect 7938 2906 8096 2940
tri 8096 2906 8250 3060 sw
tri 8334 2906 8488 3060 ne
rect 8488 2940 8490 3060
rect 8610 2940 8646 3060
rect 8488 2906 8646 2940
tri 8646 2906 8800 3060 sw
tri 8884 2906 9038 3060 ne
rect 9038 2940 9040 3060
rect 9160 2940 9196 3060
rect 9038 2906 9196 2940
tri 9196 2906 9350 3060 sw
tri 9434 2906 9588 3060 ne
rect 9588 2940 9590 3060
rect 9710 2940 9746 3060
rect 9588 2906 9746 2940
tri 9746 2906 9900 3060 sw
tri 9984 2906 10138 3060 ne
rect 10138 2940 10140 3060
rect 10260 2940 10296 3060
rect 10138 2906 10296 2940
tri 10296 2906 10450 3060 sw
tri 10534 2906 10688 3060 ne
rect 10688 2940 10690 3060
rect 10810 2940 10846 3060
rect 10688 2906 10846 2940
tri 10846 2906 11000 3060 sw
tri 11084 2906 11238 3060 ne
rect 11238 2940 11240 3060
rect 11360 2940 11396 3060
rect 11238 2906 11396 2940
tri 11396 2906 11550 3060 sw
tri 11634 2906 11788 3060 ne
rect 11788 2940 11790 3060
rect 11910 2940 11946 3060
rect 11788 2906 11946 2940
tri 11946 2906 12100 3060 sw
tri 12184 2906 12338 3060 ne
rect 12338 2940 12340 3060
rect 12460 2940 12496 3060
rect 12338 2906 12496 2940
tri 12496 2906 12650 3060 sw
tri 12734 2906 12888 3060 ne
rect 12888 2940 12890 3060
rect 13010 2940 13046 3060
rect 12888 2906 13046 2940
tri 13046 2906 13200 3060 sw
tri 13284 2906 13438 3060 ne
rect 13438 2940 13440 3060
rect 13560 2958 13596 3060
tri 13596 2958 13698 3060 sw
rect 13560 2940 14275 2958
rect 13438 2906 14275 2940
rect -156 2750 0 2906
tri 0 2750 156 2906 sw
tri 238 2750 394 2906 ne
rect 394 2750 550 2906
tri 550 2750 706 2906 sw
tri 788 2750 944 2906 ne
rect 944 2750 1100 2906
tri 1100 2750 1256 2906 sw
tri 1338 2750 1494 2906 ne
rect 1494 2750 1650 2906
tri 1650 2750 1806 2906 sw
tri 1888 2750 2044 2906 ne
rect 2044 2750 2200 2906
tri 2200 2750 2356 2906 sw
tri 2438 2750 2594 2906 ne
rect 2594 2750 2750 2906
tri 2750 2750 2906 2906 sw
tri 2988 2750 3144 2906 ne
rect 3144 2750 3300 2906
tri 3300 2750 3456 2906 sw
tri 3538 2750 3694 2906 ne
rect 3694 2750 3850 2906
tri 3850 2750 4006 2906 sw
tri 4088 2750 4244 2906 ne
rect 4244 2750 4400 2906
tri 4400 2750 4556 2906 sw
tri 4638 2750 4794 2906 ne
rect 4794 2750 4950 2906
tri 4950 2750 5106 2906 sw
tri 5188 2750 5344 2906 ne
rect 5344 2750 5500 2906
tri 5500 2750 5656 2906 sw
tri 5738 2750 5894 2906 ne
rect 5894 2750 6050 2906
tri 6050 2750 6206 2906 sw
tri 6288 2750 6444 2906 ne
rect 6444 2750 6600 2906
tri 6600 2750 6756 2906 sw
tri 6838 2750 6994 2906 ne
rect 6994 2750 7150 2906
tri 7150 2750 7306 2906 sw
tri 7388 2750 7544 2906 ne
rect 7544 2750 7700 2906
tri 7700 2750 7856 2906 sw
tri 7938 2750 8094 2906 ne
rect 8094 2750 8250 2906
tri 8250 2750 8406 2906 sw
tri 8488 2750 8644 2906 ne
rect 8644 2750 8800 2906
tri 8800 2750 8956 2906 sw
tri 9038 2750 9194 2906 ne
rect 9194 2750 9350 2906
tri 9350 2750 9506 2906 sw
tri 9588 2750 9744 2906 ne
rect 9744 2750 9900 2906
tri 9900 2750 10056 2906 sw
tri 10138 2750 10294 2906 ne
rect 10294 2750 10450 2906
tri 10450 2750 10606 2906 sw
tri 10688 2750 10844 2906 ne
rect 10844 2750 11000 2906
tri 11000 2750 11156 2906 sw
tri 11238 2750 11394 2906 ne
rect 11394 2750 11550 2906
tri 11550 2750 11706 2906 sw
tri 11788 2750 11944 2906 ne
rect 11944 2750 12100 2906
tri 12100 2750 12256 2906 sw
tri 12338 2750 12494 2906 ne
rect 12494 2750 12650 2906
tri 12650 2750 12806 2906 sw
tri 12888 2750 13044 2906 ne
rect 13044 2750 13200 2906
tri 13200 2750 13356 2906 sw
tri 13438 2750 13594 2906 ne
rect 13594 2750 14275 2906
rect -2525 2647 -394 2750
tri -394 2647 -291 2750 sw
tri -156 2647 -53 2750 ne
rect -53 2647 156 2750
tri 156 2647 259 2750 sw
tri 394 2647 497 2750 ne
rect 497 2647 706 2750
tri 706 2647 809 2750 sw
tri 944 2647 1047 2750 ne
rect 1047 2647 1256 2750
tri 1256 2647 1359 2750 sw
tri 1494 2647 1597 2750 ne
rect 1597 2647 1806 2750
tri 1806 2647 1909 2750 sw
tri 2044 2647 2147 2750 ne
rect 2147 2647 2356 2750
tri 2356 2647 2459 2750 sw
tri 2594 2647 2697 2750 ne
rect 2697 2647 2906 2750
tri 2906 2647 3009 2750 sw
tri 3144 2647 3247 2750 ne
rect 3247 2647 3456 2750
tri 3456 2647 3559 2750 sw
tri 3694 2647 3797 2750 ne
rect 3797 2647 4006 2750
tri 4006 2647 4109 2750 sw
tri 4244 2647 4347 2750 ne
rect 4347 2647 4556 2750
tri 4556 2647 4659 2750 sw
tri 4794 2647 4897 2750 ne
rect 4897 2647 5106 2750
tri 5106 2647 5209 2750 sw
tri 5344 2647 5447 2750 ne
rect 5447 2647 5656 2750
tri 5656 2647 5759 2750 sw
tri 5894 2647 5997 2750 ne
rect 5997 2647 6206 2750
tri 6206 2647 6309 2750 sw
tri 6444 2647 6547 2750 ne
rect 6547 2647 6756 2750
tri 6756 2647 6859 2750 sw
tri 6994 2647 7097 2750 ne
rect 7097 2647 7306 2750
tri 7306 2647 7409 2750 sw
tri 7544 2647 7647 2750 ne
rect 7647 2647 7856 2750
tri 7856 2647 7959 2750 sw
tri 8094 2647 8197 2750 ne
rect 8197 2647 8406 2750
tri 8406 2647 8509 2750 sw
tri 8644 2647 8747 2750 ne
rect 8747 2647 8956 2750
tri 8956 2647 9059 2750 sw
tri 9194 2647 9297 2750 ne
rect 9297 2647 9506 2750
tri 9506 2647 9609 2750 sw
tri 9744 2647 9847 2750 ne
rect 9847 2647 10056 2750
tri 10056 2647 10159 2750 sw
tri 10294 2647 10397 2750 ne
rect 10397 2647 10606 2750
tri 10606 2647 10709 2750 sw
tri 10844 2647 10947 2750 ne
rect 10947 2647 11156 2750
tri 11156 2647 11259 2750 sw
tri 11394 2647 11497 2750 ne
rect 11497 2647 11706 2750
tri 11706 2647 11809 2750 sw
tri 11944 2647 12047 2750 ne
rect 12047 2647 12256 2750
tri 12256 2647 12359 2750 sw
tri 12494 2647 12597 2750 ne
rect 12597 2647 12806 2750
tri 12806 2647 12909 2750 sw
tri 13044 2647 13147 2750 ne
rect 13147 2647 13356 2750
tri 13356 2647 13459 2750 sw
tri 13594 2647 13697 2750 ne
rect 13697 2647 14275 2750
rect -2525 2510 -291 2647
tri -291 2510 -154 2647 sw
tri -53 2510 84 2647 ne
rect 84 2510 259 2647
tri 259 2510 396 2647 sw
tri 497 2510 634 2647 ne
rect 634 2510 809 2647
tri 809 2510 946 2647 sw
tri 1047 2510 1184 2647 ne
rect 1184 2510 1359 2647
tri 1359 2510 1496 2647 sw
tri 1597 2510 1734 2647 ne
rect 1734 2510 1909 2647
tri 1909 2510 2046 2647 sw
tri 2147 2510 2284 2647 ne
rect 2284 2510 2459 2647
tri 2459 2510 2596 2647 sw
tri 2697 2510 2834 2647 ne
rect 2834 2510 3009 2647
tri 3009 2510 3146 2647 sw
tri 3247 2510 3384 2647 ne
rect 3384 2510 3559 2647
tri 3559 2510 3696 2647 sw
tri 3797 2510 3934 2647 ne
rect 3934 2510 4109 2647
tri 4109 2510 4246 2647 sw
tri 4347 2510 4484 2647 ne
rect 4484 2510 4659 2647
tri 4659 2510 4796 2647 sw
tri 4897 2510 5034 2647 ne
rect 5034 2510 5209 2647
tri 5209 2510 5346 2647 sw
tri 5447 2510 5584 2647 ne
rect 5584 2510 5759 2647
tri 5759 2510 5896 2647 sw
tri 5997 2510 6134 2647 ne
rect 6134 2510 6309 2647
tri 6309 2510 6446 2647 sw
tri 6547 2510 6684 2647 ne
rect 6684 2510 6859 2647
tri 6859 2510 6996 2647 sw
tri 7097 2510 7234 2647 ne
rect 7234 2510 7409 2647
tri 7409 2510 7546 2647 sw
tri 7647 2510 7784 2647 ne
rect 7784 2510 7959 2647
tri 7959 2510 8096 2647 sw
tri 8197 2510 8334 2647 ne
rect 8334 2510 8509 2647
tri 8509 2510 8646 2647 sw
tri 8747 2510 8884 2647 ne
rect 8884 2510 9059 2647
tri 9059 2510 9196 2647 sw
tri 9297 2510 9434 2647 ne
rect 9434 2510 9609 2647
tri 9609 2510 9746 2647 sw
tri 9847 2510 9984 2647 ne
rect 9984 2510 10159 2647
tri 10159 2510 10296 2647 sw
tri 10397 2510 10534 2647 ne
rect 10534 2510 10709 2647
tri 10709 2510 10846 2647 sw
tri 10947 2510 11084 2647 ne
rect 11084 2510 11259 2647
tri 11259 2510 11396 2647 sw
tri 11497 2510 11634 2647 ne
rect 11634 2510 11809 2647
tri 11809 2510 11946 2647 sw
tri 12047 2510 12184 2647 ne
rect 12184 2510 12359 2647
tri 12359 2510 12496 2647 sw
tri 12597 2510 12734 2647 ne
rect 12734 2510 12909 2647
tri 12909 2510 13046 2647 sw
tri 13147 2510 13284 2647 ne
rect 13284 2510 13459 2647
tri 13459 2510 13596 2647 sw
rect -2525 2492 -310 2510
rect -2525 1703 -1525 2492
tri -448 2390 -346 2492 ne
rect -346 2390 -310 2492
rect -190 2390 -154 2510
rect -1025 2200 -447 2253
tri -447 2200 -394 2253 sw
tri -346 2200 -156 2390 ne
rect -156 2356 -154 2390
tri -154 2356 0 2510 sw
tri 84 2356 238 2510 ne
rect 238 2390 240 2510
rect 360 2390 396 2510
rect 238 2356 396 2390
tri 396 2356 550 2510 sw
tri 634 2356 788 2510 ne
rect 788 2390 790 2510
rect 910 2390 946 2510
rect 788 2356 946 2390
tri 946 2356 1100 2510 sw
tri 1184 2356 1338 2510 ne
rect 1338 2390 1340 2510
rect 1460 2390 1496 2510
rect 1338 2356 1496 2390
tri 1496 2356 1650 2510 sw
tri 1734 2356 1888 2510 ne
rect 1888 2390 1890 2510
rect 2010 2390 2046 2510
rect 1888 2356 2046 2390
tri 2046 2356 2200 2510 sw
tri 2284 2356 2438 2510 ne
rect 2438 2390 2440 2510
rect 2560 2390 2596 2510
rect 2438 2356 2596 2390
tri 2596 2356 2750 2510 sw
tri 2834 2356 2988 2510 ne
rect 2988 2390 2990 2510
rect 3110 2390 3146 2510
rect 2988 2356 3146 2390
tri 3146 2356 3300 2510 sw
tri 3384 2356 3538 2510 ne
rect 3538 2390 3540 2510
rect 3660 2390 3696 2510
rect 3538 2356 3696 2390
tri 3696 2356 3850 2510 sw
tri 3934 2356 4088 2510 ne
rect 4088 2390 4090 2510
rect 4210 2390 4246 2510
rect 4088 2356 4246 2390
tri 4246 2356 4400 2510 sw
tri 4484 2356 4638 2510 ne
rect 4638 2390 4640 2510
rect 4760 2390 4796 2510
rect 4638 2356 4796 2390
tri 4796 2356 4950 2510 sw
tri 5034 2356 5188 2510 ne
rect 5188 2390 5190 2510
rect 5310 2390 5346 2510
rect 5188 2356 5346 2390
tri 5346 2356 5500 2510 sw
tri 5584 2356 5738 2510 ne
rect 5738 2390 5740 2510
rect 5860 2390 5896 2510
rect 5738 2356 5896 2390
tri 5896 2356 6050 2510 sw
tri 6134 2356 6288 2510 ne
rect 6288 2390 6290 2510
rect 6410 2390 6446 2510
rect 6288 2356 6446 2390
tri 6446 2356 6600 2510 sw
tri 6684 2356 6838 2510 ne
rect 6838 2390 6840 2510
rect 6960 2390 6996 2510
rect 6838 2356 6996 2390
tri 6996 2356 7150 2510 sw
tri 7234 2356 7388 2510 ne
rect 7388 2390 7390 2510
rect 7510 2390 7546 2510
rect 7388 2356 7546 2390
tri 7546 2356 7700 2510 sw
tri 7784 2356 7938 2510 ne
rect 7938 2390 7940 2510
rect 8060 2390 8096 2510
rect 7938 2356 8096 2390
tri 8096 2356 8250 2510 sw
tri 8334 2356 8488 2510 ne
rect 8488 2390 8490 2510
rect 8610 2390 8646 2510
rect 8488 2356 8646 2390
tri 8646 2356 8800 2510 sw
tri 8884 2356 9038 2510 ne
rect 9038 2390 9040 2510
rect 9160 2390 9196 2510
rect 9038 2356 9196 2390
tri 9196 2356 9350 2510 sw
tri 9434 2356 9588 2510 ne
rect 9588 2390 9590 2510
rect 9710 2390 9746 2510
rect 9588 2356 9746 2390
tri 9746 2356 9900 2510 sw
tri 9984 2356 10138 2510 ne
rect 10138 2390 10140 2510
rect 10260 2390 10296 2510
rect 10138 2356 10296 2390
tri 10296 2356 10450 2510 sw
tri 10534 2356 10688 2510 ne
rect 10688 2390 10690 2510
rect 10810 2390 10846 2510
rect 10688 2356 10846 2390
tri 10846 2356 11000 2510 sw
tri 11084 2356 11238 2510 ne
rect 11238 2390 11240 2510
rect 11360 2390 11396 2510
rect 11238 2356 11396 2390
tri 11396 2356 11550 2510 sw
tri 11634 2356 11788 2510 ne
rect 11788 2390 11790 2510
rect 11910 2390 11946 2510
rect 11788 2356 11946 2390
tri 11946 2356 12100 2510 sw
tri 12184 2356 12338 2510 ne
rect 12338 2390 12340 2510
rect 12460 2390 12496 2510
rect 12338 2356 12496 2390
tri 12496 2356 12650 2510 sw
tri 12734 2356 12888 2510 ne
rect 12888 2390 12890 2510
rect 13010 2390 13046 2510
rect 12888 2356 13046 2390
tri 13046 2356 13200 2510 sw
tri 13284 2356 13438 2510 ne
rect 13438 2390 13440 2510
rect 13560 2408 13596 2510
tri 13596 2408 13698 2510 sw
rect 14775 2408 15775 3197
rect 13560 2390 15775 2408
rect 13438 2356 15775 2390
rect -156 2200 0 2356
tri 0 2200 156 2356 sw
tri 238 2200 394 2356 ne
rect 394 2200 550 2356
tri 550 2200 706 2356 sw
tri 788 2200 944 2356 ne
rect 944 2200 1100 2356
tri 1100 2200 1256 2356 sw
tri 1338 2200 1494 2356 ne
rect 1494 2200 1650 2356
tri 1650 2200 1806 2356 sw
tri 1888 2200 2044 2356 ne
rect 2044 2200 2200 2356
tri 2200 2200 2356 2356 sw
tri 2438 2200 2594 2356 ne
rect 2594 2200 2750 2356
tri 2750 2200 2906 2356 sw
tri 2988 2200 3144 2356 ne
rect 3144 2200 3300 2356
tri 3300 2200 3456 2356 sw
tri 3538 2200 3694 2356 ne
rect 3694 2200 3850 2356
tri 3850 2200 4006 2356 sw
tri 4088 2200 4244 2356 ne
rect 4244 2200 4400 2356
tri 4400 2200 4556 2356 sw
tri 4638 2200 4794 2356 ne
rect 4794 2200 4950 2356
tri 4950 2200 5106 2356 sw
tri 5188 2200 5344 2356 ne
rect 5344 2200 5500 2356
tri 5500 2200 5656 2356 sw
tri 5738 2200 5894 2356 ne
rect 5894 2200 6050 2356
tri 6050 2200 6206 2356 sw
tri 6288 2200 6444 2356 ne
rect 6444 2200 6600 2356
tri 6600 2200 6756 2356 sw
tri 6838 2200 6994 2356 ne
rect 6994 2200 7150 2356
tri 7150 2200 7306 2356 sw
tri 7388 2200 7544 2356 ne
rect 7544 2200 7700 2356
tri 7700 2200 7856 2356 sw
tri 7938 2200 8094 2356 ne
rect 8094 2200 8250 2356
tri 8250 2200 8406 2356 sw
tri 8488 2200 8644 2356 ne
rect 8644 2200 8800 2356
tri 8800 2200 8956 2356 sw
tri 9038 2200 9194 2356 ne
rect 9194 2200 9350 2356
tri 9350 2200 9506 2356 sw
tri 9588 2200 9744 2356 ne
rect 9744 2200 9900 2356
tri 9900 2200 10056 2356 sw
tri 10138 2200 10294 2356 ne
rect 10294 2200 10450 2356
tri 10450 2200 10606 2356 sw
tri 10688 2200 10844 2356 ne
rect 10844 2200 11000 2356
tri 11000 2200 11156 2356 sw
tri 11238 2200 11394 2356 ne
rect 11394 2200 11550 2356
tri 11550 2200 11706 2356 sw
tri 11788 2200 11944 2356 ne
rect 11944 2200 12100 2356
tri 12100 2200 12256 2356 sw
tri 12338 2200 12494 2356 ne
rect 12494 2200 12650 2356
tri 12650 2200 12806 2356 sw
tri 12888 2200 13044 2356 ne
rect 13044 2200 13200 2356
tri 13200 2200 13356 2356 sw
tri 13438 2200 13594 2356 ne
rect 13594 2200 15775 2356
rect -1025 2097 -394 2200
tri -394 2097 -291 2200 sw
tri -156 2097 -53 2200 ne
rect -53 2097 156 2200
tri 156 2097 259 2200 sw
tri 394 2097 497 2200 ne
rect 497 2097 706 2200
tri 706 2097 809 2200 sw
tri 944 2097 1047 2200 ne
rect 1047 2097 1256 2200
tri 1256 2097 1359 2200 sw
tri 1494 2097 1597 2200 ne
rect 1597 2097 1806 2200
tri 1806 2097 1909 2200 sw
tri 2044 2097 2147 2200 ne
rect 2147 2097 2356 2200
tri 2356 2097 2459 2200 sw
tri 2594 2097 2697 2200 ne
rect 2697 2097 2906 2200
tri 2906 2097 3009 2200 sw
tri 3144 2097 3247 2200 ne
rect 3247 2097 3456 2200
tri 3456 2097 3559 2200 sw
tri 3694 2097 3797 2200 ne
rect 3797 2097 4006 2200
tri 4006 2097 4109 2200 sw
tri 4244 2097 4347 2200 ne
rect 4347 2097 4556 2200
tri 4556 2097 4659 2200 sw
tri 4794 2097 4897 2200 ne
rect 4897 2097 5106 2200
tri 5106 2097 5209 2200 sw
tri 5344 2097 5447 2200 ne
rect 5447 2097 5656 2200
tri 5656 2097 5759 2200 sw
tri 5894 2097 5997 2200 ne
rect 5997 2097 6206 2200
tri 6206 2097 6309 2200 sw
tri 6444 2097 6547 2200 ne
rect 6547 2097 6756 2200
tri 6756 2097 6859 2200 sw
tri 6994 2097 7097 2200 ne
rect 7097 2097 7306 2200
tri 7306 2097 7409 2200 sw
tri 7544 2097 7647 2200 ne
rect 7647 2097 7856 2200
tri 7856 2097 7959 2200 sw
tri 8094 2097 8197 2200 ne
rect 8197 2097 8406 2200
tri 8406 2097 8509 2200 sw
tri 8644 2097 8747 2200 ne
rect 8747 2097 8956 2200
tri 8956 2097 9059 2200 sw
tri 9194 2097 9297 2200 ne
rect 9297 2097 9506 2200
tri 9506 2097 9609 2200 sw
tri 9744 2097 9847 2200 ne
rect 9847 2097 10056 2200
tri 10056 2097 10159 2200 sw
tri 10294 2097 10397 2200 ne
rect 10397 2097 10606 2200
tri 10606 2097 10709 2200 sw
tri 10844 2097 10947 2200 ne
rect 10947 2097 11156 2200
tri 11156 2097 11259 2200 sw
tri 11394 2097 11497 2200 ne
rect 11497 2097 11706 2200
tri 11706 2097 11809 2200 sw
tri 11944 2097 12047 2200 ne
rect 12047 2097 12256 2200
tri 12256 2097 12359 2200 sw
tri 12494 2097 12597 2200 ne
rect 12597 2097 12806 2200
tri 12806 2097 12909 2200 sw
tri 13044 2097 13147 2200 ne
rect 13147 2097 13356 2200
tri 13356 2097 13459 2200 sw
tri 13594 2097 13697 2200 ne
rect 13697 2097 15775 2200
rect -1025 1960 -291 2097
tri -291 1960 -154 2097 sw
tri -53 1960 84 2097 ne
rect 84 1960 259 2097
tri 259 1960 396 2097 sw
tri 497 1960 634 2097 ne
rect 634 1960 809 2097
tri 809 1960 946 2097 sw
tri 1047 1960 1184 2097 ne
rect 1184 1960 1359 2097
tri 1359 1960 1496 2097 sw
tri 1597 1960 1734 2097 ne
rect 1734 1960 1909 2097
tri 1909 1960 2046 2097 sw
tri 2147 1960 2284 2097 ne
rect 2284 1960 2459 2097
tri 2459 1960 2596 2097 sw
tri 2697 1960 2834 2097 ne
rect 2834 1960 3009 2097
tri 3009 1960 3146 2097 sw
tri 3247 1960 3384 2097 ne
rect 3384 1960 3559 2097
tri 3559 1960 3696 2097 sw
tri 3797 1960 3934 2097 ne
rect 3934 1960 4109 2097
tri 4109 1960 4246 2097 sw
tri 4347 1960 4484 2097 ne
rect 4484 1960 4659 2097
tri 4659 1960 4796 2097 sw
tri 4897 1960 5034 2097 ne
rect 5034 1960 5209 2097
tri 5209 1960 5346 2097 sw
tri 5447 1960 5584 2097 ne
rect 5584 1960 5759 2097
tri 5759 1960 5896 2097 sw
tri 5997 1960 6134 2097 ne
rect 6134 1960 6309 2097
tri 6309 1960 6446 2097 sw
tri 6547 1960 6684 2097 ne
rect 6684 1960 6859 2097
tri 6859 1960 6996 2097 sw
tri 7097 1960 7234 2097 ne
rect 7234 1960 7409 2097
tri 7409 1960 7546 2097 sw
tri 7647 1960 7784 2097 ne
rect 7784 1960 7959 2097
tri 7959 1960 8096 2097 sw
tri 8197 1960 8334 2097 ne
rect 8334 1960 8509 2097
tri 8509 1960 8646 2097 sw
tri 8747 1960 8884 2097 ne
rect 8884 1960 9059 2097
tri 9059 1960 9196 2097 sw
tri 9297 1960 9434 2097 ne
rect 9434 1960 9609 2097
tri 9609 1960 9746 2097 sw
tri 9847 1960 9984 2097 ne
rect 9984 1960 10159 2097
tri 10159 1960 10296 2097 sw
tri 10397 1960 10534 2097 ne
rect 10534 1960 10709 2097
tri 10709 1960 10846 2097 sw
tri 10947 1960 11084 2097 ne
rect 11084 1960 11259 2097
tri 11259 1960 11396 2097 sw
tri 11497 1960 11634 2097 ne
rect 11634 1960 11809 2097
tri 11809 1960 11946 2097 sw
tri 12047 1960 12184 2097 ne
rect 12184 1960 12359 2097
tri 12359 1960 12496 2097 sw
tri 12597 1960 12734 2097 ne
rect 12734 1960 12909 2097
tri 12909 1960 13046 2097 sw
tri 13147 1960 13284 2097 ne
rect 13284 1960 13459 2097
tri 13459 1960 13596 2097 sw
rect -1025 1942 -310 1960
tri -448 1840 -346 1942 ne
rect -346 1840 -310 1942
rect -190 1840 -154 1960
rect -2525 1650 -447 1703
tri -447 1650 -394 1703 sw
tri -346 1650 -156 1840 ne
rect -156 1806 -154 1840
tri -154 1806 0 1960 sw
tri 84 1806 238 1960 ne
rect 238 1840 240 1960
rect 360 1840 396 1960
rect 238 1806 396 1840
tri 396 1806 550 1960 sw
tri 634 1806 788 1960 ne
rect 788 1840 790 1960
rect 910 1840 946 1960
rect 788 1806 946 1840
tri 946 1806 1100 1960 sw
tri 1184 1806 1338 1960 ne
rect 1338 1840 1340 1960
rect 1460 1840 1496 1960
rect 1338 1806 1496 1840
tri 1496 1806 1650 1960 sw
tri 1734 1806 1888 1960 ne
rect 1888 1840 1890 1960
rect 2010 1840 2046 1960
rect 1888 1806 2046 1840
tri 2046 1806 2200 1960 sw
tri 2284 1806 2438 1960 ne
rect 2438 1840 2440 1960
rect 2560 1840 2596 1960
rect 2438 1806 2596 1840
tri 2596 1806 2750 1960 sw
tri 2834 1806 2988 1960 ne
rect 2988 1840 2990 1960
rect 3110 1840 3146 1960
rect 2988 1806 3146 1840
tri 3146 1806 3300 1960 sw
tri 3384 1806 3538 1960 ne
rect 3538 1840 3540 1960
rect 3660 1840 3696 1960
rect 3538 1806 3696 1840
tri 3696 1806 3850 1960 sw
tri 3934 1806 4088 1960 ne
rect 4088 1840 4090 1960
rect 4210 1840 4246 1960
rect 4088 1806 4246 1840
tri 4246 1806 4400 1960 sw
tri 4484 1806 4638 1960 ne
rect 4638 1840 4640 1960
rect 4760 1840 4796 1960
rect 4638 1806 4796 1840
tri 4796 1806 4950 1960 sw
tri 5034 1806 5188 1960 ne
rect 5188 1840 5190 1960
rect 5310 1840 5346 1960
rect 5188 1806 5346 1840
tri 5346 1806 5500 1960 sw
tri 5584 1806 5738 1960 ne
rect 5738 1840 5740 1960
rect 5860 1840 5896 1960
rect 5738 1806 5896 1840
tri 5896 1806 6050 1960 sw
tri 6134 1806 6288 1960 ne
rect 6288 1840 6290 1960
rect 6410 1840 6446 1960
rect 6288 1806 6446 1840
tri 6446 1806 6600 1960 sw
tri 6684 1806 6838 1960 ne
rect 6838 1840 6840 1960
rect 6960 1840 6996 1960
rect 6838 1806 6996 1840
tri 6996 1806 7150 1960 sw
tri 7234 1806 7388 1960 ne
rect 7388 1840 7390 1960
rect 7510 1840 7546 1960
rect 7388 1806 7546 1840
tri 7546 1806 7700 1960 sw
tri 7784 1806 7938 1960 ne
rect 7938 1840 7940 1960
rect 8060 1840 8096 1960
rect 7938 1806 8096 1840
tri 8096 1806 8250 1960 sw
tri 8334 1806 8488 1960 ne
rect 8488 1840 8490 1960
rect 8610 1840 8646 1960
rect 8488 1806 8646 1840
tri 8646 1806 8800 1960 sw
tri 8884 1806 9038 1960 ne
rect 9038 1840 9040 1960
rect 9160 1840 9196 1960
rect 9038 1806 9196 1840
tri 9196 1806 9350 1960 sw
tri 9434 1806 9588 1960 ne
rect 9588 1840 9590 1960
rect 9710 1840 9746 1960
rect 9588 1806 9746 1840
tri 9746 1806 9900 1960 sw
tri 9984 1806 10138 1960 ne
rect 10138 1840 10140 1960
rect 10260 1840 10296 1960
rect 10138 1806 10296 1840
tri 10296 1806 10450 1960 sw
tri 10534 1806 10688 1960 ne
rect 10688 1840 10690 1960
rect 10810 1840 10846 1960
rect 10688 1806 10846 1840
tri 10846 1806 11000 1960 sw
tri 11084 1806 11238 1960 ne
rect 11238 1840 11240 1960
rect 11360 1840 11396 1960
rect 11238 1806 11396 1840
tri 11396 1806 11550 1960 sw
tri 11634 1806 11788 1960 ne
rect 11788 1840 11790 1960
rect 11910 1840 11946 1960
rect 11788 1806 11946 1840
tri 11946 1806 12100 1960 sw
tri 12184 1806 12338 1960 ne
rect 12338 1840 12340 1960
rect 12460 1840 12496 1960
rect 12338 1806 12496 1840
tri 12496 1806 12650 1960 sw
tri 12734 1806 12888 1960 ne
rect 12888 1840 12890 1960
rect 13010 1840 13046 1960
rect 12888 1806 13046 1840
tri 13046 1806 13200 1960 sw
tri 13284 1806 13438 1960 ne
rect 13438 1840 13440 1960
rect 13560 1858 13596 1960
tri 13596 1858 13698 1960 sw
rect 13560 1840 14275 1858
rect 13438 1806 14275 1840
rect -156 1650 0 1806
tri 0 1650 156 1806 sw
tri 238 1650 394 1806 ne
rect 394 1650 550 1806
tri 550 1650 706 1806 sw
tri 788 1650 944 1806 ne
rect 944 1650 1100 1806
tri 1100 1650 1256 1806 sw
tri 1338 1650 1494 1806 ne
rect 1494 1650 1650 1806
tri 1650 1650 1806 1806 sw
tri 1888 1650 2044 1806 ne
rect 2044 1650 2200 1806
tri 2200 1650 2356 1806 sw
tri 2438 1650 2594 1806 ne
rect 2594 1650 2750 1806
tri 2750 1650 2906 1806 sw
tri 2988 1650 3144 1806 ne
rect 3144 1650 3300 1806
tri 3300 1650 3456 1806 sw
tri 3538 1650 3694 1806 ne
rect 3694 1650 3850 1806
tri 3850 1650 4006 1806 sw
tri 4088 1650 4244 1806 ne
rect 4244 1650 4400 1806
tri 4400 1650 4556 1806 sw
tri 4638 1650 4794 1806 ne
rect 4794 1650 4950 1806
tri 4950 1650 5106 1806 sw
tri 5188 1650 5344 1806 ne
rect 5344 1650 5500 1806
tri 5500 1650 5656 1806 sw
tri 5738 1650 5894 1806 ne
rect 5894 1650 6050 1806
tri 6050 1650 6206 1806 sw
tri 6288 1650 6444 1806 ne
rect 6444 1650 6600 1806
tri 6600 1650 6756 1806 sw
tri 6838 1650 6994 1806 ne
rect 6994 1650 7150 1806
tri 7150 1650 7306 1806 sw
tri 7388 1650 7544 1806 ne
rect 7544 1650 7700 1806
tri 7700 1650 7856 1806 sw
tri 7938 1650 8094 1806 ne
rect 8094 1650 8250 1806
tri 8250 1650 8406 1806 sw
tri 8488 1650 8644 1806 ne
rect 8644 1650 8800 1806
tri 8800 1650 8956 1806 sw
tri 9038 1650 9194 1806 ne
rect 9194 1650 9350 1806
tri 9350 1650 9506 1806 sw
tri 9588 1650 9744 1806 ne
rect 9744 1650 9900 1806
tri 9900 1650 10056 1806 sw
tri 10138 1650 10294 1806 ne
rect 10294 1650 10450 1806
tri 10450 1650 10606 1806 sw
tri 10688 1650 10844 1806 ne
rect 10844 1650 11000 1806
tri 11000 1650 11156 1806 sw
tri 11238 1650 11394 1806 ne
rect 11394 1650 11550 1806
tri 11550 1650 11706 1806 sw
tri 11788 1650 11944 1806 ne
rect 11944 1650 12100 1806
tri 12100 1650 12256 1806 sw
tri 12338 1650 12494 1806 ne
rect 12494 1650 12650 1806
tri 12650 1650 12806 1806 sw
tri 12888 1650 13044 1806 ne
rect 13044 1650 13200 1806
tri 13200 1650 13356 1806 sw
tri 13438 1650 13594 1806 ne
rect 13594 1650 14275 1806
rect -2525 1547 -394 1650
tri -394 1547 -291 1650 sw
tri -156 1547 -53 1650 ne
rect -53 1547 156 1650
tri 156 1547 259 1650 sw
tri 394 1547 497 1650 ne
rect 497 1547 706 1650
tri 706 1547 809 1650 sw
tri 944 1547 1047 1650 ne
rect 1047 1547 1256 1650
tri 1256 1547 1359 1650 sw
tri 1494 1547 1597 1650 ne
rect 1597 1547 1806 1650
tri 1806 1547 1909 1650 sw
tri 2044 1547 2147 1650 ne
rect 2147 1547 2356 1650
tri 2356 1547 2459 1650 sw
tri 2594 1547 2697 1650 ne
rect 2697 1547 2906 1650
tri 2906 1547 3009 1650 sw
tri 3144 1547 3247 1650 ne
rect 3247 1547 3456 1650
tri 3456 1547 3559 1650 sw
tri 3694 1547 3797 1650 ne
rect 3797 1547 4006 1650
tri 4006 1547 4109 1650 sw
tri 4244 1547 4347 1650 ne
rect 4347 1547 4556 1650
tri 4556 1547 4659 1650 sw
tri 4794 1547 4897 1650 ne
rect 4897 1547 5106 1650
tri 5106 1547 5209 1650 sw
tri 5344 1547 5447 1650 ne
rect 5447 1547 5656 1650
tri 5656 1547 5759 1650 sw
tri 5894 1547 5997 1650 ne
rect 5997 1547 6206 1650
tri 6206 1547 6309 1650 sw
tri 6444 1547 6547 1650 ne
rect 6547 1547 6756 1650
tri 6756 1547 6859 1650 sw
tri 6994 1547 7097 1650 ne
rect 7097 1547 7306 1650
tri 7306 1547 7409 1650 sw
tri 7544 1547 7647 1650 ne
rect 7647 1547 7856 1650
tri 7856 1547 7959 1650 sw
tri 8094 1547 8197 1650 ne
rect 8197 1547 8406 1650
tri 8406 1547 8509 1650 sw
tri 8644 1547 8747 1650 ne
rect 8747 1547 8956 1650
tri 8956 1547 9059 1650 sw
tri 9194 1547 9297 1650 ne
rect 9297 1547 9506 1650
tri 9506 1547 9609 1650 sw
tri 9744 1547 9847 1650 ne
rect 9847 1547 10056 1650
tri 10056 1547 10159 1650 sw
tri 10294 1547 10397 1650 ne
rect 10397 1547 10606 1650
tri 10606 1547 10709 1650 sw
tri 10844 1547 10947 1650 ne
rect 10947 1547 11156 1650
tri 11156 1547 11259 1650 sw
tri 11394 1547 11497 1650 ne
rect 11497 1547 11706 1650
tri 11706 1547 11809 1650 sw
tri 11944 1547 12047 1650 ne
rect 12047 1547 12256 1650
tri 12256 1547 12359 1650 sw
tri 12494 1547 12597 1650 ne
rect 12597 1547 12806 1650
tri 12806 1547 12909 1650 sw
tri 13044 1547 13147 1650 ne
rect 13147 1547 13356 1650
tri 13356 1547 13459 1650 sw
tri 13594 1547 13697 1650 ne
rect 13697 1547 14275 1650
rect -2525 1410 -291 1547
tri -291 1410 -154 1547 sw
tri -53 1410 84 1547 ne
rect 84 1410 259 1547
tri 259 1410 396 1547 sw
tri 497 1410 634 1547 ne
rect 634 1410 809 1547
tri 809 1410 946 1547 sw
tri 1047 1410 1184 1547 ne
rect 1184 1410 1359 1547
tri 1359 1410 1496 1547 sw
tri 1597 1410 1734 1547 ne
rect 1734 1410 1909 1547
tri 1909 1410 2046 1547 sw
tri 2147 1410 2284 1547 ne
rect 2284 1410 2459 1547
tri 2459 1410 2596 1547 sw
tri 2697 1410 2834 1547 ne
rect 2834 1410 3009 1547
tri 3009 1410 3146 1547 sw
tri 3247 1410 3384 1547 ne
rect 3384 1410 3559 1547
tri 3559 1410 3696 1547 sw
tri 3797 1410 3934 1547 ne
rect 3934 1410 4109 1547
tri 4109 1410 4246 1547 sw
tri 4347 1410 4484 1547 ne
rect 4484 1410 4659 1547
tri 4659 1410 4796 1547 sw
tri 4897 1410 5034 1547 ne
rect 5034 1410 5209 1547
tri 5209 1410 5346 1547 sw
tri 5447 1410 5584 1547 ne
rect 5584 1410 5759 1547
tri 5759 1410 5896 1547 sw
tri 5997 1410 6134 1547 ne
rect 6134 1410 6309 1547
tri 6309 1410 6446 1547 sw
tri 6547 1410 6684 1547 ne
rect 6684 1410 6859 1547
tri 6859 1410 6996 1547 sw
tri 7097 1410 7234 1547 ne
rect 7234 1410 7409 1547
tri 7409 1410 7546 1547 sw
tri 7647 1410 7784 1547 ne
rect 7784 1410 7959 1547
tri 7959 1410 8096 1547 sw
tri 8197 1410 8334 1547 ne
rect 8334 1410 8509 1547
tri 8509 1410 8646 1547 sw
tri 8747 1410 8884 1547 ne
rect 8884 1410 9059 1547
tri 9059 1410 9196 1547 sw
tri 9297 1410 9434 1547 ne
rect 9434 1410 9609 1547
tri 9609 1410 9746 1547 sw
tri 9847 1410 9984 1547 ne
rect 9984 1410 10159 1547
tri 10159 1410 10296 1547 sw
tri 10397 1410 10534 1547 ne
rect 10534 1410 10709 1547
tri 10709 1410 10846 1547 sw
tri 10947 1410 11084 1547 ne
rect 11084 1410 11259 1547
tri 11259 1410 11396 1547 sw
tri 11497 1410 11634 1547 ne
rect 11634 1410 11809 1547
tri 11809 1410 11946 1547 sw
tri 12047 1410 12184 1547 ne
rect 12184 1410 12359 1547
tri 12359 1410 12496 1547 sw
tri 12597 1410 12734 1547 ne
rect 12734 1410 12909 1547
tri 12909 1410 13046 1547 sw
tri 13147 1410 13284 1547 ne
rect 13284 1410 13459 1547
tri 13459 1410 13596 1547 sw
rect -2525 1392 -310 1410
rect -2525 603 -1525 1392
tri -448 1290 -346 1392 ne
rect -346 1290 -310 1392
rect -190 1290 -154 1410
rect -1025 1100 -447 1153
tri -447 1100 -394 1153 sw
tri -346 1100 -156 1290 ne
rect -156 1256 -154 1290
tri -154 1256 0 1410 sw
tri 84 1256 238 1410 ne
rect 238 1290 240 1410
rect 360 1290 396 1410
rect 238 1256 396 1290
tri 396 1256 550 1410 sw
tri 634 1256 788 1410 ne
rect 788 1290 790 1410
rect 910 1290 946 1410
rect 788 1256 946 1290
tri 946 1256 1100 1410 sw
tri 1184 1256 1338 1410 ne
rect 1338 1290 1340 1410
rect 1460 1290 1496 1410
rect 1338 1256 1496 1290
tri 1496 1256 1650 1410 sw
tri 1734 1256 1888 1410 ne
rect 1888 1290 1890 1410
rect 2010 1290 2046 1410
rect 1888 1256 2046 1290
tri 2046 1256 2200 1410 sw
tri 2284 1256 2438 1410 ne
rect 2438 1290 2440 1410
rect 2560 1290 2596 1410
rect 2438 1256 2596 1290
tri 2596 1256 2750 1410 sw
tri 2834 1256 2988 1410 ne
rect 2988 1290 2990 1410
rect 3110 1290 3146 1410
rect 2988 1256 3146 1290
tri 3146 1256 3300 1410 sw
tri 3384 1256 3538 1410 ne
rect 3538 1290 3540 1410
rect 3660 1290 3696 1410
rect 3538 1256 3696 1290
tri 3696 1256 3850 1410 sw
tri 3934 1256 4088 1410 ne
rect 4088 1290 4090 1410
rect 4210 1290 4246 1410
rect 4088 1256 4246 1290
tri 4246 1256 4400 1410 sw
tri 4484 1256 4638 1410 ne
rect 4638 1290 4640 1410
rect 4760 1290 4796 1410
rect 4638 1256 4796 1290
tri 4796 1256 4950 1410 sw
tri 5034 1256 5188 1410 ne
rect 5188 1290 5190 1410
rect 5310 1290 5346 1410
rect 5188 1256 5346 1290
tri 5346 1256 5500 1410 sw
tri 5584 1256 5738 1410 ne
rect 5738 1290 5740 1410
rect 5860 1290 5896 1410
rect 5738 1256 5896 1290
tri 5896 1256 6050 1410 sw
tri 6134 1256 6288 1410 ne
rect 6288 1290 6290 1410
rect 6410 1290 6446 1410
rect 6288 1256 6446 1290
tri 6446 1256 6600 1410 sw
tri 6684 1256 6838 1410 ne
rect 6838 1290 6840 1410
rect 6960 1290 6996 1410
rect 6838 1256 6996 1290
tri 6996 1256 7150 1410 sw
tri 7234 1256 7388 1410 ne
rect 7388 1290 7390 1410
rect 7510 1290 7546 1410
rect 7388 1256 7546 1290
tri 7546 1256 7700 1410 sw
tri 7784 1256 7938 1410 ne
rect 7938 1290 7940 1410
rect 8060 1290 8096 1410
rect 7938 1256 8096 1290
tri 8096 1256 8250 1410 sw
tri 8334 1256 8488 1410 ne
rect 8488 1290 8490 1410
rect 8610 1290 8646 1410
rect 8488 1256 8646 1290
tri 8646 1256 8800 1410 sw
tri 8884 1256 9038 1410 ne
rect 9038 1290 9040 1410
rect 9160 1290 9196 1410
rect 9038 1256 9196 1290
tri 9196 1256 9350 1410 sw
tri 9434 1256 9588 1410 ne
rect 9588 1290 9590 1410
rect 9710 1290 9746 1410
rect 9588 1256 9746 1290
tri 9746 1256 9900 1410 sw
tri 9984 1256 10138 1410 ne
rect 10138 1290 10140 1410
rect 10260 1290 10296 1410
rect 10138 1256 10296 1290
tri 10296 1256 10450 1410 sw
tri 10534 1256 10688 1410 ne
rect 10688 1290 10690 1410
rect 10810 1290 10846 1410
rect 10688 1256 10846 1290
tri 10846 1256 11000 1410 sw
tri 11084 1256 11238 1410 ne
rect 11238 1290 11240 1410
rect 11360 1290 11396 1410
rect 11238 1256 11396 1290
tri 11396 1256 11550 1410 sw
tri 11634 1256 11788 1410 ne
rect 11788 1290 11790 1410
rect 11910 1290 11946 1410
rect 11788 1256 11946 1290
tri 11946 1256 12100 1410 sw
tri 12184 1256 12338 1410 ne
rect 12338 1290 12340 1410
rect 12460 1290 12496 1410
rect 12338 1256 12496 1290
tri 12496 1256 12650 1410 sw
tri 12734 1256 12888 1410 ne
rect 12888 1290 12890 1410
rect 13010 1290 13046 1410
rect 12888 1256 13046 1290
tri 13046 1256 13200 1410 sw
tri 13284 1256 13438 1410 ne
rect 13438 1290 13440 1410
rect 13560 1308 13596 1410
tri 13596 1308 13698 1410 sw
rect 14775 1308 15775 2097
rect 13560 1290 15775 1308
rect 13438 1256 15775 1290
rect -156 1100 0 1256
tri 0 1100 156 1256 sw
tri 238 1100 394 1256 ne
rect 394 1100 550 1256
tri 550 1100 706 1256 sw
tri 788 1100 944 1256 ne
rect 944 1100 1100 1256
tri 1100 1100 1256 1256 sw
tri 1338 1100 1494 1256 ne
rect 1494 1100 1650 1256
tri 1650 1100 1806 1256 sw
tri 1888 1100 2044 1256 ne
rect 2044 1100 2200 1256
tri 2200 1100 2356 1256 sw
tri 2438 1100 2594 1256 ne
rect 2594 1100 2750 1256
tri 2750 1100 2906 1256 sw
tri 2988 1100 3144 1256 ne
rect 3144 1100 3300 1256
tri 3300 1100 3456 1256 sw
tri 3538 1100 3694 1256 ne
rect 3694 1100 3850 1256
tri 3850 1100 4006 1256 sw
tri 4088 1100 4244 1256 ne
rect 4244 1100 4400 1256
tri 4400 1100 4556 1256 sw
tri 4638 1100 4794 1256 ne
rect 4794 1100 4950 1256
tri 4950 1100 5106 1256 sw
tri 5188 1100 5344 1256 ne
rect 5344 1100 5500 1256
tri 5500 1100 5656 1256 sw
tri 5738 1100 5894 1256 ne
rect 5894 1100 6050 1256
tri 6050 1100 6206 1256 sw
tri 6288 1100 6444 1256 ne
rect 6444 1100 6600 1256
tri 6600 1100 6756 1256 sw
tri 6838 1100 6994 1256 ne
rect 6994 1100 7150 1256
tri 7150 1100 7306 1256 sw
tri 7388 1100 7544 1256 ne
rect 7544 1100 7700 1256
tri 7700 1100 7856 1256 sw
tri 7938 1100 8094 1256 ne
rect 8094 1100 8250 1256
tri 8250 1100 8406 1256 sw
tri 8488 1100 8644 1256 ne
rect 8644 1100 8800 1256
tri 8800 1100 8956 1256 sw
tri 9038 1100 9194 1256 ne
rect 9194 1100 9350 1256
tri 9350 1100 9506 1256 sw
tri 9588 1100 9744 1256 ne
rect 9744 1100 9900 1256
tri 9900 1100 10056 1256 sw
tri 10138 1100 10294 1256 ne
rect 10294 1100 10450 1256
tri 10450 1100 10606 1256 sw
tri 10688 1100 10844 1256 ne
rect 10844 1100 11000 1256
tri 11000 1100 11156 1256 sw
tri 11238 1100 11394 1256 ne
rect 11394 1100 11550 1256
tri 11550 1100 11706 1256 sw
tri 11788 1100 11944 1256 ne
rect 11944 1100 12100 1256
tri 12100 1100 12256 1256 sw
tri 12338 1100 12494 1256 ne
rect 12494 1100 12650 1256
tri 12650 1100 12806 1256 sw
tri 12888 1100 13044 1256 ne
rect 13044 1100 13200 1256
tri 13200 1100 13356 1256 sw
tri 13438 1100 13594 1256 ne
rect 13594 1100 15775 1256
rect -1025 997 -394 1100
tri -394 997 -291 1100 sw
tri -156 997 -53 1100 ne
rect -53 997 156 1100
tri 156 997 259 1100 sw
tri 394 997 497 1100 ne
rect 497 997 706 1100
tri 706 997 809 1100 sw
tri 944 997 1047 1100 ne
rect 1047 997 1256 1100
tri 1256 997 1359 1100 sw
tri 1494 997 1597 1100 ne
rect 1597 997 1806 1100
tri 1806 997 1909 1100 sw
tri 2044 997 2147 1100 ne
rect 2147 997 2356 1100
tri 2356 997 2459 1100 sw
tri 2594 997 2697 1100 ne
rect 2697 997 2906 1100
tri 2906 997 3009 1100 sw
tri 3144 997 3247 1100 ne
rect 3247 997 3456 1100
tri 3456 997 3559 1100 sw
tri 3694 997 3797 1100 ne
rect 3797 997 4006 1100
tri 4006 997 4109 1100 sw
tri 4244 997 4347 1100 ne
rect 4347 997 4556 1100
tri 4556 997 4659 1100 sw
tri 4794 997 4897 1100 ne
rect 4897 997 5106 1100
tri 5106 997 5209 1100 sw
tri 5344 997 5447 1100 ne
rect 5447 997 5656 1100
tri 5656 997 5759 1100 sw
tri 5894 997 5997 1100 ne
rect 5997 997 6206 1100
tri 6206 997 6309 1100 sw
tri 6444 997 6547 1100 ne
rect 6547 997 6756 1100
tri 6756 997 6859 1100 sw
tri 6994 997 7097 1100 ne
rect 7097 997 7306 1100
tri 7306 997 7409 1100 sw
tri 7544 997 7647 1100 ne
rect 7647 997 7856 1100
tri 7856 997 7959 1100 sw
tri 8094 997 8197 1100 ne
rect 8197 997 8406 1100
tri 8406 997 8509 1100 sw
tri 8644 997 8747 1100 ne
rect 8747 997 8956 1100
tri 8956 997 9059 1100 sw
tri 9194 997 9297 1100 ne
rect 9297 997 9506 1100
tri 9506 997 9609 1100 sw
tri 9744 997 9847 1100 ne
rect 9847 997 10056 1100
tri 10056 997 10159 1100 sw
tri 10294 997 10397 1100 ne
rect 10397 997 10606 1100
tri 10606 997 10709 1100 sw
tri 10844 997 10947 1100 ne
rect 10947 997 11156 1100
tri 11156 997 11259 1100 sw
tri 11394 997 11497 1100 ne
rect 11497 997 11706 1100
tri 11706 997 11809 1100 sw
tri 11944 997 12047 1100 ne
rect 12047 997 12256 1100
tri 12256 997 12359 1100 sw
tri 12494 997 12597 1100 ne
rect 12597 997 12806 1100
tri 12806 997 12909 1100 sw
tri 13044 997 13147 1100 ne
rect 13147 997 13356 1100
tri 13356 997 13459 1100 sw
tri 13594 997 13697 1100 ne
rect 13697 997 15775 1100
rect -1025 860 -291 997
tri -291 860 -154 997 sw
tri -53 860 84 997 ne
rect 84 860 259 997
tri 259 860 396 997 sw
tri 497 860 634 997 ne
rect 634 860 809 997
tri 809 860 946 997 sw
tri 1047 860 1184 997 ne
rect 1184 860 1359 997
tri 1359 860 1496 997 sw
tri 1597 860 1734 997 ne
rect 1734 860 1909 997
tri 1909 860 2046 997 sw
tri 2147 860 2284 997 ne
rect 2284 860 2459 997
tri 2459 860 2596 997 sw
tri 2697 860 2834 997 ne
rect 2834 860 3009 997
tri 3009 860 3146 997 sw
tri 3247 860 3384 997 ne
rect 3384 860 3559 997
tri 3559 860 3696 997 sw
tri 3797 860 3934 997 ne
rect 3934 860 4109 997
tri 4109 860 4246 997 sw
tri 4347 860 4484 997 ne
rect 4484 860 4659 997
tri 4659 860 4796 997 sw
tri 4897 860 5034 997 ne
rect 5034 860 5209 997
tri 5209 860 5346 997 sw
tri 5447 860 5584 997 ne
rect 5584 860 5759 997
tri 5759 860 5896 997 sw
tri 5997 860 6134 997 ne
rect 6134 860 6309 997
tri 6309 860 6446 997 sw
tri 6547 860 6684 997 ne
rect 6684 860 6859 997
tri 6859 860 6996 997 sw
tri 7097 860 7234 997 ne
rect 7234 860 7409 997
tri 7409 860 7546 997 sw
tri 7647 860 7784 997 ne
rect 7784 860 7959 997
tri 7959 860 8096 997 sw
tri 8197 860 8334 997 ne
rect 8334 860 8509 997
tri 8509 860 8646 997 sw
tri 8747 860 8884 997 ne
rect 8884 860 9059 997
tri 9059 860 9196 997 sw
tri 9297 860 9434 997 ne
rect 9434 860 9609 997
tri 9609 860 9746 997 sw
tri 9847 860 9984 997 ne
rect 9984 860 10159 997
tri 10159 860 10296 997 sw
tri 10397 860 10534 997 ne
rect 10534 860 10709 997
tri 10709 860 10846 997 sw
tri 10947 860 11084 997 ne
rect 11084 860 11259 997
tri 11259 860 11396 997 sw
tri 11497 860 11634 997 ne
rect 11634 860 11809 997
tri 11809 860 11946 997 sw
tri 12047 860 12184 997 ne
rect 12184 860 12359 997
tri 12359 860 12496 997 sw
tri 12597 860 12734 997 ne
rect 12734 860 12909 997
tri 12909 860 13046 997 sw
tri 13147 860 13284 997 ne
rect 13284 860 13459 997
tri 13459 860 13596 997 sw
rect -1025 842 -310 860
tri -448 740 -346 842 ne
rect -346 740 -310 842
rect -190 740 -154 860
rect -2525 550 -447 603
tri -447 550 -394 603 sw
tri -346 550 -156 740 ne
rect -156 706 -154 740
tri -154 706 0 860 sw
tri 84 706 238 860 ne
rect 238 740 240 860
rect 360 740 396 860
rect 238 706 396 740
tri 396 706 550 860 sw
tri 634 706 788 860 ne
rect 788 740 790 860
rect 910 740 946 860
rect 788 706 946 740
tri 946 706 1100 860 sw
tri 1184 706 1338 860 ne
rect 1338 740 1340 860
rect 1460 740 1496 860
rect 1338 706 1496 740
tri 1496 706 1650 860 sw
tri 1734 706 1888 860 ne
rect 1888 740 1890 860
rect 2010 740 2046 860
rect 1888 706 2046 740
tri 2046 706 2200 860 sw
tri 2284 706 2438 860 ne
rect 2438 740 2440 860
rect 2560 740 2596 860
rect 2438 706 2596 740
tri 2596 706 2750 860 sw
tri 2834 706 2988 860 ne
rect 2988 740 2990 860
rect 3110 740 3146 860
rect 2988 706 3146 740
tri 3146 706 3300 860 sw
tri 3384 706 3538 860 ne
rect 3538 740 3540 860
rect 3660 740 3696 860
rect 3538 706 3696 740
tri 3696 706 3850 860 sw
tri 3934 706 4088 860 ne
rect 4088 740 4090 860
rect 4210 740 4246 860
rect 4088 706 4246 740
tri 4246 706 4400 860 sw
tri 4484 706 4638 860 ne
rect 4638 740 4640 860
rect 4760 740 4796 860
rect 4638 706 4796 740
tri 4796 706 4950 860 sw
tri 5034 706 5188 860 ne
rect 5188 740 5190 860
rect 5310 740 5346 860
rect 5188 706 5346 740
tri 5346 706 5500 860 sw
tri 5584 706 5738 860 ne
rect 5738 740 5740 860
rect 5860 740 5896 860
rect 5738 706 5896 740
tri 5896 706 6050 860 sw
tri 6134 706 6288 860 ne
rect 6288 740 6290 860
rect 6410 740 6446 860
rect 6288 706 6446 740
tri 6446 706 6600 860 sw
tri 6684 706 6838 860 ne
rect 6838 740 6840 860
rect 6960 740 6996 860
rect 6838 706 6996 740
tri 6996 706 7150 860 sw
tri 7234 706 7388 860 ne
rect 7388 740 7390 860
rect 7510 740 7546 860
rect 7388 706 7546 740
tri 7546 706 7700 860 sw
tri 7784 706 7938 860 ne
rect 7938 740 7940 860
rect 8060 740 8096 860
rect 7938 706 8096 740
tri 8096 706 8250 860 sw
tri 8334 706 8488 860 ne
rect 8488 740 8490 860
rect 8610 740 8646 860
rect 8488 706 8646 740
tri 8646 706 8800 860 sw
tri 8884 706 9038 860 ne
rect 9038 740 9040 860
rect 9160 740 9196 860
rect 9038 706 9196 740
tri 9196 706 9350 860 sw
tri 9434 706 9588 860 ne
rect 9588 740 9590 860
rect 9710 740 9746 860
rect 9588 706 9746 740
tri 9746 706 9900 860 sw
tri 9984 706 10138 860 ne
rect 10138 740 10140 860
rect 10260 740 10296 860
rect 10138 706 10296 740
tri 10296 706 10450 860 sw
tri 10534 706 10688 860 ne
rect 10688 740 10690 860
rect 10810 740 10846 860
rect 10688 706 10846 740
tri 10846 706 11000 860 sw
tri 11084 706 11238 860 ne
rect 11238 740 11240 860
rect 11360 740 11396 860
rect 11238 706 11396 740
tri 11396 706 11550 860 sw
tri 11634 706 11788 860 ne
rect 11788 740 11790 860
rect 11910 740 11946 860
rect 11788 706 11946 740
tri 11946 706 12100 860 sw
tri 12184 706 12338 860 ne
rect 12338 740 12340 860
rect 12460 740 12496 860
rect 12338 706 12496 740
tri 12496 706 12650 860 sw
tri 12734 706 12888 860 ne
rect 12888 740 12890 860
rect 13010 740 13046 860
rect 12888 706 13046 740
tri 13046 706 13200 860 sw
tri 13284 706 13438 860 ne
rect 13438 740 13440 860
rect 13560 758 13596 860
tri 13596 758 13698 860 sw
rect 13560 740 14275 758
rect 13438 706 14275 740
rect -156 550 0 706
tri 0 550 156 706 sw
tri 238 550 394 706 ne
rect 394 550 550 706
tri 550 550 706 706 sw
tri 788 550 944 706 ne
rect 944 550 1100 706
tri 1100 550 1256 706 sw
tri 1338 550 1494 706 ne
rect 1494 550 1650 706
tri 1650 550 1806 706 sw
tri 1888 550 2044 706 ne
rect 2044 550 2200 706
tri 2200 550 2356 706 sw
tri 2438 550 2594 706 ne
rect 2594 550 2750 706
tri 2750 550 2906 706 sw
tri 2988 550 3144 706 ne
rect 3144 550 3300 706
tri 3300 550 3456 706 sw
tri 3538 550 3694 706 ne
rect 3694 550 3850 706
tri 3850 550 4006 706 sw
tri 4088 550 4244 706 ne
rect 4244 550 4400 706
tri 4400 550 4556 706 sw
tri 4638 550 4794 706 ne
rect 4794 550 4950 706
tri 4950 550 5106 706 sw
tri 5188 550 5344 706 ne
rect 5344 550 5500 706
tri 5500 550 5656 706 sw
tri 5738 550 5894 706 ne
rect 5894 550 6050 706
tri 6050 550 6206 706 sw
tri 6288 550 6444 706 ne
rect 6444 550 6600 706
tri 6600 550 6756 706 sw
tri 6838 550 6994 706 ne
rect 6994 550 7150 706
tri 7150 550 7306 706 sw
tri 7388 550 7544 706 ne
rect 7544 550 7700 706
tri 7700 550 7856 706 sw
tri 7938 550 8094 706 ne
rect 8094 550 8250 706
tri 8250 550 8406 706 sw
tri 8488 550 8644 706 ne
rect 8644 550 8800 706
tri 8800 550 8956 706 sw
tri 9038 550 9194 706 ne
rect 9194 550 9350 706
tri 9350 550 9506 706 sw
tri 9588 550 9744 706 ne
rect 9744 550 9900 706
tri 9900 550 10056 706 sw
tri 10138 550 10294 706 ne
rect 10294 550 10450 706
tri 10450 550 10606 706 sw
tri 10688 550 10844 706 ne
rect 10844 550 11000 706
tri 11000 550 11156 706 sw
tri 11238 550 11394 706 ne
rect 11394 550 11550 706
tri 11550 550 11706 706 sw
tri 11788 550 11944 706 ne
rect 11944 550 12100 706
tri 12100 550 12256 706 sw
tri 12338 550 12494 706 ne
rect 12494 550 12650 706
tri 12650 550 12806 706 sw
tri 12888 550 13044 706 ne
rect 13044 550 13200 706
tri 13200 550 13356 706 sw
tri 13438 550 13594 706 ne
rect 13594 550 14275 706
rect -2525 447 -394 550
tri -394 447 -291 550 sw
tri -156 447 -53 550 ne
rect -53 447 156 550
tri 156 447 259 550 sw
tri 394 447 497 550 ne
rect 497 447 706 550
tri 706 447 809 550 sw
tri 944 447 1047 550 ne
rect 1047 447 1256 550
tri 1256 447 1359 550 sw
tri 1494 447 1597 550 ne
rect 1597 447 1806 550
tri 1806 447 1909 550 sw
tri 2044 447 2147 550 ne
rect 2147 447 2356 550
tri 2356 447 2459 550 sw
tri 2594 447 2697 550 ne
rect 2697 447 2906 550
tri 2906 447 3009 550 sw
tri 3144 447 3247 550 ne
rect 3247 447 3456 550
tri 3456 447 3559 550 sw
tri 3694 447 3797 550 ne
rect 3797 447 4006 550
tri 4006 447 4109 550 sw
tri 4244 447 4347 550 ne
rect 4347 447 4556 550
tri 4556 447 4659 550 sw
tri 4794 447 4897 550 ne
rect 4897 447 5106 550
tri 5106 447 5209 550 sw
tri 5344 447 5447 550 ne
rect 5447 447 5656 550
tri 5656 447 5759 550 sw
tri 5894 447 5997 550 ne
rect 5997 447 6206 550
tri 6206 447 6309 550 sw
tri 6444 447 6547 550 ne
rect 6547 447 6756 550
tri 6756 447 6859 550 sw
tri 6994 447 7097 550 ne
rect 7097 447 7306 550
tri 7306 447 7409 550 sw
tri 7544 447 7647 550 ne
rect 7647 447 7856 550
tri 7856 447 7959 550 sw
tri 8094 447 8197 550 ne
rect 8197 447 8406 550
tri 8406 447 8509 550 sw
tri 8644 447 8747 550 ne
rect 8747 447 8956 550
tri 8956 447 9059 550 sw
tri 9194 447 9297 550 ne
rect 9297 447 9506 550
tri 9506 447 9609 550 sw
tri 9744 447 9847 550 ne
rect 9847 447 10056 550
tri 10056 447 10159 550 sw
tri 10294 447 10397 550 ne
rect 10397 447 10606 550
tri 10606 447 10709 550 sw
tri 10844 447 10947 550 ne
rect 10947 447 11156 550
tri 11156 447 11259 550 sw
tri 11394 447 11497 550 ne
rect 11497 447 11706 550
tri 11706 447 11809 550 sw
tri 11944 447 12047 550 ne
rect 12047 447 12256 550
tri 12256 447 12359 550 sw
tri 12494 447 12597 550 ne
rect 12597 447 12806 550
tri 12806 447 12909 550 sw
tri 13044 447 13147 550 ne
rect 13147 447 13356 550
tri 13356 447 13459 550 sw
tri 13594 447 13697 550 ne
rect 13697 447 14275 550
rect -2525 310 -291 447
tri -291 310 -154 447 sw
tri -53 310 84 447 ne
rect 84 310 259 447
tri 259 310 396 447 sw
tri 497 310 634 447 ne
rect 634 310 809 447
tri 809 310 946 447 sw
tri 1047 310 1184 447 ne
rect 1184 310 1359 447
tri 1359 310 1496 447 sw
tri 1597 310 1734 447 ne
rect 1734 310 1909 447
tri 1909 310 2046 447 sw
tri 2147 310 2284 447 ne
rect 2284 310 2459 447
tri 2459 310 2596 447 sw
tri 2697 310 2834 447 ne
rect 2834 310 3009 447
tri 3009 310 3146 447 sw
tri 3247 310 3384 447 ne
rect 3384 310 3559 447
tri 3559 310 3696 447 sw
tri 3797 310 3934 447 ne
rect 3934 310 4109 447
tri 4109 310 4246 447 sw
tri 4347 310 4484 447 ne
rect 4484 310 4659 447
tri 4659 310 4796 447 sw
tri 4897 310 5034 447 ne
rect 5034 310 5209 447
tri 5209 310 5346 447 sw
tri 5447 310 5584 447 ne
rect 5584 310 5759 447
tri 5759 310 5896 447 sw
tri 5997 310 6134 447 ne
rect 6134 310 6309 447
tri 6309 310 6446 447 sw
tri 6547 310 6684 447 ne
rect 6684 310 6859 447
tri 6859 310 6996 447 sw
tri 7097 310 7234 447 ne
rect 7234 310 7409 447
tri 7409 310 7546 447 sw
tri 7647 310 7784 447 ne
rect 7784 310 7959 447
tri 7959 310 8096 447 sw
tri 8197 310 8334 447 ne
rect 8334 310 8509 447
tri 8509 310 8646 447 sw
tri 8747 310 8884 447 ne
rect 8884 310 9059 447
tri 9059 310 9196 447 sw
tri 9297 310 9434 447 ne
rect 9434 310 9609 447
tri 9609 310 9746 447 sw
tri 9847 310 9984 447 ne
rect 9984 310 10159 447
tri 10159 310 10296 447 sw
tri 10397 310 10534 447 ne
rect 10534 310 10709 447
tri 10709 310 10846 447 sw
tri 10947 310 11084 447 ne
rect 11084 310 11259 447
tri 11259 310 11396 447 sw
tri 11497 310 11634 447 ne
rect 11634 310 11809 447
tri 11809 310 11946 447 sw
tri 12047 310 12184 447 ne
rect 12184 310 12359 447
tri 12359 310 12496 447 sw
tri 12597 310 12734 447 ne
rect 12734 310 12909 447
tri 12909 310 13046 447 sw
tri 13147 310 13284 447 ne
rect 13284 310 13459 447
tri 13459 310 13596 447 sw
rect -2525 292 -310 310
rect -2525 -575 -1525 292
tri -448 190 -346 292 ne
rect -346 190 -310 292
rect -190 190 -154 310
rect -1025 0 -447 53
tri -447 0 -394 53 sw
tri -346 0 -156 190 ne
rect -156 156 -154 190
tri -154 156 0 310 sw
tri 84 156 238 310 ne
rect 238 190 240 310
rect 360 190 396 310
rect 238 156 396 190
tri 396 156 550 310 sw
tri 634 156 788 310 ne
rect 788 190 790 310
rect 910 190 946 310
rect 788 156 946 190
tri 946 156 1100 310 sw
tri 1184 156 1338 310 ne
rect 1338 190 1340 310
rect 1460 190 1496 310
rect 1338 156 1496 190
tri 1496 156 1650 310 sw
tri 1734 156 1888 310 ne
rect 1888 190 1890 310
rect 2010 190 2046 310
rect 1888 156 2046 190
tri 2046 156 2200 310 sw
tri 2284 156 2438 310 ne
rect 2438 190 2440 310
rect 2560 190 2596 310
rect 2438 156 2596 190
tri 2596 156 2750 310 sw
tri 2834 156 2988 310 ne
rect 2988 190 2990 310
rect 3110 190 3146 310
rect 2988 156 3146 190
tri 3146 156 3300 310 sw
tri 3384 156 3538 310 ne
rect 3538 190 3540 310
rect 3660 190 3696 310
rect 3538 156 3696 190
tri 3696 156 3850 310 sw
tri 3934 156 4088 310 ne
rect 4088 190 4090 310
rect 4210 190 4246 310
rect 4088 156 4246 190
tri 4246 156 4400 310 sw
tri 4484 156 4638 310 ne
rect 4638 190 4640 310
rect 4760 190 4796 310
rect 4638 156 4796 190
tri 4796 156 4950 310 sw
tri 5034 156 5188 310 ne
rect 5188 190 5190 310
rect 5310 190 5346 310
rect 5188 156 5346 190
tri 5346 156 5500 310 sw
tri 5584 156 5738 310 ne
rect 5738 190 5740 310
rect 5860 190 5896 310
rect 5738 156 5896 190
tri 5896 156 6050 310 sw
tri 6134 156 6288 310 ne
rect 6288 190 6290 310
rect 6410 190 6446 310
rect 6288 156 6446 190
tri 6446 156 6600 310 sw
tri 6684 156 6838 310 ne
rect 6838 190 6840 310
rect 6960 190 6996 310
rect 6838 156 6996 190
tri 6996 156 7150 310 sw
tri 7234 156 7388 310 ne
rect 7388 190 7390 310
rect 7510 190 7546 310
rect 7388 156 7546 190
tri 7546 156 7700 310 sw
tri 7784 156 7938 310 ne
rect 7938 190 7940 310
rect 8060 190 8096 310
rect 7938 156 8096 190
tri 8096 156 8250 310 sw
tri 8334 156 8488 310 ne
rect 8488 190 8490 310
rect 8610 190 8646 310
rect 8488 156 8646 190
tri 8646 156 8800 310 sw
tri 8884 156 9038 310 ne
rect 9038 190 9040 310
rect 9160 190 9196 310
rect 9038 156 9196 190
tri 9196 156 9350 310 sw
tri 9434 156 9588 310 ne
rect 9588 190 9590 310
rect 9710 190 9746 310
rect 9588 156 9746 190
tri 9746 156 9900 310 sw
tri 9984 156 10138 310 ne
rect 10138 190 10140 310
rect 10260 190 10296 310
rect 10138 156 10296 190
tri 10296 156 10450 310 sw
tri 10534 156 10688 310 ne
rect 10688 190 10690 310
rect 10810 190 10846 310
rect 10688 156 10846 190
tri 10846 156 11000 310 sw
tri 11084 156 11238 310 ne
rect 11238 190 11240 310
rect 11360 190 11396 310
rect 11238 156 11396 190
tri 11396 156 11550 310 sw
tri 11634 156 11788 310 ne
rect 11788 190 11790 310
rect 11910 190 11946 310
rect 11788 156 11946 190
tri 11946 156 12100 310 sw
tri 12184 156 12338 310 ne
rect 12338 190 12340 310
rect 12460 190 12496 310
rect 12338 156 12496 190
tri 12496 156 12650 310 sw
tri 12734 156 12888 310 ne
rect 12888 190 12890 310
rect 13010 190 13046 310
rect 12888 156 13046 190
tri 13046 156 13200 310 sw
tri 13284 156 13438 310 ne
rect 13438 190 13440 310
rect 13560 208 13596 310
tri 13596 208 13698 310 sw
rect 14775 208 15775 997
rect 13560 190 15775 208
rect 13438 156 15775 190
rect -156 0 0 156
tri 0 0 156 156 sw
tri 238 0 394 156 ne
rect 394 0 550 156
tri 550 0 706 156 sw
tri 788 0 944 156 ne
rect 944 0 1100 156
tri 1100 0 1256 156 sw
tri 1338 0 1494 156 ne
rect 1494 0 1650 156
tri 1650 0 1806 156 sw
tri 1888 0 2044 156 ne
rect 2044 0 2200 156
tri 2200 0 2356 156 sw
tri 2438 0 2594 156 ne
rect 2594 0 2750 156
tri 2750 0 2906 156 sw
tri 2988 0 3144 156 ne
rect 3144 0 3300 156
tri 3300 0 3456 156 sw
tri 3538 0 3694 156 ne
rect 3694 0 3850 156
tri 3850 0 4006 156 sw
tri 4088 0 4244 156 ne
rect 4244 0 4400 156
tri 4400 0 4556 156 sw
tri 4638 0 4794 156 ne
rect 4794 0 4950 156
tri 4950 0 5106 156 sw
tri 5188 0 5344 156 ne
rect 5344 0 5500 156
tri 5500 0 5656 156 sw
tri 5738 0 5894 156 ne
rect 5894 0 6050 156
tri 6050 0 6206 156 sw
tri 6288 0 6444 156 ne
rect 6444 0 6600 156
tri 6600 0 6756 156 sw
tri 6838 0 6994 156 ne
rect 6994 0 7150 156
tri 7150 0 7306 156 sw
tri 7388 0 7544 156 ne
rect 7544 0 7700 156
tri 7700 0 7856 156 sw
tri 7938 0 8094 156 ne
rect 8094 0 8250 156
tri 8250 0 8406 156 sw
tri 8488 0 8644 156 ne
rect 8644 0 8800 156
tri 8800 0 8956 156 sw
tri 9038 0 9194 156 ne
rect 9194 0 9350 156
tri 9350 0 9506 156 sw
tri 9588 0 9744 156 ne
rect 9744 0 9900 156
tri 9900 0 10056 156 sw
tri 10138 0 10294 156 ne
rect 10294 0 10450 156
tri 10450 0 10606 156 sw
tri 10688 0 10844 156 ne
rect 10844 0 11000 156
tri 11000 0 11156 156 sw
tri 11238 0 11394 156 ne
rect 11394 0 11550 156
tri 11550 0 11706 156 sw
tri 11788 0 11944 156 ne
rect 11944 0 12100 156
tri 12100 0 12256 156 sw
tri 12338 0 12494 156 ne
rect 12494 0 12650 156
tri 12650 0 12806 156 sw
tri 12888 0 13044 156 ne
rect 13044 0 13200 156
tri 13200 0 13356 156 sw
tri 13438 0 13594 156 ne
rect 13594 0 15775 156
rect -1025 -103 -394 0
tri -394 -103 -291 0 sw
tri -156 -103 -53 0 ne
rect -53 -103 156 0
rect -1025 -240 -291 -103
tri -291 -240 -154 -103 sw
tri -53 -240 84 -103 ne
rect 84 -238 156 -103
tri 156 -238 394 0 sw
tri 394 -238 632 0 ne
rect 632 -238 706 0
tri 706 -238 944 0 sw
tri 944 -238 1182 0 ne
rect 1182 -238 1256 0
tri 1256 -238 1494 0 sw
tri 1494 -238 1732 0 ne
rect 1732 -238 1806 0
tri 1806 -238 2044 0 sw
tri 2044 -238 2282 0 ne
rect 2282 -238 2356 0
tri 2356 -238 2594 0 sw
tri 2594 -238 2832 0 ne
rect 2832 -238 2906 0
tri 2906 -238 3144 0 sw
tri 3144 -238 3382 0 ne
rect 3382 -238 3456 0
tri 3456 -238 3694 0 sw
tri 3694 -238 3932 0 ne
rect 3932 -238 4006 0
tri 4006 -238 4244 0 sw
tri 4244 -238 4482 0 ne
rect 4482 -238 4556 0
tri 4556 -238 4794 0 sw
tri 4794 -238 5032 0 ne
rect 5032 -238 5106 0
tri 5106 -238 5344 0 sw
tri 5344 -238 5582 0 ne
rect 5582 -238 5656 0
tri 5656 -238 5894 0 sw
tri 5894 -238 6132 0 ne
rect 6132 -238 6206 0
tri 6206 -238 6444 0 sw
tri 6444 -238 6682 0 ne
rect 6682 -238 6756 0
tri 6756 -238 6994 0 sw
tri 6994 -238 7232 0 ne
rect 7232 -238 7306 0
tri 7306 -238 7544 0 sw
tri 7544 -238 7782 0 ne
rect 7782 -238 7856 0
tri 7856 -238 8094 0 sw
tri 8094 -238 8332 0 ne
rect 8332 -238 8406 0
tri 8406 -238 8644 0 sw
tri 8644 -238 8882 0 ne
rect 8882 -238 8956 0
tri 8956 -238 9194 0 sw
tri 9194 -238 9432 0 ne
rect 9432 -238 9506 0
tri 9506 -238 9744 0 sw
tri 9744 -238 9982 0 ne
rect 9982 -238 10056 0
tri 10056 -238 10294 0 sw
tri 10294 -238 10532 0 ne
rect 10532 -238 10606 0
tri 10606 -238 10844 0 sw
tri 10844 -238 11082 0 ne
rect 11082 -238 11156 0
tri 11156 -238 11394 0 sw
tri 11394 -238 11632 0 ne
rect 11632 -238 11706 0
tri 11706 -238 11944 0 sw
tri 11944 -238 12182 0 ne
rect 12182 -238 12256 0
tri 12256 -238 12494 0 sw
tri 12494 -238 12732 0 ne
rect 12732 -238 12806 0
tri 12806 -238 13044 0 sw
tri 13044 -156 13200 0 ne
rect 13200 -103 13356 0
tri 13356 -103 13459 0 sw
tri 13594 -103 13697 0 ne
rect 13697 -103 15775 0
rect 13200 -156 13459 -103
rect 84 -240 394 -238
rect -1025 -258 -310 -240
tri -448 -360 -346 -258 ne
rect -346 -360 -310 -258
rect -190 -360 -154 -240
tri -346 -498 -208 -360 ne
rect -208 -394 -154 -360
tri -154 -394 0 -240 sw
tri 84 -394 238 -240 ne
rect 238 -360 240 -240
rect 360 -360 394 -240
rect 238 -394 394 -360
tri 394 -394 550 -238 sw
tri 632 -259 653 -238 ne
rect 653 -240 944 -238
rect 653 -259 790 -240
rect -208 -497 0 -394
tri 0 -497 103 -394 sw
rect -208 -1575 103 -497
tri 238 -498 342 -394 ne
rect 342 -497 550 -394
tri 550 -497 653 -394 sw
tri 653 -396 790 -259 ne
rect 910 -360 944 -240
rect 790 -394 944 -360
tri 944 -394 1100 -238 sw
tri 1182 -394 1338 -238 ne
rect 1338 -240 1494 -238
rect 1338 -360 1340 -240
rect 1460 -360 1494 -240
rect 1338 -394 1494 -360
tri 1494 -394 1650 -238 sw
tri 1732 -259 1753 -238 ne
rect 1753 -240 2044 -238
rect 1753 -259 1890 -240
rect 790 -396 1100 -394
rect 342 -1075 653 -497
tri 790 -498 892 -396 ne
rect 892 -497 1100 -396
tri 1100 -497 1203 -394 sw
rect 892 -1575 1203 -497
tri 1338 -498 1442 -394 ne
rect 1442 -497 1650 -394
tri 1650 -497 1753 -394 sw
tri 1753 -396 1890 -259 ne
rect 2010 -360 2044 -240
rect 1890 -394 2044 -360
tri 2044 -394 2200 -238 sw
tri 2282 -259 2303 -238 ne
rect 2303 -240 2594 -238
rect 2303 -259 2440 -240
rect 1890 -396 2200 -394
rect 1442 -1075 1753 -497
tri 1890 -498 1992 -396 ne
rect 1992 -497 2200 -396
tri 2200 -497 2303 -394 sw
tri 2303 -396 2440 -259 ne
rect 2560 -360 2594 -240
rect 2440 -394 2594 -360
tri 2594 -394 2750 -238 sw
tri 2832 -394 2988 -238 ne
rect 2988 -240 3144 -238
rect 2988 -360 2990 -240
rect 3110 -360 3144 -240
rect 2988 -394 3144 -360
tri 3144 -394 3300 -238 sw
tri 3382 -259 3403 -238 ne
rect 3403 -240 3694 -238
rect 3403 -259 3540 -240
rect 2440 -396 2750 -394
rect 1992 -1575 2303 -497
tri 2440 -498 2542 -396 ne
rect 2542 -497 2750 -396
tri 2750 -497 2853 -394 sw
rect 2542 -1075 2853 -497
tri 2988 -498 3092 -394 ne
rect 3092 -497 3300 -394
tri 3300 -497 3403 -394 sw
tri 3403 -396 3540 -259 ne
rect 3660 -360 3694 -240
rect 3540 -394 3694 -360
tri 3694 -394 3850 -238 sw
tri 3932 -259 3953 -238 ne
rect 3953 -240 4244 -238
rect 3953 -259 4090 -240
rect 3540 -396 3850 -394
rect 3092 -1575 3403 -497
tri 3540 -498 3642 -396 ne
rect 3642 -497 3850 -396
tri 3850 -497 3953 -394 sw
tri 3953 -396 4090 -259 ne
rect 4210 -360 4244 -240
rect 4090 -394 4244 -360
tri 4244 -394 4400 -238 sw
tri 4482 -394 4638 -238 ne
rect 4638 -240 4794 -238
rect 4638 -360 4640 -240
rect 4760 -360 4794 -240
rect 4638 -394 4794 -360
tri 4794 -394 4950 -238 sw
tri 5032 -259 5053 -238 ne
rect 5053 -240 5344 -238
rect 5053 -259 5190 -240
rect 4090 -396 4400 -394
rect 3642 -1075 3953 -497
tri 4090 -498 4192 -396 ne
rect 4192 -497 4400 -396
tri 4400 -497 4503 -394 sw
rect 4192 -1575 4503 -497
tri 4638 -498 4742 -394 ne
rect 4742 -497 4950 -394
tri 4950 -497 5053 -394 sw
tri 5053 -396 5190 -259 ne
rect 5310 -360 5344 -240
rect 5190 -394 5344 -360
tri 5344 -394 5500 -238 sw
tri 5582 -259 5603 -238 ne
rect 5603 -240 5894 -238
rect 5603 -259 5740 -240
rect 5190 -396 5500 -394
rect 4742 -1075 5053 -497
tri 5190 -498 5292 -396 ne
rect 5292 -497 5500 -396
tri 5500 -497 5603 -394 sw
tri 5603 -396 5740 -259 ne
rect 5860 -360 5894 -240
rect 5740 -394 5894 -360
tri 5894 -394 6050 -238 sw
tri 6132 -394 6288 -238 ne
rect 6288 -240 6444 -238
rect 6288 -360 6290 -240
rect 6410 -360 6444 -240
rect 6288 -394 6444 -360
tri 6444 -394 6600 -238 sw
tri 6682 -259 6703 -238 ne
rect 6703 -240 6994 -238
rect 6703 -259 6840 -240
rect 5740 -396 6050 -394
rect 5292 -1575 5603 -497
tri 5740 -498 5842 -396 ne
rect 5842 -497 6050 -396
tri 6050 -497 6153 -394 sw
rect 5842 -1075 6153 -497
tri 6288 -498 6392 -394 ne
rect 6392 -497 6600 -394
tri 6600 -497 6703 -394 sw
tri 6703 -396 6840 -259 ne
rect 6960 -360 6994 -240
rect 6840 -394 6994 -360
tri 6994 -394 7150 -238 sw
tri 7232 -259 7253 -238 ne
rect 7253 -240 7544 -238
rect 7253 -259 7390 -240
rect 6840 -396 7150 -394
rect 6392 -1575 6703 -497
tri 6840 -498 6942 -396 ne
rect 6942 -497 7150 -396
tri 7150 -497 7253 -394 sw
tri 7253 -396 7390 -259 ne
rect 7510 -360 7544 -240
rect 7390 -394 7544 -360
tri 7544 -394 7700 -238 sw
tri 7782 -394 7938 -238 ne
rect 7938 -240 8094 -238
rect 7938 -360 7940 -240
rect 8060 -360 8094 -240
rect 7938 -394 8094 -360
tri 8094 -394 8250 -238 sw
tri 8332 -259 8353 -238 ne
rect 8353 -240 8644 -238
rect 8353 -259 8490 -240
rect 7390 -396 7700 -394
rect 6942 -1075 7253 -497
tri 7390 -498 7492 -396 ne
rect 7492 -497 7700 -396
tri 7700 -497 7803 -394 sw
rect 7492 -1575 7803 -497
tri 7938 -498 8042 -394 ne
rect 8042 -497 8250 -394
tri 8250 -497 8353 -394 sw
tri 8353 -396 8490 -259 ne
rect 8610 -360 8644 -240
rect 8490 -394 8644 -360
tri 8644 -394 8800 -238 sw
tri 8882 -259 8903 -238 ne
rect 8903 -240 9194 -238
rect 8903 -259 9040 -240
rect 8490 -396 8800 -394
rect 8042 -1075 8353 -497
tri 8490 -498 8592 -396 ne
rect 8592 -497 8800 -396
tri 8800 -497 8903 -394 sw
tri 8903 -396 9040 -259 ne
rect 9160 -360 9194 -240
rect 9040 -394 9194 -360
tri 9194 -394 9350 -238 sw
tri 9432 -394 9588 -238 ne
rect 9588 -240 9744 -238
rect 9588 -360 9590 -240
rect 9710 -360 9744 -240
rect 9588 -394 9744 -360
tri 9744 -394 9900 -238 sw
tri 9982 -259 10003 -238 ne
rect 10003 -240 10294 -238
rect 10003 -259 10140 -240
rect 9040 -396 9350 -394
rect 8592 -1575 8903 -497
tri 9040 -498 9142 -396 ne
rect 9142 -497 9350 -396
tri 9350 -497 9453 -394 sw
rect 9142 -1075 9453 -497
tri 9588 -498 9692 -394 ne
rect 9692 -497 9900 -394
tri 9900 -497 10003 -394 sw
tri 10003 -396 10140 -259 ne
rect 10260 -360 10294 -240
rect 10140 -394 10294 -360
tri 10294 -394 10450 -238 sw
tri 10532 -259 10553 -238 ne
rect 10553 -240 10844 -238
rect 10553 -259 10690 -240
rect 10140 -396 10450 -394
rect 9692 -1575 10003 -497
tri 10140 -498 10242 -396 ne
rect 10242 -497 10450 -396
tri 10450 -497 10553 -394 sw
tri 10553 -396 10690 -259 ne
rect 10810 -360 10844 -240
rect 10690 -394 10844 -360
tri 10844 -394 11000 -238 sw
tri 11082 -394 11238 -238 ne
rect 11238 -240 11394 -238
rect 11238 -360 11240 -240
rect 11360 -360 11394 -240
rect 11238 -394 11394 -360
tri 11394 -394 11550 -238 sw
tri 11632 -259 11653 -238 ne
rect 11653 -240 11944 -238
rect 11653 -259 11790 -240
rect 10690 -396 11000 -394
rect 10242 -1075 10553 -497
tri 10690 -498 10792 -396 ne
rect 10792 -497 11000 -396
tri 11000 -497 11103 -394 sw
rect 10792 -1575 11103 -497
tri 11238 -498 11342 -394 ne
rect 11342 -497 11550 -394
tri 11550 -497 11653 -394 sw
tri 11653 -396 11790 -259 ne
rect 11910 -360 11944 -240
rect 11790 -394 11944 -360
tri 11944 -394 12100 -238 sw
tri 12182 -259 12203 -238 ne
rect 12203 -240 12494 -238
rect 12203 -259 12340 -240
rect 11790 -396 12100 -394
rect 11342 -1075 11653 -497
tri 11790 -498 11892 -396 ne
rect 11892 -497 12100 -396
tri 12100 -497 12203 -394 sw
tri 12203 -396 12340 -259 ne
rect 12460 -360 12494 -240
rect 12340 -394 12494 -360
tri 12494 -394 12650 -238 sw
tri 12732 -394 12888 -238 ne
rect 12888 -240 13044 -238
rect 12888 -360 12890 -240
rect 13010 -360 13044 -240
rect 12888 -394 13044 -360
tri 13044 -394 13200 -238 sw
tri 13200 -394 13438 -156 ne
rect 13438 -240 13459 -156
tri 13459 -240 13596 -103 sw
rect 13438 -360 13440 -240
rect 13560 -342 13596 -240
tri 13596 -342 13698 -240 sw
rect 13560 -360 14275 -342
rect 13438 -394 14275 -360
rect 12340 -396 12650 -394
rect 11892 -1575 12203 -497
tri 12340 -498 12442 -396 ne
rect 12442 -497 12650 -396
tri 12650 -497 12753 -394 sw
rect 12442 -1075 12753 -497
tri 12888 -498 12992 -394 ne
rect 12992 -497 13200 -394
tri 13200 -497 13303 -394 sw
rect 12992 -1575 13303 -497
tri 13438 -498 13542 -394 ne
rect 13542 -653 14275 -394
rect 13542 -1075 13853 -653
rect 14775 -1575 15775 -103
rect -525 -2575 15775 -1575
<< labels >>
rlabel via1 -525 -575 -525 -575 1 G
rlabel metal5 15300 -575 15300 -575 1 S
rlabel metal5 -1750 14850 -1750 14850 1 D
rlabel viali -2350 -2250 -2350 -2250 1 PW
<< end >>

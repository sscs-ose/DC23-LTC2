* NGSPICE file created from TOP_CHILE_OPEN_LDO_pex.ext - technology: gf180mcuD

.subckt TOP_CHILE_OPEN_LDO_pex iref vin_p vss feedback ref out vdd
X0 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X3 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X4 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X5 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X6 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X7 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X8 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X9 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X10 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X11 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X12 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X13 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X14 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X15 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X16 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X17 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X18 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X19 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X20 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X21 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X22 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X23 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X24 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X25 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X26 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X27 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X28 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X29 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X30 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X31 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X32 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X33 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X34 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X35 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X36 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X37 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X38 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X39 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X40 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X41 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X42 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X43 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X44 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X45 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X46 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X47 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X48 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X49 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X50 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X51 a_313621_76595# a_315421_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X52 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X53 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X54 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X55 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X56 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X57 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X58 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X59 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X60 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X61 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X62 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X63 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=3.2335p ps=9.38u w=4.38u l=0.5u
X64 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X65 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X66 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X67 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X68 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X69 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=33.475p ps=0.14433m w=2.5u l=1u
X70 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X71 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X72 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X73 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X74 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X75 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X76 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X77 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X78 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X79 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X80 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X81 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X82 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X83 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X84 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X85 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X86 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X87 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X88 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X89 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X90 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X91 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X92 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X93 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X94 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X95 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X96 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X97 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X98 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X99 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X100 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X101 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X102 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X103 a_325921_73601# vss vss vss nfet_03v3 ad=1.3p pd=5.52u as=3.075p ps=11.23u w=5u l=1u
X104 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X105 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X106 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X107 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X108 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X109 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X110 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X111 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X112 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X113 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X114 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X115 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X116 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X117 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X118 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X119 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X120 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X121 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X122 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X123 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X124 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X125 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X126 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X127 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X128 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X129 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X130 vss iref open_ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X131 vdd vdd vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.366214n ps=0.01721 w=25u l=1u
X132 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X133 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X134 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X135 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X136 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X137 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X138 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X139 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X140 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X141 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X142 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X143 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X144 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X145 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X146 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X147 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X148 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X149 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X150 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X151 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X152 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X153 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X154 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X155 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X156 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X157 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X158 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X159 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X160 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X161 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X162 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X163 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X164 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X165 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X166 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X167 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X168 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X169 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X170 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X171 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X172 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X173 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X174 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X175 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X176 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X177 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X178 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X179 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X180 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X181 a_311821_76595# a_312421_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X182 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X183 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X184 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X185 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X186 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X187 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X188 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X189 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X190 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X191 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X192 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X193 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=3.2335p pd=9.38u as=3.8988p ps=13.77u w=4.38u l=0.5u
X194 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X195 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X196 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X197 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X198 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X199 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X200 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X201 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X202 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X203 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X204 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X205 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X206 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X207 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X208 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X209 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X210 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=2.6079p ps=9.38u w=4.38u l=0.5u
X211 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X212 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X213 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X214 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X215 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X216 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X217 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X218 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X219 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X220 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X221 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X222 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X223 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X224 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X225 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=2.6079p pd=9.38u as=4.814p ps=13.61u w=4.38u l=0.5u
X226 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X227 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X228 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X229 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X230 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X231 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X232 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X233 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=2.6079p ps=9.38u w=4.38u l=0.5u
X234 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X235 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X236 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X237 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X238 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X239 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X240 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X241 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X242 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X243 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X244 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X245 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X246 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X247 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X248 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X249 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X250 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X251 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X252 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X253 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X254 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X255 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X256 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X257 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X258 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X259 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X260 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X261 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X262 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X263 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X264 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X265 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X266 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X267 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X268 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X269 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X270 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X271 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X272 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X273 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X274 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X275 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X276 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X277 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X278 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X279 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X280 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X281 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X282 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X283 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X284 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X285 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X286 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X287 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X288 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X289 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X290 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X291 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=3.2335p pd=9.38u as=3.8988p ps=13.77u w=4.38u l=0.5u
X292 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X293 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X294 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X295 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X296 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X297 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X298 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X299 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X300 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X301 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X302 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X303 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X304 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X305 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X306 a_316021_76595# a_317221_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X307 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X308 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X309 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X310 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X311 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X312 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X313 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X314 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X315 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X316 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X317 vss iref iref vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X318 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X319 a_327783_76034# a_327175_76034# vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X320 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X321 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X322 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X323 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X324 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X325 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X326 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X327 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X328 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X329 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X330 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X331 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X332 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X333 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X334 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X335 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X336 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X337 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X338 vss vss vss ppolyf_u_1k r_width=1u r_length=5u
X339 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X340 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X341 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X342 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X343 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X344 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X345 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X346 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X347 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X348 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X349 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X350 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X351 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X352 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X353 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X354 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X355 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X356 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X357 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X358 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X359 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X360 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X361 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X362 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X363 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X364 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X365 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X366 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X367 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X368 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X369 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X370 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X371 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X372 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X373 vdd a_327783_76034# open_ldo_0.ota_0.vout vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X374 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X375 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X376 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X377 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X378 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X379 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X380 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X381 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X382 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X383 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X384 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X385 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X386 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X387 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X388 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X389 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X390 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X391 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X392 vss iref open_ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X393 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X394 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X395 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X396 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X397 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X398 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X399 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X400 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X401 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X402 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X403 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X404 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X405 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X406 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X407 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X408 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X409 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X410 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X411 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X412 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X413 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X414 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X415 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X416 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X417 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X418 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X419 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X420 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X421 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X422 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X423 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X424 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X425 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X426 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X427 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X428 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X429 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X430 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X431 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X432 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X433 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X434 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X435 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X436 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X437 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X438 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X439 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X440 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X441 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X442 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X443 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X444 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X445 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X446 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X447 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X448 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X449 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X450 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X451 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X452 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X453 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X454 vss iref a_325921_73601# vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X455 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X456 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X457 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X458 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X459 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X460 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X461 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X462 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X463 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X464 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X465 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X466 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X467 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X468 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X469 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X470 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X471 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X472 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X473 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X474 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X475 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X476 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X477 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X478 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X479 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X480 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X481 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X482 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X483 a_314221_76595# a_312421_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X484 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X485 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X486 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X487 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X488 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X489 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X490 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X491 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X492 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X493 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X494 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X495 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X496 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X497 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X498 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X499 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X500 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X501 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X502 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X503 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X504 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X505 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X506 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X507 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X508 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X509 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X510 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X511 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X512 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X513 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X514 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X515 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X516 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X517 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X518 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X519 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X520 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X521 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X522 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X523 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X524 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X525 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X526 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X527 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X528 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X529 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X530 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X531 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X532 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X533 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X534 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X535 vdd a_327783_76034# open_ldo_0.ota_0.vout vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X536 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X537 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X538 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X539 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X540 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X541 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X542 a_327783_76034# vin_p a_325921_73601# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X543 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X544 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X545 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X546 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X547 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X548 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X549 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X550 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X551 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X552 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X553 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X554 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X555 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X556 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X557 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X558 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X559 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X560 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X561 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X562 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X563 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X564 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X565 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X566 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X567 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X568 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X569 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X570 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X571 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X572 vss iref open_ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X573 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X574 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X575 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X576 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X577 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X578 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X579 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X580 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X581 a_311221_76595# a_310621_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X582 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X583 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X584 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X585 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X586 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X587 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X588 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X589 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X590 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X591 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X592 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X593 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X594 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X595 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X596 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X597 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X598 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X599 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X600 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X601 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X602 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X603 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X604 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X605 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X606 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X607 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X608 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X609 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X610 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X611 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X612 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X613 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X614 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X615 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X616 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X617 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X618 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X619 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X620 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X621 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X622 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X623 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X624 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X625 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X626 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X627 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X628 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X629 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X630 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X631 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X632 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X633 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X634 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X635 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X636 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X637 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X638 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X639 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X640 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X641 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X642 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X643 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X644 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X645 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X646 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X647 a_327175_76034# a_327175_76034# vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X648 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X649 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X650 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X651 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X652 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X653 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X654 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X655 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X656 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X657 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X658 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X659 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X660 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X661 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X662 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X663 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X664 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X665 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X666 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X667 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X668 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X669 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X670 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X671 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X672 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X673 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X674 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X675 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X676 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X677 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X678 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X679 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X680 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X681 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X682 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X683 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X684 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X685 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X686 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X687 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X688 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X689 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X690 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X691 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X692 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X693 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X694 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X695 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X696 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X697 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X698 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X699 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X700 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X701 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X702 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X703 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X704 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X705 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X706 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X707 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X708 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X709 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X710 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X711 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X712 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X713 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X714 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X715 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X716 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X717 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X718 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X719 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X720 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X721 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X722 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X723 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X724 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X725 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X726 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X727 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X728 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X729 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X730 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X731 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X732 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X733 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X734 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X735 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X736 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X737 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X738 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X739 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X740 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X741 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X742 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X743 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X744 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X745 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X746 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X747 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X748 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X749 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X750 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X751 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X752 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X753 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X754 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X755 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X756 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X757 a_316021_76595# a_315421_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X758 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X759 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X760 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X761 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X762 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X763 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X764 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X765 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X766 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X767 a_331573_72398# a_332701_72398# vss ppolyf_u_1k r_width=1u r_length=5u
X768 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X769 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X770 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X771 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X772 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X773 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X774 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X775 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X776 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X777 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X778 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X779 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X780 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X781 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X782 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X783 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X784 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X785 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X786 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X787 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X788 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X789 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X790 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X791 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X792 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X793 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X794 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X795 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X796 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X797 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X798 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X799 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X800 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X801 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X802 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X803 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X804 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X805 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X806 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X807 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X808 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X809 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X810 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X811 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X812 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X813 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X814 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X815 out a_308821_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X816 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X817 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X818 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X819 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X820 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X821 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X822 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X823 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X824 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X825 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X826 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X827 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X828 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X829 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X830 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X831 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X832 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X833 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X834 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X835 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X836 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X837 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X838 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X839 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X840 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X841 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X842 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X843 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X844 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X845 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X846 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X847 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X848 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X849 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X850 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X851 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X852 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X853 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X854 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X855 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X856 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X857 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X858 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X859 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X860 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X861 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X862 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X863 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X864 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X865 vss iref open_ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X866 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X867 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X868 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X869 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X870 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X871 a_311221_76595# a_313021_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X872 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=2.6079p pd=9.38u as=4.814p ps=13.61u w=4.38u l=0.5u
X873 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X874 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X875 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X876 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X877 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X878 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X879 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X880 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X881 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X882 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X883 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X884 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X885 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X886 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X887 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X888 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X889 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X890 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X891 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X892 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X893 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X894 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X895 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X896 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X897 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X898 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X899 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X900 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X901 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X902 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X903 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X904 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X905 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X906 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X907 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X908 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X909 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X910 open_ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X911 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X912 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X913 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X914 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X915 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X916 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X917 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X918 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X919 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X920 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X921 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X922 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X923 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X924 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X925 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X926 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X927 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X928 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X929 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X930 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X931 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X932 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X933 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X934 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X935 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X936 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X937 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X938 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X939 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X940 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X941 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X942 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X943 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X944 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X945 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X946 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X947 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X948 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X949 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X950 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X951 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X952 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X953 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X954 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X955 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X956 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X957 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X958 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X959 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X960 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X961 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X962 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X963 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X964 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X965 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X966 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X967 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X968 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X969 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X970 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X971 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X972 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X973 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X974 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X975 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X976 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X977 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X978 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X979 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X980 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X981 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X982 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X983 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X984 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X985 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X986 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X987 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X988 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X989 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X990 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X991 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X992 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X993 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X994 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X995 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X996 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X997 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X998 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X999 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1000 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1001 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1002 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1003 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1004 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1005 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1006 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1007 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1008 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1009 vss a_310021_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1010 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1011 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1012 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1013 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1014 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1015 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1016 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1017 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1018 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1019 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1020 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1021 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1022 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1023 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1024 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1025 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1026 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1027 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1028 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1029 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1030 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1031 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1032 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1033 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1034 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1035 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1036 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1037 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1038 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1039 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1040 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1041 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1042 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1043 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1044 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1045 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1046 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1047 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1048 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1049 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1050 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1051 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1052 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1053 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1054 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1055 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1056 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1057 a_331573_72398# a_327783_76034# vss ppolyf_u_1k r_width=1u r_length=5u
X1058 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1059 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1060 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1061 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1062 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1063 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1064 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1065 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1066 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1067 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1068 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1069 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1070 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1071 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1072 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1073 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1074 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1075 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1076 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1077 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1078 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1079 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1080 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1081 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1082 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1083 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1084 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1085 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1086 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1087 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1088 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1089 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1090 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1091 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1092 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1093 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1094 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1095 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1096 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1097 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1098 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1099 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1100 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1101 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1102 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1103 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1104 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1105 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1106 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1107 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1108 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1109 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1110 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1111 open_ldo_0.ota_0.vout a_327783_76034# vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X1112 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1113 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1114 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1115 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1116 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1117 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1118 vdd vdd vdd vdd pfet_03v3 ad=3.25p pd=11.299999u as=0 ps=0 w=5u l=1u
X1119 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1120 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1121 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1122 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1123 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1124 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1125 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1126 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1127 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1128 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1129 open_ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1130 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1131 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1132 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1133 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1134 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1135 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1136 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1137 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1138 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1139 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1140 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1141 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1142 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1143 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1144 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1145 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1146 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1147 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1148 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1149 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1150 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1151 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1152 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1153 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1154 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1155 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1156 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1157 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1158 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1159 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1160 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1161 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1162 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1163 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1164 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1165 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1166 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1167 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1168 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1169 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1170 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1171 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1172 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1173 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1174 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1175 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1176 open_ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1177 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1178 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1179 a_327175_76034# ref a_325921_73601# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1180 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1181 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1182 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1183 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1184 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1185 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1186 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1187 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1188 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1189 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1190 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1191 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1192 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1193 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1194 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1195 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1196 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1197 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1198 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1199 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1200 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1201 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1202 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1203 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1204 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1205 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1206 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1207 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1208 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1209 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1210 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1211 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1212 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1213 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1214 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1215 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1216 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1217 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1218 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1219 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1220 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1221 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1222 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1223 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1224 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1225 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1226 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1227 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1228 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1229 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1230 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1231 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1232 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1233 feedback a_317221_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1234 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1235 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1236 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1237 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1238 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1239 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1240 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1241 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1242 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1243 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1244 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1245 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=0 ps=0 w=2.5u l=1u
X1246 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1247 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1248 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1249 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1250 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1251 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1252 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1253 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1254 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1255 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1256 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1257 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1258 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1259 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1260 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1261 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1262 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1263 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1264 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1265 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1266 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1267 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1268 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1269 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1270 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1271 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1272 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1273 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1274 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1275 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1276 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1277 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1278 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1279 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1280 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1281 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1282 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1283 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1284 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1285 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1286 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1287 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1288 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1289 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1290 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1291 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1292 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1293 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1294 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1295 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1296 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1297 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1298 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1299 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1300 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1301 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1302 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1303 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1304 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1305 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1306 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1307 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1308 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1309 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1310 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1311 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1312 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1313 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1314 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1315 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1316 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1317 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1318 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1319 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1320 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1321 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1322 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1323 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1324 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1325 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1326 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1327 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1328 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1329 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1330 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1331 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1332 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1333 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1334 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1335 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1336 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1337 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1338 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1339 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1340 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1341 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1342 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1343 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1344 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1345 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1346 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1347 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1348 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1349 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1350 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1351 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1352 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1353 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1354 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1355 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1356 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1357 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1358 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1359 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1360 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1361 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1362 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1363 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1364 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1365 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1366 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1367 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1368 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1369 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1370 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1371 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1372 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1373 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1374 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1375 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1376 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1377 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1378 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1379 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1380 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1381 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1382 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1383 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1384 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1385 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1386 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1387 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1388 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1389 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1390 vdd vdd vdd vdd pfet_03v3 ad=1.3p pd=5.52u as=0 ps=0 w=5u l=1u
X1391 a_314221_76595# a_314821_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1392 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1393 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1394 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1395 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1396 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1397 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1398 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1399 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1400 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1401 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1402 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1403 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1404 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1405 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1406 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1407 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1408 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1409 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1410 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1411 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1412 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1413 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1414 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1415 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1416 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1417 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1418 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1419 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1420 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1421 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1422 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1423 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1424 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1425 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1426 open_ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1427 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1428 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1429 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1430 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1431 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1432 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1433 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1434 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1435 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1436 open_ldo_0.ota_0.vout a_327783_76034# vdd vdd pfet_03v3 ad=6.5p pd=25.519999u as=6.5p ps=25.519999u w=25u l=1u
X1437 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1438 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1439 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1440 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1441 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1442 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1443 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1444 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1445 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1446 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1447 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1448 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1449 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1450 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1451 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1452 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1453 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1454 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1455 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1456 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1457 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1458 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1459 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1460 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1461 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1462 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1463 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1464 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1465 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1466 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1467 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1468 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1469 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1470 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1471 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1472 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1473 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1474 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1475 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1476 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1477 vss vss vss ppolyf_u_1k r_width=1u r_length=5u
X1478 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1479 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1480 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1481 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1482 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1483 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1484 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1485 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1486 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1487 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1488 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1489 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1490 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1491 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1492 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1493 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1494 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1495 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1496 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1497 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1498 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1499 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1500 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1501 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1502 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1503 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1504 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1505 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1506 a_309421_76595# a_308821_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1507 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1508 iref iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1509 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1510 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1511 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1512 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1513 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1514 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1515 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1516 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1517 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1518 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1519 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1520 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1521 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1522 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1523 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1524 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1525 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1526 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1527 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1528 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1529 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1530 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1531 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1532 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1533 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1534 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1535 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1536 a_311821_76595# a_310021_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1537 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1538 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1539 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1540 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1541 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1542 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1543 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1544 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1545 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1546 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1547 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1548 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1549 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1550 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1551 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1552 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1553 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1554 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1555 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1556 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1557 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1558 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1559 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1560 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1561 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1562 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1563 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1564 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1565 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1566 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1567 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1568 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1569 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1570 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1571 a_325921_73601# iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1572 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1573 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1574 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1575 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1576 open_ldo_0.ota_0.vout a_332701_72398# cap_mim_2f0_m4m5_noshield c_width=22u c_length=22u
X1577 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1578 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1579 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1580 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1581 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1582 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1583 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1584 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1585 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1586 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1587 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1588 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1589 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1590 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1591 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1592 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1593 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1594 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1595 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1596 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1597 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1598 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1599 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1600 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1601 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1602 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1603 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1604 a_325921_73601# vin_p a_327783_76034# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1605 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1606 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1607 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1608 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1609 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1610 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1611 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1612 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1613 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1614 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1615 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1616 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1617 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1618 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1619 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1620 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1621 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1622 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1623 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1624 open_ldo_0.ota_0.vout iref vss vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1625 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=0 ps=0 w=2.5u l=1u
X1626 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1627 vdd a_327175_76034# a_327175_76034# vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1628 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1629 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1630 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1631 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1632 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1633 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1634 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1635 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1636 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1637 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1638 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1639 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1640 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1641 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1642 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1643 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1644 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1645 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1646 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1647 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1648 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1649 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1650 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1651 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1652 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1653 feedback a_314821_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1654 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1655 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1656 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1657 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1658 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1659 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1660 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1661 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1662 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1663 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1664 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1665 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1666 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1667 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1668 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1669 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1670 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1671 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1672 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1673 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1674 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1675 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1676 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1677 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1678 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1679 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1680 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1681 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1682 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1683 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1684 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1685 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1686 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1687 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1688 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1689 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1690 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1691 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1692 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1693 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1694 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1695 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1696 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1697 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1698 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1699 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1700 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1701 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1702 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1703 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1704 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1705 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1706 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1707 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1708 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1709 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1710 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1711 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1712 vss vss vss vss nfet_03v3 ad=0.65p pd=3.02u as=0 ps=0 w=2.5u l=1u
X1713 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1714 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1715 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1716 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1717 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1718 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1719 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1720 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1721 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1722 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1723 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1724 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1725 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1726 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1727 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1728 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1729 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1730 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1731 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1732 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1733 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1734 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1735 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1736 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1737 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1738 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1739 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1740 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1741 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1742 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1743 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1744 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1745 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1746 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1747 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1748 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1749 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1750 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1751 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1752 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1753 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1754 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1755 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1756 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1757 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1758 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1759 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1760 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1761 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1762 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1763 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1764 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1765 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1766 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1767 vss vss vss vss nfet_03v3 ad=1.525p pd=6.22u as=0 ps=0 w=2.5u l=1u
X1768 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1769 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1770 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1771 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1772 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1773 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1774 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1775 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1776 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1777 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1778 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1779 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1780 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1781 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1782 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1783 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1784 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1785 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1786 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1787 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1788 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1789 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1790 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1791 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1792 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1793 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1794 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1795 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1796 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1797 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1798 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1799 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1800 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1801 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1802 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1803 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1804 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1805 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1806 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1807 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1808 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1809 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1810 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1811 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1812 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1813 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1814 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1815 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1816 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1817 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1818 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1819 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1820 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1821 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1822 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1823 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1824 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1825 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1826 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1827 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1828 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1829 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1830 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1831 a_313621_76595# a_313021_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1832 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1833 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1834 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1835 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1836 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1837 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1838 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1839 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1840 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1841 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1842 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1843 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1844 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1845 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1846 vdd a_327175_76034# a_327783_76034# vdd pfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X1847 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1848 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1849 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1850 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1851 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1852 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1853 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1854 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1855 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1856 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1857 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1858 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1859 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1860 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1861 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1862 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1863 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1864 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1865 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1866 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1867 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1868 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1869 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1870 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1871 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1872 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1873 vdd vdd vdd vdd pfet_03v3 ad=16.25p pd=51.3u as=0 ps=0 w=25u l=1u
X1874 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1875 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1876 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1877 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1878 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1879 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1880 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1881 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1882 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1883 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1884 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1885 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1886 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1887 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1888 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1889 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1890 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1891 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1892 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1893 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1894 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1895 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1896 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1897 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1898 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1899 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1900 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1901 vss vss vss ppolyf_u_1k r_width=1u r_length=20u
X1902 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1903 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1904 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1905 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1906 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1907 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1908 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1909 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1910 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1911 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1912 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1913 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1914 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1915 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1916 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1917 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1918 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1919 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1920 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1921 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1922 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1923 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1924 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1925 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1926 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1927 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1928 a_309421_76595# a_310621_72467# vss ppolyf_u_1k r_width=1u r_length=20u
X1929 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1930 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1931 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1932 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1933 vss vss vss ppolyf_u_1k r_width=1u r_length=20u
X1934 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1935 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1936 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1937 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1938 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1939 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1940 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1941 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1942 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1943 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1944 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1945 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1946 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1947 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1948 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1949 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1950 vss vss a_325921_73601# vss nfet_03v3 ad=3.05p pd=11.219999u as=1.3p ps=5.52u w=5u l=1u
X1951 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1952 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1953 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1954 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1955 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1956 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1957 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1958 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1959 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1960 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1961 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=3.2335p ps=9.38u w=4.38u l=0.5u
X1962 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1963 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1964 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1965 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1966 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X1967 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1968 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1969 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1970 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1971 vss iref open_ldo_0.ota_0.vout vss nfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=1u
X1972 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1973 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1974 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1975 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1976 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1977 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1978 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1979 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1980 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1981 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1982 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1983 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X1984 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1985 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1986 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1987 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1988 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X1989 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1990 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1991 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1992 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1993 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1994 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X1995 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X1996 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1997 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1998 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X1999 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2000 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2001 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2002 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2003 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2004 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=4.814p ps=13.61u w=4.38u l=0.5u
X2005 a_325921_73601# ref a_327175_76034# vss nfet_03v3 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=1u
X2006 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2007 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2008 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2009 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2010 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2011 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2012 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2013 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2014 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2015 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2016 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2017 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=3.8988p pd=13.77u as=6.322p ps=16.92u w=4.38u l=0.5u
X2018 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2019 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2020 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2021 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2022 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2023 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2024 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2025 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X2026 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2027 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2028 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2029 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=4.814p pd=13.61u as=3.8988p ps=13.77u w=4.38u l=0.5u
X2030 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2031 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2032 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2033 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2034 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2035 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2036 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=4.814p ps=13.61u w=4.38u l=0.5u
X2037 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2038 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2039 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2040 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2041 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2042 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2043 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2044 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2045 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2046 out open_ldo_0.ota_0.vout vdd vdd pfet_03v3 ad=5.163599p pd=17.56u as=6.322p ps=16.92u w=4.38u l=0.5u
X2047 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
X2048 vdd open_ldo_0.ota_0.vout out vdd pfet_03v3 ad=6.322p pd=16.92u as=5.163599p ps=17.56u w=4.38u l=0.5u
C0 a_325921_73601# iref 0.215656f
C1 vdd feedback 11.426401f
C2 m1_317211_77525# feedback 0.137209f
C3 a_313621_76595# a_316021_76595# 0.14109f
C4 a_332701_72398# iref 0.573472f
C5 vdd ref 12.195901f
C6 open_ldo_0.ota_0.vout iref 3.66853f
C7 a_325921_73601# a_327783_76034# 0.434752f
C8 a_325921_73601# vin_p 0.967832f
C9 a_313021_72467# a_312421_72467# 0.864964f
C10 open_ldo_0.ota_0.vout out 1.31128p
C11 a_317221_72467# a_314821_72467# 0.120932f
C12 a_327783_76034# vin_p 1.10184f
C13 a_325921_73601# a_327175_76034# 0.216749f
C14 a_332701_72398# a_327783_76034# 0.332743f
C15 open_ldo_0.ota_0.vout a_327783_76034# 3.13106f
C16 a_332701_72398# open_ldo_0.ota_0.vout 2.737f
C17 a_311221_76595# a_311821_76595# 0.802011f
C18 a_327783_76034# a_327175_76034# 1.10962f
C19 a_309421_76595# a_311221_76595# 0.14109f
C20 a_327175_76034# vin_p 0.389594f
C21 vdd iref 3.26831f
C22 a_313621_76595# a_314221_76595# 0.802011f
C23 vdd out 2.35665p
C24 a_313621_76595# a_311221_76595# 0.14109f
C25 a_310021_72467# a_312421_72467# 0.14109f
C26 ref iref 2.99563f
C27 out feedback 0.411961f
C28 a_327783_76034# vdd 9.13877f
C29 a_308821_72467# vdd 0.121652f
C30 vdd vin_p 8.31014f
C31 a_325921_73601# ref 2.366f
C32 a_310021_72467# a_310621_72467# 0.864964f
C33 a_332701_72398# vdd 0.494722f
C34 open_ldo_0.ota_0.vout vdd 1.77216p
C35 feedback vin_p 0.211703f
C36 a_316021_76595# feedback 0.600659f
C37 ref vin_p 1.26274f
C38 a_327175_76034# vdd 3.02748f
C39 a_332701_72398# ref 0.423289f
C40 open_ldo_0.ota_0.vout ref 0.134195f
C41 a_309421_76595# out 0.120238f
C42 a_308821_72467# a_310021_72467# 0.120932f
C43 a_314821_72467# a_312421_72467# 0.14109f
C44 a_327175_76034# ref 1.05237f
C45 a_315421_72467# a_314821_72467# 0.864964f
C46 iref vss 29.6738f
C47 vin_p vss 13.0541f
C48 ref vss 12.4705f
C49 feedback vss 16.2747f
C50 out vss 0.153743p
C51 vdd vss 33.3066p
C52 m1_318411_71393# vss 0.237793f $ **FLOATING
C53 m1_316611_71393# vss 0.193159f $ **FLOATING
C54 m1_314811_71393# vss 0.192608f $ **FLOATING
C55 m1_314211_71393# vss 0.193159f $ **FLOATING
C56 m1_312411_71393# vss 0.192608f $ **FLOATING
C57 m1_311811_71393# vss 0.193159f $ **FLOATING
C58 m1_310011_71393# vss 0.192608f $ **FLOATING
C59 m1_308211_71393# vss 0.217848f $ **FLOATING
C60 m1_318411_71793# vss 0.269211f $ **FLOATING
C61 m1_308211_71793# vss 0.248714f $ **FLOATING
C62 m1_318411_77125# vss 0.290611f $ **FLOATING
C63 m1_308211_77125# vss 0.270516f $ **FLOATING
C64 m1_318411_77525# vss 0.222777f $ **FLOATING
C65 m1_317211_77525# vss 0.177465f $ **FLOATING
C66 m1_316011_77525# vss 0.205536f $ **FLOATING
C67 m1_315411_77525# vss 0.205536f $ **FLOATING
C68 m1_313611_77525# vss 0.205536f $ **FLOATING
C69 m1_313011_77525# vss 0.205536f $ **FLOATING
C70 m1_311211_77525# vss 0.205536f $ **FLOATING
C71 m1_310611_77525# vss 0.269682f $ **FLOATING
C72 m1_309411_77525# vss 0.267473f $ **FLOATING
C73 m1_308211_77525# vss 0.227432f $ **FLOATING
C74 a_332701_72398# vss 2.96596f
C75 a_331573_72398# vss 1.30142f
C76 a_327783_76034# vss 4.70165f
C77 a_327175_76034# vss 2.39286f
C78 a_325921_73601# vss 3.68453f
C79 a_317221_72467# vss 1.84846f
C80 a_316021_76595# vss 2.16602f
C81 a_315421_72467# vss 1.55755f
C82 a_314821_72467# vss 1.94527f
C83 a_314221_76595# vss 1.80662f
C84 a_313621_76595# vss 2.46883f
C85 a_313021_72467# vss 1.56132f
C86 a_312421_72467# vss 1.93093f
C87 a_311821_76595# vss 1.81178f
C88 a_311221_76595# vss 2.46883f
C89 a_310621_72467# vss 1.55755f
C90 a_310021_72467# vss 1.94527f
C91 a_309421_76595# vss 2.67953f
C92 a_308821_72467# vss 1.81856f
C93 open_ldo_0.ota_0.vout vss 0.130198p
.ends


* Extracted by KLayout with GF180MCU LVS runset on : 16/01/2024 03:17

.SUBCKT waffle-12x12
M$1 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$2 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$3 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$4 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$5 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$6 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$7 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$8 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$9 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$10 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$11 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$12 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$13 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$14 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$15 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$16 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$17 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$18 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$19 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$20 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$21 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$22 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$23 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$24 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$25 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$26 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$27 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$28 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$29 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$30 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$31 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$32 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$33 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$34 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$35 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$36 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$37 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$38 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$39 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$40 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$41 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$42 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$43 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$44 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$45 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$46 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$47 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$48 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$49 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$50 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$51 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$52 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$53 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$54 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$55 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$56 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$57 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$58 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$59 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$60 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$61 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$62 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$63 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$64 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$65 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$66 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$67 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$68 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$69 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$70 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$71 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$72 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$73 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$74 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$75 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$76 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$77 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$78 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=5.5934P PS=9.39333333333U
+ PD=16.02U
M$79 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$80 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$81 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$82 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$83 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$84 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=5.5934P PS=9.39333333333U
+ PD=16.02U
M$85 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$86 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$87 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$88 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$89 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$90 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$91 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$92 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$93 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$94 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$95 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$96 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$97 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$98 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$99 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$100 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$101 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$102 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$103 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$104 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$105 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$106 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$107 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$108 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$109 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$110 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$111 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$112 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$113 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$114 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$115 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$116 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$117 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$118 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$119 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$120 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$121 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$122 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.33125P AD=4.15233333333P PS=9.38U
+ PD=10.8733333333U
M$123 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$124 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$125 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$126 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$127 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$128 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$129 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$130 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$131 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$132 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$133 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$134 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.33125P AD=4.15233333333P PS=9.38U
+ PD=10.8733333333U
M$135 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$136 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$137 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$138 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$139 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$140 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$141 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$142 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$143 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$144 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$145 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$146 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$147 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$148 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$149 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$150 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$151 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$152 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$153 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$154 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$155 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$156 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$157 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$158 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$159 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$160 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$161 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$162 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$163 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$164 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$165 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$166 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$167 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$168 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$169 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$170 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$171 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$172 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$173 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$174 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$175 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$176 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$177 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$178 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$179 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$180 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$181 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$182 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$183 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$184 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$185 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$186 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=5.5934P PS=9.39333333333U
+ PD=16.02U
M$187 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=5.5934P PS=9.39333333333U
+ PD=16.02U
M$188 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$189 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$190 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$191 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$192 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$193 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$194 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$195 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$196 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$197 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$198 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$199 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$200 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$201 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$202 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$203 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$204 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$205 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$206 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$207 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$208 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$209 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$210 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$211 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$212 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$213 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.33125P AD=4.15233333333P PS=9.38U
+ PD=10.8733333333U
M$214 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$215 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$216 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$217 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$218 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$219 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$220 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$221 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$222 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$223 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$224 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$225 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$226 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$227 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$228 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$229 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$230 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$231 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$232 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$233 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$234 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$235 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$236 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$237 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$238 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$239 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$240 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$241 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$242 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$243 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$244 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$245 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$246 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$247 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$248 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$249 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$250 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=3.4318P PS=9.39333333333U
+ PD=8.3U
M$251 S G D D pfet_03v3 L=0.5U W=4.38U AS=4.15233333333P AD=1.3923P
+ PS=10.8733333333U PD=9.42U
M$252 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.33125P AD=4.15233333333P PS=9.38U
+ PD=10.8733333333U
M$253 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
M$254 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$255 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$256 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$257 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$258 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$259 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$260 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=4.15233333333P PS=9.42U
+ PD=10.8733333333U
M$261 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$262 S G D D pfet_03v3 L=0.5U W=4.38U AS=3.4318P AD=1.3923P PS=8.3U PD=9.42U
M$263 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3923P AD=3.4318P PS=9.42U PD=8.3U
M$264 D G S D pfet_03v3 L=0.5U W=4.38U AS=1.3516P AD=4.15233333333P
+ PS=9.39333333333U PD=10.8733333333U
.ENDS waffle-12x12

* Extracted by KLayout with GF180MCU LVS runset on : 24/12/2023 05:15

* cell resistor
* pin OUT,VDD,VSS
* pin gf180mcu_gnd
.SUBCKT resistor OUT|VDD|VSS gf180mcu_gnd
* device instance $1 r0 *1 10,0.5 ppolyf_u
R$1 OUT|VDD|VSS OUT|VDD|VSS gf180mcu_gnd 388.888888889 ppolyf_u L=20U W=18U
.ENDS resistor

* NGSPICE file created from gf180mcu_fd_io__asig_5p0_gab.ext - technology: gf180mcuC

.subckt gf180mcu_fd_io__asig_5p0_gab VSS VDD ASIG5V DVSS DVDD
X0 DVDD.t1 DVSS.t36 cap_nmos_06v0 c_width=15u c_length=15u
X1 DVDD.t2 DVSS.t35 cap_nmos_06v0 c_width=15u c_length=15u
X2 DVDD.t3 DVSS.t34 cap_nmos_06v0 c_width=15u c_length=15u
X3 DVDD.t4 DVSS.t33 cap_nmos_06v0 c_width=15u c_length=15u
X4 DVDD.t5 DVSS.t32 cap_nmos_06v0 c_width=15u c_length=15u
D0 DVSS.t3 DVDD.t6 diode_nd2ps_06v0 pj=82u area=40p
X5 DVDD.t7 DVSS.t31 cap_nmos_06v0 c_width=15u c_length=15u
X6 DVDD.t8 DVSS.t30 cap_nmos_06v0 c_width=15u c_length=15u
X7 DVDD.t9 DVSS.t29 cap_nmos_06v0 c_width=15u c_length=15u
X8 DVDD.t10 DVSS.t28 cap_nmos_06v0 c_width=15u c_length=15u
X9 DVDD.t11 DVSS.t27 cap_nmos_06v0 c_width=15u c_length=15u
X10 DVDD.t12 DVSS.t26 cap_nmos_06v0 c_width=15u c_length=15u
X11 DVDD.t13 DVSS.t25 cap_nmos_06v0 c_width=15u c_length=15u
X12 DVDD.t14 DVSS.t24 cap_nmos_06v0 c_width=15u c_length=15u
X13 DVDD.t15 DVSS.t23 cap_nmos_06v0 c_width=15u c_length=15u
X14 DVDD.t16 DVSS.t22 cap_nmos_06v0 c_width=15u c_length=15u
D1 DVSS.t37 ASIG5V.t0 diode_nd2ps_06v0 pj=0.106m area=0.15n
X15 DVDD.t17 DVSS.t21 cap_nmos_06v0 c_width=15u c_length=15u
X16 DVDD.t18 DVSS.t20 cap_nmos_06v0 c_width=15u c_length=15u
X17 DVDD.t19 DVSS.t19 cap_nmos_06v0 c_width=15u c_length=15u
D2 DVSS.t37 ASIG5V.t1 diode_nd2ps_06v0 pj=0.106m area=0.15n
D3 ASIG5V.t2 DVDD.t0 diode_pd2nw_06v0 pj=0.106m area=0.15n
X18 DVDD.t20 DVSS.t18 cap_nmos_06v0 c_width=15u c_length=15u
X19 DVDD.t21 DVSS.t17 cap_nmos_06v0 c_width=15u c_length=15u
D4 ASIG5V.t3 DVDD.t0 diode_pd2nw_06v0 pj=0.106m area=0.15n
D5 DVSS.t37 ASIG5V.t4 diode_nd2ps_06v0 pj=0.106m area=0.15n
X20 DVDD.t22 DVSS.t16 cap_nmos_06v0 c_width=15u c_length=15u
D6 ASIG5V.t5 DVDD.t0 diode_pd2nw_06v0 pj=0.106m area=0.15n
X21 DVDD.t23 DVSS.t15 cap_nmos_06v0 c_width=15u c_length=15u
X22 DVDD.t24 DVSS.t14 cap_nmos_06v0 c_width=15u c_length=15u
D7 DVSS.t3 DVDD.t25 diode_nd2ps_06v0 pj=82u area=40p
X23 DVDD.t26 DVSS.t13 cap_nmos_06v0 c_width=15u c_length=15u
X24 DVDD.t27 DVSS.t12 cap_nmos_06v0 c_width=15u c_length=15u
X25 DVDD.t28 DVSS.t11 cap_nmos_06v0 c_width=15u c_length=15u
X26 DVDD.t29 DVSS.t10 cap_nmos_06v0 c_width=15u c_length=15u
X27 DVDD.t30 DVSS.t9 cap_nmos_06v0 c_width=15u c_length=15u
D8 DVSS.t3 DVDD.t31 diode_nd2ps_06v0 pj=82u area=40p
X28 DVDD.t32 DVSS.t8 cap_nmos_06v0 c_width=15u c_length=15u
D9 DVSS.t37 ASIG5V.t6 diode_nd2ps_06v0 pj=0.106m area=0.15n
X29 DVDD.t33 DVSS.t7 cap_nmos_06v0 c_width=15u c_length=15u
X30 DVDD.t34 DVSS.t6 cap_nmos_06v0 c_width=15u c_length=15u
X31 DVDD.t35 DVSS.t5 cap_nmos_06v0 c_width=15u c_length=15u
X32 DVDD.t36 DVSS.t4 cap_nmos_06v0 c_width=15u c_length=15u
D10 DVSS.t3 DVDD.t37 diode_nd2ps_06v0 pj=82u area=40p
D11 ASIG5V.t7 DVDD.t0 diode_pd2nw_06v0 pj=0.106m area=0.15n
X33 DVDD.t38 DVSS.t2 cap_nmos_06v0 c_width=15u c_length=15u
X34 DVDD.t39 DVSS.t1 cap_nmos_06v0 c_width=15u c_length=15u
X35 DVDD.t40 DVSS.t0 cap_nmos_06v0 c_width=15u c_length=15u
R0 DVDD.n2024 DVDD.n2023 47.4925
R1 DVDD.n2055 DVDD.n2054 47.4925
R2 DVDD.n2156 DVDD.n2155 47.4925
R3 DVDD.n2209 DVDD.n2208 47.4925
R4 DVDD.n2232 DVDD.n2231 47.4925
R5 DVDD.n18931 DVDD.n18930 47.4925
R6 DVDD.n7100 DVDD.n7099 47.4925
R7 DVDD.n7033 DVDD.n7032 47.4925
R8 DVDD.n6938 DVDD.n6937 47.4925
R9 DVDD.n6943 DVDD.n6942 47.4925
R10 DVDD.n6786 DVDD.n6785 47.4925
R11 DVDD.n6802 DVDD.n6801 47.4925
R12 DVDD.n6520 DVDD.n6519 47.4925
R13 DVDD.n6553 DVDD.n6552 47.4925
R14 DVDD.n1859 DVDD.n1858 47.4925
R15 DVDD.n1862 DVDD.n1861 47.4925
R16 DVDD.n3925 DVDD.n3924 47.4925
R17 DVDD.n3930 DVDD.n3929 47.4925
R18 DVDD.n19833 DVDD.n19832 47.4925
R19 DVDD.n19802 DVDD.n19801 47.4925
R20 DVDD.n19988 DVDD.n19987 47.4925
R21 DVDD.n19935 DVDD.n19934 47.4925
R22 DVDD.n19049 DVDD.n19048 47.4925
R23 DVDD.n20011 DVDD.n20010 47.4925
R24 DVDD.n4613 DVDD.n4612 47.4925
R25 DVDD.n3879 DVDD.n3878 47.4925
R26 DVDD.n4717 DVDD.n4716 47.4925
R27 DVDD.n4712 DVDD.n4711 47.4925
R28 DVDD.n4839 DVDD.n4838 47.4925
R29 DVDD.n4823 DVDD.n4822 47.4925
R30 DVDD.n5144 DVDD.n5143 47.4925
R31 DVDD.n5111 DVDD.n5110 47.4925
R32 DVDD.n19640 DVDD.n19639 47.4925
R33 DVDD.n19637 DVDD.n19636 47.4925
R34 DVDD.n5235 DVDD.n5234 47.4925
R35 DVDD.n5230 DVDD.n5229 47.4925
R36 DVDD.n7742 DVDD.n7741 8.0005
R37 DVDD.n7744 DVDD.n7743 8.0005
R38 DVDD.n18282 DVDD.n18281 8.0005
R39 DVDD.n18284 DVDD.n18283 8.0005
R40 DVDD.n17172 DVDD.n17171 6.3005
R41 DVDD.n11203 DVDD.n11202 6.3005
R42 DVDD.n12916 DVDD.n12874 6.3005
R43 DVDD.n9023 DVDD.n8981 6.3005
R44 DVDD.n17290 DVDD.n17289 6.3005
R45 DVDD.n17288 DVDD.n17287 6.3005
R46 DVDD.n13905 DVDD.n13904 6.3005
R47 DVDD.n13907 DVDD.n13906 6.3005
R48 DVDD.n17585 DVDD.n17584 6.3005
R49 DVDD.n14206 DVDD.n14205 6.3005
R50 DVDD.n17666 DVDD.n17665 6.3005
R51 DVDD.n14293 DVDD.n14292 6.3005
R52 DVDD.n14296 DVDD.n14295 6.3005
R53 DVDD.n14295 DVDD.n14294 6.3005
R54 DVDD.n17669 DVDD.n17668 6.3005
R55 DVDD.n17668 DVDD.n17667 6.3005
R56 DVDD.n13911 DVDD.n13910 4.5005
R57 DVDD.n17294 DVDD.n17293 4.5005
R58 DVDD.n17673 DVDD.n17672 4.5005
R59 DVDD.n14300 DVDD.n14299 4.5005
R60 DVDD.n7766 DVDD 4.0005
R61 DVDD.n18285 DVDD 4.0005
R62 DVDD.n9815 DVDD.n9814 3.81094
R63 DVDD.n1545 DVDD.n1544 3.81094
R64 DVDD.n1674 DVDD.n959 3.81094
R65 DVDD.n11541 DVDD.n11418 3.81094
R66 DVDD.n9958 DVDD.n9957 3.81094
R67 DVDD.n3320 DVDD.n3319 3.81094
R68 DVDD.n1283 DVDD.n1121 3.81094
R69 DVDD.n11916 DVDD.n11915 3.81094
R70 DVDD.n12323 DVDD.n11306 3.81094
R71 DVDD.n7162 DVDD.n7161 3.81094
R72 DVDD.n18287 DVDD.n18286 3.81094
R73 DVDD.n3157 DVDD.n3031 3.81094
R74 DVDD.n9519 DVDD.n9518 3.81094
R75 DVDD.n1012 DVDD.n1011 3.81093
R76 DVDD.n1733 DVDD.n1732 3.81093
R77 DVDD.n1089 DVDD.n1088 3.81093
R78 DVDD.n11423 DVDD.n11422 3.81093
R79 DVDD.n1123 DVDD.n1122 3.81093
R80 DVDD.n7768 DVDD.n7767 3.80354
R81 DVDD.n3452 DVDD.n3451 3.80354
R82 DVDD.n3575 DVDD.n3574 3.80354
R83 DVDD.n3674 DVDD.n3673 3.80354
R84 DVDD.n2916 DVDD.n2915 3.80354
R85 DVDD.n3001 DVDD.n3000 3.80353
R86 DVDD.t19 DVDD.n7766 3.6505
R87 DVDD.n7767 DVDD.t19 3.6505
R88 DVDD.n18776 DVDD.t4 3.6505
R89 DVDD.n3451 DVDD.t14 3.6505
R90 DVDD.n3574 DVDD.t38 3.6505
R91 DVDD.n7161 DVDD.t11 3.6505
R92 DVDD.n7815 DVDD.t20 3.6505
R93 DVDD.n7935 DVDD.t35 3.6505
R94 DVDD.n8361 DVDD.t16 3.6505
R95 DVDD.n2054 DVDD.t29 3.6505
R96 DVDD.n2208 DVDD.t23 3.6505
R97 DVDD.n2231 DVDD.t24 3.6505
R98 DVDD.n7099 DVDD.t34 3.6505
R99 DVDD.n6937 DVDD.t27 3.6505
R100 DVDD.n6785 DVDD.t3 3.6505
R101 DVDD.n6552 DVDD.t22 3.6505
R102 DVDD.n1858 DVDD.t26 3.6505
R103 DVDD.n3924 DVDD.t30 3.6505
R104 DVDD.n19832 DVDD.t15 3.6505
R105 DVDD.n19987 DVDD.t39 3.6505
R106 DVDD.n20010 DVDD.t2 3.6505
R107 DVDD.n3878 DVDD.t17 3.6505
R108 DVDD.n4711 DVDD.t8 3.6505
R109 DVDD.n4822 DVDD.t21 3.6505
R110 DVDD.n5143 DVDD.t36 3.6505
R111 DVDD.n19636 DVDD.t10 3.6505
R112 DVDD.n5229 DVDD.t13 3.6505
R113 DVDD.n1544 DVDD.t7 3.6505
R114 DVDD.n959 DVDD.t32 3.6505
R115 DVDD.n1732 DVDD.t33 3.6505
R116 DVDD.n11422 DVDD.t40 3.6505
R117 DVDD.t12 DVDD.n18285 3.6505
R118 DVDD.n18286 DVDD.t12 3.6505
R119 DVDD.n11915 DVDD.t18 3.6505
R120 DVDD.n1122 DVDD.t1 3.6505
R121 DVDD.n11306 DVDD.t28 3.6505
R122 DVDD.n11299 DVDD.t5 3.6505
R123 DVDD.n3031 DVDD.t9 3.6505
R124 DVDD.n2054 DVDD.n2053 3.62748
R125 DVDD.n2208 DVDD.n2207 3.62748
R126 DVDD.n18930 DVDD.n18929 3.62748
R127 DVDD.n7032 DVDD.n7031 3.62748
R128 DVDD.n6942 DVDD.n6941 3.62748
R129 DVDD.n6801 DVDD.n6800 3.62748
R130 DVDD.n6552 DVDD.n6551 3.62748
R131 DVDD.n1861 DVDD.n1860 3.62748
R132 DVDD.n3929 DVDD.n3928 3.62748
R133 DVDD.n19832 DVDD.n19831 3.62748
R134 DVDD.n19987 DVDD.n19986 3.62748
R135 DVDD.n19048 DVDD.n19047 3.62748
R136 DVDD.n4612 DVDD.n4611 3.62748
R137 DVDD.n4716 DVDD.n4715 3.62748
R138 DVDD.n4838 DVDD.n4837 3.62748
R139 DVDD.n5143 DVDD.n5142 3.62748
R140 DVDD.n19639 DVDD.n19638 3.62748
R141 DVDD.n5234 DVDD.n5233 3.62748
R142 DVDD.n2023 DVDD.n2022 3.62747
R143 DVDD.n2155 DVDD.n2154 3.62747
R144 DVDD.n2231 DVDD.n2230 3.62747
R145 DVDD.n7099 DVDD.n7098 3.62747
R146 DVDD.n6937 DVDD.n6936 3.62747
R147 DVDD.n6785 DVDD.n6784 3.62747
R148 DVDD.n6519 DVDD.n6518 3.62747
R149 DVDD.n1858 DVDD.n1857 3.62747
R150 DVDD.n3924 DVDD.n3923 3.62747
R151 DVDD.n19801 DVDD.n19800 3.62747
R152 DVDD.n19934 DVDD.n19933 3.62747
R153 DVDD.n20010 DVDD.n20009 3.62747
R154 DVDD.n3878 DVDD.n3877 3.62747
R155 DVDD.n4711 DVDD.n4710 3.62747
R156 DVDD.n4822 DVDD.n4821 3.62747
R157 DVDD.n5110 DVDD.n5109 3.62747
R158 DVDD.n19636 DVDD.n19635 3.62747
R159 DVDD.n5229 DVDD.n5228 3.62747
R160 DVDD.n18777 DVDD.n18776 3.1796
R161 DVDD.n13889 DVDD.n13888 3.1505
R162 DVDD.n4241 DVDD.n4240 3.1505
R163 DVDD.n13885 DVDD.n13884 3.1505
R164 DVDD.n5799 DVDD.n5798 3.1505
R165 DVDD.n4230 DVDD.n4229 3.1505
R166 DVDD.n4222 DVDD.n4221 3.1505
R167 DVDD.n4226 DVDD.n4225 3.1505
R168 DVDD.n5801 DVDD.n5800 3.1505
R169 DVDD.n5791 DVDD.n5790 3.1505
R170 DVDD.n5793 DVDD.n5792 3.1505
R171 DVDD.n17269 DVDD.n17268 3.1505
R172 DVDD.n17280 DVDD.n17279 3.1505
R173 DVDD.n17276 DVDD.n17275 3.1505
R174 DVDD.n17272 DVDD.n17271 3.1505
R175 DVDD.n17284 DVDD.n17283 3.1505
R176 DVDD.n13893 DVDD.n13892 3.1505
R177 DVDD.n13897 DVDD.n13896 3.1505
R178 DVDD.n13901 DVDD.n13900 3.1505
R179 DVDD.n17406 DVDD.n17405 3.1505
R180 DVDD.n14000 DVDD.n13999 3.1505
R181 DVDD.n17239 DVDD.n17238 3.1505
R182 DVDD.n14089 DVDD.n14088 3.1505
R183 DVDD.n14209 DVDD.n14208 3.1505
R184 DVDD.n14208 DVDD.n14207 3.1505
R185 DVDD.n17588 DVDD.n17587 3.1505
R186 DVDD.n17587 DVDD.n17586 3.1505
R187 DVDD.n17592 DVDD.n17591 3.1505
R188 DVDD.n17650 DVDD.n17649 3.1505
R189 DVDD.n17654 DVDD.n17653 3.1505
R190 DVDD.n17658 DVDD.n17657 3.1505
R191 DVDD.n17662 DVDD.n17661 3.1505
R192 DVDD.n14289 DVDD.n14288 3.1505
R193 DVDD.n14285 DVDD.n14284 3.1505
R194 DVDD.n14281 DVDD.n14280 3.1505
R195 DVDD.n14277 DVDD.n14276 3.1505
R196 DVDD.n14273 DVDD.n14272 3.1505
R197 DVDD.n4174 DVDD.n4173 3.1505
R198 DVDD.n4170 DVDD.n4169 3.1505
R199 DVDD.n4339 DVDD.n4338 3.1505
R200 DVDD.n4343 DVDD.n4342 3.1505
R201 DVDD.n5785 DVDD.n5784 3.1505
R202 DVDD.n5781 DVDD.n5780 3.1505
R203 DVDD.n5777 DVDD.n5776 3.1505
R204 DVDD.n5773 DVDD.n5772 3.1505
R205 DVDD.n17647 DVDD.n17646 3.1505
R206 DVDD.n19430 DVDD.n19429 3.10835
R207 DVDD.n13224 DVDD.n13223 3.10835
R208 DVDD.n11341 DVDD.n11340 3.10835
R209 DVDD.n11338 DVDD.n11337 3.10835
R210 DVDD.n11300 DVDD.n11299 3.10835
R211 DVDD.n9313 DVDD.n9312 3.1048
R212 DVDD.n7816 DVDD.n7815 3.1048
R213 DVDD.n7936 DVDD.n7935 3.1048
R214 DVDD.n8362 DVDD.n8361 3.1048
R215 DVDD.n14141 DVDD.n14140 2.83716
R216 DVDD.n14255 DVDD.n14254 2.53461
R217 DVDD.n17264 DVDD.n17263 2.49083
R218 DVDD.n13916 DVDD.n13915 2.49083
R219 DVDD.n17642 DVDD.n17641 2.49083
R220 DVDD.n14305 DVDD.n14304 2.49083
R221 DVDD.n17623 DVDD.n17622 2.47025
R222 DVDD.n6110 DVDD.n6109 2.25096
R223 DVDD.n12740 DVDD.n12465 2.25096
R224 DVDD.n6122 DVDD.n4068 2.25096
R225 DVDD.n8824 DVDD.n8490 2.25096
R226 DVDD.n14431 DVDD.n11207 2.25095
R227 DVDD.n12758 DVDD.n12458 2.25091
R228 DVDD.n5576 DVDD.n5575 2.25073
R229 DVDD.n5623 DVDD.n5622 2.25073
R230 DVDD.n5669 DVDD.n5668 2.25073
R231 DVDD.n12850 DVDD.n12417 2.25073
R232 DVDD.n12813 DVDD.n12437 2.25073
R233 DVDD.n12777 DVDD.n12450 2.25073
R234 DVDD.n6230 DVDD.n4038 2.25073
R235 DVDD.n6192 DVDD.n4048 2.25073
R236 DVDD.n6154 DVDD.n4058 2.25073
R237 DVDD.n8932 DVDD.n8437 2.25073
R238 DVDD.n8894 DVDD.n8456 2.25073
R239 DVDD.n8856 DVDD.n8474 2.25073
R240 DVDD.n4505 DVDD.n4504 2.25073
R241 DVDD.n6092 DVDD.n5707 2.25069
R242 DVDD.n4542 DVDD.n4075 2.25069
R243 DVDD.n8809 DVDD.n8497 2.25069
R244 DVDD.n14449 DVDD.n11198 2.2505
R245 DVDD.n14449 DVDD.n14439 2.2505
R246 DVDD.n14449 DVDD.n14448 2.2505
R247 DVDD.n6017 DVDD.n5998 2.2505
R248 DVDD.n6017 DVDD.n6007 2.2505
R249 DVDD.n5307 DVDD.n5306 2.2505
R250 DVDD.n4747 DVDD.n4746 2.2505
R251 DVDD.n4652 DVDD.n4651 2.2505
R252 DVDD.n3887 DVDD.n3884 2.2505
R253 DVDD.n19992 DVDD.n19991 2.2505
R254 DVDD.n19837 DVDD.n19836 2.2505
R255 DVDD.n6017 DVDD.n6010 2.2505
R256 DVDD.n6017 DVDD.n6016 2.2505
R257 DVDD.n6040 DVDD.n6039 2.2505
R258 DVDD.n6069 DVDD.n6068 2.2505
R259 DVDD.n13151 DVDD.n13150 2.2505
R260 DVDD.n11573 DVDD.n11572 2.2505
R261 DVDD.n18331 DVDD.n18330 2.2505
R262 DVDD.n1680 DVDD.n1679 2.2505
R263 DVDD.n1539 DVDD.n1538 2.2505
R264 DVDD.n12668 DVDD.n12484 2.2505
R265 DVDD.n12668 DVDD.n12661 2.2505
R266 DVDD.n12668 DVDD.n12475 2.2505
R267 DVDD.n12668 DVDD.n12667 2.2505
R268 DVDD.n17282 DVDD.n17281 2.2505
R269 DVDD.n5803 DVDD.n5802 2.2505
R270 DVDD.n5789 DVDD.n5788 2.2505
R271 DVDD.n5795 DVDD.n5794 2.2505
R272 DVDD.n5813 DVDD.n5811 2.2505
R273 DVDD.n5797 DVDD.n5796 2.2505
R274 DVDD.n17278 DVDD.n17277 2.2505
R275 DVDD.n17274 DVDD.n17273 2.2505
R276 DVDD.n17270 DVDD.n17267 2.2505
R277 DVDD.n17286 DVDD.n17285 2.2505
R278 DVDD.n17818 DVDD.n17185 2.2505
R279 DVDD.n17818 DVDD.n17817 2.2505
R280 DVDD.n17818 DVDD.n17170 2.2505
R281 DVDD.n14005 DVDD.n14004 2.2505
R282 DVDD.n17411 DVDD.n17410 2.2505
R283 DVDD.n14094 DVDD.n14093 2.2505
R284 DVDD.n17244 DVDD.n17243 2.2505
R285 DVDD.n14215 DVDD.n14214 2.2505
R286 DVDD.n14214 DVDD.n14213 2.2505
R287 DVDD.n17594 DVDD.n17593 2.2505
R288 DVDD.n17648 DVDD.n17645 2.2505
R289 DVDD.n17652 DVDD.n17651 2.2505
R290 DVDD.n17656 DVDD.n17655 2.2505
R291 DVDD.n17660 DVDD.n17659 2.2505
R292 DVDD.n17664 DVDD.n17663 2.2505
R293 DVDD.n5783 DVDD.n5782 2.2505
R294 DVDD.n5787 DVDD.n5786 2.2505
R295 DVDD.n5775 DVDD.n5774 2.2505
R296 DVDD.n5779 DVDD.n5778 2.2505
R297 DVDD.n5875 DVDD.n5874 2.2505
R298 DVDD.n4345 DVDD.n4344 2.2505
R299 DVDD.n4468 DVDD.n4109 2.2505
R300 DVDD.n4468 DVDD.n4100 2.2505
R301 DVDD.n4491 DVDD.n4490 2.2505
R302 DVDD.n6453 DVDD.n4001 2.2505
R303 DVDD.n6973 DVDD.n6972 2.2505
R304 DVDD.n7108 DVDD.n7105 2.2505
R305 DVDD.n7072 DVDD.n7071 2.2505
R306 DVDD.n2213 DVDD.n2212 2.2505
R307 DVDD.n2059 DVDD.n2058 2.2505
R308 DVDD.n4468 DVDD.n4461 2.2505
R309 DVDD.n4468 DVDD.n4467 2.2505
R310 DVDD.n4172 DVDD.n4171 2.2505
R311 DVDD.n4176 DVDD.n4175 2.2505
R312 DVDD.n4168 DVDD.n4167 2.2505
R313 DVDD.n4341 DVDD.n4340 2.2505
R314 DVDD.n4519 DVDD.n4518 2.2505
R315 DVDD.n4232 DVDD.n4231 2.2505
R316 DVDD.n4220 DVDD.n4219 2.2505
R317 DVDD.n4228 DVDD.n4227 2.2505
R318 DVDD.n4224 DVDD.n4223 2.2505
R319 DVDD.n4243 DVDD.n4242 2.2505
R320 DVDD.n8754 DVDD.n8732 2.2505
R321 DVDD.n8754 DVDD.n8735 2.2505
R322 DVDD.n9240 DVDD.n9239 2.2505
R323 DVDD.n3569 DVDD.n3568 2.2505
R324 DVDD.n3458 DVDD.n3457 2.2505
R325 DVDD.n9990 DVDD.n9989 2.2505
R326 DVDD.n8754 DVDD.n8744 2.2505
R327 DVDD.n8754 DVDD.n8753 2.2505
R328 DVDD.n14291 DVDD.n14290 2.2505
R329 DVDD.n14287 DVDD.n14286 2.2505
R330 DVDD.n14283 DVDD.n14282 2.2505
R331 DVDD.n14279 DVDD.n14278 2.2505
R332 DVDD.n14275 DVDD.n14274 2.2505
R333 DVDD.n13891 DVDD.n13890 2.2505
R334 DVDD.n13895 DVDD.n13894 2.2505
R335 DVDD.n13899 DVDD.n13898 2.2505
R336 DVDD.n13903 DVDD.n13902 2.2505
R337 DVDD.n13887 DVDD.n13886 2.2505
R338 DVDD.n10053 DVDD.n7155 2.2505
R339 DVDD.n5814 DVDD.n5813 2.25042
R340 DVDD.n5816 DVDD.n5795 2.25042
R341 DVDD.n5880 DVDD.n5779 2.25042
R342 DVDD.n5878 DVDD.n5787 2.25042
R343 DVDD.n4244 DVDD.n4243 2.25042
R344 DVDD.n4246 DVDD.n4228 2.25042
R345 DVDD.n4346 DVDD.n4345 2.25042
R346 DVDD.n4334 DVDD.n4176 2.25042
R347 DVDD.n6070 DVDD.n5723 2.25038
R348 DVDD.n4520 DVDD.n4094 2.25038
R349 DVDD.n5578 DVDD.n4600 2.25034
R350 DVDD.n12848 DVDD.n12426 2.25034
R351 DVDD.n6228 DVDD.n4046 2.25034
R352 DVDD.n8930 DVDD.n8446 2.25034
R353 DVDD.n5625 DVDD.n4585 2.25025
R354 DVDD.n12811 DVDD.n12445 2.25025
R355 DVDD.n6190 DVDD.n4056 2.25025
R356 DVDD.n8892 DVDD.n8464 2.25025
R357 DVDD.n5671 DVDD.n4570 2.25016
R358 DVDD.n12726 DVDD.n12472 2.25016
R359 DVDD.n12775 DVDD.n12774 2.25016
R360 DVDD.n6152 DVDD.n4066 2.25016
R361 DVDD.n8854 DVDD.n8482 2.25016
R362 DVDD.n6107 DVDD.n6106 2.25011
R363 DVDD.n12738 DVDD.n12737 2.25011
R364 DVDD.n6120 DVDD.n6119 2.25011
R365 DVDD.n8822 DVDD.n8821 2.25011
R366 DVDD.n5809 DVDD.n5803 2.24737
R367 DVDD.n5876 DVDD.n5875 2.24737
R368 DVDD.n4238 DVDD.n4232 2.24737
R369 DVDD.n12919 DVDD.n12918 2.1005
R370 DVDD.n12918 DVDD.n12917 2.1005
R371 DVDD.n9026 DVDD.n9025 2.1005
R372 DVDD.n9025 DVDD.n9024 2.1005
R373 DVDD.n9034 DVDD.n9033 2.1005
R374 DVDD.n9033 DVDD.n9032 2.1005
R375 DVDD.n8979 DVDD.n8978 2.1005
R376 DVDD.n8978 DVDD.n8977 2.1005
R377 DVDD.n8973 DVDD.n8972 2.1005
R378 DVDD.n8972 DVDD.n8971 2.1005
R379 DVDD.n8965 DVDD.n8964 2.1005
R380 DVDD.n8964 DVDD.n8963 2.1005
R381 DVDD.n8957 DVDD.n8956 2.1005
R382 DVDD.n8956 DVDD.n8955 2.1005
R383 DVDD.n4032 DVDD.n4031 2.1005
R384 DVDD.n4031 DVDD.n4030 2.1005
R385 DVDD.n4023 DVDD.n4022 2.1005
R386 DVDD.n4022 DVDD.n4021 2.1005
R387 DVDD.n4017 DVDD.n4016 2.1005
R388 DVDD.n4016 DVDD.n4015 2.1005
R389 DVDD.n4009 DVDD.n4008 2.1005
R390 DVDD.n4008 DVDD.n4007 2.1005
R391 DVDD.n5537 DVDD.n5536 2.1005
R392 DVDD.n5536 DVDD.n5535 2.1005
R393 DVDD.n5525 DVDD.n5524 2.1005
R394 DVDD.n5524 DVDD.n5523 2.1005
R395 DVDD.n5519 DVDD.n5518 2.1005
R396 DVDD.n5518 DVDD.n5517 2.1005
R397 DVDD.n5511 DVDD.n5510 2.1005
R398 DVDD.n5510 DVDD.n5509 2.1005
R399 DVDD.n12940 DVDD.n12939 2.1005
R400 DVDD.n12939 DVDD.n12938 2.1005
R401 DVDD.n12927 DVDD.n12926 2.1005
R402 DVDD.n12926 DVDD.n12925 2.1005
R403 DVDD.n12935 DVDD.n12934 2.1005
R404 DVDD.n12934 DVDD.n12933 2.1005
R405 DVDD.n12954 DVDD.n12953 2.1005
R406 DVDD.n12953 DVDD.n12952 2.1005
R407 DVDD.n12946 DVDD.n12945 2.1005
R408 DVDD.n12945 DVDD.n12944 2.1005
R409 DVDD.n12915 DVDD.n12914 2.1005
R410 DVDD.n12914 DVDD.n12913 2.1005
R411 DVDD.n8992 DVDD.n8991 2.1005
R412 DVDD.n8991 DVDD.n8990 2.1005
R413 DVDD.n9014 DVDD.n9013 2.1005
R414 DVDD.n9013 DVDD.n9012 2.1005
R415 DVDD.n9022 DVDD.n9021 2.1005
R416 DVDD.n9021 DVDD.n9020 2.1005
R417 DVDD.n9006 DVDD.n9005 2.1005
R418 DVDD.n9005 DVDD.n9004 2.1005
R419 DVDD.n9000 DVDD.n8999 2.1005
R420 DVDD.n8999 DVDD.n8998 2.1005
R421 DVDD.n8984 DVDD.n8983 2.1005
R422 DVDD.n8983 DVDD.n8982 2.1005
R423 DVDD.n4500 DVDD.n4499 2.1005
R424 DVDD.n4499 DVDD.n4498 2.1005
R425 DVDD.n5715 DVDD.n5714 2.1005
R426 DVDD.n5714 DVDD.n5713 2.1005
R427 DVDD.n6057 DVDD.n6056 2.1005
R428 DVDD.n6056 DVDD.n6055 2.1005
R429 DVDD.n4086 DVDD.n4085 2.1005
R430 DVDD.n4085 DVDD.n4084 2.1005
R431 DVDD.n4515 DVDD.n4514 2.1005
R432 DVDD.n4514 DVDD.n4513 2.1005
R433 DVDD.n4090 DVDD.n4089 2.1005
R434 DVDD.n4089 DVDD.n4088 2.1005
R435 DVDD.n6065 DVDD.n6064 2.1005
R436 DVDD.n6064 DVDD.n6063 2.1005
R437 DVDD.n5719 DVDD.n5718 2.1005
R438 DVDD.n5718 DVDD.n5717 2.1005
R439 DVDD.n12881 DVDD.n12880 2.1005
R440 DVDD.n12880 DVDD.n12879 2.1005
R441 DVDD.n12895 DVDD.n12894 2.1005
R442 DVDD.n12894 DVDD.n12893 2.1005
R443 DVDD.n12907 DVDD.n12906 2.1005
R444 DVDD.n12906 DVDD.n12905 2.1005
R445 DVDD.n12899 DVDD.n12898 2.1005
R446 DVDD.n12898 DVDD.n12897 2.1005
R447 DVDD.n12887 DVDD.n12886 2.1005
R448 DVDD.n12886 DVDD.n12885 2.1005
R449 DVDD.n17389 DVDD.n17388 2.1005
R450 DVDD.n17381 DVDD.n17380 2.1005
R451 DVDD.n17377 DVDD.n17376 2.1005
R452 DVDD.n17373 DVDD.n17372 2.1005
R453 DVDD.n17369 DVDD.n17368 2.1005
R454 DVDD.n4212 DVDD.n4211 2.1005
R455 DVDD.n4216 DVDD.n4215 2.1005
R456 DVDD.n4256 DVDD.n4255 2.1005
R457 DVDD.n4260 DVDD.n4259 2.1005
R458 DVDD.n13979 DVDD.n13978 2.1005
R459 DVDD.n13983 DVDD.n13982 2.1005
R460 DVDD.n13987 DVDD.n13986 2.1005
R461 DVDD.n13991 DVDD.n13990 2.1005
R462 DVDD.n13995 DVDD.n13994 2.1005
R463 DVDD.n17397 DVDD.n17396 2.1005
R464 DVDD.n17401 DVDD.n17400 2.1005
R465 DVDD.n17393 DVDD.n17392 2.1005
R466 DVDD.n17385 DVDD.n17384 2.1005
R467 DVDD.n17234 DVDD.n17233 2.1005
R468 DVDD.n17230 DVDD.n17229 2.1005
R469 DVDD.n17226 DVDD.n17225 2.1005
R470 DVDD.n17222 DVDD.n17221 2.1005
R471 DVDD.n17218 DVDD.n17217 2.1005
R472 DVDD.n17214 DVDD.n17213 2.1005
R473 DVDD.n17210 DVDD.n17209 2.1005
R474 DVDD.n17206 DVDD.n17205 2.1005
R475 DVDD.n17202 DVDD.n17201 2.1005
R476 DVDD.n4200 DVDD.n4199 2.1005
R477 DVDD.n4204 DVDD.n4203 2.1005
R478 DVDD.n4281 DVDD.n4280 2.1005
R479 DVDD.n4285 DVDD.n4284 2.1005
R480 DVDD.n14068 DVDD.n14067 2.1005
R481 DVDD.n14072 DVDD.n14071 2.1005
R482 DVDD.n14076 DVDD.n14075 2.1005
R483 DVDD.n14080 DVDD.n14079 2.1005
R484 DVDD.n14084 DVDD.n14083 2.1005
R485 DVDD.n14182 DVDD.n14181 2.1005
R486 DVDD.n14201 DVDD.n14200 2.1005
R487 DVDD.n14200 DVDD.n14199 2.1005
R488 DVDD.n14195 DVDD.n14194 2.1005
R489 DVDD.n14194 DVDD.n14193 2.1005
R490 DVDD.n14189 DVDD.n14188 2.1005
R491 DVDD.n14188 DVDD.n14187 2.1005
R492 DVDD.n14183 DVDD.n14182 2.1005
R493 DVDD.n14177 DVDD.n14176 2.1005
R494 DVDD.n14176 DVDD.n14175 2.1005
R495 DVDD.n4315 DVDD.n4314 2.1005
R496 DVDD.n4314 DVDD.n4313 2.1005
R497 DVDD.n4307 DVDD.n4306 2.1005
R498 DVDD.n4306 DVDD.n4305 2.1005
R499 DVDD.n4193 DVDD.n4192 2.1005
R500 DVDD.n4192 DVDD.n4191 2.1005
R501 DVDD.n4185 DVDD.n4184 2.1005
R502 DVDD.n4184 DVDD.n4183 2.1005
R503 DVDD.n17550 DVDD.n17549 2.1005
R504 DVDD.n17549 DVDD.n17548 2.1005
R505 DVDD.n17554 DVDD.n17553 2.1005
R506 DVDD.n17553 DVDD.n17552 2.1005
R507 DVDD.n17558 DVDD.n17557 2.1005
R508 DVDD.n17557 DVDD.n17556 2.1005
R509 DVDD.n17562 DVDD.n17561 2.1005
R510 DVDD.n17561 DVDD.n17560 2.1005
R511 DVDD.n17566 DVDD.n17565 2.1005
R512 DVDD.n17565 DVDD.n17564 2.1005
R513 DVDD.n17570 DVDD.n17569 2.1005
R514 DVDD.n17569 DVDD.n17568 2.1005
R515 DVDD.n17574 DVDD.n17573 2.1005
R516 DVDD.n17573 DVDD.n17572 2.1005
R517 DVDD.n17578 DVDD.n17577 2.1005
R518 DVDD.n17577 DVDD.n17576 2.1005
R519 DVDD.n17582 DVDD.n17581 2.1005
R520 DVDD.n17581 DVDD.n17580 2.1005
R521 DVDD.n14220 DVDD.n14218 1.6285
R522 DVDD.n17516 DVDD.n17514 1.62213
R523 DVDD.n17182 DVDD.n17181 1.5755
R524 DVDD.n17181 DVDD.n17180 1.5755
R525 DVDD.n17811 DVDD.n17810 1.5755
R526 DVDD.n17810 DVDD.n17809 1.5755
R527 DVDD.n17814 DVDD.n17813 1.5755
R528 DVDD.n17813 DVDD.n17812 1.5755
R529 DVDD.n12478 DVDD.n12477 1.5755
R530 DVDD.n12477 DVDD.n12476 1.5755
R531 DVDD.n12481 DVDD.n12480 1.5755
R532 DVDD.n12480 DVDD.n12479 1.5755
R533 DVDD.n12658 DVDD.n12657 1.5755
R534 DVDD.n12657 DVDD.n12656 1.5755
R535 DVDD.n12664 DVDD.n12663 1.5755
R536 DVDD.n12663 DVDD.n12662 1.5755
R537 DVDD.n6001 DVDD.n6000 1.5755
R538 DVDD.n6000 DVDD.n5999 1.5755
R539 DVDD.n6004 DVDD.n6003 1.5755
R540 DVDD.n6003 DVDD.n6002 1.5755
R541 DVDD.n5995 DVDD.n5994 1.5755
R542 DVDD.n5994 DVDD.n5993 1.5755
R543 DVDD.n6013 DVDD.n6012 1.5755
R544 DVDD.n6012 DVDD.n6011 1.5755
R545 DVDD.n4106 DVDD.n4105 1.5755
R546 DVDD.n4105 DVDD.n4104 1.5755
R547 DVDD.n4458 DVDD.n4457 1.5755
R548 DVDD.n4457 DVDD.n4456 1.5755
R549 DVDD.n4097 DVDD.n4096 1.5755
R550 DVDD.n4096 DVDD.n4095 1.5755
R551 DVDD.n4464 DVDD.n4463 1.5755
R552 DVDD.n4463 DVDD.n4462 1.5755
R553 DVDD.n8738 DVDD.n8737 1.5755
R554 DVDD.n8737 DVDD.n8736 1.5755
R555 DVDD.n8741 DVDD.n8740 1.5755
R556 DVDD.n8740 DVDD.n8739 1.5755
R557 DVDD.n8747 DVDD.n8746 1.5755
R558 DVDD.n8746 DVDD.n8745 1.5755
R559 DVDD.n8750 DVDD.n8749 1.5755
R560 DVDD.n8749 DVDD.n8748 1.5755
R561 DVDD.n14436 DVDD.n14435 1.5755
R562 DVDD.n14435 DVDD.n14434 1.5755
R563 DVDD.n14442 DVDD.n14441 1.5755
R564 DVDD.n14441 DVDD.n14440 1.5755
R565 DVDD.n14445 DVDD.n14444 1.5755
R566 DVDD.n14444 DVDD.n14443 1.5755
R567 DVDD.n5916 DVDD.n5915 1.5755
R568 DVDD.n5915 DVDD.n5914 1.5755
R569 DVDD.n5906 DVDD.n5905 1.5755
R570 DVDD.n5905 DVDD.n5904 1.5755
R571 DVDD.n5910 DVDD.n5909 1.5755
R572 DVDD.n5909 DVDD.n5908 1.5755
R573 DVDD.n5898 DVDD.n5897 1.5755
R574 DVDD.n5897 DVDD.n5896 1.5755
R575 DVDD.n17705 DVDD.n17704 1.5755
R576 DVDD.n17704 DVDD.n17703 1.5755
R577 DVDD.n17711 DVDD.n17710 1.5755
R578 DVDD.n17710 DVDD.n17709 1.5755
R579 DVDD.n17732 DVDD.n17731 1.5755
R580 DVDD.n17731 DVDD.n17730 1.5755
R581 DVDD.n17726 DVDD.n17725 1.5755
R582 DVDD.n17725 DVDD.n17724 1.5755
R583 DVDD.n17720 DVDD.n17719 1.5755
R584 DVDD.n17719 DVDD.n17718 1.5755
R585 DVDD.n17714 DVDD.n17713 1.5755
R586 DVDD.n17713 DVDD.n17712 1.5755
R587 DVDD.n5892 DVDD.n5891 1.5755
R588 DVDD.n5891 DVDD.n5890 1.5755
R589 DVDD.n4361 DVDD.n4360 1.5755
R590 DVDD.n4360 DVDD.n4359 1.5755
R591 DVDD.n4373 DVDD.n4372 1.5755
R592 DVDD.n4372 DVDD.n4371 1.5755
R593 DVDD.n4367 DVDD.n4366 1.5755
R594 DVDD.n4366 DVDD.n4365 1.5755
R595 DVDD.n8629 DVDD.n8628 1.5755
R596 DVDD.n8628 DVDD.n8627 1.5755
R597 DVDD.n8635 DVDD.n8634 1.5755
R598 DVDD.n8634 DVDD.n8633 1.5755
R599 DVDD.n8647 DVDD.n8646 1.5755
R600 DVDD.n8646 DVDD.n8645 1.5755
R601 DVDD.n8641 DVDD.n8640 1.5755
R602 DVDD.n8640 DVDD.n8639 1.5755
R603 DVDD.n14330 DVDD.n14329 1.5755
R604 DVDD.n14329 DVDD.n14328 1.5755
R605 DVDD.n14352 DVDD.n14351 1.5755
R606 DVDD.n14351 DVDD.n14350 1.5755
R607 DVDD.n14346 DVDD.n14345 1.5755
R608 DVDD.n14345 DVDD.n14344 1.5755
R609 DVDD.n14340 DVDD.n14339 1.5755
R610 DVDD.n14339 DVDD.n14338 1.5755
R611 DVDD.n14102 DVDD.n14101 1.5755
R612 DVDD.n17192 DVDD.n17191 1.5755
R613 DVDD.n19054 DVDD.n19053 1.5005
R614 DVDD.n20050 DVDD.n20049 1.5005
R615 DVDD.n4899 DVDD.n4898 1.5005
R616 DVDD.n5163 DVDD.n5162 1.5005
R617 DVDD.n5533 DVDD.n5532 1.5005
R618 DVDD.n5532 DVDD.n5531 1.5005
R619 DVDD.n5541 DVDD.n5540 1.5005
R620 DVDD.n5540 DVDD.n5539 1.5005
R621 DVDD.n5522 DVDD.n5521 1.5005
R622 DVDD.n5521 DVDD.n5520 1.5005
R623 DVDD.n5515 DVDD.n5514 1.5005
R624 DVDD.n5514 DVDD.n5513 1.5005
R625 DVDD.n5507 DVDD.n5506 1.5005
R626 DVDD.n5506 DVDD.n5505 1.5005
R627 DVDD.n6039 DVDD.n6038 1.5005
R628 DVDD.n6038 DVDD.n6037 1.5005
R629 DVDD.n6061 DVDD.n6060 1.5005
R630 DVDD.n6060 DVDD.n6059 1.5005
R631 DVDD.n6068 DVDD.n6067 1.5005
R632 DVDD.n6067 DVDD.n6066 1.5005
R633 DVDD.n5723 DVDD.n5722 1.5005
R634 DVDD.n5722 DVDD.n5721 1.5005
R635 DVDD.n5711 DVDD.n5710 1.5005
R636 DVDD.n5710 DVDD.n5709 1.5005
R637 DVDD.n12911 DVDD.n12910 1.5005
R638 DVDD.n1723 DVDD.n1722 1.5005
R639 DVDD.n19436 DVDD.n19435 1.5005
R640 DVDD.n11854 DVDD.n11853 1.5005
R641 DVDD.n12344 DVDD.n12343 1.5005
R642 DVDD.n12931 DVDD.n12930 1.5005
R643 DVDD.n12930 DVDD.n12929 1.5005
R644 DVDD.n12957 DVDD.n12956 1.5005
R645 DVDD.n12956 DVDD.n12955 1.5005
R646 DVDD.n12950 DVDD.n12949 1.5005
R647 DVDD.n12949 DVDD.n12948 1.5005
R648 DVDD.n12942 DVDD.n12937 1.5005
R649 DVDD.n12937 DVDD.n12936 1.5005
R650 DVDD.n12910 DVDD.n12909 1.5005
R651 DVDD.n12903 DVDD.n12902 1.5005
R652 DVDD.n12902 DVDD.n12901 1.5005
R653 DVDD.n12896 DVDD.n12876 1.5005
R654 DVDD.n12876 DVDD.n12875 1.5005
R655 DVDD.n12891 DVDD.n12890 1.5005
R656 DVDD.n12890 DVDD.n12889 1.5005
R657 DVDD.n12883 DVDD.n12878 1.5005
R658 DVDD.n12878 DVDD.n12877 1.5005
R659 DVDD.n12923 DVDD.n12922 1.5005
R660 DVDD.n12922 DVDD.n12921 1.5005
R661 DVDD.n17379 DVDD.n17378 1.5005
R662 DVDD.n17375 DVDD.n17374 1.5005
R663 DVDD.n17371 DVDD.n17370 1.5005
R664 DVDD.n17367 DVDD.n17366 1.5005
R665 DVDD.n17403 DVDD.n17402 1.5005
R666 DVDD.n17399 DVDD.n17398 1.5005
R667 DVDD.n17395 DVDD.n17394 1.5005
R668 DVDD.n17391 DVDD.n17390 1.5005
R669 DVDD.n17387 DVDD.n17386 1.5005
R670 DVDD.n17383 DVDD.n17382 1.5005
R671 DVDD.n17236 DVDD.n17235 1.5005
R672 DVDD.n17232 DVDD.n17231 1.5005
R673 DVDD.n17228 DVDD.n17227 1.5005
R674 DVDD.n17224 DVDD.n17223 1.5005
R675 DVDD.n17220 DVDD.n17219 1.5005
R676 DVDD.n17216 DVDD.n17215 1.5005
R677 DVDD.n17212 DVDD.n17211 1.5005
R678 DVDD.n17208 DVDD.n17207 1.5005
R679 DVDD.n17204 DVDD.n17203 1.5005
R680 DVDD.n17200 DVDD.n17199 1.5005
R681 DVDD.n17547 DVDD.n17546 1.5005
R682 DVDD.n17546 DVDD.n17545 1.5005
R683 DVDD.n17551 DVDD.n17544 1.5005
R684 DVDD.n17544 DVDD.n17543 1.5005
R685 DVDD.n17555 DVDD.n17542 1.5005
R686 DVDD.n17542 DVDD.n17541 1.5005
R687 DVDD.n17559 DVDD.n17540 1.5005
R688 DVDD.n17540 DVDD.n17539 1.5005
R689 DVDD.n17563 DVDD.n17538 1.5005
R690 DVDD.n17538 DVDD.n17537 1.5005
R691 DVDD.n17567 DVDD.n17536 1.5005
R692 DVDD.n17536 DVDD.n17535 1.5005
R693 DVDD.n17571 DVDD.n17534 1.5005
R694 DVDD.n17534 DVDD.n17533 1.5005
R695 DVDD.n17575 DVDD.n17532 1.5005
R696 DVDD.n17532 DVDD.n17531 1.5005
R697 DVDD.n17579 DVDD.n17530 1.5005
R698 DVDD.n17530 DVDD.n17529 1.5005
R699 DVDD.n17583 DVDD.n17528 1.5005
R700 DVDD.n17528 DVDD.n17527 1.5005
R701 DVDD.n2271 DVDD.n2270 1.5005
R702 DVDD.n18946 DVDD.n18935 1.5005
R703 DVDD.n6862 DVDD.n6861 1.5005
R704 DVDD.n6572 DVDD.n6571 1.5005
R705 DVDD.n4210 DVDD.n4209 1.5005
R706 DVDD.n4218 DVDD.n4217 1.5005
R707 DVDD.n4214 DVDD.n4213 1.5005
R708 DVDD.n4262 DVDD.n4261 1.5005
R709 DVDD.n4258 DVDD.n4257 1.5005
R710 DVDD.n4198 DVDD.n4197 1.5005
R711 DVDD.n4206 DVDD.n4205 1.5005
R712 DVDD.n4202 DVDD.n4201 1.5005
R713 DVDD.n4287 DVDD.n4286 1.5005
R714 DVDD.n4283 DVDD.n4282 1.5005
R715 DVDD.n4312 DVDD.n4311 1.5005
R716 DVDD.n4311 DVDD.n4310 1.5005
R717 DVDD.n4316 DVDD.n4309 1.5005
R718 DVDD.n4309 DVDD.n4308 1.5005
R719 DVDD.n4190 DVDD.n4189 1.5005
R720 DVDD.n4189 DVDD.n4188 1.5005
R721 DVDD.n4194 DVDD.n4187 1.5005
R722 DVDD.n4187 DVDD.n4186 1.5005
R723 DVDD.n4182 DVDD.n4181 1.5005
R724 DVDD.n4181 DVDD.n4180 1.5005
R725 DVDD.n4028 DVDD.n4027 1.5005
R726 DVDD.n4027 DVDD.n4026 1.5005
R727 DVDD.n4036 DVDD.n4035 1.5005
R728 DVDD.n4035 DVDD.n4034 1.5005
R729 DVDD.n4020 DVDD.n4019 1.5005
R730 DVDD.n4019 DVDD.n4018 1.5005
R731 DVDD.n4013 DVDD.n4012 1.5005
R732 DVDD.n4012 DVDD.n4011 1.5005
R733 DVDD.n4005 DVDD.n4004 1.5005
R734 DVDD.n4004 DVDD.n4003 1.5005
R735 DVDD.n4504 DVDD.n4503 1.5005
R736 DVDD.n4503 DVDD.n4502 1.5005
R737 DVDD.n4518 DVDD.n4517 1.5005
R738 DVDD.n4517 DVDD.n4516 1.5005
R739 DVDD.n4094 DVDD.n4093 1.5005
R740 DVDD.n4093 DVDD.n4092 1.5005
R741 DVDD.n4082 DVDD.n4081 1.5005
R742 DVDD.n4081 DVDD.n4080 1.5005
R743 DVDD.n4490 DVDD.n4488 1.5005
R744 DVDD.n4488 DVDD.n4487 1.5005
R745 DVDD.n9753 DVDD.n9752 1.5005
R746 DVDD.n9540 DVDD.n9539 1.5005
R747 DVDD.n13981 DVDD.n13980 1.5005
R748 DVDD.n13985 DVDD.n13984 1.5005
R749 DVDD.n13989 DVDD.n13988 1.5005
R750 DVDD.n13993 DVDD.n13992 1.5005
R751 DVDD.n13997 DVDD.n13996 1.5005
R752 DVDD.n14070 DVDD.n14069 1.5005
R753 DVDD.n14074 DVDD.n14073 1.5005
R754 DVDD.n14078 DVDD.n14077 1.5005
R755 DVDD.n14082 DVDD.n14081 1.5005
R756 DVDD.n14086 DVDD.n14085 1.5005
R757 DVDD.n14204 DVDD.n14203 1.5005
R758 DVDD.n14203 DVDD.n14202 1.5005
R759 DVDD.n14198 DVDD.n14197 1.5005
R760 DVDD.n14197 DVDD.n14196 1.5005
R761 DVDD.n14192 DVDD.n14191 1.5005
R762 DVDD.n14191 DVDD.n14190 1.5005
R763 DVDD.n14186 DVDD.n14185 1.5005
R764 DVDD.n14185 DVDD.n14184 1.5005
R765 DVDD.n14180 DVDD.n14179 1.5005
R766 DVDD.n14179 DVDD.n14178 1.5005
R767 DVDD.n9030 DVDD.n9029 1.5005
R768 DVDD.n9029 DVDD.n9028 1.5005
R769 DVDD.n9038 DVDD.n9037 1.5005
R770 DVDD.n9037 DVDD.n9036 1.5005
R771 DVDD.n8976 DVDD.n8975 1.5005
R772 DVDD.n8975 DVDD.n8974 1.5005
R773 DVDD.n8969 DVDD.n8968 1.5005
R774 DVDD.n8968 DVDD.n8967 1.5005
R775 DVDD.n8961 DVDD.n8960 1.5005
R776 DVDD.n8960 DVDD.n8959 1.5005
R777 DVDD.n9018 DVDD.n9017 1.5005
R778 DVDD.n9017 DVDD.n9016 1.5005
R779 DVDD.n9010 DVDD.n9009 1.5005
R780 DVDD.n9009 DVDD.n9008 1.5005
R781 DVDD.n9003 DVDD.n9002 1.5005
R782 DVDD.n9002 DVDD.n9001 1.5005
R783 DVDD.n8996 DVDD.n8995 1.5005
R784 DVDD.n8995 DVDD.n8994 1.5005
R785 DVDD.n8988 DVDD.n8987 1.5005
R786 DVDD.n8987 DVDD.n8986 1.5005
R787 DVDD.n18783 DVDD.n18782 1.5005
R788 DVDD.n3715 DVDD.n3714 1.5005
R789 DVDD.n4265 DVDD.n4218 1.50017
R790 DVDD.n4290 DVDD.n4206 1.50017
R791 DVDD.n4319 DVDD.n4194 1.50017
R792 DVDD.n4263 DVDD.n4262 1.50013
R793 DVDD.n4288 DVDD.n4287 1.50013
R794 DVDD.n4317 DVDD.n4316 1.50013
R795 DVDD.n5542 DVDD.n5541 1.49676
R796 DVDD.n6253 DVDD.n4036 1.49676
R797 DVDD.n13975 DVDD.n13974 1.39476
R798 DVDD.n13971 DVDD.n13970 1.39476
R799 DVDD.n13955 DVDD.n13954 1.39476
R800 DVDD.n13946 DVDD.n13943 1.39476
R801 DVDD.n13939 DVDD.n13938 1.39476
R802 DVDD.n13934 DVDD.n13933 1.39476
R803 DVDD.n13929 DVDD.n13928 1.39476
R804 DVDD.n13924 DVDD.n13922 1.39476
R805 DVDD.n17253 DVDD.n17252 1.39476
R806 DVDD.n17249 DVDD.n17248 1.39476
R807 DVDD.n17448 DVDD.n17447 1.39476
R808 DVDD.n17439 DVDD.n17438 1.39476
R809 DVDD.n17432 DVDD.n17431 1.39476
R810 DVDD.n17427 DVDD.n17426 1.39476
R811 DVDD.n17422 DVDD.n17421 1.39476
R812 DVDD.n17352 DVDD.n17351 1.39476
R813 DVDD.n17348 DVDD.n17347 1.39476
R814 DVDD.n17332 DVDD.n17331 1.39476
R815 DVDD.n17323 DVDD.n17320 1.39476
R816 DVDD.n17316 DVDD.n17315 1.39476
R817 DVDD.n17311 DVDD.n17310 1.39476
R818 DVDD.n17306 DVDD.n17305 1.39476
R819 DVDD.n17301 DVDD.n17300 1.39476
R820 DVDD.n14167 DVDD.n14166 1.39476
R821 DVDD.n14170 DVDD.n14169 1.39476
R822 DVDD.n14150 DVDD.n14149 1.39476
R823 DVDD.n14142 DVDD.n14138 1.39476
R824 DVDD.n14134 DVDD.n14133 1.39476
R825 DVDD.n14128 DVDD.n14127 1.39476
R826 DVDD.n14124 DVDD.n14123 1.39476
R827 DVDD.n14115 DVDD.n14114 1.39476
R828 DVDD.n14111 DVDD.n14110 1.39476
R829 DVDD.n14052 DVDD.n14051 1.39476
R830 DVDD.n14043 DVDD.n14040 1.39476
R831 DVDD.n14036 DVDD.n14035 1.39476
R832 DVDD.n14031 DVDD.n14030 1.39476
R833 DVDD.n14026 DVDD.n14025 1.39476
R834 DVDD.n17681 DVDD.n17679 1.39476
R835 DVDD.n17681 DVDD.n17680 1.39476
R836 DVDD.n17636 DVDD.n17635 1.39476
R837 DVDD.n17631 DVDD.n17630 1.39476
R838 DVDD.n17623 DVDD.n17618 1.39476
R839 DVDD.n17623 DVDD.n17619 1.39476
R840 DVDD.n17613 DVDD.n17612 1.39476
R841 DVDD.n17608 DVDD.n17607 1.39476
R842 DVDD.n17603 DVDD.n17602 1.39476
R843 DVDD.n17511 DVDD.n17510 1.39476
R844 DVDD.n17507 DVDD.n17506 1.39476
R845 DVDD.n17491 DVDD.n17490 1.39476
R846 DVDD.n17482 DVDD.n17481 1.39476
R847 DVDD.n17475 DVDD.n17474 1.39476
R848 DVDD.n17470 DVDD.n17469 1.39476
R849 DVDD.n17465 DVDD.n17464 1.39476
R850 DVDD.n14314 DVDD.n14312 1.39476
R851 DVDD.n14314 DVDD.n14313 1.39476
R852 DVDD.n14268 DVDD.n14267 1.39476
R853 DVDD.n14263 DVDD.n14262 1.39476
R854 DVDD.n14255 DVDD.n14251 1.39476
R855 DVDD.n14255 DVDD.n14252 1.39476
R856 DVDD.n14246 DVDD.n14245 1.39476
R857 DVDD.n14241 DVDD.n14240 1.39476
R858 DVDD.n14237 DVDD.n14236 1.39476
R859 DVDD.n13930 DVDD.n13929 1.313
R860 DVDD.n13935 DVDD.n13934 1.313
R861 DVDD.n13940 DVDD.n13939 1.313
R862 DVDD.n13951 DVDD.n13950 1.313
R863 DVDD.n13956 DVDD.n13955 1.313
R864 DVDD.n13972 DVDD.n13971 1.313
R865 DVDD.n13976 DVDD.n13975 1.313
R866 DVDD.n17302 DVDD.n17301 1.313
R867 DVDD.n17258 DVDD.n17186 1.313
R868 DVDD.n14315 DVDD.n14314 1.313
R869 DVDD.n13925 DVDD.n13924 1.313
R870 DVDD.n17418 DVDD.n17417 1.313
R871 DVDD.n17423 DVDD.n17422 1.313
R872 DVDD.n17428 DVDD.n17427 1.313
R873 DVDD.n17433 DVDD.n17432 1.313
R874 DVDD.n17444 DVDD.n17443 1.313
R875 DVDD.n17449 DVDD.n17448 1.313
R876 DVDD.n17250 DVDD.n17249 1.313
R877 DVDD.n17254 DVDD.n17253 1.313
R878 DVDD.n17307 DVDD.n17306 1.313
R879 DVDD.n17312 DVDD.n17311 1.313
R880 DVDD.n17317 DVDD.n17316 1.313
R881 DVDD.n17328 DVDD.n17327 1.313
R882 DVDD.n17333 DVDD.n17332 1.313
R883 DVDD.n17349 DVDD.n17348 1.313
R884 DVDD.n17353 DVDD.n17352 1.313
R885 DVDD.n14116 DVDD.n14115 1.313
R886 DVDD.n14112 DVDD.n14111 1.313
R887 DVDD.n14053 DVDD.n14052 1.313
R888 DVDD.n14048 DVDD.n14047 1.313
R889 DVDD.n14037 DVDD.n14036 1.313
R890 DVDD.n14032 DVDD.n14031 1.313
R891 DVDD.n14027 DVDD.n14026 1.313
R892 DVDD.n14022 DVDD.n14021 1.313
R893 DVDD.n17466 DVDD.n17465 1.313
R894 DVDD.n17471 DVDD.n17470 1.313
R895 DVDD.n17476 DVDD.n17475 1.313
R896 DVDD.n17487 DVDD.n17486 1.313
R897 DVDD.n17492 DVDD.n17491 1.313
R898 DVDD.n17508 DVDD.n17507 1.313
R899 DVDD.n17512 DVDD.n17511 1.313
R900 DVDD.n14238 DVDD.n14237 1.313
R901 DVDD.n14243 DVDD.n14241 1.313
R902 DVDD.n14248 DVDD.n14246 1.313
R903 DVDD.n14260 DVDD.n14258 1.313
R904 DVDD.n14265 DVDD.n14263 1.313
R905 DVDD.n14270 DVDD.n14268 1.313
R906 DVDD.n14233 DVDD.n14165 1.313
R907 DVDD.n14173 DVDD.n14167 1.313
R908 DVDD.n14171 DVDD.n14170 1.313
R909 DVDD.n14152 DVDD.n14150 1.313
R910 DVDD.n14147 DVDD.n14146 1.313
R911 DVDD.n14135 DVDD.n14134 1.313
R912 DVDD.n14130 DVDD.n14128 1.313
R913 DVDD.n14125 DVDD.n14124 1.313
R914 DVDD.n14120 DVDD.n14066 1.313
R915 DVDD.n17605 DVDD.n17603 1.313
R916 DVDD.n17610 DVDD.n17608 1.313
R917 DVDD.n17615 DVDD.n17613 1.313
R918 DVDD.n17628 DVDD.n17626 1.313
R919 DVDD.n17633 DVDD.n17631 1.313
R920 DVDD.n17638 DVDD.n17636 1.313
R921 DVDD.n17683 DVDD.n17681 1.313
R922 DVDD.n17600 DVDD.n17599 1.313
R923 DVDD.n6117 DVDD.t25 1.30762
R924 DVDD.n4572 DVDD.t37 1.30762
R925 DVDD.n4587 DVDD.t31 1.30762
R926 DVDD.n4557 DVDD.t6 1.30762
R927 DVDD.n14254 DVDD.n14253 1.23378
R928 DVDD.n2755 DVDD.n2754 1.19477
R929 DVDD.n791 DVDD.n790 1.19477
R930 DVDD.n14813 DVDD.n14812 1.19194
R931 DVDD.n18225 DVDD.n18224 1.19194
R932 DVDD.n14439 DVDD.n14438 1.1255
R933 DVDD.n14438 DVDD.n14437 1.1255
R934 DVDD.n11198 DVDD.n11197 1.1255
R935 DVDD.n11197 DVDD.n11196 1.1255
R936 DVDD.n14448 DVDD.n14447 1.1255
R937 DVDD.n14447 DVDD.n14446 1.1255
R938 DVDD.n11201 DVDD.n11200 1.1255
R939 DVDD.n11200 DVDD.n11199 1.1255
R940 DVDD.n14355 DVDD.n14354 1.1255
R941 DVDD.n14354 DVDD.n14353 1.1255
R942 DVDD.n14349 DVDD.n14348 1.1255
R943 DVDD.n14348 DVDD.n14347 1.1255
R944 DVDD.n14343 DVDD.n14342 1.1255
R945 DVDD.n14342 DVDD.n14341 1.1255
R946 DVDD.n14337 DVDD.n14336 1.1255
R947 DVDD.n14336 DVDD.n14335 1.1255
R948 DVDD.n5919 DVDD.n5918 1.1255
R949 DVDD.n6007 DVDD.n6006 1.1255
R950 DVDD.n6006 DVDD.n6005 1.1255
R951 DVDD.n6010 DVDD.n6009 1.1255
R952 DVDD.n6009 DVDD.n6008 1.1255
R953 DVDD.n5998 DVDD.n5997 1.1255
R954 DVDD.n5997 DVDD.n5996 1.1255
R955 DVDD.n6016 DVDD.n6015 1.1255
R956 DVDD.n6015 DVDD.n6014 1.1255
R957 DVDD.n5907 DVDD.n5900 1.1255
R958 DVDD.n5900 DVDD.n5899 1.1255
R959 DVDD.n5913 DVDD.n5912 1.1255
R960 DVDD.n5912 DVDD.n5911 1.1255
R961 DVDD.n5918 DVDD.n5917 1.1255
R962 DVDD.n5903 DVDD.n5902 1.1255
R963 DVDD.n5902 DVDD.n5901 1.1255
R964 DVDD.n12484 DVDD.n12483 1.1255
R965 DVDD.n12483 DVDD.n12482 1.1255
R966 DVDD.n12661 DVDD.n12660 1.1255
R967 DVDD.n12660 DVDD.n12659 1.1255
R968 DVDD.n12475 DVDD.n12474 1.1255
R969 DVDD.n12474 DVDD.n12473 1.1255
R970 DVDD.n17723 DVDD.n17722 1.1255
R971 DVDD.n17722 DVDD.n17721 1.1255
R972 DVDD.n17717 DVDD.n17716 1.1255
R973 DVDD.n17716 DVDD.n17715 1.1255
R974 DVDD.n5889 DVDD.n5888 1.1255
R975 DVDD.n5888 DVDD.n5887 1.1255
R976 DVDD.n5895 DVDD.n5894 1.1255
R977 DVDD.n5894 DVDD.n5893 1.1255
R978 DVDD.n12667 DVDD.n12666 1.1255
R979 DVDD.n12666 DVDD.n12665 1.1255
R980 DVDD.n17179 DVDD.n17178 1.1255
R981 DVDD.n17178 DVDD.n17177 1.1255
R982 DVDD.n17185 DVDD.n17184 1.1255
R983 DVDD.n17184 DVDD.n17183 1.1255
R984 DVDD.n17817 DVDD.n17816 1.1255
R985 DVDD.n17816 DVDD.n17815 1.1255
R986 DVDD.n17170 DVDD.n17169 1.1255
R987 DVDD.n17169 DVDD.n17168 1.1255
R988 DVDD.n17702 DVDD.n17701 1.1255
R989 DVDD.n17701 DVDD.n17700 1.1255
R990 DVDD.n17708 DVDD.n17707 1.1255
R991 DVDD.n17707 DVDD.n17706 1.1255
R992 DVDD.n17735 DVDD.n17734 1.1255
R993 DVDD.n17734 DVDD.n17733 1.1255
R994 DVDD.n17729 DVDD.n17728 1.1255
R995 DVDD.n17728 DVDD.n17727 1.1255
R996 DVDD.n14014 DVDD.n14013 1.1255
R997 DVDD.n17361 DVDD.n17360 1.1255
R998 DVDD.n14226 DVDD.n14225 1.1255
R999 DVDD.n14225 DVDD.n14224 1.1255
R1000 DVDD.n17522 DVDD.n17521 1.1255
R1001 DVDD.n17521 DVDD.n17520 1.1255
R1002 DVDD.n4109 DVDD.n4108 1.1255
R1003 DVDD.n4108 DVDD.n4107 1.1255
R1004 DVDD.n4461 DVDD.n4460 1.1255
R1005 DVDD.n4460 DVDD.n4459 1.1255
R1006 DVDD.n4100 DVDD.n4099 1.1255
R1007 DVDD.n4099 DVDD.n4098 1.1255
R1008 DVDD.n4467 DVDD.n4466 1.1255
R1009 DVDD.n4466 DVDD.n4465 1.1255
R1010 DVDD.n4358 DVDD.n4357 1.1255
R1011 DVDD.n4357 DVDD.n4356 1.1255
R1012 DVDD.n4376 DVDD.n4375 1.1255
R1013 DVDD.n4375 DVDD.n4374 1.1255
R1014 DVDD.n4370 DVDD.n4369 1.1255
R1015 DVDD.n4369 DVDD.n4368 1.1255
R1016 DVDD.n4364 DVDD.n4363 1.1255
R1017 DVDD.n4363 DVDD.n4362 1.1255
R1018 DVDD.n3447 DVDD.n3446 1.1255
R1019 DVDD.n7790 DVDD.n7789 1.1255
R1020 DVDD.n3580 DVDD.n3579 1.1255
R1021 DVDD.n3669 DVDD.n3668 1.1255
R1022 DVDD.n18644 DVDD.n18643 1.1255
R1023 DVDD.n18741 DVDD.n18740 1.1255
R1024 DVDD.n8735 DVDD.n8734 1.1255
R1025 DVDD.n8734 DVDD.n8733 1.1255
R1026 DVDD.n8744 DVDD.n8743 1.1255
R1027 DVDD.n8743 DVDD.n8742 1.1255
R1028 DVDD.n8732 DVDD.n8731 1.1255
R1029 DVDD.n8731 DVDD.n8730 1.1255
R1030 DVDD.n8753 DVDD.n8752 1.1255
R1031 DVDD.n8752 DVDD.n8751 1.1255
R1032 DVDD.n8632 DVDD.n8631 1.1255
R1033 DVDD.n8631 DVDD.n8630 1.1255
R1034 DVDD.n8650 DVDD.n8649 1.1255
R1035 DVDD.n8649 DVDD.n8648 1.1255
R1036 DVDD.n8644 DVDD.n8643 1.1255
R1037 DVDD.n8643 DVDD.n8642 1.1255
R1038 DVDD.n8638 DVDD.n8637 1.1255
R1039 DVDD.n8637 DVDD.n8636 1.1255
R1040 DVDD.n17405 DVDD.n17404 1.12437
R1041 DVDD.n17238 DVDD.n17237 1.12437
R1042 DVDD.n17587 DVDD.n17585 1.12437
R1043 DVDD.n12958 DVDD.n12957 1.12142
R1044 DVDD.n9039 DVDD.n9038 1.12142
R1045 DVDD.n2736 DVDD.n2713 1.12072
R1046 DVDD.n15388 DVDD.n15387 1.12072
R1047 DVDD.n2777 DVDD.n2501 1.12072
R1048 DVDD.n15518 DVDD.n15517 1.12072
R1049 DVDD.n17736 DVDD.n17735 1.12072
R1050 DVDD.n774 DVDD.n753 1.12072
R1051 DVDD.n18211 DVDD.n10733 1.12072
R1052 DVDD.n811 DVDD.n524 1.12072
R1053 DVDD.n18093 DVDD.n17167 1.12072
R1054 DVDD.n4377 DVDD.n4376 1.12072
R1055 DVDD.n4401 DVDD.n4166 1.12072
R1056 DVDD.n13729 DVDD.n13728 1.12072
R1057 DVDD.n5942 DVDD.n5771 1.12072
R1058 DVDD.n14380 DVDD.n13880 1.12072
R1059 DVDD.n12605 DVDD.n12504 1.12072
R1060 DVDD.n8675 DVDD.n8548 1.12072
R1061 DVDD.n8651 DVDD.n8650 1.12072
R1062 DVDD.n14356 DVDD.n14355 1.12053
R1063 DVDD.n5920 DVDD.n5919 1.12053
R1064 DVDD.n16068 DVDD.n16067 1.12038
R1065 DVDD.n15693 DVDD.n15692 1.12038
R1066 DVDD.n13999 DVDD.n13998 1.10854
R1067 DVDD.n14088 DVDD.n14087 1.10854
R1068 DVDD.n14208 DVDD.n14206 1.10854
R1069 DVDD.n13947 DVDD.n13946 1.08671
R1070 DVDD.n17324 DVDD.n17323 1.08671
R1071 DVDD.n17440 DVDD.n17439 1.08671
R1072 DVDD.n14044 DVDD.n14043 1.08671
R1073 DVDD.n17483 DVDD.n17482 1.08671
R1074 DVDD.n14256 DVDD.n14255 1.08671
R1075 DVDD.n14143 DVDD.n14142 1.08671
R1076 DVDD.n17624 DVDD.n17623 1.08671
R1077 DVDD.t25 DVDD 1.0505
R1078 DVDD DVDD.t6 1.0505
R1079 DVDD DVDD.t37 1.0505
R1080 DVDD DVDD.t31 1.0505
R1081 DVDD.t0 DVDD.n4177 1.0505
R1082 DVDD.n4337 DVDD.n4336 1.0505
R1083 DVDD.n14013 DVDD.n14012 0.981907
R1084 DVDD.n14100 DVDD.n14099 0.981907
R1085 DVDD.n14225 DVDD.n14223 0.981907
R1086 DVDD.n17360 DVDD.n17359 0.966078
R1087 DVDD.n17190 DVDD.n17189 0.966078
R1088 DVDD.n17521 DVDD.n17519 0.966078
R1089 DVDD.n17361 DVDD.n17356 0.879031
R1090 DVDD.n17522 DVDD.n17516 0.879031
R1091 DVDD.n14014 DVDD.n14009 0.875231
R1092 DVDD.n14226 DVDD.n14220 0.875231
R1093 DVDD.n15993 DVDD.n15992 0.858403
R1094 DVDD.n5529 DVDD.n5528 0.788
R1095 DVDD.n5528 DVDD.n5527 0.788
R1096 DVDD.n4078 DVDD.n4077 0.788
R1097 DVDD.n4077 DVDD.n4076 0.788
R1098 DVDD.n4208 DVDD.n4207 0.788
R1099 DVDD.n4196 DVDD.n4195 0.788
R1100 DVDD.n4179 DVDD.n4178 0.788
R1101 DVDD.n4178 DVDD.t0 0.788
R1102 DVDD.n17194 DVDD.n17193 0.766594
R1103 DVDD.n14104 DVDD.n14103 0.762133
R1104 DVDD.n9392 DVDD.n9391 0.75203
R1105 DVDD.n13303 DVDD.n13302 0.75203
R1106 DVDD.n9887 DVDD.n9886 0.75167
R1107 DVDD.n11988 DVDD.n11987 0.75167
R1108 DVDD.n9485 DVDD.n9484 0.75158
R1109 DVDD.n12290 DVDD.n12289 0.75158
R1110 DVDD.n11514 DVDD.n11513 0.7505
R1111 DVDD.n18267 DVDD.n18266 0.7505
R1112 DVDD.n19416 DVDD.n19415 0.7505
R1113 DVDD.n1670 DVDD.n1669 0.7505
R1114 DVDD.n1550 DVDD.n1549 0.7505
R1115 DVDD.n1782 DVDD.n1781 0.7505
R1116 DVDD.n19106 DVDD.n19105 0.7505
R1117 DVDD.n17462 DVDD.n17258 0.7505
R1118 DVDD.n13936 DVDD.n13935 0.7505
R1119 DVDD.n13941 DVDD.n13940 0.7505
R1120 DVDD.n13948 DVDD.n13947 0.7505
R1121 DVDD.n13952 DVDD.n13951 0.7505
R1122 DVDD.n13957 DVDD.n13956 0.7505
R1123 DVDD.n13926 DVDD.n13925 0.7505
R1124 DVDD.n13931 DVDD.n13930 0.7505
R1125 DVDD.n17419 DVDD.n17418 0.7505
R1126 DVDD.n17424 DVDD.n17423 0.7505
R1127 DVDD.n17429 DVDD.n17428 0.7505
R1128 DVDD.n17434 DVDD.n17433 0.7505
R1129 DVDD.n17441 DVDD.n17440 0.7505
R1130 DVDD.n17445 DVDD.n17444 0.7505
R1131 DVDD.n17450 DVDD.n17449 0.7505
R1132 DVDD.n17303 DVDD.n17302 0.7505
R1133 DVDD.n17308 DVDD.n17307 0.7505
R1134 DVDD.n17313 DVDD.n17312 0.7505
R1135 DVDD.n17318 DVDD.n17317 0.7505
R1136 DVDD.n17325 DVDD.n17324 0.7505
R1137 DVDD.n17329 DVDD.n17328 0.7505
R1138 DVDD.n17334 DVDD.n17333 0.7505
R1139 DVDD.n14054 DVDD.n14053 0.7505
R1140 DVDD.n14049 DVDD.n14048 0.7505
R1141 DVDD.n14045 DVDD.n14044 0.7505
R1142 DVDD.n14038 DVDD.n14037 0.7505
R1143 DVDD.n14033 DVDD.n14032 0.7505
R1144 DVDD.n14028 DVDD.n14027 0.7505
R1145 DVDD.n14023 DVDD.n14022 0.7505
R1146 DVDD.n17467 DVDD.n17466 0.7505
R1147 DVDD.n17472 DVDD.n17471 0.7505
R1148 DVDD.n17477 DVDD.n17476 0.7505
R1149 DVDD.n17484 DVDD.n17483 0.7505
R1150 DVDD.n17488 DVDD.n17487 0.7505
R1151 DVDD.n17493 DVDD.n17492 0.7505
R1152 DVDD.n14239 DVDD.n14238 0.7505
R1153 DVDD.n14244 DVDD.n14243 0.7505
R1154 DVDD.n14249 DVDD.n14248 0.7505
R1155 DVDD.n14257 DVDD.n14256 0.7505
R1156 DVDD.n14261 DVDD.n14260 0.7505
R1157 DVDD.n14266 DVDD.n14265 0.7505
R1158 DVDD.n14271 DVDD.n14270 0.7505
R1159 DVDD.n14316 DVDD.n14315 0.7505
R1160 DVDD.n14234 DVDD.n14233 0.7505
R1161 DVDD.n14153 DVDD.n14152 0.7505
R1162 DVDD.n14148 DVDD.n14147 0.7505
R1163 DVDD.n14144 DVDD.n14143 0.7505
R1164 DVDD.n14136 DVDD.n14135 0.7505
R1165 DVDD.n14131 DVDD.n14130 0.7505
R1166 DVDD.n14126 DVDD.n14125 0.7505
R1167 DVDD.n14121 DVDD.n14120 0.7505
R1168 DVDD.n17606 DVDD.n17605 0.7505
R1169 DVDD.n17611 DVDD.n17610 0.7505
R1170 DVDD.n17616 DVDD.n17615 0.7505
R1171 DVDD.n17625 DVDD.n17624 0.7505
R1172 DVDD.n17629 DVDD.n17628 0.7505
R1173 DVDD.n17634 DVDD.n17633 0.7505
R1174 DVDD.n17639 DVDD.n17638 0.7505
R1175 DVDD.n17684 DVDD.n17683 0.7505
R1176 DVDD.n17601 DVDD.n17600 0.7505
R1177 DVDD.n18858 DVDD.n18857 0.7505
R1178 DVDD.n9930 DVDD.n9929 0.7505
R1179 DVDD.n3325 DVDD.n3324 0.7505
R1180 DVDD.n18357 DVDD.n18356 0.7505
R1181 DVDD.n7134 DVDD.n7133 0.7505
R1182 DVDD.n7691 DVDD.n7690 0.7505
R1183 DVDD.n18668 DVDD.n18667 0.7505
R1184 DVDD.n18586 DVDD.n18585 0.7505
R1185 DVDD.n18601 DVDD.n18600 0.7505
R1186 DVDD.n18616 DVDD.n18615 0.7505
R1187 DVDD.n18632 DVDD.n18631 0.7505
R1188 DVDD.n18649 DVDD.n18648 0.7505
R1189 DVDD.n18736 DVDD.n18735 0.7505
R1190 DVDD.n18725 DVDD.n18724 0.7505
R1191 DVDD.n18710 DVDD.n18709 0.7505
R1192 DVDD.n18696 DVDD.n18695 0.7505
R1193 DVDD.n18467 DVDD.n18466 0.7505
R1194 DVDD.n18395 DVDD.n18394 0.7505
R1195 DVDD.n12919 DVDD.n12916 0.662783
R1196 DVDD.n12916 DVDD.n12915 0.662783
R1197 DVDD.n9026 DVDD.n9023 0.662538
R1198 DVDD.n9023 DVDD.n9022 0.662538
R1199 DVDD.n17173 DVDD.n17172 0.643962
R1200 DVDD.n11204 DVDD.n11203 0.643769
R1201 DVDD.n4610 DVDD.n4609 0.643357
R1202 DVDD.n18333 DVDD.n3888 0.643357
R1203 DVDD.n20215 DVDD.n20079 0.643357
R1204 DVDD.n20211 DVDD.n20210 0.643357
R1205 DVDD.n20117 DVDD.n20116 0.643357
R1206 DVDD.n19464 DVDD.n19081 0.643357
R1207 DVDD.n18333 DVDD.n18332 0.643357
R1208 DVDD.n20215 DVDD.n293 0.643357
R1209 DVDD.n19464 DVDD.n19463 0.643357
R1210 DVDD.n18333 DVDD.n7109 0.643357
R1211 DVDD.n7074 DVDD.n7073 0.643357
R1212 DVDD.n20215 DVDD.n2300 0.643357
R1213 DVDD.n19596 DVDD.n19595 0.643357
R1214 DVDD.n19502 DVDD.n19501 0.643357
R1215 DVDD.n19464 DVDD.n18973 0.643357
R1216 DVDD.n19464 DVDD.n18810 0.643357
R1217 DVDD.n20215 DVDD.n3779 0.643357
R1218 DVDD.n18333 DVDD.n10054 0.643357
R1219 DVDD.n14790 DVDD.n14771 0.643357
R1220 DVDD.n18449 DVDD.n18448 0.643357
R1221 DVDD.n13924 DVDD.n13923 0.637389
R1222 DVDD.n17417 DVDD.n17416 0.637389
R1223 DVDD.n4103 DVDD.n4102 0.6305
R1224 DVDD.n4102 DVDD.n4101 0.6305
R1225 DVDD.n4355 DVDD.n4354 0.6305
R1226 DVDD.n4354 DVDD.n4353 0.6305
R1227 DVDD.n3157 DVDD.n3156 0.628944
R1228 DVDD.n13945 DVDD.n13944 0.628675
R1229 DVDD.n13946 DVDD.n13945 0.628675
R1230 DVDD.n17437 DVDD.n17436 0.628675
R1231 DVDD.n17439 DVDD.n17437 0.628675
R1232 DVDD.n17322 DVDD.n17321 0.628675
R1233 DVDD.n17323 DVDD.n17322 0.628675
R1234 DVDD.n14042 DVDD.n14041 0.628675
R1235 DVDD.n14043 DVDD.n14042 0.628675
R1236 DVDD.n17480 DVDD.n17479 0.628675
R1237 DVDD.n17482 DVDD.n17480 0.628675
R1238 DVDD.n14141 DVDD.n14139 0.628675
R1239 DVDD.n14142 DVDD.n14141 0.628675
R1240 DVDD.n1241 DVDD.n1123 0.626961
R1241 DVDD.n2024 DVDD 0.608566
R1242 DVDD.n2156 DVDD 0.608566
R1243 DVDD.n2232 DVDD 0.608566
R1244 DVDD.n6938 DVDD 0.608566
R1245 DVDD.n6786 DVDD 0.608566
R1246 DVDD.n6520 DVDD 0.608566
R1247 DVDD.n1859 DVDD 0.608566
R1248 DVDD.n3925 DVDD 0.608566
R1249 DVDD.n19802 DVDD 0.608566
R1250 DVDD.n19935 DVDD 0.608566
R1251 DVDD.n20011 DVDD 0.608566
R1252 DVDD.n4712 DVDD 0.608566
R1253 DVDD.n4823 DVDD 0.608566
R1254 DVDD.n5111 DVDD 0.608566
R1255 DVDD.n19637 DVDD 0.608566
R1256 DVDD.n5230 DVDD 0.608566
R1257 DVDD.n2055 DVDD 0.608476
R1258 DVDD.n2209 DVDD 0.608476
R1259 DVDD.n18931 DVDD 0.608476
R1260 DVDD.n7033 DVDD 0.608476
R1261 DVDD.n6943 DVDD 0.608476
R1262 DVDD.n6802 DVDD 0.608476
R1263 DVDD.n6553 DVDD 0.608476
R1264 DVDD.n1862 DVDD 0.608476
R1265 DVDD.n3930 DVDD 0.608476
R1266 DVDD.n19833 DVDD 0.608476
R1267 DVDD.n19988 DVDD 0.608476
R1268 DVDD.n19049 DVDD 0.608476
R1269 DVDD.n4613 DVDD 0.608476
R1270 DVDD.n4717 DVDD 0.608476
R1271 DVDD.n4839 DVDD 0.608476
R1272 DVDD.n5144 DVDD 0.608476
R1273 DVDD.n19640 DVDD 0.608476
R1274 DVDD.n5235 DVDD 0.608476
R1275 DVDD DVDD.n7097 0.608386
R1276 DVDD DVDD.n3876 0.608386
R1277 DVDD DVDD.n7765 0.606676
R1278 DVDD DVDD.n18775 0.606676
R1279 DVDD.n9886 DVDD 0.606676
R1280 DVDD.n9485 DVDD 0.606676
R1281 DVDD.n9391 DVDD 0.606676
R1282 DVDD.n9314 DVDD 0.606676
R1283 DVDD DVDD.n19428 0.606676
R1284 DVDD DVDD.n18277 0.606676
R1285 DVDD.n11987 DVDD 0.606676
R1286 DVDD.n12290 DVDD 0.606676
R1287 DVDD.n13225 DVDD 0.606676
R1288 DVDD.n13302 DVDD 0.606676
R1289 DVDD.n17293 DVDD.n17292 0.594352
R1290 DVDD.n13910 DVDD.n13909 0.594352
R1291 DVDD.n17672 DVDD.n17671 0.594352
R1292 DVDD.n14299 DVDD.n14298 0.594352
R1293 DVDD.n7163 DVDD.n7162 0.578545
R1294 DVDD.n1013 DVDD.n1012 0.578545
R1295 DVDD.n1734 DVDD.n1733 0.578545
R1296 DVDD.n1089 DVDD.n1087 0.578544
R1297 DVDD.n11424 DVDD.n11423 0.578544
R1298 DVDD.n9816 DVDD.n9815 0.57846
R1299 DVDD.n9958 DVDD.n9956 0.57846
R1300 DVDD.n1546 DVDD.n1545 0.57846
R1301 DVDD.n1674 DVDD.n1673 0.57846
R1302 DVDD.n11541 DVDD.n11540 0.57846
R1303 DVDD.n3321 DVDD.n3320 0.57846
R1304 DVDD.n11917 DVDD.n11916 0.57846
R1305 DVDD.n1283 DVDD.n1282 0.57846
R1306 DVDD.n12323 DVDD.n12322 0.57846
R1307 DVDD.n18287 DVDD.n10125 0.578459
R1308 DVDD.n9519 DVDD.n9517 0.578459
R1309 DVDD.n3674 DVDD.n3672 0.577423
R1310 DVDD.n2916 DVDD.n2914 0.577423
R1311 DVDD.n3002 DVDD.n3001 0.577423
R1312 DVDD.n3576 DVDD.n3575 0.577338
R1313 DVDD.n3452 DVDD.n3450 0.577338
R1314 DVDD.n7769 DVDD.n7768 0.577338
R1315 DVDD.n7817 DVDD.n7816 0.563519
R1316 DVDD.n7936 DVDD.n7934 0.563519
R1317 DVDD.n8363 DVDD.n8362 0.563519
R1318 DVDD.n9313 DVDD.n9311 0.56343
R1319 DVDD.n11342 DVDD.n11341 0.563421
R1320 DVDD.n11338 DVDD.n11336 0.563421
R1321 DVDD.n11301 DVDD.n11300 0.563421
R1322 DVDD.n19431 DVDD.n19430 0.563333
R1323 DVDD.n13224 DVDD.n13222 0.563333
R1324 DVDD.n18266 DVDD.n18265 0.563
R1325 DVDD.n19415 DVDD.n19414 0.563
R1326 DVDD.n18333 DVDD.n10102 0.563
R1327 DVDD.n18238 DVDD.n18237 0.563
R1328 DVDD.n249 DVDD.n248 0.563
R1329 DVDD.n20215 DVDD.n843 0.563
R1330 DVDD.n161 DVDD.n160 0.563
R1331 DVDD.n19464 DVDD.n19180 0.563
R1332 DVDD.n18333 DVDD.n10070 0.563
R1333 DVDD.n14800 DVDD.n14799 0.563
R1334 DVDD.n18682 DVDD.n18681 0.563
R1335 DVDD.n18580 DVDD.n18579 0.563
R1336 DVDD.n20215 DVDD.n2811 0.563
R1337 DVDD.n19464 DVDD.n18484 0.563
R1338 DVDD.n3651 DVDD.n3650 0.563
R1339 DVDD.n18778 DVDD.n18777 0.561353
R1340 DVDD.n1783 DVDD.n1782 0.5005
R1341 DVDD DVDD.n6111 0.5
R1342 DVDD DVDD.n6116 0.5
R1343 DVDD.n4565 DVDD 0.5
R1344 DVDD DVDD.n4564 0.5
R1345 DVDD.n4580 DVDD 0.5
R1346 DVDD DVDD.n4579 0.5
R1347 DVDD.n4595 DVDD 0.5
R1348 DVDD DVDD.n4594 0.5
R1349 DVDD.n5813 DVDD.n5812 0.455365
R1350 DVDD.n4345 DVDD.n4337 0.455365
R1351 DVDD.n3274 DVDD.n3158 0.446103
R1352 DVDD.n1328 DVDD.n1120 0.44482
R1353 DVDD.n14012 DVDD.n14010 0.439434
R1354 DVDD.n13922 DVDD.n13921 0.439434
R1355 DVDD.n17189 DVDD.n17187 0.439434
R1356 DVDD.n17359 DVDD.n17357 0.439434
R1357 DVDD.n17359 DVDD.n17358 0.439434
R1358 DVDD.n17300 DVDD.n17299 0.439434
R1359 DVDD.n14223 DVDD.n14221 0.439434
R1360 DVDD.n14099 DVDD.n14097 0.439434
R1361 DVDD.n14099 DVDD.n14098 0.439434
R1362 DVDD.n14012 DVDD.n14011 0.439434
R1363 DVDD.n17679 DVDD.n17678 0.439434
R1364 DVDD.n17519 DVDD.n17517 0.439434
R1365 DVDD.n17519 DVDD.n17518 0.439434
R1366 DVDD.n17189 DVDD.n17188 0.439434
R1367 DVDD.n14312 DVDD.n14311 0.439434
R1368 DVDD.n14223 DVDD.n14222 0.439434
R1369 DVDD.n5701 DVDD.n5700 0.4091
R1370 DVDD.n8484 DVDD.n8483 0.4091
R1371 DVDD.n12453 DVDD.n12452 0.4091
R1372 DVDD.n4061 DVDD.n4060 0.4091
R1373 DVDD.n12440 DVDD.n12439 0.4091
R1374 DVDD.n4051 DVDD.n4050 0.4091
R1375 DVDD.n12421 DVDD.n12420 0.4091
R1376 DVDD.n4041 DVDD.n4040 0.4091
R1377 DVDD.n7160 DVDD.n7159 0.404524
R1378 DVDD.n9960 DVDD.n9959 0.404438
R1379 DVDD.n9813 DVDD.n9812 0.404438
R1380 DVDD.n9521 DVDD.n9520 0.404438
R1381 DVDD.n3318 DVDD.n3317 0.404438
R1382 DVDD.n1091 DVDD.n1090 0.403241
R1383 DVDD.n1010 DVDD.n1009 0.403241
R1384 DVDD.n1731 DVDD.n1730 0.403241
R1385 DVDD.n11421 DVDD.n11420 0.403241
R1386 DVDD.n1543 DVDD.n1542 0.403154
R1387 DVDD.n1676 DVDD.n1675 0.403154
R1388 DVDD.n11543 DVDD.n11542 0.403154
R1389 DVDD.n18289 DVDD.n18288 0.403154
R1390 DVDD.n11914 DVDD.n11913 0.403154
R1391 DVDD.n1285 DVDD.n1284 0.403154
R1392 DVDD.n12325 DVDD.n12324 0.403154
R1393 DVDD.n14358 DVDD.n14357 0.396996
R1394 DVDD.n5922 DVDD.n5921 0.396996
R1395 DVDD.n12585 DVDD.n12584 0.396996
R1396 DVDD.n17738 DVDD.n17737 0.396996
R1397 DVDD.n4379 DVDD.n4378 0.396996
R1398 DVDD.n8653 DVDD.n8652 0.396996
R1399 DVDD.n15278 DVDD.n15274 0.382213
R1400 DVDD.n18282 DVDD.n18280 0.378092
R1401 DVDD.n3443 DVDD.n3442 0.37805
R1402 DVDD.n3584 DVDD.n3583 0.37805
R1403 DVDD.n15278 DVDD.n15277 0.3755
R1404 DVDD.n15282 DVDD.n15281 0.3755
R1405 DVDD.n15286 DVDD.n15285 0.3755
R1406 DVDD.n15135 DVDD.n15130 0.3755
R1407 DVDD.n15288 DVDD.n15287 0.3755
R1408 DVDD.n3676 DVDD.n3675 0.375019
R1409 DVDD.n2999 DVDD.n2998 0.375019
R1410 DVDD.n2918 DVDD.n2917 0.375019
R1411 DVDD.n7736 DVDD.n7735 0.374932
R1412 DVDD.n3454 DVDD.n3453 0.374932
R1413 DVDD.n3573 DVDD.n3572 0.374932
R1414 DVDD.n17622 DVDD.n17621 0.37479
R1415 DVDD.n17270 DVDD.n17269 0.373473
R1416 DVDD.n13887 DVDD.n13885 0.373473
R1417 DVDD.n17648 DVDD.n17647 0.373473
R1418 DVDD.n14275 DVDD.n14273 0.373473
R1419 DVDD.n3329 DVDD.n3328 0.372367
R1420 DVDD.n7811 DVDD.n7810 0.37102
R1421 DVDD.n17410 DVDD.n17409 0.36457
R1422 DVDD.n14004 DVDD.n14003 0.36457
R1423 DVDD.n17243 DVDD.n17242 0.36457
R1424 DVDD.n14093 DVDD.n14092 0.36457
R1425 DVDD.n17593 DVDD.n17592 0.36457
R1426 DVDD.n14214 DVDD.n14212 0.36457
R1427 DVDD.n7742 DVDD.n7740 0.348975
R1428 DVDD.n13692 DVDD.n13691 0.345264
R1429 DVDD.n14399 DVDD.n14398 0.345264
R1430 DVDD.n5959 DVDD.n5958 0.345264
R1431 DVDD.n12622 DVDD.n12621 0.345264
R1432 DVDD.n17775 DVDD.n17774 0.345264
R1433 DVDD.n4420 DVDD.n4419 0.345264
R1434 DVDD.n8694 DVDD.n8693 0.345264
R1435 DVDD.n2796 DVDD.n2795 0.344378
R1436 DVDD.n828 DVDD.n827 0.344378
R1437 DVDD.n15504 DVDD.n15503 0.340657
R1438 DVDD.n18107 DVDD.n18106 0.340657
R1439 DVDD.n15274 DVDD.n15273 0.323092
R1440 DVDD.n19684 DVDD.n19683 0.308636
R1441 DVDD.n1329 DVDD.n1328 0.308636
R1442 DVDD.n1906 DVDD.n1905 0.308636
R1443 DVDD.n3274 DVDD.n3273 0.308636
R1444 DVDD.n5530 DVDD.n5529 0.271967
R1445 DVDD.n4079 DVDD.n4078 0.271967
R1446 DVDD.n4198 DVDD.n4196 0.269064
R1447 DVDD.n4210 DVDD.n4208 0.269064
R1448 DVDD.n4182 DVDD.n4179 0.269064
R1449 DVDD.n17622 DVDD.n17620 0.267993
R1450 DVDD.n13905 DVDD.n13903 0.264014
R1451 DVDD.n14293 DVDD.n14291 0.264014
R1452 DVDD.n17288 DVDD.n17286 0.263608
R1453 DVDD.n17666 DVDD.n17664 0.263608
R1454 DVDD.n17192 DVDD.n17190 0.253766
R1455 DVDD.n17291 DVDD.n17290 0.249014
R1456 DVDD.n13908 DVDD.n13907 0.249014
R1457 DVDD.n17670 DVDD.n17669 0.249014
R1458 DVDD.n14297 DVDD.n14296 0.249014
R1459 DVDD.n14102 DVDD.n14100 0.237937
R1460 DVDD.n13915 DVDD.n13914 0.23535
R1461 DVDD.n17263 DVDD.n17262 0.23535
R1462 DVDD.n14304 DVDD.n14303 0.23535
R1463 DVDD.n17641 DVDD.n17640 0.23535
R1464 DVDD.n3675 DVDD 0.234468
R1465 DVDD DVDD.n2999 0.234468
R1466 DVDD.n2917 DVDD 0.234468
R1467 DVDD DVDD.n7736 0.234465
R1468 DVDD.n3453 DVDD 0.234465
R1469 DVDD DVDD.n3573 0.234465
R1470 DVDD.n2487 DVDD.n2486 0.2255
R1471 DVDD.n2484 DVDD.n2483 0.2255
R1472 DVDD.n2482 DVDD.n2481 0.2255
R1473 DVDD.n2475 DVDD.n2474 0.2255
R1474 DVDD.n2467 DVDD.n2466 0.2255
R1475 DVDD.n2464 DVDD.n2463 0.2255
R1476 DVDD.n2462 DVDD.n2461 0.2255
R1477 DVDD.n2460 DVDD.n2459 0.2255
R1478 DVDD.n2458 DVDD.n2457 0.2255
R1479 DVDD.n2497 DVDD.n2496 0.2255
R1480 DVDD.n2498 DVDD.n2497 0.2255
R1481 DVDD.n2449 DVDD.n2447 0.2255
R1482 DVDD.n2450 DVDD.n2449 0.2255
R1483 DVDD.n2425 DVDD.n2424 0.2255
R1484 DVDD.n2419 DVDD.n2418 0.2255
R1485 DVDD.n2415 DVDD.n2414 0.2255
R1486 DVDD.n2413 DVDD.n2412 0.2255
R1487 DVDD.n2411 DVDD.n2410 0.2255
R1488 DVDD.n2409 DVDD.n2408 0.2255
R1489 DVDD.n2407 DVDD.n2406 0.2255
R1490 DVDD.n2405 DVDD.n2404 0.2255
R1491 DVDD.n2403 DVDD.n2402 0.2255
R1492 DVDD.n2393 DVDD.n2392 0.2255
R1493 DVDD.n2385 DVDD.n2384 0.2255
R1494 DVDD.n2378 DVDD.n2377 0.2255
R1495 DVDD.n2372 DVDD.n2371 0.2255
R1496 DVDD.n2370 DVDD.n2369 0.2255
R1497 DVDD.n2368 DVDD.n2367 0.2255
R1498 DVDD.n2366 DVDD.n2365 0.2255
R1499 DVDD.n2364 DVDD.n2363 0.2255
R1500 DVDD.n2362 DVDD.n2361 0.2255
R1501 DVDD.n2360 DVDD.n2359 0.2255
R1502 DVDD.n2358 DVDD.n2357 0.2255
R1503 DVDD.n2356 DVDD.n2355 0.2255
R1504 DVDD.n2354 DVDD.n2353 0.2255
R1505 DVDD.n2352 DVDD.n2351 0.2255
R1506 DVDD.n2350 DVDD.n2349 0.2255
R1507 DVDD.n2348 DVDD.n2347 0.2255
R1508 DVDD.n2342 DVDD.n2341 0.2255
R1509 DVDD.n2334 DVDD.n2333 0.2255
R1510 DVDD.n2327 DVDD.n2326 0.2255
R1511 DVDD.n2317 DVDD.n2316 0.2255
R1512 DVDD.n2315 DVDD.n2314 0.2255
R1513 DVDD.n2313 DVDD.n2312 0.2255
R1514 DVDD.n2311 DVDD.n2310 0.2255
R1515 DVDD.n2309 DVDD.n2308 0.2255
R1516 DVDD.n2307 DVDD.n2306 0.2255
R1517 DVDD.n2305 DVDD.n2304 0.2255
R1518 DVDD.n2303 DVDD.n2302 0.2255
R1519 DVDD.n416 DVDD.n415 0.2255
R1520 DVDD.n418 DVDD.n417 0.2255
R1521 DVDD.n420 DVDD.n419 0.2255
R1522 DVDD.n422 DVDD.n421 0.2255
R1523 DVDD.n424 DVDD.n423 0.2255
R1524 DVDD.n426 DVDD.n425 0.2255
R1525 DVDD.n428 DVDD.n427 0.2255
R1526 DVDD.n430 DVDD.n429 0.2255
R1527 DVDD.n398 DVDD.n397 0.2255
R1528 DVDD.n405 DVDD.n404 0.2255
R1529 DVDD.n413 DVDD.n412 0.2255
R1530 DVDD.n523 DVDD.n522 0.2255
R1531 DVDD.n520 DVDD.n519 0.2255
R1532 DVDD.n518 DVDD.n517 0.2255
R1533 DVDD.n516 DVDD.n515 0.2255
R1534 DVDD.n514 DVDD.n513 0.2255
R1535 DVDD.n512 DVDD.n511 0.2255
R1536 DVDD.n510 DVDD.n509 0.2255
R1537 DVDD.n508 DVDD.n507 0.2255
R1538 DVDD.n506 DVDD.n505 0.2255
R1539 DVDD.n504 DVDD.n503 0.2255
R1540 DVDD.n495 DVDD.n494 0.2255
R1541 DVDD.n486 DVDD.n485 0.2255
R1542 DVDD.n481 DVDD.n480 0.2255
R1543 DVDD.n478 DVDD.n477 0.2255
R1544 DVDD.n476 DVDD.n475 0.2255
R1545 DVDD.n474 DVDD.n473 0.2255
R1546 DVDD.n470 DVDD.n469 0.2255
R1547 DVDD.n468 DVDD.n467 0.2255
R1548 DVDD.n466 DVDD.n465 0.2255
R1549 DVDD.n464 DVDD.n463 0.2255
R1550 DVDD.n462 DVDD.n461 0.2255
R1551 DVDD.n460 DVDD.n459 0.2255
R1552 DVDD.n458 DVDD.n457 0.2255
R1553 DVDD.n456 DVDD.n455 0.2255
R1554 DVDD.n454 DVDD.n453 0.2255
R1555 DVDD.n449 DVDD.n448 0.2255
R1556 DVDD.n440 DVDD.n439 0.2255
R1557 DVDD.n435 DVDD.n434 0.2255
R1558 DVDD.n752 DVDD.n646 0.2255
R1559 DVDD.n2689 DVDD.n2651 0.2255
R1560 DVDD.n2699 DVDD.n2698 0.2255
R1561 DVDD.n2696 DVDD.n2695 0.2255
R1562 DVDD.n629 DVDD.n628 0.2255
R1563 DVDD.n636 DVDD.n635 0.2255
R1564 DVDD.n644 DVDD.n643 0.2255
R1565 DVDD.n750 DVDD.n749 0.2255
R1566 DVDD.n748 DVDD.n747 0.2255
R1567 DVDD.n746 DVDD.n745 0.2255
R1568 DVDD.n744 DVDD.n743 0.2255
R1569 DVDD.n742 DVDD.n741 0.2255
R1570 DVDD.n740 DVDD.n739 0.2255
R1571 DVDD.n738 DVDD.n737 0.2255
R1572 DVDD.n736 DVDD.n735 0.2255
R1573 DVDD.n734 DVDD.n733 0.2255
R1574 DVDD.n727 DVDD.n726 0.2255
R1575 DVDD.n718 DVDD.n717 0.2255
R1576 DVDD.n713 DVDD.n712 0.2255
R1577 DVDD.n710 DVDD.n709 0.2255
R1578 DVDD.n708 DVDD.n707 0.2255
R1579 DVDD.n706 DVDD.n705 0.2255
R1580 DVDD.n704 DVDD.n703 0.2255
R1581 DVDD.n702 DVDD.n701 0.2255
R1582 DVDD.n700 DVDD.n699 0.2255
R1583 DVDD.n696 DVDD.n695 0.2255
R1584 DVDD.n694 DVDD.n693 0.2255
R1585 DVDD.n692 DVDD.n691 0.2255
R1586 DVDD.n690 DVDD.n689 0.2255
R1587 DVDD.n688 DVDD.n687 0.2255
R1588 DVDD.n686 DVDD.n685 0.2255
R1589 DVDD.n681 DVDD.n680 0.2255
R1590 DVDD.n672 DVDD.n671 0.2255
R1591 DVDD.n667 DVDD.n666 0.2255
R1592 DVDD.n662 DVDD.n661 0.2255
R1593 DVDD.n658 DVDD.n657 0.2255
R1594 DVDD.n656 DVDD.n655 0.2255
R1595 DVDD.n654 DVDD.n653 0.2255
R1596 DVDD.n652 DVDD.n651 0.2255
R1597 DVDD.n650 DVDD.n649 0.2255
R1598 DVDD.n648 DVDD.n647 0.2255
R1599 DVDD.n2503 DVDD.n2502 0.2255
R1600 DVDD.n2505 DVDD.n2504 0.2255
R1601 DVDD.n2507 DVDD.n2506 0.2255
R1602 DVDD.n2511 DVDD.n2510 0.2255
R1603 DVDD.n2513 DVDD.n2512 0.2255
R1604 DVDD.n2515 DVDD.n2514 0.2255
R1605 DVDD.n2517 DVDD.n2516 0.2255
R1606 DVDD.n2525 DVDD.n2524 0.2255
R1607 DVDD.n2532 DVDD.n2531 0.2255
R1608 DVDD.n2540 DVDD.n2539 0.2255
R1609 DVDD.n2546 DVDD.n2545 0.2255
R1610 DVDD.n2548 DVDD.n2547 0.2255
R1611 DVDD.n2550 DVDD.n2549 0.2255
R1612 DVDD.n2552 DVDD.n2551 0.2255
R1613 DVDD.n2554 DVDD.n2553 0.2255
R1614 DVDD.n2556 DVDD.n2555 0.2255
R1615 DVDD.n2558 DVDD.n2557 0.2255
R1616 DVDD.n2560 DVDD.n2559 0.2255
R1617 DVDD.n2564 DVDD.n2563 0.2255
R1618 DVDD.n2566 DVDD.n2565 0.2255
R1619 DVDD.n2568 DVDD.n2567 0.2255
R1620 DVDD.n2570 DVDD.n2569 0.2255
R1621 DVDD.n2576 DVDD.n2575 0.2255
R1622 DVDD.n2583 DVDD.n2582 0.2255
R1623 DVDD.n2591 DVDD.n2590 0.2255
R1624 DVDD.n2599 DVDD.n2598 0.2255
R1625 DVDD.n2601 DVDD.n2600 0.2255
R1626 DVDD.n2603 DVDD.n2602 0.2255
R1627 DVDD.n2605 DVDD.n2604 0.2255
R1628 DVDD.n2607 DVDD.n2606 0.2255
R1629 DVDD.n2609 DVDD.n2608 0.2255
R1630 DVDD.n2611 DVDD.n2610 0.2255
R1631 DVDD.n2613 DVDD.n2612 0.2255
R1632 DVDD.n2615 DVDD.n2614 0.2255
R1633 DVDD.n2621 DVDD.n2620 0.2255
R1634 DVDD.n2645 DVDD.n2644 0.2255
R1635 DVDD.n2646 DVDD.n2645 0.2255
R1636 DVDD.n2709 DVDD.n2708 0.2255
R1637 DVDD.n2710 DVDD.n2709 0.2255
R1638 DVDD.n2656 DVDD.n2655 0.2255
R1639 DVDD.n2658 DVDD.n2657 0.2255
R1640 DVDD.n2660 DVDD.n2659 0.2255
R1641 DVDD.n2662 DVDD.n2661 0.2255
R1642 DVDD.n2665 DVDD.n2664 0.2255
R1643 DVDD.n2673 DVDD.n2672 0.2255
R1644 DVDD.n2682 DVDD.n2681 0.2255
R1645 DVDD.n13832 DVDD.n13831 0.2255
R1646 DVDD.n13835 DVDD.n13834 0.2255
R1647 DVDD.n5727 DVDD.n5726 0.2255
R1648 DVDD.n5731 DVDD.n5730 0.2255
R1649 DVDD.n5733 DVDD.n5732 0.2255
R1650 DVDD.n5737 DVDD.n5736 0.2255
R1651 DVDD.n5744 DVDD.n5743 0.2255
R1652 DVDD.n5769 DVDD.n5768 0.2255
R1653 DVDD.n5763 DVDD.n5762 0.2255
R1654 DVDD.n5760 DVDD.n5759 0.2255
R1655 DVDD.n5758 DVDD.n5757 0.2255
R1656 DVDD.n5756 DVDD.n5755 0.2255
R1657 DVDD.n5752 DVDD.n5751 0.2255
R1658 DVDD.n4115 DVDD.n4114 0.2255
R1659 DVDD.n4119 DVDD.n4118 0.2255
R1660 DVDD.n4123 DVDD.n4122 0.2255
R1661 DVDD.n4127 DVDD.n4126 0.2255
R1662 DVDD.n4134 DVDD.n4133 0.2255
R1663 DVDD.n4164 DVDD.n4163 0.2255
R1664 DVDD.n4156 DVDD.n4155 0.2255
R1665 DVDD.n4143 DVDD.n4142 0.2255
R1666 DVDD.n4139 DVDD.n4138 0.2255
R1667 DVDD.n8499 DVDD.n8498 0.2255
R1668 DVDD.n8503 DVDD.n8502 0.2255
R1669 DVDD.n8509 DVDD.n8508 0.2255
R1670 DVDD.n8516 DVDD.n8515 0.2255
R1671 DVDD.n8546 DVDD.n8545 0.2255
R1672 DVDD.n8538 DVDD.n8537 0.2255
R1673 DVDD.n8527 DVDD.n8526 0.2255
R1674 DVDD.n8525 DVDD.n8524 0.2255
R1675 DVDD.n8523 DVDD.n8522 0.2255
R1676 DVDD.n8519 DVDD.n8518 0.2255
R1677 DVDD.n11209 DVDD.n11208 0.2255
R1678 DVDD.n11211 DVDD.n11210 0.2255
R1679 DVDD.n11218 DVDD.n11217 0.2255
R1680 DVDD.n13878 DVDD.n13877 0.2255
R1681 DVDD.n13870 DVDD.n13869 0.2255
R1682 DVDD.n13859 DVDD.n13858 0.2255
R1683 DVDD.n13857 DVDD.n13856 0.2255
R1684 DVDD.n13855 DVDD.n13854 0.2255
R1685 DVDD.n13849 DVDD.n13848 0.2255
R1686 DVDD.n13842 DVDD.n13841 0.2255
R1687 DVDD.n12941 DVDD.n12940 0.222565
R1688 DVDD.n8958 DVDD.n8957 0.222565
R1689 DVDD.n12882 DVDD.n12881 0.222565
R1690 DVDD.n8985 DVDD.n8984 0.222565
R1691 DVDD.n4109 DVDD.n4103 0.222038
R1692 DVDD.n4358 DVDD.n4355 0.222038
R1693 DVDD.n17220 DVDD.n17218 0.220713
R1694 DVDD.n17218 DVDD.n17216 0.220713
R1695 DVDD.n14070 DVDD.n14068 0.220713
R1696 DVDD.n17387 DVDD.n17385 0.220713
R1697 DVDD.n17385 DVDD.n17383 0.220713
R1698 DVDD.n13981 DVDD.n13979 0.220713
R1699 DVDD.n17567 DVDD.n17566 0.220713
R1700 DVDD.n17566 DVDD.n17563 0.220713
R1701 DVDD.n14180 DVDD.n14177 0.220713
R1702 DVDD.n14323 DVDD.n14322 0.21611
R1703 DVDD.n17691 DVDD.n17690 0.21611
R1704 DVDD.n5882 DVDD.n5881 0.208315
R1705 DVDD.n12578 DVDD.n12577 0.208315
R1706 DVDD.n4348 DVDD.n4347 0.208315
R1707 DVDD.n8622 DVDD.n8621 0.208315
R1708 DVDD.n1090 DVDD 0.206051
R1709 DVDD DVDD.n1010 0.206051
R1710 DVDD DVDD.n1731 0.206051
R1711 DVDD DVDD.n11421 0.206051
R1712 DVDD DVDD.n1120 0.206051
R1713 DVDD DVDD.n1543 0.206049
R1714 DVDD.n1675 DVDD 0.206049
R1715 DVDD.n11542 DVDD 0.206049
R1716 DVDD.n18288 DVDD 0.206049
R1717 DVDD DVDD.n11914 0.206049
R1718 DVDD.n1284 DVDD 0.206049
R1719 DVDD.n12324 DVDD 0.206049
R1720 DVDD DVDD.n7160 0.204759
R1721 DVDD.n3158 DVDD 0.204759
R1722 DVDD.n9959 DVDD 0.204756
R1723 DVDD DVDD.n9813 0.204756
R1724 DVDD.n9520 DVDD 0.204756
R1725 DVDD DVDD.n3318 0.204756
R1726 DVDD.n5852 DVDD.n5851 0.202291
R1727 DVDD.n5835 DVDD.n5834 0.202291
R1728 DVDD.n12550 DVDD.n12549 0.202291
R1729 DVDD.n12533 DVDD.n12532 0.202291
R1730 DVDD.n4298 DVDD.n4297 0.202291
R1731 DVDD.n4273 DVDD.n4272 0.202291
R1732 DVDD.n8594 DVDD.n8593 0.202291
R1733 DVDD.n8577 DVDD.n8576 0.202291
R1734 DVDD.n5869 DVDD.n5868 0.200343
R1735 DVDD.n12567 DVDD.n12566 0.200343
R1736 DVDD.n4327 DVDD.n4326 0.200343
R1737 DVDD.n8611 DVDD.n8610 0.200343
R1738 DVDD.n5818 DVDD.n5817 0.200165
R1739 DVDD.n12516 DVDD.n12515 0.200165
R1740 DVDD.n4248 DVDD.n4247 0.200165
R1741 DVDD.n8560 DVDD.n8559 0.200165
R1742 DVDD DVDD.n7744 0.196382
R1743 DVDD.n6007 DVDD.n6001 0.183192
R1744 DVDD.n4467 DVDD.n4464 0.183192
R1745 DVDD.n5898 DVDD.n5895 0.183192
R1746 DVDD.n5919 DVDD.n5898 0.183192
R1747 DVDD.n8632 DVDD.n8629 0.183192
R1748 DVDD.n9903 DVDD.n9902 0.173278
R1749 DVDD DVDD.n18284 0.167265
R1750 DVDD.n14091 DVDD.n14090 0.164223
R1751 DVDD.n14002 DVDD.n14001 0.164223
R1752 DVDD.n14211 DVDD.n14210 0.164223
R1753 DVDD.n17241 DVDD.n17240 0.163984
R1754 DVDD.n17408 DVDD.n17407 0.163984
R1755 DVDD.n17590 DVDD.n17589 0.163984
R1756 DVDD.n14089 DVDD.n14086 0.156085
R1757 DVDD.n14000 DVDD.n13997 0.156085
R1758 DVDD.n14209 DVDD.n14204 0.156085
R1759 DVDD.n19771 DVDD.n19770 0.155874
R1760 DVDD.n19841 DVDD.n19840 0.155874
R1761 DVDD.n19996 DVDD.n19995 0.155874
R1762 DVDD.n4707 DVDD.n4706 0.155874
R1763 DVDD.n1416 DVDD.n1415 0.155874
R1764 DVDD.n1535 DVDD.n1534 0.155874
R1765 DVDD.n1684 DVDD.n1683 0.155874
R1766 DVDD.n11414 DVDD.n11413 0.155874
R1767 DVDD.n1993 DVDD.n1992 0.155874
R1768 DVDD.n2063 DVDD.n2062 0.155874
R1769 DVDD.n2217 DVDD.n2216 0.155874
R1770 DVDD.n6977 DVDD.n6976 0.155874
R1771 DVDD.n3187 DVDD.n3186 0.155874
R1772 DVDD.n3462 DVDD.n3461 0.155874
R1773 DVDD.n3565 DVDD.n3564 0.155874
R1774 DVDD.n9994 DVDD.n9993 0.155874
R1775 DVDD.n17239 DVDD.n17236 0.155846
R1776 DVDD.n17406 DVDD.n17403 0.155846
R1777 DVDD.n17588 DVDD.n17583 0.155846
R1778 DVDD.n1149 DVDD.n1148 0.149142
R1779 DVDD.n1554 DVDD.n1553 0.149142
R1780 DVDD.n1666 DVDD.n1665 0.149142
R1781 DVDD.n11470 DVDD.n11469 0.149142
R1782 DVDD.n3156 DVDD.n3120 0.141056
R1783 DVDD.n18392 DVDD.n18391 0.14
R1784 DVDD.n15939 DVDD.n15938 0.133067
R1785 DVDD.n12484 DVDD.n12478 0.128577
R1786 DVDD.n8753 DVDD.n8750 0.128577
R1787 DVDD.n17729 DVDD.n17726 0.128577
R1788 DVDD.n17726 DVDD.n17723 0.128577
R1789 DVDD.n14355 DVDD.n14330 0.128577
R1790 DVDD.n1241 DVDD.n1240 0.121593
R1791 DVDD.n7297 DVDD 0.114903
R1792 DVDD DVDD.n0 0.114226
R1793 DVDD DVDD.n7664 0.11306
R1794 DVDD.n7587 DVDD.n7583 0.112722
R1795 DVDD.n16352 DVDD.n16351 0.110256
R1796 DVDD.n16363 DVDD.n16362 0.110256
R1797 DVDD.n16329 DVDD.n16328 0.110256
R1798 DVDD.n16276 DVDD.n16275 0.110256
R1799 DVDD.n16267 DVDD.n16266 0.110256
R1800 DVDD.n16158 DVDD.n16157 0.110256
R1801 DVDD.n16149 DVDD.n16148 0.110256
R1802 DVDD.n16948 DVDD.n16947 0.110256
R1803 DVDD.n17006 DVDD.n17005 0.110256
R1804 DVDD.n11159 DVDD.n11158 0.110256
R1805 DVDD.n11147 DVDD.n11146 0.110256
R1806 DVDD.n16523 DVDD.n16522 0.110256
R1807 DVDD.n17164 DVDD.n17163 0.110256
R1808 DVDD.n17117 DVDD.n17116 0.110256
R1809 DVDD.n17067 DVDD.n17066 0.110256
R1810 DVDD.n11016 DVDD.n11015 0.110256
R1811 DVDD.n11024 DVDD.n11023 0.110256
R1812 DVDD.n11072 DVDD.n11071 0.110256
R1813 DVDD.n11079 DVDD.n11078 0.110256
R1814 DVDD.n15530 DVDD.n15529 0.110256
R1815 DVDD.n15524 DVDD.n15523 0.110256
R1816 DVDD.n11193 DVDD.n11192 0.110256
R1817 DVDD.n7543 DVDD.n7539 0.110054
R1818 DVDD.n12 DVDD.n8 0.109536
R1819 DVDD.n94 DVDD.n90 0.109536
R1820 DVDD.n40 DVDD.n36 0.109536
R1821 DVDD.n7189 DVDD.n7185 0.109536
R1822 DVDD.n20230 DVDD.n20226 0.109536
R1823 DVDD.n7689 DVDD.n7688 0.109536
R1824 DVDD.n7185 DVDD.n7184 0.108841
R1825 DVDD.n7690 DVDD.n7689 0.107849
R1826 DVDD.n7595 DVDD.n7594 0.107643
R1827 DVDD.n7597 DVDD.n7596 0.107643
R1828 DVDD.n7591 DVDD.n7590 0.107643
R1829 DVDD.n7587 DVDD.n7586 0.107643
R1830 DVDD.n7406 DVDD.n7405 0.107643
R1831 DVDD.n7402 DVDD.n7401 0.107643
R1832 DVDD.n7398 DVDD.n7397 0.107643
R1833 DVDD.n7394 DVDD.n7393 0.107643
R1834 DVDD.n7418 DVDD.n7417 0.107643
R1835 DVDD.n7422 DVDD.n7421 0.107643
R1836 DVDD.n7426 DVDD.n7425 0.107643
R1837 DVDD.n7380 DVDD.n7379 0.107643
R1838 DVDD.n7376 DVDD.n7375 0.107643
R1839 DVDD.n7372 DVDD.n7371 0.107643
R1840 DVDD.n7368 DVDD.n7367 0.107643
R1841 DVDD.n7364 DVDD.n7363 0.107643
R1842 DVDD.n7360 DVDD.n7359 0.107643
R1843 DVDD.n7356 DVDD.n7355 0.107643
R1844 DVDD.n108 DVDD.n107 0.107643
R1845 DVDD.n24 DVDD.n23 0.107643
R1846 DVDD.n20 DVDD.n19 0.107643
R1847 DVDD.n16 DVDD.n15 0.107643
R1848 DVDD.n7384 DVDD.n7383 0.107643
R1849 DVDD.n7386 DVDD.n7385 0.107643
R1850 DVDD.n7410 DVDD.n7409 0.107643
R1851 DVDD.n12 DVDD.n11 0.107643
R1852 DVDD.n7414 DVDD.n7413 0.107643
R1853 DVDD.n7390 DVDD.n7389 0.107643
R1854 DVDD.n7553 DVDD.n7552 0.107643
R1855 DVDD.n7551 DVDD.n7550 0.107643
R1856 DVDD.n7547 DVDD.n7546 0.107643
R1857 DVDD.n7543 DVDD.n7542 0.107643
R1858 DVDD.n7454 DVDD.n7453 0.107643
R1859 DVDD.n7450 DVDD.n7449 0.107643
R1860 DVDD.n7446 DVDD.n7445 0.107643
R1861 DVDD.n7442 DVDD.n7441 0.107643
R1862 DVDD.n7466 DVDD.n7465 0.107643
R1863 DVDD.n62 DVDD.n61 0.107643
R1864 DVDD.n66 DVDD.n65 0.107643
R1865 DVDD.n70 DVDD.n69 0.107643
R1866 DVDD.n74 DVDD.n73 0.107643
R1867 DVDD.n78 DVDD.n77 0.107643
R1868 DVDD.n82 DVDD.n81 0.107643
R1869 DVDD.n86 DVDD.n85 0.107643
R1870 DVDD.n88 DVDD.n87 0.107643
R1871 DVDD.n106 DVDD.n105 0.107643
R1872 DVDD.n102 DVDD.n101 0.107643
R1873 DVDD.n98 DVDD.n97 0.107643
R1874 DVDD.n58 DVDD.n57 0.107643
R1875 DVDD.n54 DVDD.n53 0.107643
R1876 DVDD.n94 DVDD.n93 0.107643
R1877 DVDD.n7474 DVDD.n7473 0.107643
R1878 DVDD.n7470 DVDD.n7469 0.107643
R1879 DVDD.n7462 DVDD.n7461 0.107643
R1880 DVDD.n7458 DVDD.n7457 0.107643
R1881 DVDD.n7438 DVDD.n7437 0.107643
R1882 DVDD.n7199 DVDD.n7198 0.107643
R1883 DVDD.n7193 DVDD.n7192 0.107643
R1884 DVDD.n7197 DVDD.n7196 0.107643
R1885 DVDD.n7503 DVDD.n7502 0.107643
R1886 DVDD.n7507 DVDD.n7506 0.107643
R1887 DVDD.n7499 DVDD.n7498 0.107643
R1888 DVDD.n7253 DVDD.n7252 0.107643
R1889 DVDD.n7249 DVDD.n7248 0.107643
R1890 DVDD.n7245 DVDD.n7244 0.107643
R1891 DVDD.n7241 DVDD.n7240 0.107643
R1892 DVDD.n7237 DVDD.n7236 0.107643
R1893 DVDD.n7233 DVDD.n7232 0.107643
R1894 DVDD.n7229 DVDD.n7228 0.107643
R1895 DVDD.n34 DVDD.n33 0.107643
R1896 DVDD.n52 DVDD.n51 0.107643
R1897 DVDD.n48 DVDD.n47 0.107643
R1898 DVDD.n44 DVDD.n43 0.107643
R1899 DVDD.n7259 DVDD.n7258 0.107643
R1900 DVDD.n7257 DVDD.n7256 0.107643
R1901 DVDD.n7479 DVDD.n7478 0.107643
R1902 DVDD.n7483 DVDD.n7482 0.107643
R1903 DVDD.n40 DVDD.n39 0.107643
R1904 DVDD.n7487 DVDD.n7486 0.107643
R1905 DVDD.n7491 DVDD.n7490 0.107643
R1906 DVDD.n7511 DVDD.n7510 0.107643
R1907 DVDD.n7495 DVDD.n7494 0.107643
R1908 DVDD.n7189 DVDD.n7188 0.107643
R1909 DVDD.n7623 DVDD.n7512 0.107643
R1910 DVDD.n15342 DVDD.n15341 0.107643
R1911 DVDD.n15352 DVDD.n15351 0.107643
R1912 DVDD.n15361 DVDD.n15360 0.107643
R1913 DVDD.n15368 DVDD.n15367 0.107643
R1914 DVDD.n15370 DVDD.n15369 0.107643
R1915 DVDD.n15372 DVDD.n15371 0.107643
R1916 DVDD.n15374 DVDD.n15373 0.107643
R1917 DVDD.n15376 DVDD.n15375 0.107643
R1918 DVDD.n15384 DVDD.n15383 0.107643
R1919 DVDD.n15326 DVDD.n15325 0.107643
R1920 DVDD.n15325 DVDD.n15324 0.107643
R1921 DVDD.n15320 DVDD.n15319 0.107643
R1922 DVDD.n15313 DVDD.n15312 0.107643
R1923 DVDD.n15073 DVDD.n15072 0.107643
R1924 DVDD.n15071 DVDD.n15070 0.107643
R1925 DVDD.n15069 DVDD.n15068 0.107643
R1926 DVDD.n15067 DVDD.n15066 0.107643
R1927 DVDD.n15065 DVDD.n15064 0.107643
R1928 DVDD.n15063 DVDD.n15062 0.107643
R1929 DVDD.n15061 DVDD.n15060 0.107643
R1930 DVDD.n15059 DVDD.n15058 0.107643
R1931 DVDD.n15052 DVDD.n15051 0.107643
R1932 DVDD.n15043 DVDD.n15042 0.107643
R1933 DVDD.n15035 DVDD.n15034 0.107643
R1934 DVDD.n15028 DVDD.n15027 0.107643
R1935 DVDD.n15026 DVDD.n15025 0.107643
R1936 DVDD.n15024 DVDD.n15023 0.107643
R1937 DVDD.n14975 DVDD.n14974 0.107643
R1938 DVDD.n14966 DVDD.n14965 0.107643
R1939 DVDD.n10353 DVDD.n10352 0.107643
R1940 DVDD.n10358 DVDD.n10357 0.107643
R1941 DVDD.n10360 DVDD.n10359 0.107643
R1942 DVDD.n10362 DVDD.n10361 0.107643
R1943 DVDD.n10364 DVDD.n10363 0.107643
R1944 DVDD.n10366 DVDD.n10365 0.107643
R1945 DVDD.n10373 DVDD.n10372 0.107643
R1946 DVDD.n10381 DVDD.n10380 0.107643
R1947 DVDD.n10732 DVDD.n10731 0.107643
R1948 DVDD.n10539 DVDD.n10538 0.107643
R1949 DVDD.n10537 DVDD.n10536 0.107643
R1950 DVDD.n10535 DVDD.n10534 0.107643
R1951 DVDD.n10533 DVDD.n10532 0.107643
R1952 DVDD.n10531 DVDD.n10530 0.107643
R1953 DVDD.n10529 DVDD.n10528 0.107643
R1954 DVDD.n10527 DVDD.n10526 0.107643
R1955 DVDD.n10525 DVDD.n10524 0.107643
R1956 DVDD.n10523 DVDD.n10522 0.107643
R1957 DVDD.n10516 DVDD.n10515 0.107643
R1958 DVDD.n10507 DVDD.n10506 0.107643
R1959 DVDD.n10501 DVDD.n10500 0.107643
R1960 DVDD.n10498 DVDD.n10497 0.107643
R1961 DVDD.n10496 DVDD.n10495 0.107643
R1962 DVDD.n10445 DVDD.n10444 0.107643
R1963 DVDD.n10436 DVDD.n10435 0.107643
R1964 DVDD.n10425 DVDD.n10424 0.107643
R1965 DVDD.n14936 DVDD.n14935 0.107643
R1966 DVDD.n14950 DVDD.n14949 0.107643
R1967 DVDD.n10337 DVDD.n10336 0.107643
R1968 DVDD.n10347 DVDD.n10346 0.107643
R1969 DVDD.n15912 DVDD.n15911 0.107643
R1970 DVDD.n15917 DVDD.n15916 0.107643
R1971 DVDD.n15918 DVDD.n15917 0.107643
R1972 DVDD.n15793 DVDD.n15792 0.107643
R1973 DVDD.n15804 DVDD.n15803 0.107643
R1974 DVDD.n15813 DVDD.n15812 0.107643
R1975 DVDD.n15816 DVDD.n15815 0.107643
R1976 DVDD.n15820 DVDD.n15819 0.107643
R1977 DVDD.n15822 DVDD.n15821 0.107643
R1978 DVDD.n15824 DVDD.n15823 0.107643
R1979 DVDD.n15826 DVDD.n15825 0.107643
R1980 DVDD.n15828 DVDD.n15827 0.107643
R1981 DVDD.n15832 DVDD.n15831 0.107643
R1982 DVDD.n15834 DVDD.n15833 0.107643
R1983 DVDD.n15836 DVDD.n15835 0.107643
R1984 DVDD.n15838 DVDD.n15837 0.107643
R1985 DVDD.n15847 DVDD.n15846 0.107643
R1986 DVDD.n15856 DVDD.n15855 0.107643
R1987 DVDD.n15867 DVDD.n15866 0.107643
R1988 DVDD.n15875 DVDD.n15874 0.107643
R1989 DVDD.n15877 DVDD.n15876 0.107643
R1990 DVDD.n15879 DVDD.n15878 0.107643
R1991 DVDD.n15885 DVDD.n15884 0.107643
R1992 DVDD.n15887 DVDD.n15886 0.107643
R1993 DVDD.n15889 DVDD.n15888 0.107643
R1994 DVDD.n15891 DVDD.n15890 0.107643
R1995 DVDD.n16112 DVDD.n16111 0.107643
R1996 DVDD.n16104 DVDD.n16103 0.107643
R1997 DVDD.n16096 DVDD.n16095 0.107643
R1998 DVDD.n16088 DVDD.n16087 0.107643
R1999 DVDD.n16086 DVDD.n16085 0.107643
R2000 DVDD.n16084 DVDD.n16083 0.107643
R2001 DVDD.n16082 DVDD.n16081 0.107643
R2002 DVDD.n16074 DVDD.n16073 0.107643
R2003 DVDD.n16556 DVDD.n16555 0.107643
R2004 DVDD.n16563 DVDD.n16562 0.107643
R2005 DVDD.n16571 DVDD.n16570 0.107643
R2006 DVDD.n16576 DVDD.n16575 0.107643
R2007 DVDD.n16692 DVDD.n16691 0.107643
R2008 DVDD.n16686 DVDD.n16685 0.107643
R2009 DVDD.n16684 DVDD.n16683 0.107643
R2010 DVDD.n16682 DVDD.n16681 0.107643
R2011 DVDD.n16678 DVDD.n16677 0.107643
R2012 DVDD.n16676 DVDD.n16675 0.107643
R2013 DVDD.n16669 DVDD.n16668 0.107643
R2014 DVDD.n16658 DVDD.n16657 0.107643
R2015 DVDD.n16650 DVDD.n16649 0.107643
R2016 DVDD.n16645 DVDD.n16644 0.107643
R2017 DVDD.n16643 DVDD.n16642 0.107643
R2018 DVDD.n16641 DVDD.n16640 0.107643
R2019 DVDD.n16637 DVDD.n16636 0.107643
R2020 DVDD.n16635 DVDD.n16634 0.107643
R2021 DVDD.n16631 DVDD.n16630 0.107643
R2022 DVDD.n16629 DVDD.n16628 0.107643
R2023 DVDD.n16625 DVDD.n16624 0.107643
R2024 DVDD.n16623 DVDD.n16622 0.107643
R2025 DVDD.n16619 DVDD.n16618 0.107643
R2026 DVDD.n16612 DVDD.n16611 0.107643
R2027 DVDD.n16601 DVDD.n16600 0.107643
R2028 DVDD.n16593 DVDD.n16592 0.107643
R2029 DVDD.n16588 DVDD.n16587 0.107643
R2030 DVDD.n16586 DVDD.n16585 0.107643
R2031 DVDD.n16584 DVDD.n16583 0.107643
R2032 DVDD.n16582 DVDD.n16581 0.107643
R2033 DVDD.n16580 DVDD.n16579 0.107643
R2034 DVDD.n16578 DVDD.n16577 0.107643
R2035 DVDD.n15757 DVDD.n15756 0.107643
R2036 DVDD.n15761 DVDD.n15760 0.107643
R2037 DVDD.n15763 DVDD.n15762 0.107643
R2038 DVDD.n15769 DVDD.n15768 0.107643
R2039 DVDD.n15771 DVDD.n15770 0.107643
R2040 DVDD.n15773 DVDD.n15772 0.107643
R2041 DVDD.n15775 DVDD.n15774 0.107643
R2042 DVDD.n15784 DVDD.n15783 0.107643
R2043 DVDD.n16814 DVDD.n16813 0.107643
R2044 DVDD.n16812 DVDD.n16811 0.107643
R2045 DVDD.n16810 DVDD.n16809 0.107643
R2046 DVDD.n16808 DVDD.n16807 0.107643
R2047 DVDD.n16806 DVDD.n16805 0.107643
R2048 DVDD.n16791 DVDD.n16790 0.107643
R2049 DVDD.n16781 DVDD.n16780 0.107643
R2050 DVDD.n16773 DVDD.n16772 0.107643
R2051 DVDD.n16768 DVDD.n16767 0.107643
R2052 DVDD.n16766 DVDD.n16765 0.107643
R2053 DVDD.n16764 DVDD.n16763 0.107643
R2054 DVDD.n16762 DVDD.n16761 0.107643
R2055 DVDD.n16760 DVDD.n16759 0.107643
R2056 DVDD.n16758 DVDD.n16757 0.107643
R2057 DVDD.n16756 DVDD.n16755 0.107643
R2058 DVDD.n16754 DVDD.n16753 0.107643
R2059 DVDD.n16752 DVDD.n16751 0.107643
R2060 DVDD.n16748 DVDD.n16747 0.107643
R2061 DVDD.n16914 DVDD.n16913 0.107643
R2062 DVDD.n16904 DVDD.n16903 0.107643
R2063 DVDD.n16896 DVDD.n16895 0.107643
R2064 DVDD.n16891 DVDD.n16890 0.107643
R2065 DVDD.n16887 DVDD.n16886 0.107643
R2066 DVDD.n16881 DVDD.n16880 0.107643
R2067 DVDD.n16177 DVDD.n16176 0.107643
R2068 DVDD.n16179 DVDD.n16178 0.107643
R2069 DVDD.n16187 DVDD.n16186 0.107643
R2070 DVDD.n16189 DVDD.n16188 0.107643
R2071 DVDD.n16191 DVDD.n16190 0.107643
R2072 DVDD.n16193 DVDD.n16192 0.107643
R2073 DVDD.n16195 DVDD.n16194 0.107643
R2074 DVDD.n16205 DVDD.n16204 0.107643
R2075 DVDD.n16214 DVDD.n16213 0.107643
R2076 DVDD.n16224 DVDD.n16223 0.107643
R2077 DVDD.n16231 DVDD.n16230 0.107643
R2078 DVDD.n15538 DVDD.n15537 0.107643
R2079 DVDD.n15544 DVDD.n15543 0.107643
R2080 DVDD.n15546 DVDD.n15545 0.107643
R2081 DVDD.n15548 DVDD.n15547 0.107643
R2082 DVDD.n15550 DVDD.n15549 0.107643
R2083 DVDD.n15552 DVDD.n15551 0.107643
R2084 DVDD.n15556 DVDD.n15555 0.107643
R2085 DVDD.n15558 DVDD.n15557 0.107643
R2086 DVDD.n15560 DVDD.n15559 0.107643
R2087 DVDD.n15570 DVDD.n15569 0.107643
R2088 DVDD.n15579 DVDD.n15578 0.107643
R2089 DVDD.n15589 DVDD.n15588 0.107643
R2090 DVDD.n15596 DVDD.n15595 0.107643
R2091 DVDD.n15598 DVDD.n15597 0.107643
R2092 DVDD.n15602 DVDD.n15601 0.107643
R2093 DVDD.n15604 DVDD.n15603 0.107643
R2094 DVDD.n15606 DVDD.n15605 0.107643
R2095 DVDD.n15608 DVDD.n15607 0.107643
R2096 DVDD.n15610 DVDD.n15609 0.107643
R2097 DVDD.n15612 DVDD.n15611 0.107643
R2098 DVDD.n15752 DVDD.n15751 0.107643
R2099 DVDD.n15744 DVDD.n15743 0.107643
R2100 DVDD.n15737 DVDD.n15736 0.107643
R2101 DVDD.n15729 DVDD.n15728 0.107643
R2102 DVDD.n15727 DVDD.n15726 0.107643
R2103 DVDD.n15725 DVDD.n15724 0.107643
R2104 DVDD.n15723 DVDD.n15722 0.107643
R2105 DVDD.n15716 DVDD.n15715 0.107643
R2106 DVDD.n15707 DVDD.n15706 0.107643
R2107 DVDD.n15708 DVDD.n15707 0.107643
R2108 DVDD.n15699 DVDD.n15698 0.107643
R2109 DVDD.n16725 DVDD.n16724 0.107643
R2110 DVDD.n16732 DVDD.n16731 0.107643
R2111 DVDD.n16739 DVDD.n16738 0.107643
R2112 DVDD.n16744 DVDD.n16743 0.107643
R2113 DVDD.n16380 DVDD.n16376 0.107643
R2114 DVDD.n16381 DVDD.n16380 0.107643
R2115 DVDD.n16340 DVDD.n16339 0.107643
R2116 DVDD.n16337 DVDD.n16336 0.107643
R2117 DVDD.n16335 DVDD.n16334 0.107643
R2118 DVDD.n16311 DVDD.n16310 0.107643
R2119 DVDD.n16309 DVDD.n16308 0.107643
R2120 DVDD.n16307 DVDD.n16306 0.107643
R2121 DVDD.n16305 DVDD.n16304 0.107643
R2122 DVDD.n16303 DVDD.n16302 0.107643
R2123 DVDD.n16301 DVDD.n16300 0.107643
R2124 DVDD.n16299 DVDD.n16298 0.107643
R2125 DVDD.n16295 DVDD.n16294 0.107643
R2126 DVDD.n16258 DVDD.n16257 0.107643
R2127 DVDD.n16256 DVDD.n16255 0.107643
R2128 DVDD.n16254 DVDD.n16253 0.107643
R2129 DVDD.n16252 DVDD.n16251 0.107643
R2130 DVDD.n16250 DVDD.n16249 0.107643
R2131 DVDD.n16248 DVDD.n16247 0.107643
R2132 DVDD.n16246 DVDD.n16245 0.107643
R2133 DVDD.n16244 DVDD.n16243 0.107643
R2134 DVDD.n16240 DVDD.n16239 0.107643
R2135 DVDD.n16238 DVDD.n16237 0.107643
R2136 DVDD.n16236 DVDD.n16235 0.107643
R2137 DVDD.n16175 DVDD.n16174 0.107643
R2138 DVDD.n16138 DVDD.n16137 0.107643
R2139 DVDD.n16136 DVDD.n16135 0.107643
R2140 DVDD.n16134 DVDD.n16133 0.107643
R2141 DVDD.n16130 DVDD.n16129 0.107643
R2142 DVDD.n16128 DVDD.n16127 0.107643
R2143 DVDD.n16126 DVDD.n16125 0.107643
R2144 DVDD.n16120 DVDD.n16119 0.107643
R2145 DVDD.n16925 DVDD.n16924 0.107643
R2146 DVDD.n16929 DVDD.n16928 0.107643
R2147 DVDD.n16931 DVDD.n16930 0.107643
R2148 DVDD.n16933 DVDD.n16932 0.107643
R2149 DVDD.n16991 DVDD.n16990 0.107643
R2150 DVDD.n16989 DVDD.n16988 0.107643
R2151 DVDD.n16987 DVDD.n16986 0.107643
R2152 DVDD.n16985 DVDD.n16984 0.107643
R2153 DVDD.n16983 DVDD.n16982 0.107643
R2154 DVDD.n16981 DVDD.n16980 0.107643
R2155 DVDD.n16979 DVDD.n16978 0.107643
R2156 DVDD.n16977 DVDD.n16976 0.107643
R2157 DVDD.n16975 DVDD.n16974 0.107643
R2158 DVDD.n16973 DVDD.n16972 0.107643
R2159 DVDD.n16965 DVDD.n16964 0.107643
R2160 DVDD.n16940 DVDD.n16939 0.107643
R2161 DVDD.n16993 DVDD.n16992 0.107643
R2162 DVDD.n16998 DVDD.n16997 0.107643
R2163 DVDD.n16879 DVDD.n16878 0.107643
R2164 DVDD.n16858 DVDD.n16857 0.107643
R2165 DVDD.n17041 DVDD.n17040 0.107643
R2166 DVDD.n17039 DVDD.n17038 0.107643
R2167 DVDD.n17035 DVDD.n17034 0.107643
R2168 DVDD.n17033 DVDD.n17032 0.107643
R2169 DVDD.n17031 DVDD.n17030 0.107643
R2170 DVDD.n17025 DVDD.n17024 0.107643
R2171 DVDD.n11185 DVDD.n11184 0.107643
R2172 DVDD.n11183 DVDD.n11182 0.107643
R2173 DVDD.n11181 DVDD.n11180 0.107643
R2174 DVDD.n11179 DVDD.n11178 0.107643
R2175 DVDD.n11177 DVDD.n11176 0.107643
R2176 DVDD.n11144 DVDD.n11143 0.107643
R2177 DVDD.n11142 DVDD.n11141 0.107643
R2178 DVDD.n16516 DVDD.n16515 0.107643
R2179 DVDD.n17158 DVDD.n17157 0.107643
R2180 DVDD.n17150 DVDD.n17149 0.107643
R2181 DVDD.n17148 DVDD.n17147 0.107643
R2182 DVDD.n17146 DVDD.n17145 0.107643
R2183 DVDD.n17144 DVDD.n17143 0.107643
R2184 DVDD.n17142 DVDD.n17141 0.107643
R2185 DVDD.n17138 DVDD.n17137 0.107643
R2186 DVDD.n17134 DVDD.n17133 0.107643
R2187 DVDD.n17112 DVDD.n17111 0.107643
R2188 DVDD.n17109 DVDD.n17108 0.107643
R2189 DVDD.n17107 DVDD.n17106 0.107643
R2190 DVDD.n17103 DVDD.n17102 0.107643
R2191 DVDD.n17101 DVDD.n17100 0.107643
R2192 DVDD.n17097 DVDD.n17096 0.107643
R2193 DVDD.n17095 DVDD.n17094 0.107643
R2194 DVDD.n17093 DVDD.n17092 0.107643
R2195 DVDD.n17089 DVDD.n17088 0.107643
R2196 DVDD.n17087 DVDD.n17086 0.107643
R2197 DVDD.n17062 DVDD.n17061 0.107643
R2198 DVDD.n17057 DVDD.n17056 0.107643
R2199 DVDD.n17055 DVDD.n17054 0.107643
R2200 DVDD.n17053 DVDD.n17052 0.107643
R2201 DVDD.n17051 DVDD.n17050 0.107643
R2202 DVDD.n17047 DVDD.n17046 0.107643
R2203 DVDD.n17045 DVDD.n17044 0.107643
R2204 DVDD.n10992 DVDD.n10991 0.107643
R2205 DVDD.n10996 DVDD.n10995 0.107643
R2206 DVDD.n10998 DVDD.n10997 0.107643
R2207 DVDD.n11000 DVDD.n10999 0.107643
R2208 DVDD.n11002 DVDD.n11001 0.107643
R2209 DVDD.n11004 DVDD.n11003 0.107643
R2210 DVDD.n11006 DVDD.n11005 0.107643
R2211 DVDD.n11008 DVDD.n11007 0.107643
R2212 DVDD.n11039 DVDD.n11038 0.107643
R2213 DVDD.n11045 DVDD.n11044 0.107643
R2214 DVDD.n11047 DVDD.n11046 0.107643
R2215 DVDD.n11049 DVDD.n11048 0.107643
R2216 DVDD.n11051 DVDD.n11050 0.107643
R2217 DVDD.n11053 DVDD.n11052 0.107643
R2218 DVDD.n11055 DVDD.n11054 0.107643
R2219 DVDD.n11057 DVDD.n11056 0.107643
R2220 DVDD.n11059 DVDD.n11058 0.107643
R2221 DVDD.n11061 DVDD.n11060 0.107643
R2222 DVDD.n11063 DVDD.n11062 0.107643
R2223 DVDD.n11065 DVDD.n11064 0.107643
R2224 DVDD.n11096 DVDD.n11095 0.107643
R2225 DVDD.n11098 DVDD.n11097 0.107643
R2226 DVDD.n11100 DVDD.n11099 0.107643
R2227 DVDD.n11102 DVDD.n11101 0.107643
R2228 DVDD.n11104 DVDD.n11103 0.107643
R2229 DVDD.n11106 DVDD.n11105 0.107643
R2230 DVDD.n11108 DVDD.n11107 0.107643
R2231 DVDD.n11110 DVDD.n11109 0.107643
R2232 DVDD.n11123 DVDD.n11122 0.107643
R2233 DVDD.n7684 DVDD.n7683 0.107643
R2234 DVDD.n7676 DVDD.n7675 0.107643
R2235 DVDD.n7680 DVDD.n7679 0.107643
R2236 DVDD.n7688 DVDD.n7687 0.107643
R2237 DVDD.n7306 DVDD.n7305 0.107643
R2238 DVDD.n7322 DVDD.n7321 0.107643
R2239 DVDD.n7318 DVDD.n7317 0.107643
R2240 DVDD.n7314 DVDD.n7313 0.107643
R2241 DVDD.n7310 DVDD.n7309 0.107643
R2242 DVDD.n7334 DVDD.n7333 0.107643
R2243 DVDD.n7338 DVDD.n7337 0.107643
R2244 DVDD.n7342 DVDD.n7341 0.107643
R2245 DVDD.n20252 DVDD.n20251 0.107643
R2246 DVDD.n20256 DVDD.n20255 0.107643
R2247 DVDD.n20260 DVDD.n20259 0.107643
R2248 DVDD.n20264 DVDD.n20263 0.107643
R2249 DVDD.n20268 DVDD.n20267 0.107643
R2250 DVDD.n20272 DVDD.n20271 0.107643
R2251 DVDD.n20276 DVDD.n20275 0.107643
R2252 DVDD.n20340 DVDD.n20339 0.107643
R2253 DVDD.n20242 DVDD.n20241 0.107643
R2254 DVDD.n20238 DVDD.n20237 0.107643
R2255 DVDD.n20234 DVDD.n20233 0.107643
R2256 DVDD.n20248 DVDD.n20247 0.107643
R2257 DVDD.n20244 DVDD.n20243 0.107643
R2258 DVDD.n7330 DVDD.n7329 0.107643
R2259 DVDD.n7326 DVDD.n7325 0.107643
R2260 DVDD.n20230 DVDD.n20229 0.107643
R2261 DVDD.n7297 DVDD.n7204 0.107557
R2262 DVDD.n20216 DVDD.n20215 0.0993568
R2263 DVDD.n7539 DVDD.n7538 0.0989868
R2264 DVDD.n7598 DVDD 0.0970016
R2265 DVDD.n7583 DVDD.n7582 0.0969425
R2266 DVDD DVDD.n0 0.0938784
R2267 DVDD.n374 DVDD.n373 0.0929542
R2268 DVDD.n605 DVDD.n604 0.0929542
R2269 DVDD.n13736 DVDD.n13735 0.0929542
R2270 DVDD.n9027 DVDD.n9026 0.092212
R2271 DVDD.n9022 DVDD.n9019 0.092212
R2272 DVDD.n12920 DVDD.n12919 0.0919674
R2273 DVDD.n12915 DVDD.n12912 0.0919674
R2274 DVDD.n20341 DVDD.n20216 0.0916836
R2275 DVDD.n7674 DVDD.n7598 0.0908035
R2276 DVDD.n2690 DVDD 0.0894467
R2277 DVDD.n10330 DVDD.n10329 0.0889932
R2278 DVDD DVDD.n7302 0.0870792
R2279 DVDD DVDD.n11224 0.0817673
R2280 DVDD.n373 DVDD.n372 0.0800338
R2281 DVDD.n604 DVDD.n603 0.0800338
R2282 DVDD.n13737 DVDD.n13736 0.0800338
R2283 DVDD.n2485 DVDD 0.0786244
R2284 DVDD.n4777 DVDD.n4776 0.0763268
R2285 DVDD.n11603 DVDD.n11602 0.0763268
R2286 DVDD.n6907 DVDD.n6906 0.0763268
R2287 DVDD.n7859 DVDD.n7858 0.0763268
R2288 DVDD.n11487 DVDD.n11486 0.0729606
R2289 DVDD.n2691 DVDD.n2690 0.0715072
R2290 DVDD.n14009 DVDD.n14008 0.0709162
R2291 DVDD.n14220 DVDD.n14219 0.0709162
R2292 DVDD.n16349 DVDD 0.0661438
R2293 DVDD.n7744 DVDD.n7742 0.0640294
R2294 DVDD.n18284 DVDD.n18282 0.0640294
R2295 DVDD.n17356 DVDD.n17355 0.0624362
R2296 DVDD.n17516 DVDD.n17515 0.0624362
R2297 DVDD.n14103 DVDD.n14102 0.061834
R2298 DVDD.n15463 DVDD.n15462 0.0617992
R2299 DVDD.n18144 DVDD.n18143 0.0617992
R2300 DVDD.n10329 DVDD.n10328 0.0617844
R2301 DVDD.n13530 DVDD.n13529 0.0584331
R2302 DVDD.n14591 DVDD.n14590 0.0584331
R2303 DVDD.n17951 DVDD.n17950 0.0584331
R2304 DVDD.n13611 DVDD.n13610 0.0582559
R2305 DVDD.n14673 DVDD.n14672 0.0582559
R2306 DVDD.n14503 DVDD.n14502 0.0582559
R2307 DVDD.n5695 DVDD.n5694 0.0582559
R2308 DVDD.n12746 DVDD.n12745 0.0582559
R2309 DVDD.n18029 DVDD.n18028 0.0582559
R2310 DVDD.n17870 DVDD.n17869 0.0582559
R2311 DVDD.n6128 DVDD.n6127 0.0582559
R2312 DVDD.n8830 DVDD.n8829 0.0582559
R2313 DVDD.n16832 DVDD.n16820 0.0580122
R2314 DVDD.n16488 DVDD.n16476 0.0580122
R2315 DVDD.n17290 DVDD.n17288 0.0576622
R2316 DVDD.n13907 DVDD.n13905 0.0576622
R2317 DVDD.n17669 DVDD.n17666 0.0576622
R2318 DVDD.n14296 DVDD.n14293 0.0576622
R2319 DVDD.n2485 DVDD 0.0567182
R2320 DVDD.n11224 DVDD 0.0567182
R2321 DVDD.n3333 DVDD.n3332 0.0563
R2322 DVDD.n3334 DVDD.n3333 0.0563
R2323 DVDD.n3335 DVDD.n3334 0.0563
R2324 DVDD.n3336 DVDD.n3335 0.0563
R2325 DVDD.n3337 DVDD.n3336 0.0563
R2326 DVDD.n3338 DVDD.n3337 0.0563
R2327 DVDD.n3339 DVDD.n3338 0.0563
R2328 DVDD.n3340 DVDD.n3339 0.0563
R2329 DVDD.n3341 DVDD.n3340 0.0563
R2330 DVDD.n3342 DVDD.n3341 0.0563
R2331 DVDD.n3343 DVDD.n3342 0.0563
R2332 DVDD.n3344 DVDD.n3343 0.0563
R2333 DVDD.n3345 DVDD.n3344 0.0563
R2334 DVDD.n3346 DVDD.n3345 0.0563
R2335 DVDD.n3347 DVDD.n3346 0.0563
R2336 DVDD.n3348 DVDD.n3347 0.0563
R2337 DVDD.n3349 DVDD.n3348 0.0563
R2338 DVDD.n3350 DVDD.n3349 0.0563
R2339 DVDD.n3351 DVDD.n3350 0.0563
R2340 DVDD.n3352 DVDD.n3351 0.0563
R2341 DVDD.n3353 DVDD.n3352 0.0563
R2342 DVDD.n3354 DVDD.n3353 0.0563
R2343 DVDD.n3446 DVDD.n3354 0.0563
R2344 DVDD.n3439 DVDD.n3438 0.0563
R2345 DVDD.n3438 DVDD.n3437 0.0563
R2346 DVDD.n3437 DVDD.n3436 0.0563
R2347 DVDD.n3436 DVDD.n3435 0.0563
R2348 DVDD.n3435 DVDD.n3434 0.0563
R2349 DVDD.n3434 DVDD.n3433 0.0563
R2350 DVDD.n3358 DVDD.n3357 0.0563
R2351 DVDD.n3357 DVDD.n3356 0.0563
R2352 DVDD.n3356 DVDD.n3355 0.0563
R2353 DVDD.n3355 DVDD.n2866 0.0563
R2354 DVDD.n3580 DVDD.n2866 0.0563
R2355 DVDD.n7791 DVDD.n7790 0.0563
R2356 DVDD.n7792 DVDD.n7791 0.0563
R2357 DVDD.n7793 DVDD.n7792 0.0563
R2358 DVDD.n7794 DVDD.n7793 0.0563
R2359 DVDD.n7795 DVDD.n7794 0.0563
R2360 DVDD.n7796 DVDD.n7795 0.0563
R2361 DVDD.n7797 DVDD.n7796 0.0563
R2362 DVDD.n7798 DVDD.n7797 0.0563
R2363 DVDD.n7799 DVDD.n7798 0.0563
R2364 DVDD.n7800 DVDD.n7799 0.0563
R2365 DVDD.n7801 DVDD.n7800 0.0563
R2366 DVDD.n7802 DVDD.n7801 0.0563
R2367 DVDD.n7803 DVDD.n7802 0.0563
R2368 DVDD.n7804 DVDD.n7803 0.0563
R2369 DVDD.n7805 DVDD.n7804 0.0563
R2370 DVDD.n7806 DVDD.n7805 0.0563
R2371 DVDD.n7807 DVDD.n7806 0.0563
R2372 DVDD.n17193 DVDD.n17192 0.0555679
R2373 DVDD.n19316 DVDD.n19315 0.0554213
R2374 DVDD.n16349 DVDD.n16345 0.0532076
R2375 DVDD.n7662 DVDD.n7660 0.052798
R2376 DVDD.n2022 DVDD 0.0502899
R2377 DVDD.n2154 DVDD 0.0502899
R2378 DVDD.n2230 DVDD 0.0502899
R2379 DVDD.n7098 DVDD 0.0502899
R2380 DVDD.n6936 DVDD 0.0502899
R2381 DVDD.n6784 DVDD 0.0502899
R2382 DVDD.n6518 DVDD 0.0502899
R2383 DVDD.n1857 DVDD 0.0502899
R2384 DVDD.n3923 DVDD 0.0502899
R2385 DVDD.n19800 DVDD 0.0502899
R2386 DVDD.n19933 DVDD 0.0502899
R2387 DVDD.n20009 DVDD 0.0502899
R2388 DVDD.n3877 DVDD 0.0502899
R2389 DVDD.n4710 DVDD 0.0502899
R2390 DVDD.n4821 DVDD 0.0502899
R2391 DVDD.n5109 DVDD 0.0502899
R2392 DVDD.n19635 DVDD 0.0502899
R2393 DVDD.n5228 DVDD 0.0502899
R2394 DVDD.n2053 DVDD 0.0502827
R2395 DVDD.n2207 DVDD 0.0502827
R2396 DVDD.n18929 DVDD 0.0502827
R2397 DVDD.n7031 DVDD 0.0502827
R2398 DVDD.n6941 DVDD 0.0502827
R2399 DVDD.n6800 DVDD 0.0502827
R2400 DVDD.n6551 DVDD 0.0502827
R2401 DVDD.n1860 DVDD 0.0502827
R2402 DVDD.n3928 DVDD 0.0502827
R2403 DVDD.n19831 DVDD 0.0502827
R2404 DVDD.n19986 DVDD 0.0502827
R2405 DVDD.n19047 DVDD 0.0502827
R2406 DVDD.n4611 DVDD 0.0502827
R2407 DVDD.n4715 DVDD 0.0502827
R2408 DVDD.n4837 DVDD 0.0502827
R2409 DVDD.n5142 DVDD 0.0502827
R2410 DVDD.n19638 DVDD 0.0502827
R2411 DVDD.n5233 DVDD 0.0502827
R2412 DVDD.n18346 DVDD.n18345 0.04775
R2413 DVDD.n20338 DVDD.n20302 0.047668
R2414 DVDD.n7301 DVDD.n7300 0.047612
R2415 DVDD.n10469 DVDD.n10468 0.0475895
R2416 DVDD.n7790 DVDD.n7693 0.0473
R2417 DVDD.n3446 DVDD.n3445 0.04685
R2418 DVDD.n3581 DVDD.n3580 0.04685
R2419 DVDD.n7808 DVDD.n7807 0.04685
R2420 DVDD.n3332 DVDD.n3331 0.0464
R2421 DVDD.n3440 DVDD.n3439 0.0464
R2422 DVDD.n3668 DVDD.n3586 0.0464
R2423 DVDD.n18645 DVDD.n18644 0.0464
R2424 DVDD.n18777 DVDD 0.0463897
R2425 DVDD.n10469 DVDD.n10467 0.0463522
R2426 DVDD.n7301 DVDD.n7299 0.0462939
R2427 DVDD.n7662 DVDD.n7661 0.0457907
R2428 DVDD.n20338 DVDD.n20337 0.0457773
R2429 DVDD.n3359 DVDD.n3358 0.0455
R2430 DVDD.n16707 DVDD.n16706 0.0452896
R2431 DVDD.n1905 DVDD.n1904 0.0448795
R2432 DVDD.n19683 DVDD.n19682 0.0448795
R2433 DVDD.n1328 DVDD.n1327 0.0448795
R2434 DVDD.n3275 DVDD.n3274 0.0448795
R2435 DVDD.n11341 DVDD 0.0446291
R2436 DVDD DVDD.n11338 0.0446291
R2437 DVDD.n11300 DVDD 0.0446291
R2438 DVDD.n19430 DVDD 0.0446286
R2439 DVDD DVDD.n13224 0.0446286
R2440 DVDD.n7816 DVDD 0.0445411
R2441 DVDD DVDD.n7936 0.0445411
R2442 DVDD.n8362 DVDD 0.0445411
R2443 DVDD DVDD.n9313 0.0445405
R2444 DVDD.n16489 DVDD.n16488 0.0433911
R2445 DVDD.n16833 DVDD.n16832 0.0433911
R2446 DVDD.n16538 DVDD.n16537 0.0433911
R2447 DVDD.n3433 DVDD.n3432 0.0428
R2448 DVDD.n11140 DVDD 0.0423002
R2449 DVDD.n1905 DVDD.n1859 0.0420792
R2450 DVDD.n19683 DVDD.n19637 0.0420792
R2451 DVDD.n3668 DVDD.n3667 0.0419
R2452 DVDD.n18349 DVDD.n18348 0.04055
R2453 DVDD.n18740 DVDD.n18739 0.0392
R2454 DVDD.n15915 DVDD.n15914 0.0384256
R2455 DVDD.n15339 DVDD 0.0373056
R2456 DVDD.n1242 DVDD.n1241 0.0356325
R2457 DVDD.n18343 DVDD.n18342 0.03515
R2458 DVDD.n3036 DVDD.n3035 0.0349444
R2459 DVDD.n3035 DVDD.n3034 0.0349444
R2460 DVDD.n3034 DVDD.n3033 0.0349444
R2461 DVDD.n3033 DVDD.n3032 0.0349444
R2462 DVDD.n3032 DVDD.n3028 0.0349444
R2463 DVDD.n3325 DVDD.n3028 0.0349444
R2464 DVDD.n11140 DVDD.n11139 0.0346544
R2465 DVDD.n13736 DVDD.n11266 0.0333127
R2466 DVDD.n373 DVDD.n304 0.0333127
R2467 DVDD.n604 DVDD.n535 0.0333127
R2468 DVDD.n3156 DVDD.n3155 0.033206
R2469 DVDD.n15339 DVDD 0.03312
R2470 DVDD.n15914 DVDD 0.03312
R2471 DVDD.n7216 DVDD.n7215 0.0324667
R2472 DVDD.n10693 DVDD.n10692 0.0324667
R2473 DVDD.n7626 DVDD.n7625 0.0322741
R2474 DVDD.n20314 DVDD.n20313 0.0322741
R2475 DVDD.n15075 DVDD.n15074 0.0322733
R2476 DVDD.n7287 DVDD.n7286 0.0322733
R2477 DVDD.n7650 DVDD.n7649 0.0321049
R2478 DVDD.n20292 DVDD.n20291 0.0321049
R2479 DVDD.n3426 DVDD.n3425 0.032
R2480 DVDD.n3419 DVDD.n3418 0.032
R2481 DVDD.n3413 DVDD.n3412 0.032
R2482 DVDD.n3406 DVDD.n3405 0.032
R2483 DVDD.n3399 DVDD.n3398 0.032
R2484 DVDD.n3393 DVDD.n3392 0.032
R2485 DVDD.n3387 DVDD.n3386 0.032
R2486 DVDD.n3380 DVDD.n3379 0.032
R2487 DVDD.n3373 DVDD.n3372 0.032
R2488 DVDD.n3366 DVDD.n3365 0.032
R2489 DVDD.n3661 DVDD.n3660 0.032
R2490 DVDD.n3654 DVDD.n3653 0.032
R2491 DVDD.n3606 DVDD.n3605 0.032
R2492 DVDD.n3599 DVDD.n3598 0.032
R2493 DVDD.n3592 DVDD.n3591 0.032
R2494 DVDD.n18430 DVDD.n18429 0.032
R2495 DVDD.n18446 DVDD.n18445 0.032
R2496 DVDD.n14748 DVDD.n14747 0.032
R2497 DVDD.n14753 DVDD.n14752 0.032
R2498 DVDD.n14769 DVDD.n14768 0.032
R2499 DVDD.n14762 DVDD.n14761 0.032
R2500 DVDD.n9471 DVDD.n9470 0.0306622
R2501 DVDD.n9470 DVDD.n9469 0.0306622
R2502 DVDD.n9469 DVDD.n9468 0.0306622
R2503 DVDD.n9468 DVDD.n9467 0.0306622
R2504 DVDD.n9467 DVDD.n9466 0.0306622
R2505 DVDD.n9466 DVDD.n9465 0.0306622
R2506 DVDD.n9465 DVDD.n9464 0.0306622
R2507 DVDD.n9464 DVDD.n9463 0.0306622
R2508 DVDD.n9463 DVDD.n9462 0.0306622
R2509 DVDD.n9462 DVDD.n9461 0.0306622
R2510 DVDD.n9461 DVDD.n9460 0.0306622
R2511 DVDD.n9460 DVDD.n9459 0.0306622
R2512 DVDD.n9459 DVDD.n9458 0.0306622
R2513 DVDD.n9458 DVDD.n9457 0.0306622
R2514 DVDD.n8099 DVDD.n8098 0.0306622
R2515 DVDD.n9929 DVDD.n9928 0.0306622
R2516 DVDD.n9928 DVDD.n9927 0.0306622
R2517 DVDD.n9927 DVDD.n9926 0.0306622
R2518 DVDD.n9926 DVDD.n9925 0.0306622
R2519 DVDD.n9925 DVDD.n9924 0.0306622
R2520 DVDD.n9924 DVDD.n9923 0.0306622
R2521 DVDD.n9923 DVDD.n9922 0.0306622
R2522 DVDD.n9922 DVDD.n9921 0.0306622
R2523 DVDD.n9921 DVDD.n9920 0.0306622
R2524 DVDD.n9920 DVDD.n9919 0.0306622
R2525 DVDD.n9919 DVDD.n9918 0.0306622
R2526 DVDD.n9918 DVDD.n9917 0.0306622
R2527 DVDD.n9917 DVDD.n9916 0.0306622
R2528 DVDD.n9916 DVDD.n9915 0.0306622
R2529 DVDD.n9915 DVDD.n9914 0.0306622
R2530 DVDD.n9914 DVDD.n9913 0.0306622
R2531 DVDD.n9913 DVDD.n9912 0.0306622
R2532 DVDD.n9912 DVDD.n9911 0.0306622
R2533 DVDD.n9911 DVDD.n9910 0.0306622
R2534 DVDD.n9910 DVDD.n9909 0.0306622
R2535 DVDD.n9909 DVDD.n9908 0.0306622
R2536 DVDD.n9908 DVDD.n9907 0.0306622
R2537 DVDD.n9907 DVDD.n9906 0.0306622
R2538 DVDD.n7635 DVDD.n7634 0.03065
R2539 DVDD.n7659 DVDD.n7658 0.03065
R2540 DVDD.n20301 DVDD.n20300 0.03065
R2541 DVDD.n20323 DVDD.n20322 0.03065
R2542 DVDD.n7225 DVDD.n7224 0.030425
R2543 DVDD.n7264 DVDD.n7263 0.030425
R2544 DVDD.n7613 DVDD.n7612 0.030425
R2545 DVDD.n7640 DVDD.n7639 0.030425
R2546 DVDD.n20281 DVDD.n20280 0.030425
R2547 DVDD.n20328 DVDD.n20327 0.030425
R2548 DVDD.n15084 DVDD.n15083 0.030425
R2549 DVDD.n15089 DVDD.n15088 0.030425
R2550 DVDD.n10702 DVDD.n10701 0.030425
R2551 DVDD.n10707 DVDD.n10706 0.030425
R2552 DVDD.n7296 DVDD.n7295 0.030425
R2553 DVDD.n7277 DVDD.n7276 0.030425
R2554 DVDD.n8296 DVDD.n8295 0.0304189
R2555 DVDD.n8297 DVDD.n8296 0.0299324
R2556 DVDD.n6105 DVDD.n6104 0.0295115
R2557 DVDD.n12448 DVDD.n12447 0.0295115
R2558 DVDD.n4558 DVDD.n4557 0.0295115
R2559 DVDD.n8472 DVDD.n8471 0.0295115
R2560 DVDD.n12435 DVDD.n12434 0.0295115
R2561 DVDD.n5620 DVDD.n5619 0.0295115
R2562 DVDD.n4573 DVDD.n4572 0.0295115
R2563 DVDD.n8454 DVDD.n8453 0.0295115
R2564 DVDD.n12416 DVDD.n12415 0.0295115
R2565 DVDD.n4588 DVDD.n4587 0.0295115
R2566 DVDD.n8436 DVDD.n8435 0.0295115
R2567 DVDD.n3326 DVDD.n3325 0.0291111
R2568 DVDD.n8098 DVDD.n8097 0.0289595
R2569 DVDD.n15704 DVDD 0.0288569
R2570 DVDD.n9472 DVDD.n9471 0.0287162
R2571 DVDD.n18992 DVDD.n18991 0.0284
R2572 DVDD.n19152 DVDD.n19151 0.0284
R2573 DVDD.n3846 DVDD.n3845 0.0284
R2574 DVDD.n10072 DVDD.n10071 0.0284
R2575 DVDD.n131 DVDD.n130 0.0284
R2576 DVDD.n1808 DVDD.n1807 0.0284
R2577 DVDD.n10595 DVDD.n10594 0.0284
R2578 DVDD.n10614 DVDD.n10613 0.0284
R2579 DVDD.n15705 DVDD.n15704 0.0282682
R2580 DVDD.n18423 DVDD.n18422 0.02795
R2581 DVDD.n18439 DVDD.n18438 0.0275
R2582 DVDD.n3001 DVDD 0.0269933
R2583 DVDD DVDD.n3674 0.026993
R2584 DVDD DVDD.n2916 0.026993
R2585 DVDD.n3575 DVDD 0.0269892
R2586 DVDD.n7768 DVDD 0.0269892
R2587 DVDD DVDD.n3452 0.0269892
R2588 DVDD.n7610 DVDD.n7609 0.0269368
R2589 DVDD.n20325 DVDD.n20324 0.0269368
R2590 DVDD.n7261 DVDD.n7260 0.0267443
R2591 DVDD.n10704 DVDD.n10703 0.0267443
R2592 DVDD.n7637 DVDD.n7636 0.0266462
R2593 DVDD.n20278 DVDD.n20277 0.0266462
R2594 DVDD.n15086 DVDD.n15085 0.0264781
R2595 DVDD.n7274 DVDD.n7273 0.0264774
R2596 DVDD DVDD.n1089 0.0260195
R2597 DVDD.n11423 DVDD 0.0260195
R2598 DVDD.n1123 DVDD 0.0260195
R2599 DVDD.n1012 DVDD 0.0260192
R2600 DVDD.n1733 DVDD 0.0260192
R2601 DVDD DVDD.n3157 0.026019
R2602 DVDD.n7162 DVDD 0.0260187
R2603 DVDD DVDD.n18287 0.0260158
R2604 DVDD DVDD.n9519 0.0260158
R2605 DVDD.n11916 DVDD 0.0260155
R2606 DVDD DVDD.n1283 0.0260155
R2607 DVDD DVDD.n12323 0.0260155
R2608 DVDD DVDD.n9958 0.0260153
R2609 DVDD.n1545 DVDD 0.0260153
R2610 DVDD DVDD.n1674 0.0260153
R2611 DVDD DVDD.n11541 0.0260153
R2612 DVDD.n3320 DVDD 0.0260153
R2613 DVDD.n9815 DVDD 0.026015
R2614 DVDD.n9906 DVDD.n9905 0.0255541
R2615 DVDD.n9929 DVDD.n7813 0.0253108
R2616 DVDD.n12737 DVDD.n12736 0.0248
R2617 DVDD.n6106 DVDD.n6103 0.0248
R2618 DVDD.n6119 DVDD.n6118 0.0248
R2619 DVDD.n8821 DVDD.n8820 0.0248
R2620 DVDD.n12450 DVDD.n12449 0.0248
R2621 DVDD.n5668 DVDD.n5666 0.0248
R2622 DVDD.n4058 DVDD.n4057 0.0248
R2623 DVDD.n8474 DVDD.n8473 0.0248
R2624 DVDD.n12437 DVDD.n12436 0.0248
R2625 DVDD.n5622 DVDD.n5621 0.0248
R2626 DVDD.n4048 DVDD.n4047 0.0248
R2627 DVDD.n8456 DVDD.n8455 0.0248
R2628 DVDD.n5575 DVDD.n5573 0.0248
R2629 DVDD.n4038 DVDD.n4037 0.0248
R2630 DVDD.n3037 DVDD.n3036 0.024193
R2631 DVDD.n7219 DVDD.n7218 0.024125
R2632 DVDD.n7222 DVDD.n7221 0.024125
R2633 DVDD.n7270 DVDD.n7269 0.024125
R2634 DVDD.n7267 DVDD.n7266 0.024125
R2635 DVDD.n7616 DVDD.n7615 0.024125
R2636 DVDD.n7619 DVDD.n7618 0.024125
R2637 DVDD.n7632 DVDD.n7631 0.024125
R2638 DVDD.n7629 DVDD.n7628 0.024125
R2639 DVDD.n7643 DVDD.n7642 0.024125
R2640 DVDD.n7646 DVDD.n7645 0.024125
R2641 DVDD.n7656 DVDD.n7655 0.024125
R2642 DVDD.n7653 DVDD.n7652 0.024125
R2643 DVDD.n20284 DVDD.n20283 0.024125
R2644 DVDD.n20287 DVDD.n20286 0.024125
R2645 DVDD.n20298 DVDD.n20297 0.024125
R2646 DVDD.n20295 DVDD.n20294 0.024125
R2647 DVDD.n20331 DVDD.n20330 0.024125
R2648 DVDD.n20334 DVDD.n20333 0.024125
R2649 DVDD.n20320 DVDD.n20319 0.024125
R2650 DVDD.n20317 DVDD.n20316 0.024125
R2651 DVDD.n15078 DVDD.n15077 0.024125
R2652 DVDD.n15081 DVDD.n15080 0.024125
R2653 DVDD.n15095 DVDD.n15094 0.024125
R2654 DVDD.n15092 DVDD.n15091 0.024125
R2655 DVDD.n10696 DVDD.n10695 0.024125
R2656 DVDD.n10699 DVDD.n10698 0.024125
R2657 DVDD.n10713 DVDD.n10712 0.024125
R2658 DVDD.n10710 DVDD.n10709 0.024125
R2659 DVDD.n7290 DVDD.n7289 0.024125
R2660 DVDD.n7293 DVDD.n7292 0.024125
R2661 DVDD.n7283 DVDD.n7282 0.024125
R2662 DVDD.n7280 DVDD.n7279 0.024125
R2663 DVDD DVDD.n16349 0.023649
R2664 DVDD.n12463 DVDD.n12462 0.023
R2665 DVDD.n12471 DVDD.n12470 0.023
R2666 DVDD.n5705 DVDD.n5704 0.023
R2667 DVDD.n4554 DVDD.n4553 0.023
R2668 DVDD.n6113 DVDD.n6112 0.023
R2669 DVDD.n4074 DVDD.n4073 0.023
R2670 DVDD.n8488 DVDD.n8487 0.023
R2671 DVDD.n8496 DVDD.n8495 0.023
R2672 DVDD.n12772 DVDD.n12771 0.023
R2673 DVDD.n12457 DVDD.n12456 0.023
R2674 DVDD.n5663 DVDD.n5662 0.023
R2675 DVDD.n4569 DVDD.n4568 0.023
R2676 DVDD.n4561 DVDD.n4560 0.023
R2677 DVDD.n4065 DVDD.n4064 0.023
R2678 DVDD.n8469 DVDD.n8468 0.023
R2679 DVDD.n8481 DVDD.n8480 0.023
R2680 DVDD.n12432 DVDD.n12431 0.023
R2681 DVDD.n12444 DVDD.n12443 0.023
R2682 DVDD.n5617 DVDD.n5616 0.023
R2683 DVDD.n4584 DVDD.n4583 0.023
R2684 DVDD.n4576 DVDD.n4575 0.023
R2685 DVDD.n4055 DVDD.n4054 0.023
R2686 DVDD.n8451 DVDD.n8450 0.023
R2687 DVDD.n8463 DVDD.n8462 0.023
R2688 DVDD.n12413 DVDD.n12412 0.023
R2689 DVDD.n12425 DVDD.n12424 0.023
R2690 DVDD.n5570 DVDD.n5569 0.023
R2691 DVDD.n4599 DVDD.n4598 0.023
R2692 DVDD.n4591 DVDD.n4590 0.023
R2693 DVDD.n4045 DVDD.n4044 0.023
R2694 DVDD.n8433 DVDD.n8432 0.023
R2695 DVDD.n8445 DVDD.n8444 0.023
R2696 DVDD.n1158 DVDD.n1157 0.0224685
R2697 DVDD.n1157 DVDD.n1156 0.0224685
R2698 DVDD.n1156 DVDD.n1155 0.0224685
R2699 DVDD.n1155 DVDD.n1154 0.0224685
R2700 DVDD.n1154 DVDD.n1153 0.0224685
R2701 DVDD.n1153 DVDD.n1152 0.0224685
R2702 DVDD.n1145 DVDD.n1144 0.0224685
R2703 DVDD.n1144 DVDD.n1143 0.0224685
R2704 DVDD.n1143 DVDD.n1142 0.0224685
R2705 DVDD.n1142 DVDD.n1141 0.0224685
R2706 DVDD.n1141 DVDD.n1140 0.0224685
R2707 DVDD.n1140 DVDD.n1139 0.0224685
R2708 DVDD.n1139 DVDD.n1138 0.0224685
R2709 DVDD.n1138 DVDD.n1137 0.0224685
R2710 DVDD.n1137 DVDD.n1136 0.0224685
R2711 DVDD.n1136 DVDD.n1135 0.0224685
R2712 DVDD.n1135 DVDD.n1134 0.0224685
R2713 DVDD.n1134 DVDD.n1133 0.0224685
R2714 DVDD.n1133 DVDD.n1132 0.0224685
R2715 DVDD.n1132 DVDD.n1131 0.0224685
R2716 DVDD.n1131 DVDD.n1130 0.0224685
R2717 DVDD.n1130 DVDD.n1129 0.0224685
R2718 DVDD.n1129 DVDD.n1128 0.0224685
R2719 DVDD.n1128 DVDD.n1127 0.0224685
R2720 DVDD.n1127 DVDD.n1126 0.0224685
R2721 DVDD.n1126 DVDD.n1125 0.0224685
R2722 DVDD.n1125 DVDD.n1124 0.0224685
R2723 DVDD.n1124 DVDD.n1061 0.0224685
R2724 DVDD.n1550 DVDD.n1061 0.0224685
R2725 DVDD.n1558 DVDD.n1557 0.0224685
R2726 DVDD.n1559 DVDD.n1558 0.0224685
R2727 DVDD.n1560 DVDD.n1559 0.0224685
R2728 DVDD.n1561 DVDD.n1560 0.0224685
R2729 DVDD.n1562 DVDD.n1561 0.0224685
R2730 DVDD.n1563 DVDD.n1562 0.0224685
R2731 DVDD.n1643 DVDD.n1642 0.0224685
R2732 DVDD.n1644 DVDD.n1643 0.0224685
R2733 DVDD.n1645 DVDD.n1644 0.0224685
R2734 DVDD.n1646 DVDD.n1645 0.0224685
R2735 DVDD.n1669 DVDD.n1646 0.0224685
R2736 DVDD.n871 DVDD.n870 0.0224685
R2737 DVDD.n11450 DVDD.n11449 0.0224685
R2738 DVDD.n11451 DVDD.n11450 0.0224685
R2739 DVDD.n11452 DVDD.n11451 0.0224685
R2740 DVDD.n11453 DVDD.n11452 0.0224685
R2741 DVDD.n11454 DVDD.n11453 0.0224685
R2742 DVDD.n11455 DVDD.n11454 0.0224685
R2743 DVDD.n11456 DVDD.n11455 0.0224685
R2744 DVDD.n11457 DVDD.n11456 0.0224685
R2745 DVDD.n11458 DVDD.n11457 0.0224685
R2746 DVDD.n11459 DVDD.n11458 0.0224685
R2747 DVDD.n11460 DVDD.n11459 0.0224685
R2748 DVDD.n11461 DVDD.n11460 0.0224685
R2749 DVDD.n11462 DVDD.n11461 0.0224685
R2750 DVDD.n11463 DVDD.n11462 0.0224685
R2751 DVDD.n11464 DVDD.n11463 0.0224685
R2752 DVDD.n11465 DVDD.n11464 0.0224685
R2753 DVDD.n11466 DVDD.n11465 0.0224685
R2754 DVDD.n11513 DVDD.n11512 0.0224685
R2755 DVDD.n11512 DVDD.n11511 0.0224685
R2756 DVDD.n11511 DVDD.n11510 0.0224685
R2757 DVDD.n11510 DVDD.n11509 0.0224685
R2758 DVDD.n11509 DVDD.n11508 0.0224685
R2759 DVDD.n11508 DVDD.n11507 0.0224685
R2760 DVDD.n11507 DVDD.n11506 0.0224685
R2761 DVDD.n11506 DVDD.n11505 0.0224685
R2762 DVDD.n11505 DVDD.n11504 0.0224685
R2763 DVDD.n11504 DVDD.n11503 0.0224685
R2764 DVDD.n11503 DVDD.n11502 0.0224685
R2765 DVDD.n11502 DVDD.n11501 0.0224685
R2766 DVDD.n11501 DVDD.n11500 0.0224685
R2767 DVDD.n11500 DVDD.n11499 0.0224685
R2768 DVDD.n11499 DVDD.n11498 0.0224685
R2769 DVDD.n11498 DVDD.n11497 0.0224685
R2770 DVDD.n11497 DVDD.n11496 0.0224685
R2771 DVDD.n11496 DVDD.n11495 0.0224685
R2772 DVDD.n11495 DVDD.n11494 0.0224685
R2773 DVDD.n11494 DVDD.n11493 0.0224685
R2774 DVDD.n11493 DVDD.n11492 0.0224685
R2775 DVDD.n11492 DVDD.n11491 0.0224685
R2776 DVDD.n11491 DVDD.n11490 0.0224685
R2777 DVDD.n12158 DVDD.n12157 0.0224685
R2778 DVDD.n12276 DVDD.n12275 0.0224685
R2779 DVDD.n12275 DVDD.n12274 0.0224685
R2780 DVDD.n12274 DVDD.n12273 0.0224685
R2781 DVDD.n12273 DVDD.n12272 0.0224685
R2782 DVDD.n12272 DVDD.n12271 0.0224685
R2783 DVDD.n12271 DVDD.n12270 0.0224685
R2784 DVDD.n12270 DVDD.n12269 0.0224685
R2785 DVDD.n12269 DVDD.n12268 0.0224685
R2786 DVDD.n12268 DVDD.n12267 0.0224685
R2787 DVDD.n12267 DVDD.n12266 0.0224685
R2788 DVDD.n12266 DVDD.n12265 0.0224685
R2789 DVDD.n12265 DVDD.n12264 0.0224685
R2790 DVDD.n12264 DVDD.n12263 0.0224685
R2791 DVDD.n12263 DVDD.n12262 0.0224685
R2792 DVDD.n17513 DVDD.n17512 0.0223919
R2793 DVDD.n17512 DVDD.n17509 0.0223919
R2794 DVDD.n17509 DVDD.n17508 0.0223919
R2795 DVDD.n17508 DVDD.n17505 0.0223919
R2796 DVDD.n17492 DVDD.n17489 0.0223919
R2797 DVDD.n17487 DVDD.n17485 0.0223919
R2798 DVDD.n17483 DVDD.n17478 0.0223919
R2799 DVDD.n17476 DVDD.n17473 0.0223919
R2800 DVDD.n17471 DVDD.n17468 0.0223919
R2801 DVDD.n17466 DVDD.n17463 0.0223919
R2802 DVDD.n17258 DVDD.n17257 0.0223919
R2803 DVDD.n17354 DVDD.n17353 0.0223919
R2804 DVDD.n17353 DVDD.n17350 0.0223919
R2805 DVDD.n17350 DVDD.n17349 0.0223919
R2806 DVDD.n17349 DVDD.n17346 0.0223919
R2807 DVDD.n17333 DVDD.n17330 0.0223919
R2808 DVDD.n17328 DVDD.n17326 0.0223919
R2809 DVDD.n17324 DVDD.n17319 0.0223919
R2810 DVDD.n17317 DVDD.n17314 0.0223919
R2811 DVDD.n17312 DVDD.n17309 0.0223919
R2812 DVDD.n17307 DVDD.n17304 0.0223919
R2813 DVDD.n17302 DVDD.n17298 0.0223919
R2814 DVDD.n17286 DVDD.n17284 0.0223919
R2815 DVDD.n17284 DVDD.n17282 0.0223919
R2816 DVDD.n17282 DVDD.n17280 0.0223919
R2817 DVDD.n17280 DVDD.n17278 0.0223919
R2818 DVDD.n17278 DVDD.n17276 0.0223919
R2819 DVDD.n17276 DVDD.n17274 0.0223919
R2820 DVDD.n17274 DVDD.n17272 0.0223919
R2821 DVDD.n17272 DVDD.n17270 0.0223919
R2822 DVDD.n5799 DVDD.n5797 0.0223919
R2823 DVDD.n5803 DVDD.n5799 0.0223919
R2824 DVDD.n5803 DVDD.n5801 0.0223919
R2825 DVDD.n5791 DVDD.n5789 0.0223919
R2826 DVDD.n5795 DVDD.n5791 0.0223919
R2827 DVDD.n5795 DVDD.n5793 0.0223919
R2828 DVDD.n4243 DVDD.n4241 0.0223919
R2829 DVDD.n4232 DVDD.n4230 0.0223919
R2830 DVDD.n4222 DVDD.n4220 0.0223919
R2831 DVDD.n4228 DVDD.n4222 0.0223919
R2832 DVDD.n4228 DVDD.n4226 0.0223919
R2833 DVDD.n4226 DVDD.n4224 0.0223919
R2834 DVDD.n13889 DVDD.n13887 0.0223919
R2835 DVDD.n13891 DVDD.n13889 0.0223919
R2836 DVDD.n13893 DVDD.n13891 0.0223919
R2837 DVDD.n13895 DVDD.n13893 0.0223919
R2838 DVDD.n13897 DVDD.n13895 0.0223919
R2839 DVDD.n13899 DVDD.n13897 0.0223919
R2840 DVDD.n13901 DVDD.n13899 0.0223919
R2841 DVDD.n13903 DVDD.n13901 0.0223919
R2842 DVDD.n14117 DVDD.n14116 0.0223919
R2843 DVDD.n14116 DVDD.n14113 0.0223919
R2844 DVDD.n14113 DVDD.n14112 0.0223919
R2845 DVDD.n14112 DVDD.n14109 0.0223919
R2846 DVDD.n14053 DVDD.n14050 0.0223919
R2847 DVDD.n14048 DVDD.n14046 0.0223919
R2848 DVDD.n14044 DVDD.n14039 0.0223919
R2849 DVDD.n14037 DVDD.n14034 0.0223919
R2850 DVDD.n14032 DVDD.n14029 0.0223919
R2851 DVDD.n14027 DVDD.n14024 0.0223919
R2852 DVDD.n14022 DVDD.n14020 0.0223919
R2853 DVDD.n13977 DVDD.n13976 0.0223919
R2854 DVDD.n13976 DVDD.n13973 0.0223919
R2855 DVDD.n13973 DVDD.n13972 0.0223919
R2856 DVDD.n13972 DVDD.n13969 0.0223919
R2857 DVDD.n13956 DVDD.n13953 0.0223919
R2858 DVDD.n13951 DVDD.n13949 0.0223919
R2859 DVDD.n13947 DVDD.n13942 0.0223919
R2860 DVDD.n13940 DVDD.n13937 0.0223919
R2861 DVDD.n13935 DVDD.n13932 0.0223919
R2862 DVDD.n13930 DVDD.n13927 0.0223919
R2863 DVDD.n13925 DVDD.n13920 0.0223919
R2864 DVDD.n17255 DVDD.n17254 0.0223919
R2865 DVDD.n17254 DVDD.n17251 0.0223919
R2866 DVDD.n17251 DVDD.n17250 0.0223919
R2867 DVDD.n17250 DVDD.n17247 0.0223919
R2868 DVDD.n17449 DVDD.n17446 0.0223919
R2869 DVDD.n17444 DVDD.n17442 0.0223919
R2870 DVDD.n17440 DVDD.n17435 0.0223919
R2871 DVDD.n17433 DVDD.n17430 0.0223919
R2872 DVDD.n17428 DVDD.n17425 0.0223919
R2873 DVDD.n17423 DVDD.n17420 0.0223919
R2874 DVDD.n17418 DVDD.n17415 0.0223919
R2875 DVDD.n14315 DVDD.n14309 0.0223919
R2876 DVDD.n14315 DVDD.n14310 0.0223919
R2877 DVDD.n14270 DVDD.n14269 0.0223919
R2878 DVDD.n14265 DVDD.n14264 0.0223919
R2879 DVDD.n14260 DVDD.n14259 0.0223919
R2880 DVDD.n14256 DVDD.n14250 0.0223919
R2881 DVDD.n14248 DVDD.n14247 0.0223919
R2882 DVDD.n14243 DVDD.n14242 0.0223919
R2883 DVDD.n14238 DVDD.n14235 0.0223919
R2884 DVDD.n14233 DVDD.n14232 0.0223919
R2885 DVDD.n14174 DVDD.n14173 0.0223919
R2886 DVDD.n14173 DVDD.n14172 0.0223919
R2887 DVDD.n14172 DVDD.n14171 0.0223919
R2888 DVDD.n14171 DVDD.n14168 0.0223919
R2889 DVDD.n14152 DVDD.n14151 0.0223919
R2890 DVDD.n14147 DVDD.n14145 0.0223919
R2891 DVDD.n14143 DVDD.n14137 0.0223919
R2892 DVDD.n14135 DVDD.n14132 0.0223919
R2893 DVDD.n14130 DVDD.n14129 0.0223919
R2894 DVDD.n14125 DVDD.n14122 0.0223919
R2895 DVDD.n14120 DVDD.n14119 0.0223919
R2896 DVDD.n17683 DVDD.n17677 0.0223919
R2897 DVDD.n17683 DVDD.n17682 0.0223919
R2898 DVDD.n17638 DVDD.n17637 0.0223919
R2899 DVDD.n17633 DVDD.n17632 0.0223919
R2900 DVDD.n17628 DVDD.n17627 0.0223919
R2901 DVDD.n17624 DVDD.n17617 0.0223919
R2902 DVDD.n17615 DVDD.n17614 0.0223919
R2903 DVDD.n17610 DVDD.n17609 0.0223919
R2904 DVDD.n17605 DVDD.n17604 0.0223919
R2905 DVDD.n17600 DVDD.n17598 0.0223919
R2906 DVDD.n17664 DVDD.n17662 0.0223919
R2907 DVDD.n17662 DVDD.n17660 0.0223919
R2908 DVDD.n17660 DVDD.n17658 0.0223919
R2909 DVDD.n17658 DVDD.n17656 0.0223919
R2910 DVDD.n17656 DVDD.n17654 0.0223919
R2911 DVDD.n17654 DVDD.n17652 0.0223919
R2912 DVDD.n17652 DVDD.n17650 0.0223919
R2913 DVDD.n17650 DVDD.n17648 0.0223919
R2914 DVDD.n5779 DVDD.n5773 0.0223919
R2915 DVDD.n5779 DVDD.n5777 0.0223919
R2916 DVDD.n5777 DVDD.n5775 0.0223919
R2917 DVDD.n5787 DVDD.n5781 0.0223919
R2918 DVDD.n5787 DVDD.n5785 0.0223919
R2919 DVDD.n5785 DVDD.n5783 0.0223919
R2920 DVDD.n4345 DVDD.n4343 0.0223919
R2921 DVDD.n4343 DVDD.n4341 0.0223919
R2922 DVDD.n4341 DVDD.n4339 0.0223919
R2923 DVDD.n4170 DVDD.n4168 0.0223919
R2924 DVDD.n4176 DVDD.n4170 0.0223919
R2925 DVDD.n4176 DVDD.n4174 0.0223919
R2926 DVDD.n4174 DVDD.n4172 0.0223919
R2927 DVDD.n14277 DVDD.n14275 0.0223919
R2928 DVDD.n14279 DVDD.n14277 0.0223919
R2929 DVDD.n14281 DVDD.n14279 0.0223919
R2930 DVDD.n14283 DVDD.n14281 0.0223919
R2931 DVDD.n14285 DVDD.n14283 0.0223919
R2932 DVDD.n14287 DVDD.n14285 0.0223919
R2933 DVDD.n14289 DVDD.n14287 0.0223919
R2934 DVDD.n14291 DVDD.n14289 0.0223919
R2935 DVDD.n13372 DVDD.n13371 0.0222913
R2936 DVDD.n7302 DVDD.n7301 0.0222662
R2937 DVDD.n13371 DVDD.n13370 0.021937
R2938 DVDD.n10076 DVDD.n10075 0.021875
R2939 DVDD.n1812 DVDD.n1811 0.021875
R2940 DVDD.n18996 DVDD.n18995 0.02165
R2941 DVDD.n3842 DVDD.n3841 0.02165
R2942 DVDD.n127 DVDD.n126 0.02165
R2943 DVDD.n10599 DVDD.n10598 0.02165
R2944 DVDD.n19148 DVDD.n19147 0.021425
R2945 DVDD.n10610 DVDD.n10609 0.021425
R2946 DVDD.n12157 DVDD.n12156 0.0212283
R2947 DVDD.n12277 DVDD.n12276 0.0210512
R2948 DVDD.n19156 DVDD.n19155 0.02075
R2949 DVDD.n10618 DVDD.n10617 0.02075
R2950 DVDD.n20290 DVDD.n0 0.0205764
R2951 DVDD.n3850 DVDD.n3849 0.020525
R2952 DVDD.n135 DVDD.n134 0.020525
R2953 DVDD.n15984 DVDD.n15983 0.0202699
R2954 DVDD.n15980 DVDD.n15979 0.0202699
R2955 DVDD.n15969 DVDD.n15968 0.0202699
R2956 DVDD.n15965 DVDD.n15964 0.0202699
R2957 DVDD.n15956 DVDD.n15955 0.0202699
R2958 DVDD.n15943 DVDD.n15942 0.0202699
R2959 DVDD.n15947 DVDD.n15946 0.0202699
R2960 DVDD.n16066 DVDD.n16065 0.0202699
R2961 DVDD.n16062 DVDD.n16061 0.0202699
R2962 DVDD.n16058 DVDD.n16057 0.0202699
R2963 DVDD.n16049 DVDD.n16048 0.0202699
R2964 DVDD.n16045 DVDD.n16044 0.0202699
R2965 DVDD.n16036 DVDD.n16035 0.0202699
R2966 DVDD.n16032 DVDD.n16031 0.0202699
R2967 DVDD.n16019 DVDD.n16018 0.0202699
R2968 DVDD.n16015 DVDD.n16014 0.0202699
R2969 DVDD.n16006 DVDD.n16005 0.0202699
R2970 DVDD.n16002 DVDD.n16001 0.0202699
R2971 DVDD.n15683 DVDD.n15682 0.0202699
R2972 DVDD.n15687 DVDD.n15686 0.0202699
R2973 DVDD.n15678 DVDD.n15677 0.0202699
R2974 DVDD.n15674 DVDD.n15673 0.0202699
R2975 DVDD.n15670 DVDD.n15669 0.0202699
R2976 DVDD.n15661 DVDD.n15660 0.0202699
R2977 DVDD.n15657 DVDD.n15656 0.0202699
R2978 DVDD.n15648 DVDD.n15647 0.0202699
R2979 DVDD.n15644 DVDD.n15643 0.0202699
R2980 DVDD.n15631 DVDD.n15630 0.0202699
R2981 DVDD.n15627 DVDD.n15626 0.0202699
R2982 DVDD.n15926 DVDD.n15925 0.0202699
R2983 DVDD.n15930 DVDD.n15929 0.0202699
R2984 DVDD.n8164 DVDD.n8163 0.0202699
R2985 DVDD.n8160 DVDD.n8159 0.0202699
R2986 DVDD.n8151 DVDD.n8150 0.0202699
R2987 DVDD.n8147 DVDD.n8146 0.0202699
R2988 DVDD.n8143 DVDD.n8142 0.0202699
R2989 DVDD.n9412 DVDD.n9411 0.0202699
R2990 DVDD.n9405 DVDD.n9404 0.0202699
R2991 DVDD.n9401 DVDD.n9400 0.0202699
R2992 DVDD.n8128 DVDD.n8127 0.0202699
R2993 DVDD.n8132 DVDD.n8131 0.0202699
R2994 DVDD.n9899 DVDD.n9898 0.0202699
R2995 DVDD.n9895 DVDD.n9894 0.0202699
R2996 DVDD.n15976 DVDD.n15975 0.0200816
R2997 DVDD.n8121 DVDD.n8120 0.0200816
R2998 DVDD DVDD.n7297 0.0200421
R2999 DVDD.n10080 DVDD.n10079 0.01985
R3000 DVDD.n1816 DVDD.n1815 0.01985
R3001 DVDD.n14316 DVDD.n14271 0.0196339
R3002 DVDD.n14271 DVDD.n14266 0.0196339
R3003 DVDD.n14266 DVDD.n14261 0.0196339
R3004 DVDD.n14261 DVDD.n14257 0.0196339
R3005 DVDD.n14257 DVDD.n14249 0.0196339
R3006 DVDD.n14249 DVDD.n14244 0.0196339
R3007 DVDD.n14244 DVDD.n14239 0.0196339
R3008 DVDD.n14239 DVDD.n14234 0.0196339
R3009 DVDD.n14155 DVDD.n14154 0.0196339
R3010 DVDD.n14154 DVDD.n14153 0.0196339
R3011 DVDD.n14153 DVDD.n14148 0.0196339
R3012 DVDD.n14148 DVDD.n14144 0.0196339
R3013 DVDD.n14144 DVDD.n14136 0.0196339
R3014 DVDD.n14136 DVDD.n14131 0.0196339
R3015 DVDD.n14131 DVDD.n14126 0.0196339
R3016 DVDD.n14126 DVDD.n14121 0.0196339
R3017 DVDD.n14056 DVDD.n14055 0.0196339
R3018 DVDD.n14055 DVDD.n14054 0.0196339
R3019 DVDD.n14054 DVDD.n14049 0.0196339
R3020 DVDD.n14049 DVDD.n14045 0.0196339
R3021 DVDD.n14045 DVDD.n14038 0.0196339
R3022 DVDD.n14038 DVDD.n14033 0.0196339
R3023 DVDD.n14033 DVDD.n14028 0.0196339
R3024 DVDD.n14028 DVDD.n14023 0.0196339
R3025 DVDD.n13959 DVDD.n13958 0.0196339
R3026 DVDD.n13958 DVDD.n13957 0.0196339
R3027 DVDD.n13957 DVDD.n13952 0.0196339
R3028 DVDD.n13952 DVDD.n13948 0.0196339
R3029 DVDD.n13948 DVDD.n13941 0.0196339
R3030 DVDD.n13941 DVDD.n13936 0.0196339
R3031 DVDD.n13936 DVDD.n13931 0.0196339
R3032 DVDD.n13931 DVDD.n13926 0.0196339
R3033 DVDD.n19761 DVDD.n19760 0.0196339
R3034 DVDD.n19762 DVDD.n19761 0.0196339
R3035 DVDD.n19763 DVDD.n19762 0.0196339
R3036 DVDD.n19764 DVDD.n19763 0.0196339
R3037 DVDD.n19765 DVDD.n19764 0.0196339
R3038 DVDD.n19766 DVDD.n19765 0.0196339
R3039 DVDD.n19767 DVDD.n19766 0.0196339
R3040 DVDD.n19775 DVDD.n19774 0.0196339
R3041 DVDD.n19776 DVDD.n19775 0.0196339
R3042 DVDD.n19777 DVDD.n19776 0.0196339
R3043 DVDD.n19778 DVDD.n19777 0.0196339
R3044 DVDD.n19779 DVDD.n19778 0.0196339
R3045 DVDD.n19780 DVDD.n19779 0.0196339
R3046 DVDD.n19781 DVDD.n19780 0.0196339
R3047 DVDD.n19782 DVDD.n19781 0.0196339
R3048 DVDD.n19783 DVDD.n19782 0.0196339
R3049 DVDD.n19784 DVDD.n19783 0.0196339
R3050 DVDD.n19785 DVDD.n19784 0.0196339
R3051 DVDD.n19786 DVDD.n19785 0.0196339
R3052 DVDD.n19787 DVDD.n19786 0.0196339
R3053 DVDD.n19788 DVDD.n19787 0.0196339
R3054 DVDD.n19789 DVDD.n19788 0.0196339
R3055 DVDD.n19790 DVDD.n19789 0.0196339
R3056 DVDD.n19791 DVDD.n19790 0.0196339
R3057 DVDD.n19792 DVDD.n19791 0.0196339
R3058 DVDD.n19793 DVDD.n19792 0.0196339
R3059 DVDD.n19794 DVDD.n19793 0.0196339
R3060 DVDD.n19795 DVDD.n19794 0.0196339
R3061 DVDD.n19796 DVDD.n19795 0.0196339
R3062 DVDD.n19797 DVDD.n19796 0.0196339
R3063 DVDD.n19798 DVDD.n19797 0.0196339
R3064 DVDD.n19799 DVDD.n19798 0.0196339
R3065 DVDD.n19837 DVDD.n19799 0.0196339
R3066 DVDD.n19845 DVDD.n19844 0.0196339
R3067 DVDD.n19846 DVDD.n19845 0.0196339
R3068 DVDD.n19847 DVDD.n19846 0.0196339
R3069 DVDD.n19848 DVDD.n19847 0.0196339
R3070 DVDD.n19849 DVDD.n19848 0.0196339
R3071 DVDD.n19850 DVDD.n19849 0.0196339
R3072 DVDD.n19851 DVDD.n19850 0.0196339
R3073 DVDD.n19928 DVDD.n19927 0.0196339
R3074 DVDD.n19929 DVDD.n19928 0.0196339
R3075 DVDD.n19930 DVDD.n19929 0.0196339
R3076 DVDD.n19931 DVDD.n19930 0.0196339
R3077 DVDD.n19932 DVDD.n19931 0.0196339
R3078 DVDD.n19992 DVDD.n19932 0.0196339
R3079 DVDD.n20178 DVDD.n20177 0.0196339
R3080 DVDD.n4684 DVDD.n4683 0.0196339
R3081 DVDD.n4685 DVDD.n4684 0.0196339
R3082 DVDD.n4686 DVDD.n4685 0.0196339
R3083 DVDD.n4687 DVDD.n4686 0.0196339
R3084 DVDD.n4688 DVDD.n4687 0.0196339
R3085 DVDD.n4689 DVDD.n4688 0.0196339
R3086 DVDD.n4690 DVDD.n4689 0.0196339
R3087 DVDD.n4691 DVDD.n4690 0.0196339
R3088 DVDD.n4692 DVDD.n4691 0.0196339
R3089 DVDD.n4693 DVDD.n4692 0.0196339
R3090 DVDD.n4694 DVDD.n4693 0.0196339
R3091 DVDD.n4695 DVDD.n4694 0.0196339
R3092 DVDD.n4696 DVDD.n4695 0.0196339
R3093 DVDD.n4697 DVDD.n4696 0.0196339
R3094 DVDD.n4698 DVDD.n4697 0.0196339
R3095 DVDD.n4699 DVDD.n4698 0.0196339
R3096 DVDD.n4700 DVDD.n4699 0.0196339
R3097 DVDD.n4701 DVDD.n4700 0.0196339
R3098 DVDD.n4702 DVDD.n4701 0.0196339
R3099 DVDD.n4703 DVDD.n4702 0.0196339
R3100 DVDD.n4748 DVDD.n4747 0.0196339
R3101 DVDD.n4749 DVDD.n4748 0.0196339
R3102 DVDD.n4750 DVDD.n4749 0.0196339
R3103 DVDD.n4751 DVDD.n4750 0.0196339
R3104 DVDD.n4752 DVDD.n4751 0.0196339
R3105 DVDD.n4753 DVDD.n4752 0.0196339
R3106 DVDD.n4754 DVDD.n4753 0.0196339
R3107 DVDD.n4755 DVDD.n4754 0.0196339
R3108 DVDD.n4756 DVDD.n4755 0.0196339
R3109 DVDD.n4757 DVDD.n4756 0.0196339
R3110 DVDD.n4758 DVDD.n4757 0.0196339
R3111 DVDD.n4759 DVDD.n4758 0.0196339
R3112 DVDD.n4760 DVDD.n4759 0.0196339
R3113 DVDD.n4761 DVDD.n4760 0.0196339
R3114 DVDD.n4762 DVDD.n4761 0.0196339
R3115 DVDD.n4763 DVDD.n4762 0.0196339
R3116 DVDD.n4764 DVDD.n4763 0.0196339
R3117 DVDD.n4765 DVDD.n4764 0.0196339
R3118 DVDD.n4766 DVDD.n4765 0.0196339
R3119 DVDD.n4767 DVDD.n4766 0.0196339
R3120 DVDD.n4768 DVDD.n4767 0.0196339
R3121 DVDD.n4769 DVDD.n4768 0.0196339
R3122 DVDD.n4770 DVDD.n4769 0.0196339
R3123 DVDD.n4771 DVDD.n4770 0.0196339
R3124 DVDD.n4772 DVDD.n4771 0.0196339
R3125 DVDD.n4773 DVDD.n4772 0.0196339
R3126 DVDD.n5012 DVDD.n5011 0.0196339
R3127 DVDD.n5013 DVDD.n5012 0.0196339
R3128 DVDD.n5068 DVDD.n5067 0.0196339
R3129 DVDD.n5069 DVDD.n5068 0.0196339
R3130 DVDD.n5070 DVDD.n5069 0.0196339
R3131 DVDD.n5071 DVDD.n5070 0.0196339
R3132 DVDD.n5072 DVDD.n5071 0.0196339
R3133 DVDD.n5073 DVDD.n5072 0.0196339
R3134 DVDD.n5074 DVDD.n5073 0.0196339
R3135 DVDD.n5075 DVDD.n5074 0.0196339
R3136 DVDD.n5076 DVDD.n5075 0.0196339
R3137 DVDD.n5077 DVDD.n5076 0.0196339
R3138 DVDD.n5078 DVDD.n5077 0.0196339
R3139 DVDD.n5079 DVDD.n5078 0.0196339
R3140 DVDD.n5080 DVDD.n5079 0.0196339
R3141 DVDD.n5081 DVDD.n5080 0.0196339
R3142 DVDD.n5082 DVDD.n5081 0.0196339
R3143 DVDD.n5083 DVDD.n5082 0.0196339
R3144 DVDD.n5084 DVDD.n5083 0.0196339
R3145 DVDD.n5361 DVDD.n5360 0.0196339
R3146 DVDD.n5362 DVDD.n5361 0.0196339
R3147 DVDD.n1406 DVDD.n1405 0.0196339
R3148 DVDD.n1407 DVDD.n1406 0.0196339
R3149 DVDD.n1408 DVDD.n1407 0.0196339
R3150 DVDD.n1409 DVDD.n1408 0.0196339
R3151 DVDD.n1410 DVDD.n1409 0.0196339
R3152 DVDD.n1411 DVDD.n1410 0.0196339
R3153 DVDD.n1412 DVDD.n1411 0.0196339
R3154 DVDD.n1420 DVDD.n1419 0.0196339
R3155 DVDD.n1421 DVDD.n1420 0.0196339
R3156 DVDD.n1422 DVDD.n1421 0.0196339
R3157 DVDD.n1423 DVDD.n1422 0.0196339
R3158 DVDD.n1424 DVDD.n1423 0.0196339
R3159 DVDD.n1425 DVDD.n1424 0.0196339
R3160 DVDD.n1426 DVDD.n1425 0.0196339
R3161 DVDD.n1427 DVDD.n1426 0.0196339
R3162 DVDD.n1428 DVDD.n1427 0.0196339
R3163 DVDD.n1429 DVDD.n1428 0.0196339
R3164 DVDD.n1430 DVDD.n1429 0.0196339
R3165 DVDD.n1431 DVDD.n1430 0.0196339
R3166 DVDD.n1432 DVDD.n1431 0.0196339
R3167 DVDD.n1433 DVDD.n1432 0.0196339
R3168 DVDD.n1434 DVDD.n1433 0.0196339
R3169 DVDD.n1435 DVDD.n1434 0.0196339
R3170 DVDD.n1436 DVDD.n1435 0.0196339
R3171 DVDD.n1437 DVDD.n1436 0.0196339
R3172 DVDD.n1438 DVDD.n1437 0.0196339
R3173 DVDD.n1439 DVDD.n1438 0.0196339
R3174 DVDD.n1440 DVDD.n1439 0.0196339
R3175 DVDD.n1441 DVDD.n1440 0.0196339
R3176 DVDD.n1442 DVDD.n1441 0.0196339
R3177 DVDD.n1443 DVDD.n1442 0.0196339
R3178 DVDD.n1444 DVDD.n1443 0.0196339
R3179 DVDD.n1538 DVDD.n1444 0.0196339
R3180 DVDD.n1531 DVDD.n1530 0.0196339
R3181 DVDD.n1530 DVDD.n1529 0.0196339
R3182 DVDD.n1529 DVDD.n1528 0.0196339
R3183 DVDD.n1528 DVDD.n1527 0.0196339
R3184 DVDD.n1527 DVDD.n1526 0.0196339
R3185 DVDD.n1526 DVDD.n1525 0.0196339
R3186 DVDD.n1525 DVDD.n1524 0.0196339
R3187 DVDD.n1449 DVDD.n1448 0.0196339
R3188 DVDD.n1448 DVDD.n1447 0.0196339
R3189 DVDD.n1447 DVDD.n1446 0.0196339
R3190 DVDD.n1446 DVDD.n1445 0.0196339
R3191 DVDD.n1445 DVDD.n957 0.0196339
R3192 DVDD.n1680 DVDD.n957 0.0196339
R3193 DVDD.n256 DVDD.n255 0.0196339
R3194 DVDD.n11391 DVDD.n11390 0.0196339
R3195 DVDD.n11392 DVDD.n11391 0.0196339
R3196 DVDD.n11393 DVDD.n11392 0.0196339
R3197 DVDD.n11394 DVDD.n11393 0.0196339
R3198 DVDD.n11395 DVDD.n11394 0.0196339
R3199 DVDD.n11396 DVDD.n11395 0.0196339
R3200 DVDD.n11397 DVDD.n11396 0.0196339
R3201 DVDD.n11398 DVDD.n11397 0.0196339
R3202 DVDD.n11399 DVDD.n11398 0.0196339
R3203 DVDD.n11400 DVDD.n11399 0.0196339
R3204 DVDD.n11401 DVDD.n11400 0.0196339
R3205 DVDD.n11402 DVDD.n11401 0.0196339
R3206 DVDD.n11403 DVDD.n11402 0.0196339
R3207 DVDD.n11404 DVDD.n11403 0.0196339
R3208 DVDD.n11405 DVDD.n11404 0.0196339
R3209 DVDD.n11406 DVDD.n11405 0.0196339
R3210 DVDD.n11407 DVDD.n11406 0.0196339
R3211 DVDD.n11408 DVDD.n11407 0.0196339
R3212 DVDD.n11409 DVDD.n11408 0.0196339
R3213 DVDD.n11410 DVDD.n11409 0.0196339
R3214 DVDD.n11574 DVDD.n11573 0.0196339
R3215 DVDD.n11575 DVDD.n11574 0.0196339
R3216 DVDD.n11576 DVDD.n11575 0.0196339
R3217 DVDD.n11577 DVDD.n11576 0.0196339
R3218 DVDD.n11578 DVDD.n11577 0.0196339
R3219 DVDD.n11579 DVDD.n11578 0.0196339
R3220 DVDD.n11580 DVDD.n11579 0.0196339
R3221 DVDD.n11581 DVDD.n11580 0.0196339
R3222 DVDD.n11582 DVDD.n11581 0.0196339
R3223 DVDD.n11583 DVDD.n11582 0.0196339
R3224 DVDD.n11584 DVDD.n11583 0.0196339
R3225 DVDD.n11585 DVDD.n11584 0.0196339
R3226 DVDD.n11586 DVDD.n11585 0.0196339
R3227 DVDD.n11587 DVDD.n11586 0.0196339
R3228 DVDD.n11588 DVDD.n11587 0.0196339
R3229 DVDD.n11589 DVDD.n11588 0.0196339
R3230 DVDD.n11590 DVDD.n11589 0.0196339
R3231 DVDD.n11591 DVDD.n11590 0.0196339
R3232 DVDD.n11592 DVDD.n11591 0.0196339
R3233 DVDD.n11593 DVDD.n11592 0.0196339
R3234 DVDD.n11594 DVDD.n11593 0.0196339
R3235 DVDD.n11595 DVDD.n11594 0.0196339
R3236 DVDD.n11596 DVDD.n11595 0.0196339
R3237 DVDD.n11597 DVDD.n11596 0.0196339
R3238 DVDD.n11598 DVDD.n11597 0.0196339
R3239 DVDD.n11599 DVDD.n11598 0.0196339
R3240 DVDD.n11742 DVDD.n11741 0.0196339
R3241 DVDD.n11741 DVDD.n11740 0.0196339
R3242 DVDD.n11686 DVDD.n11685 0.0196339
R3243 DVDD.n11685 DVDD.n11684 0.0196339
R3244 DVDD.n11684 DVDD.n11683 0.0196339
R3245 DVDD.n11683 DVDD.n11682 0.0196339
R3246 DVDD.n11682 DVDD.n11681 0.0196339
R3247 DVDD.n11681 DVDD.n11680 0.0196339
R3248 DVDD.n11680 DVDD.n11679 0.0196339
R3249 DVDD.n11679 DVDD.n11678 0.0196339
R3250 DVDD.n11678 DVDD.n11677 0.0196339
R3251 DVDD.n11677 DVDD.n11676 0.0196339
R3252 DVDD.n11676 DVDD.n11675 0.0196339
R3253 DVDD.n11675 DVDD.n11674 0.0196339
R3254 DVDD.n11674 DVDD.n11673 0.0196339
R3255 DVDD.n11673 DVDD.n11672 0.0196339
R3256 DVDD.n11672 DVDD.n11671 0.0196339
R3257 DVDD.n11671 DVDD.n11670 0.0196339
R3258 DVDD.n11670 DVDD.n11669 0.0196339
R3259 DVDD.n13099 DVDD.n13098 0.0196339
R3260 DVDD.n13098 DVDD.n13097 0.0196339
R3261 DVDD.n17684 DVDD.n17639 0.0196339
R3262 DVDD.n17639 DVDD.n17634 0.0196339
R3263 DVDD.n17634 DVDD.n17629 0.0196339
R3264 DVDD.n17629 DVDD.n17625 0.0196339
R3265 DVDD.n17625 DVDD.n17616 0.0196339
R3266 DVDD.n17616 DVDD.n17611 0.0196339
R3267 DVDD.n17611 DVDD.n17606 0.0196339
R3268 DVDD.n17606 DVDD.n17601 0.0196339
R3269 DVDD.n17495 DVDD.n17494 0.0196339
R3270 DVDD.n17494 DVDD.n17493 0.0196339
R3271 DVDD.n17493 DVDD.n17488 0.0196339
R3272 DVDD.n17488 DVDD.n17484 0.0196339
R3273 DVDD.n17484 DVDD.n17477 0.0196339
R3274 DVDD.n17477 DVDD.n17472 0.0196339
R3275 DVDD.n17472 DVDD.n17467 0.0196339
R3276 DVDD.n17467 DVDD.n17462 0.0196339
R3277 DVDD.n17452 DVDD.n17451 0.0196339
R3278 DVDD.n17451 DVDD.n17450 0.0196339
R3279 DVDD.n17450 DVDD.n17445 0.0196339
R3280 DVDD.n17445 DVDD.n17441 0.0196339
R3281 DVDD.n17441 DVDD.n17434 0.0196339
R3282 DVDD.n17434 DVDD.n17429 0.0196339
R3283 DVDD.n17429 DVDD.n17424 0.0196339
R3284 DVDD.n17424 DVDD.n17419 0.0196339
R3285 DVDD.n17336 DVDD.n17335 0.0196339
R3286 DVDD.n17335 DVDD.n17334 0.0196339
R3287 DVDD.n17334 DVDD.n17329 0.0196339
R3288 DVDD.n17329 DVDD.n17325 0.0196339
R3289 DVDD.n17325 DVDD.n17318 0.0196339
R3290 DVDD.n17318 DVDD.n17313 0.0196339
R3291 DVDD.n17313 DVDD.n17308 0.0196339
R3292 DVDD.n17308 DVDD.n17303 0.0196339
R3293 DVDD.n1983 DVDD.n1982 0.0196339
R3294 DVDD.n1984 DVDD.n1983 0.0196339
R3295 DVDD.n1985 DVDD.n1984 0.0196339
R3296 DVDD.n1986 DVDD.n1985 0.0196339
R3297 DVDD.n1987 DVDD.n1986 0.0196339
R3298 DVDD.n1988 DVDD.n1987 0.0196339
R3299 DVDD.n1989 DVDD.n1988 0.0196339
R3300 DVDD.n1997 DVDD.n1996 0.0196339
R3301 DVDD.n1998 DVDD.n1997 0.0196339
R3302 DVDD.n1999 DVDD.n1998 0.0196339
R3303 DVDD.n2000 DVDD.n1999 0.0196339
R3304 DVDD.n2001 DVDD.n2000 0.0196339
R3305 DVDD.n2002 DVDD.n2001 0.0196339
R3306 DVDD.n2003 DVDD.n2002 0.0196339
R3307 DVDD.n2004 DVDD.n2003 0.0196339
R3308 DVDD.n2005 DVDD.n2004 0.0196339
R3309 DVDD.n2006 DVDD.n2005 0.0196339
R3310 DVDD.n2007 DVDD.n2006 0.0196339
R3311 DVDD.n2008 DVDD.n2007 0.0196339
R3312 DVDD.n2009 DVDD.n2008 0.0196339
R3313 DVDD.n2010 DVDD.n2009 0.0196339
R3314 DVDD.n2011 DVDD.n2010 0.0196339
R3315 DVDD.n2012 DVDD.n2011 0.0196339
R3316 DVDD.n2013 DVDD.n2012 0.0196339
R3317 DVDD.n2014 DVDD.n2013 0.0196339
R3318 DVDD.n2015 DVDD.n2014 0.0196339
R3319 DVDD.n2016 DVDD.n2015 0.0196339
R3320 DVDD.n2017 DVDD.n2016 0.0196339
R3321 DVDD.n2018 DVDD.n2017 0.0196339
R3322 DVDD.n2019 DVDD.n2018 0.0196339
R3323 DVDD.n2020 DVDD.n2019 0.0196339
R3324 DVDD.n2021 DVDD.n2020 0.0196339
R3325 DVDD.n2059 DVDD.n2021 0.0196339
R3326 DVDD.n2067 DVDD.n2066 0.0196339
R3327 DVDD.n2068 DVDD.n2067 0.0196339
R3328 DVDD.n2069 DVDD.n2068 0.0196339
R3329 DVDD.n2070 DVDD.n2069 0.0196339
R3330 DVDD.n2071 DVDD.n2070 0.0196339
R3331 DVDD.n2072 DVDD.n2071 0.0196339
R3332 DVDD.n2073 DVDD.n2072 0.0196339
R3333 DVDD.n2149 DVDD.n2148 0.0196339
R3334 DVDD.n2150 DVDD.n2149 0.0196339
R3335 DVDD.n2151 DVDD.n2150 0.0196339
R3336 DVDD.n2152 DVDD.n2151 0.0196339
R3337 DVDD.n2153 DVDD.n2152 0.0196339
R3338 DVDD.n2213 DVDD.n2153 0.0196339
R3339 DVDD.n19563 DVDD.n19562 0.0196339
R3340 DVDD.n7000 DVDD.n6999 0.0196339
R3341 DVDD.n6999 DVDD.n6998 0.0196339
R3342 DVDD.n6998 DVDD.n6997 0.0196339
R3343 DVDD.n6997 DVDD.n6996 0.0196339
R3344 DVDD.n6996 DVDD.n6995 0.0196339
R3345 DVDD.n6995 DVDD.n6994 0.0196339
R3346 DVDD.n6994 DVDD.n6993 0.0196339
R3347 DVDD.n6993 DVDD.n6992 0.0196339
R3348 DVDD.n6992 DVDD.n6991 0.0196339
R3349 DVDD.n6991 DVDD.n6990 0.0196339
R3350 DVDD.n6990 DVDD.n6989 0.0196339
R3351 DVDD.n6989 DVDD.n6988 0.0196339
R3352 DVDD.n6988 DVDD.n6987 0.0196339
R3353 DVDD.n6987 DVDD.n6986 0.0196339
R3354 DVDD.n6986 DVDD.n6985 0.0196339
R3355 DVDD.n6985 DVDD.n6984 0.0196339
R3356 DVDD.n6984 DVDD.n6983 0.0196339
R3357 DVDD.n6983 DVDD.n6982 0.0196339
R3358 DVDD.n6982 DVDD.n6981 0.0196339
R3359 DVDD.n6981 DVDD.n6980 0.0196339
R3360 DVDD.n6973 DVDD.n6935 0.0196339
R3361 DVDD.n6935 DVDD.n6934 0.0196339
R3362 DVDD.n6934 DVDD.n6933 0.0196339
R3363 DVDD.n6933 DVDD.n6932 0.0196339
R3364 DVDD.n6932 DVDD.n6931 0.0196339
R3365 DVDD.n6931 DVDD.n6930 0.0196339
R3366 DVDD.n6930 DVDD.n6929 0.0196339
R3367 DVDD.n6929 DVDD.n6928 0.0196339
R3368 DVDD.n6928 DVDD.n6927 0.0196339
R3369 DVDD.n6927 DVDD.n6926 0.0196339
R3370 DVDD.n6926 DVDD.n6925 0.0196339
R3371 DVDD.n6925 DVDD.n6924 0.0196339
R3372 DVDD.n6924 DVDD.n6923 0.0196339
R3373 DVDD.n6923 DVDD.n6922 0.0196339
R3374 DVDD.n6922 DVDD.n6921 0.0196339
R3375 DVDD.n6921 DVDD.n6920 0.0196339
R3376 DVDD.n6920 DVDD.n6919 0.0196339
R3377 DVDD.n6919 DVDD.n6918 0.0196339
R3378 DVDD.n6918 DVDD.n6917 0.0196339
R3379 DVDD.n6917 DVDD.n6916 0.0196339
R3380 DVDD.n6916 DVDD.n6915 0.0196339
R3381 DVDD.n6915 DVDD.n6914 0.0196339
R3382 DVDD.n6914 DVDD.n6913 0.0196339
R3383 DVDD.n6913 DVDD.n6912 0.0196339
R3384 DVDD.n6912 DVDD.n6911 0.0196339
R3385 DVDD.n6911 DVDD.n6910 0.0196339
R3386 DVDD.n6672 DVDD.n6671 0.0196339
R3387 DVDD.n6671 DVDD.n6670 0.0196339
R3388 DVDD.n6614 DVDD.n6613 0.0196339
R3389 DVDD.n6613 DVDD.n6612 0.0196339
R3390 DVDD.n6612 DVDD.n6611 0.0196339
R3391 DVDD.n6611 DVDD.n6610 0.0196339
R3392 DVDD.n6610 DVDD.n6609 0.0196339
R3393 DVDD.n6609 DVDD.n6608 0.0196339
R3394 DVDD.n6608 DVDD.n6607 0.0196339
R3395 DVDD.n6607 DVDD.n6606 0.0196339
R3396 DVDD.n6606 DVDD.n6605 0.0196339
R3397 DVDD.n6605 DVDD.n6604 0.0196339
R3398 DVDD.n6604 DVDD.n6603 0.0196339
R3399 DVDD.n6603 DVDD.n6602 0.0196339
R3400 DVDD.n6602 DVDD.n6601 0.0196339
R3401 DVDD.n6601 DVDD.n6600 0.0196339
R3402 DVDD.n6600 DVDD.n6599 0.0196339
R3403 DVDD.n6599 DVDD.n6598 0.0196339
R3404 DVDD.n6598 DVDD.n6597 0.0196339
R3405 DVDD.n6400 DVDD.n6399 0.0196339
R3406 DVDD.n6399 DVDD.n6398 0.0196339
R3407 DVDD.n3197 DVDD.n3196 0.0196339
R3408 DVDD.n3196 DVDD.n3195 0.0196339
R3409 DVDD.n3195 DVDD.n3194 0.0196339
R3410 DVDD.n3194 DVDD.n3193 0.0196339
R3411 DVDD.n3193 DVDD.n3192 0.0196339
R3412 DVDD.n3192 DVDD.n3191 0.0196339
R3413 DVDD.n3191 DVDD.n3190 0.0196339
R3414 DVDD.n3183 DVDD.n3182 0.0196339
R3415 DVDD.n3182 DVDD.n3181 0.0196339
R3416 DVDD.n3181 DVDD.n3180 0.0196339
R3417 DVDD.n3180 DVDD.n3179 0.0196339
R3418 DVDD.n3179 DVDD.n3178 0.0196339
R3419 DVDD.n3178 DVDD.n3177 0.0196339
R3420 DVDD.n3177 DVDD.n3176 0.0196339
R3421 DVDD.n3176 DVDD.n3175 0.0196339
R3422 DVDD.n3175 DVDD.n3174 0.0196339
R3423 DVDD.n3174 DVDD.n3173 0.0196339
R3424 DVDD.n3173 DVDD.n3172 0.0196339
R3425 DVDD.n3172 DVDD.n3171 0.0196339
R3426 DVDD.n3171 DVDD.n3170 0.0196339
R3427 DVDD.n3170 DVDD.n3169 0.0196339
R3428 DVDD.n3169 DVDD.n3168 0.0196339
R3429 DVDD.n3168 DVDD.n3167 0.0196339
R3430 DVDD.n3167 DVDD.n3166 0.0196339
R3431 DVDD.n3166 DVDD.n3165 0.0196339
R3432 DVDD.n3165 DVDD.n3164 0.0196339
R3433 DVDD.n3164 DVDD.n3163 0.0196339
R3434 DVDD.n3163 DVDD.n3162 0.0196339
R3435 DVDD.n3162 DVDD.n3161 0.0196339
R3436 DVDD.n3161 DVDD.n3160 0.0196339
R3437 DVDD.n3160 DVDD.n3159 0.0196339
R3438 DVDD.n3159 DVDD.n2969 0.0196339
R3439 DVDD.n3458 DVDD.n2969 0.0196339
R3440 DVDD.n3466 DVDD.n3465 0.0196339
R3441 DVDD.n3467 DVDD.n3466 0.0196339
R3442 DVDD.n3468 DVDD.n3467 0.0196339
R3443 DVDD.n3469 DVDD.n3468 0.0196339
R3444 DVDD.n3470 DVDD.n3469 0.0196339
R3445 DVDD.n3471 DVDD.n3470 0.0196339
R3446 DVDD.n3472 DVDD.n3471 0.0196339
R3447 DVDD.n3548 DVDD.n3547 0.0196339
R3448 DVDD.n3549 DVDD.n3548 0.0196339
R3449 DVDD.n3550 DVDD.n3549 0.0196339
R3450 DVDD.n3551 DVDD.n3550 0.0196339
R3451 DVDD.n3552 DVDD.n3551 0.0196339
R3452 DVDD.n3568 DVDD.n3552 0.0196339
R3453 DVDD.n3742 DVDD.n3741 0.0196339
R3454 DVDD.n10017 DVDD.n10016 0.0196339
R3455 DVDD.n10016 DVDD.n10015 0.0196339
R3456 DVDD.n10015 DVDD.n10014 0.0196339
R3457 DVDD.n10014 DVDD.n10013 0.0196339
R3458 DVDD.n10013 DVDD.n10012 0.0196339
R3459 DVDD.n10012 DVDD.n10011 0.0196339
R3460 DVDD.n10011 DVDD.n10010 0.0196339
R3461 DVDD.n10010 DVDD.n10009 0.0196339
R3462 DVDD.n10009 DVDD.n10008 0.0196339
R3463 DVDD.n10008 DVDD.n10007 0.0196339
R3464 DVDD.n10007 DVDD.n10006 0.0196339
R3465 DVDD.n10006 DVDD.n10005 0.0196339
R3466 DVDD.n10005 DVDD.n10004 0.0196339
R3467 DVDD.n10004 DVDD.n10003 0.0196339
R3468 DVDD.n10003 DVDD.n10002 0.0196339
R3469 DVDD.n10002 DVDD.n10001 0.0196339
R3470 DVDD.n10001 DVDD.n10000 0.0196339
R3471 DVDD.n10000 DVDD.n9999 0.0196339
R3472 DVDD.n9999 DVDD.n9998 0.0196339
R3473 DVDD.n9998 DVDD.n9997 0.0196339
R3474 DVDD.n9990 DVDD.n7156 0.0196339
R3475 DVDD.n7831 DVDD.n7156 0.0196339
R3476 DVDD.n7832 DVDD.n7831 0.0196339
R3477 DVDD.n7833 DVDD.n7832 0.0196339
R3478 DVDD.n7834 DVDD.n7833 0.0196339
R3479 DVDD.n7835 DVDD.n7834 0.0196339
R3480 DVDD.n7836 DVDD.n7835 0.0196339
R3481 DVDD.n7837 DVDD.n7836 0.0196339
R3482 DVDD.n7838 DVDD.n7837 0.0196339
R3483 DVDD.n7839 DVDD.n7838 0.0196339
R3484 DVDD.n7840 DVDD.n7839 0.0196339
R3485 DVDD.n7841 DVDD.n7840 0.0196339
R3486 DVDD.n7842 DVDD.n7841 0.0196339
R3487 DVDD.n7843 DVDD.n7842 0.0196339
R3488 DVDD.n7844 DVDD.n7843 0.0196339
R3489 DVDD.n7845 DVDD.n7844 0.0196339
R3490 DVDD.n7846 DVDD.n7845 0.0196339
R3491 DVDD.n7847 DVDD.n7846 0.0196339
R3492 DVDD.n7848 DVDD.n7847 0.0196339
R3493 DVDD.n7849 DVDD.n7848 0.0196339
R3494 DVDD.n7850 DVDD.n7849 0.0196339
R3495 DVDD.n7851 DVDD.n7850 0.0196339
R3496 DVDD.n7852 DVDD.n7851 0.0196339
R3497 DVDD.n7853 DVDD.n7852 0.0196339
R3498 DVDD.n7854 DVDD.n7853 0.0196339
R3499 DVDD.n7855 DVDD.n7854 0.0196339
R3500 DVDD.n9640 DVDD.n9639 0.0196339
R3501 DVDD.n9639 DVDD.n9638 0.0196339
R3502 DVDD.n9582 DVDD.n9581 0.0196339
R3503 DVDD.n9581 DVDD.n9580 0.0196339
R3504 DVDD.n9580 DVDD.n9579 0.0196339
R3505 DVDD.n9579 DVDD.n9578 0.0196339
R3506 DVDD.n9578 DVDD.n9577 0.0196339
R3507 DVDD.n9577 DVDD.n9576 0.0196339
R3508 DVDD.n9576 DVDD.n9575 0.0196339
R3509 DVDD.n9575 DVDD.n9574 0.0196339
R3510 DVDD.n9574 DVDD.n9573 0.0196339
R3511 DVDD.n9573 DVDD.n9572 0.0196339
R3512 DVDD.n9572 DVDD.n9571 0.0196339
R3513 DVDD.n9571 DVDD.n9570 0.0196339
R3514 DVDD.n9570 DVDD.n9569 0.0196339
R3515 DVDD.n9569 DVDD.n9568 0.0196339
R3516 DVDD.n9568 DVDD.n9567 0.0196339
R3517 DVDD.n9567 DVDD.n9566 0.0196339
R3518 DVDD.n9566 DVDD.n9565 0.0196339
R3519 DVDD.n9186 DVDD.n9185 0.0196339
R3520 DVDD.n9185 DVDD.n9184 0.0196339
R3521 DVDD.n19000 DVDD.n18999 0.019625
R3522 DVDD.n10603 DVDD.n10602 0.019625
R3523 DVDD.n17297 DVDD.n17296 0.0195541
R3524 DVDD.n17676 DVDD.n17675 0.0195541
R3525 DVDD DVDD.n7598 0.0193923
R3526 DVDD.n15973 DVDD.n15972 0.0193285
R3527 DVDD.n8124 DVDD.n8123 0.0193285
R3528 DVDD.n19768 DVDD.n19767 0.0192795
R3529 DVDD.n19838 DVDD.n19837 0.0192795
R3530 DVDD.n19993 DVDD.n19992 0.0192795
R3531 DVDD.n4704 DVDD.n4703 0.0192795
R3532 DVDD.n4774 DVDD.n4773 0.0192795
R3533 DVDD.n1413 DVDD.n1412 0.0192795
R3534 DVDD.n1538 DVDD.n1537 0.0192795
R3535 DVDD.n1681 DVDD.n1680 0.0192795
R3536 DVDD.n11411 DVDD.n11410 0.0192795
R3537 DVDD.n11600 DVDD.n11599 0.0192795
R3538 DVDD.n1990 DVDD.n1989 0.0192795
R3539 DVDD.n2060 DVDD.n2059 0.0192795
R3540 DVDD.n2214 DVDD.n2213 0.0192795
R3541 DVDD.n6980 DVDD.n6979 0.0192795
R3542 DVDD.n6910 DVDD.n6909 0.0192795
R3543 DVDD.n3190 DVDD.n3189 0.0192795
R3544 DVDD.n3459 DVDD.n3458 0.0192795
R3545 DVDD.n3568 DVDD.n3567 0.0192795
R3546 DVDD.n9997 DVDD.n9996 0.0192795
R3547 DVDD.n7856 DVDD.n7855 0.0192795
R3548 DVDD.n13919 DVDD.n13913 0.0191486
R3549 DVDD.n14308 DVDD.n14302 0.0191486
R3550 DVDD.n15951 DVDD.n15950 0.0191402
R3551 DVDD.n15691 DVDD.n15690 0.0191402
R3552 DVDD.n9408 DVDD.n9407 0.0191402
R3553 DVDD.n19313 DVDD.n19312 0.0191024
R3554 DVDD.n10160 DVDD.n10159 0.0191024
R3555 DVDD.n11483 DVDD.n11482 0.0191024
R3556 DVDD.n11479 DVDD.n11478 0.0191024
R3557 DVDD.n12187 DVDD.n12186 0.0191024
R3558 DVDD.n12191 DVDD.n12190 0.0191024
R3559 DVDD.n12217 DVDD.n12216 0.0191024
R3560 DVDD.n12210 DVDD.n12209 0.0191024
R3561 DVDD.n12206 DVDD.n12205 0.0191024
R3562 DVDD.n13508 DVDD.n13507 0.0191024
R3563 DVDD.n13512 DVDD.n13511 0.0191024
R3564 DVDD.n13521 DVDD.n13520 0.0191024
R3565 DVDD.n13525 DVDD.n13524 0.0191024
R3566 DVDD.n13534 DVDD.n13533 0.0191024
R3567 DVDD.n13538 DVDD.n13537 0.0191024
R3568 DVDD.n13545 DVDD.n13544 0.0191024
R3569 DVDD.n13549 DVDD.n13548 0.0191024
R3570 DVDD.n13553 DVDD.n13552 0.0191024
R3571 DVDD.n13560 DVDD.n13559 0.0191024
R3572 DVDD.n13564 DVDD.n13563 0.0191024
R3573 DVDD.n13573 DVDD.n13572 0.0191024
R3574 DVDD.n13577 DVDD.n13576 0.0191024
R3575 DVDD.n13587 DVDD.n13586 0.0191024
R3576 DVDD.n13591 DVDD.n13590 0.0191024
R3577 DVDD.n13600 DVDD.n13599 0.0191024
R3578 DVDD.n13604 DVDD.n13603 0.0191024
R3579 DVDD.n13615 DVDD.n13614 0.0191024
R3580 DVDD.n13619 DVDD.n13618 0.0191024
R3581 DVDD.n13626 DVDD.n13625 0.0191024
R3582 DVDD.n13630 DVDD.n13629 0.0191024
R3583 DVDD.n13634 DVDD.n13633 0.0191024
R3584 DVDD.n13641 DVDD.n13640 0.0191024
R3585 DVDD.n13645 DVDD.n13644 0.0191024
R3586 DVDD.n13654 DVDD.n13653 0.0191024
R3587 DVDD.n13658 DVDD.n13657 0.0191024
R3588 DVDD.n13668 DVDD.n13667 0.0191024
R3589 DVDD.n13672 DVDD.n13671 0.0191024
R3590 DVDD.n13681 DVDD.n13680 0.0191024
R3591 DVDD.n13685 DVDD.n13684 0.0191024
R3592 DVDD.n13699 DVDD.n13698 0.0191024
R3593 DVDD.n13703 DVDD.n13702 0.0191024
R3594 DVDD.n13723 DVDD.n13722 0.0191024
R3595 DVDD.n13719 DVDD.n13718 0.0191024
R3596 DVDD.n13712 DVDD.n13711 0.0191024
R3597 DVDD.n2718 DVDD.n2717 0.0191024
R3598 DVDD.n2727 DVDD.n2726 0.0191024
R3599 DVDD.n2731 DVDD.n2730 0.0191024
R3600 DVDD.n2738 DVDD.n2737 0.0191024
R3601 DVDD.n2742 DVDD.n2741 0.0191024
R3602 DVDD.n2746 DVDD.n2745 0.0191024
R3603 DVDD.n2759 DVDD.n2758 0.0191024
R3604 DVDD.n2768 DVDD.n2767 0.0191024
R3605 DVDD.n2772 DVDD.n2771 0.0191024
R3606 DVDD.n2779 DVDD.n2778 0.0191024
R3607 DVDD.n2783 DVDD.n2782 0.0191024
R3608 DVDD.n2787 DVDD.n2786 0.0191024
R3609 DVDD.n2799 DVDD.n2798 0.0191024
R3610 DVDD.n2805 DVDD.n2804 0.0191024
R3611 DVDD.n2808 DVDD.n2807 0.0191024
R3612 DVDD.n18579 DVDD.n18578 0.0191024
R3613 DVDD.n18576 DVDD.n18575 0.0191024
R3614 DVDD.n18573 DVDD.n18572 0.0191024
R3615 DVDD.n18675 DVDD.n18674 0.0191024
R3616 DVDD.n18678 DVDD.n18677 0.0191024
R3617 DVDD.n18481 DVDD.n18480 0.0191024
R3618 DVDD.n18478 DVDD.n18477 0.0191024
R3619 DVDD.n18472 DVDD.n18471 0.0191024
R3620 DVDD.n10058 DVDD.n10057 0.0191024
R3621 DVDD.n10064 DVDD.n10063 0.0191024
R3622 DVDD.n10067 DVDD.n10066 0.0191024
R3623 DVDD.n14801 DVDD.n14800 0.0191024
R3624 DVDD.n14804 DVDD.n14803 0.0191024
R3625 DVDD.n14807 DVDD.n14806 0.0191024
R3626 DVDD.n14817 DVDD.n14816 0.0191024
R3627 DVDD.n14821 DVDD.n14820 0.0191024
R3628 DVDD.n15390 DVDD.n15389 0.0191024
R3629 DVDD.n15394 DVDD.n15393 0.0191024
R3630 DVDD.n15398 DVDD.n15397 0.0191024
R3631 DVDD.n15407 DVDD.n15406 0.0191024
R3632 DVDD.n15411 DVDD.n15410 0.0191024
R3633 DVDD.n15420 DVDD.n15419 0.0191024
R3634 DVDD.n15424 DVDD.n15423 0.0191024
R3635 DVDD.n15437 DVDD.n15436 0.0191024
R3636 DVDD.n15441 DVDD.n15440 0.0191024
R3637 DVDD.n15450 DVDD.n15449 0.0191024
R3638 DVDD.n15454 DVDD.n15453 0.0191024
R3639 DVDD.n15472 DVDD.n15471 0.0191024
R3640 DVDD.n15476 DVDD.n15475 0.0191024
R3641 DVDD.n15487 DVDD.n15486 0.0191024
R3642 DVDD.n15491 DVDD.n15490 0.0191024
R3643 DVDD.n15500 DVDD.n15499 0.0191024
R3644 DVDD.n15508 DVDD.n15507 0.0191024
R3645 DVDD.n15512 DVDD.n15511 0.0191024
R3646 DVDD.n14737 DVDD.n14736 0.0191024
R3647 DVDD.n14733 DVDD.n14732 0.0191024
R3648 DVDD.n14724 DVDD.n14723 0.0191024
R3649 DVDD.n14720 DVDD.n14719 0.0191024
R3650 DVDD.n14713 DVDD.n14712 0.0191024
R3651 DVDD.n14709 DVDD.n14708 0.0191024
R3652 DVDD.n14705 DVDD.n14704 0.0191024
R3653 DVDD.n14696 DVDD.n14695 0.0191024
R3654 DVDD.n14692 DVDD.n14691 0.0191024
R3655 DVDD.n14683 DVDD.n14682 0.0191024
R3656 DVDD.n14679 DVDD.n14678 0.0191024
R3657 DVDD.n14669 DVDD.n14668 0.0191024
R3658 DVDD.n14665 DVDD.n14664 0.0191024
R3659 DVDD.n14654 DVDD.n14653 0.0191024
R3660 DVDD.n14650 DVDD.n14649 0.0191024
R3661 DVDD.n14641 DVDD.n14640 0.0191024
R3662 DVDD.n14637 DVDD.n14636 0.0191024
R3663 DVDD.n14630 DVDD.n14629 0.0191024
R3664 DVDD.n14626 DVDD.n14625 0.0191024
R3665 DVDD.n14622 DVDD.n14621 0.0191024
R3666 DVDD.n14613 DVDD.n14612 0.0191024
R3667 DVDD.n14609 DVDD.n14608 0.0191024
R3668 DVDD.n14600 DVDD.n14599 0.0191024
R3669 DVDD.n14596 DVDD.n14595 0.0191024
R3670 DVDD.n14592 DVDD.n14591 0.0191024
R3671 DVDD.n14587 DVDD.n14586 0.0191024
R3672 DVDD.n14583 DVDD.n14582 0.0191024
R3673 DVDD.n14576 DVDD.n14575 0.0191024
R3674 DVDD.n14572 DVDD.n14571 0.0191024
R3675 DVDD.n14568 DVDD.n14567 0.0191024
R3676 DVDD.n14559 DVDD.n14558 0.0191024
R3677 DVDD.n14555 DVDD.n14554 0.0191024
R3678 DVDD.n14546 DVDD.n14545 0.0191024
R3679 DVDD.n14542 DVDD.n14541 0.0191024
R3680 DVDD.n14529 DVDD.n14528 0.0191024
R3681 DVDD.n14525 DVDD.n14524 0.0191024
R3682 DVDD.n14516 DVDD.n14515 0.0191024
R3683 DVDD.n14512 DVDD.n14511 0.0191024
R3684 DVDD.n14499 DVDD.n14498 0.0191024
R3685 DVDD.n14495 DVDD.n14494 0.0191024
R3686 DVDD.n14488 DVDD.n14487 0.0191024
R3687 DVDD.n14484 DVDD.n14483 0.0191024
R3688 DVDD.n14480 DVDD.n14479 0.0191024
R3689 DVDD.n14471 DVDD.n14470 0.0191024
R3690 DVDD.n14467 DVDD.n14466 0.0191024
R3691 DVDD.n14458 DVDD.n14457 0.0191024
R3692 DVDD.n14454 DVDD.n14453 0.0191024
R3693 DVDD.n14412 DVDD.n14411 0.0191024
R3694 DVDD.n14408 DVDD.n14407 0.0191024
R3695 DVDD.n14390 DVDD.n14389 0.0191024
R3696 DVDD.n14386 DVDD.n14385 0.0191024
R3697 DVDD.n14375 DVDD.n14374 0.0191024
R3698 DVDD.n14371 DVDD.n14370 0.0191024
R3699 DVDD.n14362 DVDD.n14361 0.0191024
R3700 DVDD.n19774 DVDD.n19773 0.0191024
R3701 DVDD.n19844 DVDD.n19843 0.0191024
R3702 DVDD.n19999 DVDD.n19998 0.0191024
R3703 DVDD.n3859 DVDD.n3858 0.0191024
R3704 DVDD.n3865 DVDD.n3864 0.0191024
R3705 DVDD.n3868 DVDD.n3867 0.0191024
R3706 DVDD.n4747 DVDD.n4709 0.0191024
R3707 DVDD.n4781 DVDD.n4780 0.0191024
R3708 DVDD.n4785 DVDD.n4784 0.0191024
R3709 DVDD.n5047 DVDD.n5046 0.0191024
R3710 DVDD.n5051 DVDD.n5050 0.0191024
R3711 DVDD.n5205 DVDD.n5204 0.0191024
R3712 DVDD.n5212 DVDD.n5211 0.0191024
R3713 DVDD.n5216 DVDD.n5215 0.0191024
R3714 DVDD.n5220 DVDD.n5219 0.0191024
R3715 DVDD.n5474 DVDD.n5473 0.0191024
R3716 DVDD.n5478 DVDD.n5477 0.0191024
R3717 DVDD.n5487 DVDD.n5486 0.0191024
R3718 DVDD.n5491 DVDD.n5490 0.0191024
R3719 DVDD.n5548 DVDD.n5547 0.0191024
R3720 DVDD.n5552 DVDD.n5551 0.0191024
R3721 DVDD.n5559 DVDD.n5558 0.0191024
R3722 DVDD.n5597 DVDD.n5596 0.0191024
R3723 DVDD.n5601 DVDD.n5600 0.0191024
R3724 DVDD.n5648 DVDD.n5647 0.0191024
R3725 DVDD.n5652 DVDD.n5651 0.0191024
R3726 DVDD.n5688 DVDD.n5687 0.0191024
R3727 DVDD.n6084 DVDD.n6083 0.0191024
R3728 DVDD.n6080 DVDD.n6079 0.0191024
R3729 DVDD.n6076 DVDD.n6075 0.0191024
R3730 DVDD.n6026 DVDD.n6025 0.0191024
R3731 DVDD.n6022 DVDD.n6021 0.0191024
R3732 DVDD.n5970 DVDD.n5969 0.0191024
R3733 DVDD.n5966 DVDD.n5965 0.0191024
R3734 DVDD.n5952 DVDD.n5951 0.0191024
R3735 DVDD.n5948 DVDD.n5947 0.0191024
R3736 DVDD.n5937 DVDD.n5936 0.0191024
R3737 DVDD.n5933 DVDD.n5932 0.0191024
R3738 DVDD.n5926 DVDD.n5925 0.0191024
R3739 DVDD.n1419 DVDD.n1418 0.0191024
R3740 DVDD.n1532 DVDD.n1531 0.0191024
R3741 DVDD.n1687 DVDD.n1686 0.0191024
R3742 DVDD.n10106 DVDD.n10105 0.0191024
R3743 DVDD.n10112 DVDD.n10111 0.0191024
R3744 DVDD.n10115 DVDD.n10114 0.0191024
R3745 DVDD.n11573 DVDD.n11416 0.0191024
R3746 DVDD.n11607 DVDD.n11606 0.0191024
R3747 DVDD.n11611 DVDD.n11610 0.0191024
R3748 DVDD.n11707 DVDD.n11706 0.0191024
R3749 DVDD.n11703 DVDD.n11702 0.0191024
R3750 DVDD.n12385 DVDD.n12384 0.0191024
R3751 DVDD.n12392 DVDD.n12391 0.0191024
R3752 DVDD.n12396 DVDD.n12395 0.0191024
R3753 DVDD.n12400 DVDD.n12399 0.0191024
R3754 DVDD.n12989 DVDD.n12988 0.0191024
R3755 DVDD.n12985 DVDD.n12984 0.0191024
R3756 DVDD.n12976 DVDD.n12975 0.0191024
R3757 DVDD.n12972 DVDD.n12971 0.0191024
R3758 DVDD.n12869 DVDD.n12868 0.0191024
R3759 DVDD.n12865 DVDD.n12864 0.0191024
R3760 DVDD.n12858 DVDD.n12857 0.0191024
R3761 DVDD.n12830 DVDD.n12829 0.0191024
R3762 DVDD.n12826 DVDD.n12825 0.0191024
R3763 DVDD.n12789 DVDD.n12788 0.0191024
R3764 DVDD.n12785 DVDD.n12784 0.0191024
R3765 DVDD.n12753 DVDD.n12752 0.0191024
R3766 DVDD.n12716 DVDD.n12715 0.0191024
R3767 DVDD.n12712 DVDD.n12711 0.0191024
R3768 DVDD.n12708 DVDD.n12707 0.0191024
R3769 DVDD.n12677 DVDD.n12676 0.0191024
R3770 DVDD.n12673 DVDD.n12672 0.0191024
R3771 DVDD.n12633 DVDD.n12632 0.0191024
R3772 DVDD.n12629 DVDD.n12628 0.0191024
R3773 DVDD.n12615 DVDD.n12614 0.0191024
R3774 DVDD.n12611 DVDD.n12610 0.0191024
R3775 DVDD.n12600 DVDD.n12599 0.0191024
R3776 DVDD.n12596 DVDD.n12595 0.0191024
R3777 DVDD.n12589 DVDD.n12588 0.0191024
R3778 DVDD.n758 DVDD.n757 0.0191024
R3779 DVDD.n765 DVDD.n764 0.0191024
R3780 DVDD.n769 DVDD.n768 0.0191024
R3781 DVDD.n776 DVDD.n775 0.0191024
R3782 DVDD.n780 DVDD.n779 0.0191024
R3783 DVDD.n784 DVDD.n783 0.0191024
R3784 DVDD.n795 DVDD.n794 0.0191024
R3785 DVDD.n802 DVDD.n801 0.0191024
R3786 DVDD.n806 DVDD.n805 0.0191024
R3787 DVDD.n813 DVDD.n812 0.0191024
R3788 DVDD.n817 DVDD.n816 0.0191024
R3789 DVDD.n821 DVDD.n820 0.0191024
R3790 DVDD.n831 DVDD.n830 0.0191024
R3791 DVDD.n837 DVDD.n836 0.0191024
R3792 DVDD.n840 DVDD.n839 0.0191024
R3793 DVDD.n248 DVDD.n247 0.0191024
R3794 DVDD.n245 DVDD.n244 0.0191024
R3795 DVDD.n242 DVDD.n241 0.0191024
R3796 DVDD.n154 DVDD.n153 0.0191024
R3797 DVDD.n157 DVDD.n156 0.0191024
R3798 DVDD.n19177 DVDD.n19176 0.0191024
R3799 DVDD.n19174 DVDD.n19173 0.0191024
R3800 DVDD.n19168 DVDD.n19167 0.0191024
R3801 DVDD.n10090 DVDD.n10089 0.0191024
R3802 DVDD.n10096 DVDD.n10095 0.0191024
R3803 DVDD.n10099 DVDD.n10098 0.0191024
R3804 DVDD.n18237 DVDD.n18236 0.0191024
R3805 DVDD.n18234 DVDD.n18233 0.0191024
R3806 DVDD.n18231 DVDD.n18230 0.0191024
R3807 DVDD.n18221 DVDD.n18220 0.0191024
R3808 DVDD.n18217 DVDD.n18216 0.0191024
R3809 DVDD.n18210 DVDD.n18209 0.0191024
R3810 DVDD.n18206 DVDD.n18205 0.0191024
R3811 DVDD.n18202 DVDD.n18201 0.0191024
R3812 DVDD.n18195 DVDD.n18194 0.0191024
R3813 DVDD.n18191 DVDD.n18190 0.0191024
R3814 DVDD.n18182 DVDD.n18181 0.0191024
R3815 DVDD.n18178 DVDD.n18177 0.0191024
R3816 DVDD.n18168 DVDD.n18167 0.0191024
R3817 DVDD.n18164 DVDD.n18163 0.0191024
R3818 DVDD.n18155 DVDD.n18154 0.0191024
R3819 DVDD.n18151 DVDD.n18150 0.0191024
R3820 DVDD.n18137 DVDD.n18136 0.0191024
R3821 DVDD.n18133 DVDD.n18132 0.0191024
R3822 DVDD.n18122 DVDD.n18121 0.0191024
R3823 DVDD.n18118 DVDD.n18117 0.0191024
R3824 DVDD.n18111 DVDD.n18110 0.0191024
R3825 DVDD.n18103 DVDD.n18102 0.0191024
R3826 DVDD.n18099 DVDD.n18098 0.0191024
R3827 DVDD.n18088 DVDD.n18087 0.0191024
R3828 DVDD.n18084 DVDD.n18083 0.0191024
R3829 DVDD.n18077 DVDD.n18076 0.0191024
R3830 DVDD.n18073 DVDD.n18072 0.0191024
R3831 DVDD.n18066 DVDD.n18065 0.0191024
R3832 DVDD.n18062 DVDD.n18061 0.0191024
R3833 DVDD.n18058 DVDD.n18057 0.0191024
R3834 DVDD.n18051 DVDD.n18050 0.0191024
R3835 DVDD.n18047 DVDD.n18046 0.0191024
R3836 DVDD.n18038 DVDD.n18037 0.0191024
R3837 DVDD.n18034 DVDD.n18033 0.0191024
R3838 DVDD.n18025 DVDD.n18024 0.0191024
R3839 DVDD.n18021 DVDD.n18020 0.0191024
R3840 DVDD.n18010 DVDD.n18009 0.0191024
R3841 DVDD.n18006 DVDD.n18005 0.0191024
R3842 DVDD.n17999 DVDD.n17998 0.0191024
R3843 DVDD.n17995 DVDD.n17994 0.0191024
R3844 DVDD.n17988 DVDD.n17987 0.0191024
R3845 DVDD.n17984 DVDD.n17983 0.0191024
R3846 DVDD.n17980 DVDD.n17979 0.0191024
R3847 DVDD.n17973 DVDD.n17972 0.0191024
R3848 DVDD.n17969 DVDD.n17968 0.0191024
R3849 DVDD.n17960 DVDD.n17959 0.0191024
R3850 DVDD.n17956 DVDD.n17955 0.0191024
R3851 DVDD.n17952 DVDD.n17951 0.0191024
R3852 DVDD.n17947 DVDD.n17946 0.0191024
R3853 DVDD.n17943 DVDD.n17942 0.0191024
R3854 DVDD.n17936 DVDD.n17935 0.0191024
R3855 DVDD.n17932 DVDD.n17931 0.0191024
R3856 DVDD.n17928 DVDD.n17927 0.0191024
R3857 DVDD.n17921 DVDD.n17920 0.0191024
R3858 DVDD.n17917 DVDD.n17916 0.0191024
R3859 DVDD.n17908 DVDD.n17907 0.0191024
R3860 DVDD.n17904 DVDD.n17903 0.0191024
R3861 DVDD.n17894 DVDD.n17893 0.0191024
R3862 DVDD.n17890 DVDD.n17889 0.0191024
R3863 DVDD.n17881 DVDD.n17880 0.0191024
R3864 DVDD.n17877 DVDD.n17876 0.0191024
R3865 DVDD.n17866 DVDD.n17865 0.0191024
R3866 DVDD.n17862 DVDD.n17861 0.0191024
R3867 DVDD.n17855 DVDD.n17854 0.0191024
R3868 DVDD.n17851 DVDD.n17850 0.0191024
R3869 DVDD.n17847 DVDD.n17846 0.0191024
R3870 DVDD.n17840 DVDD.n17839 0.0191024
R3871 DVDD.n17836 DVDD.n17835 0.0191024
R3872 DVDD.n17827 DVDD.n17826 0.0191024
R3873 DVDD.n17823 DVDD.n17822 0.0191024
R3874 DVDD.n17786 DVDD.n17785 0.0191024
R3875 DVDD.n17782 DVDD.n17781 0.0191024
R3876 DVDD.n17768 DVDD.n17767 0.0191024
R3877 DVDD.n17764 DVDD.n17763 0.0191024
R3878 DVDD.n17753 DVDD.n17752 0.0191024
R3879 DVDD.n17749 DVDD.n17748 0.0191024
R3880 DVDD.n17742 DVDD.n17741 0.0191024
R3881 DVDD.n1996 DVDD.n1995 0.0191024
R3882 DVDD.n2066 DVDD.n2065 0.0191024
R3883 DVDD.n2220 DVDD.n2219 0.0191024
R3884 DVDD.n7080 DVDD.n7079 0.0191024
R3885 DVDD.n7086 DVDD.n7085 0.0191024
R3886 DVDD.n7089 DVDD.n7088 0.0191024
R3887 DVDD.n6974 DVDD.n6973 0.0191024
R3888 DVDD.n6903 DVDD.n6902 0.0191024
R3889 DVDD.n6899 DVDD.n6898 0.0191024
R3890 DVDD.n6637 DVDD.n6636 0.0191024
R3891 DVDD.n6633 DVDD.n6632 0.0191024
R3892 DVDD.n6477 DVDD.n6476 0.0191024
R3893 DVDD.n6470 DVDD.n6469 0.0191024
R3894 DVDD.n6466 DVDD.n6465 0.0191024
R3895 DVDD.n6462 DVDD.n6461 0.0191024
R3896 DVDD.n6285 DVDD.n6284 0.0191024
R3897 DVDD.n6281 DVDD.n6280 0.0191024
R3898 DVDD.n6272 DVDD.n6271 0.0191024
R3899 DVDD.n6268 DVDD.n6267 0.0191024
R3900 DVDD.n6248 DVDD.n6247 0.0191024
R3901 DVDD.n6244 DVDD.n6243 0.0191024
R3902 DVDD.n6237 DVDD.n6236 0.0191024
R3903 DVDD.n6208 DVDD.n6207 0.0191024
R3904 DVDD.n6204 DVDD.n6203 0.0191024
R3905 DVDD.n6166 DVDD.n6165 0.0191024
R3906 DVDD.n6162 DVDD.n6161 0.0191024
R3907 DVDD.n6137 DVDD.n6136 0.0191024
R3908 DVDD.n4534 DVDD.n4533 0.0191024
R3909 DVDD.n4530 DVDD.n4529 0.0191024
R3910 DVDD.n4526 DVDD.n4525 0.0191024
R3911 DVDD.n4477 DVDD.n4476 0.0191024
R3912 DVDD.n4473 DVDD.n4472 0.0191024
R3913 DVDD.n4433 DVDD.n4432 0.0191024
R3914 DVDD.n4429 DVDD.n4428 0.0191024
R3915 DVDD.n4411 DVDD.n4410 0.0191024
R3916 DVDD.n4407 DVDD.n4406 0.0191024
R3917 DVDD.n4396 DVDD.n4395 0.0191024
R3918 DVDD.n4392 DVDD.n4391 0.0191024
R3919 DVDD.n4383 DVDD.n4382 0.0191024
R3920 DVDD.n3184 DVDD.n3183 0.0191024
R3921 DVDD.n3465 DVDD.n3464 0.0191024
R3922 DVDD.n3562 DVDD.n3561 0.0191024
R3923 DVDD.n7138 DVDD.n7137 0.0191024
R3924 DVDD.n7144 DVDD.n7143 0.0191024
R3925 DVDD.n7147 DVDD.n7146 0.0191024
R3926 DVDD.n9991 DVDD.n9990 0.0191024
R3927 DVDD.n7863 DVDD.n7862 0.0191024
R3928 DVDD.n7867 DVDD.n7866 0.0191024
R3929 DVDD.n9605 DVDD.n9604 0.0191024
R3930 DVDD.n9601 DVDD.n9600 0.0191024
R3931 DVDD.n8406 DVDD.n8405 0.0191024
R3932 DVDD.n8413 DVDD.n8412 0.0191024
R3933 DVDD.n8417 DVDD.n8416 0.0191024
R3934 DVDD.n8421 DVDD.n8420 0.0191024
R3935 DVDD.n9071 DVDD.n9070 0.0191024
R3936 DVDD.n9067 DVDD.n9066 0.0191024
R3937 DVDD.n9058 DVDD.n9057 0.0191024
R3938 DVDD.n9054 DVDD.n9053 0.0191024
R3939 DVDD.n8950 DVDD.n8949 0.0191024
R3940 DVDD.n8946 DVDD.n8945 0.0191024
R3941 DVDD.n8939 DVDD.n8938 0.0191024
R3942 DVDD.n8910 DVDD.n8909 0.0191024
R3943 DVDD.n8906 DVDD.n8905 0.0191024
R3944 DVDD.n8868 DVDD.n8867 0.0191024
R3945 DVDD.n8864 DVDD.n8863 0.0191024
R3946 DVDD.n8839 DVDD.n8838 0.0191024
R3947 DVDD.n8801 DVDD.n8800 0.0191024
R3948 DVDD.n8797 DVDD.n8796 0.0191024
R3949 DVDD.n8793 DVDD.n8792 0.0191024
R3950 DVDD.n8763 DVDD.n8762 0.0191024
R3951 DVDD.n8759 DVDD.n8758 0.0191024
R3952 DVDD.n8707 DVDD.n8706 0.0191024
R3953 DVDD.n8703 DVDD.n8702 0.0191024
R3954 DVDD.n8685 DVDD.n8684 0.0191024
R3955 DVDD.n8681 DVDD.n8680 0.0191024
R3956 DVDD.n8670 DVDD.n8669 0.0191024
R3957 DVDD.n8666 DVDD.n8665 0.0191024
R3958 DVDD.n8657 DVDD.n8656 0.0191024
R3959 DVDD.n7664 DVDD.n7663 0.018978
R3960 DVDD.n16041 DVDD.n16040 0.0189519
R3961 DVDD.n16010 DVDD.n16009 0.0189519
R3962 DVDD.n15653 DVDD.n15652 0.0189519
R3963 DVDD.n15922 DVDD.n15921 0.0189519
R3964 DVDD.n8156 DVDD.n8155 0.0189519
R3965 DVDD.n11449 DVDD.n11448 0.0189252
R3966 DVDD.n12180 DVDD.n12179 0.0189252
R3967 DVDD.n13707 DVDD.n13706 0.0189252
R3968 DVDD.n18681 DVDD.n18680 0.0189252
R3969 DVDD.n15480 DVDD.n15479 0.0189252
R3970 DVDD.n14741 DVDD.n14740 0.0189252
R3971 DVDD.n14658 DVDD.n14657 0.0189252
R3972 DVDD.n14382 DVDD.n14381 0.0189252
R3973 DVDD.n5040 DVDD.n5039 0.0189252
R3974 DVDD.n5944 DVDD.n5943 0.0189252
R3975 DVDD.n11714 DVDD.n11713 0.0189252
R3976 DVDD.n12607 DVDD.n12606 0.0189252
R3977 DVDD.n160 DVDD.n159 0.0189252
R3978 DVDD.n18129 DVDD.n18128 0.0189252
R3979 DVDD.n18092 DVDD.n18091 0.0189252
R3980 DVDD.n18014 DVDD.n18013 0.0189252
R3981 DVDD.n17760 DVDD.n17759 0.0189252
R3982 DVDD.n6644 DVDD.n6643 0.0189252
R3983 DVDD.n4403 DVDD.n4402 0.0189252
R3984 DVDD.n9612 DVDD.n9611 0.0189252
R3985 DVDD.n8677 DVDD.n8676 0.0189252
R3986 DVDD.n16040 DVDD.n16039 0.0187636
R3987 DVDD.n16011 DVDD.n16010 0.0187636
R3988 DVDD.n15652 DVDD.n15651 0.0187636
R3989 DVDD.n15921 DVDD.n15920 0.0187636
R3990 DVDD.n8155 DVDD.n8154 0.0187636
R3991 DVDD.n1152 DVDD.n1151 0.018748
R3992 DVDD.n1551 DVDD.n1550 0.018748
R3993 DVDD.n1669 DVDD.n1668 0.018748
R3994 DVDD.n11467 DVDD.n11466 0.018748
R3995 DVDD.n11490 DVDD.n11489 0.018748
R3996 DVDD.n19160 DVDD.n19159 0.018725
R3997 DVDD.n10622 DVDD.n10621 0.018725
R3998 DVDD.n1146 DVDD.n1145 0.0185709
R3999 DVDD.n1557 DVDD.n1556 0.0185709
R4000 DVDD.n1663 DVDD.n1662 0.0185709
R4001 DVDD.n872 DVDD.n871 0.0185709
R4002 DVDD.n11513 DVDD.n11472 0.0185709
R4003 DVDD.n12462 DVDD.n12461 0.0185
R4004 DVDD.n12470 DVDD.n12469 0.0185
R4005 DVDD.n5704 DVDD.n5703 0.0185
R4006 DVDD.n4555 DVDD.n4554 0.0185
R4007 DVDD.n6114 DVDD.n6113 0.0185
R4008 DVDD.n4073 DVDD.n4072 0.0185
R4009 DVDD.n8487 DVDD.n8486 0.0185
R4010 DVDD.n8495 DVDD.n8494 0.0185
R4011 DVDD.n12773 DVDD.n12772 0.0185
R4012 DVDD.n12456 DVDD.n12455 0.0185
R4013 DVDD.n5662 DVDD.n5661 0.0185
R4014 DVDD.n4568 DVDD.n4567 0.0185
R4015 DVDD.n4562 DVDD.n4561 0.0185
R4016 DVDD.n4064 DVDD.n4063 0.0185
R4017 DVDD.n8468 DVDD.n8467 0.0185
R4018 DVDD.n8480 DVDD.n8479 0.0185
R4019 DVDD.n12431 DVDD.n12430 0.0185
R4020 DVDD.n12443 DVDD.n12442 0.0185
R4021 DVDD.n5616 DVDD.n5615 0.0185
R4022 DVDD.n4583 DVDD.n4582 0.0185
R4023 DVDD.n4577 DVDD.n4576 0.0185
R4024 DVDD.n4054 DVDD.n4053 0.0185
R4025 DVDD.n8450 DVDD.n8449 0.0185
R4026 DVDD.n8462 DVDD.n8461 0.0185
R4027 DVDD.n12412 DVDD.n12411 0.0185
R4028 DVDD.n12424 DVDD.n12423 0.0185
R4029 DVDD.n5569 DVDD.n5568 0.0185
R4030 DVDD.n4598 DVDD.n4597 0.0185
R4031 DVDD.n4592 DVDD.n4591 0.0185
R4032 DVDD.n4044 DVDD.n4043 0.0185
R4033 DVDD.n8432 DVDD.n8431 0.0185
R4034 DVDD.n8444 DVDD.n8443 0.0185
R4035 DVDD.n3854 DVDD.n3853 0.0185
R4036 DVDD.n139 DVDD.n138 0.0185
R4037 DVDD.n1642 DVDD.n1641 0.0182165
R4038 DVDD.n12183 DVDD.n12182 0.0182165
R4039 DVDD.n13727 DVDD.n13726 0.0182165
R4040 DVDD.n18484 DVDD.n18483 0.0182165
R4041 DVDD.n15483 DVDD.n15482 0.0182165
R4042 DVDD.n15516 DVDD.n15515 0.0182165
R4043 DVDD.n14661 DVDD.n14660 0.0182165
R4044 DVDD.n14379 DVDD.n14378 0.0182165
R4045 DVDD.n5043 DVDD.n5042 0.0182165
R4046 DVDD.n5941 DVDD.n5940 0.0182165
R4047 DVDD.n11711 DVDD.n11710 0.0182165
R4048 DVDD.n12604 DVDD.n12603 0.0182165
R4049 DVDD.n19180 DVDD.n19179 0.0182165
R4050 DVDD.n18126 DVDD.n18125 0.0182165
R4051 DVDD.n18095 DVDD.n18094 0.0182165
R4052 DVDD.n18017 DVDD.n18016 0.0182165
R4053 DVDD.n17757 DVDD.n17756 0.0182165
R4054 DVDD.n6641 DVDD.n6640 0.0182165
R4055 DVDD.n4400 DVDD.n4399 0.0182165
R4056 DVDD.n9609 DVDD.n9608 0.0182165
R4057 DVDD.n8674 DVDD.n8673 0.0182165
R4058 DVDD.n12213 DVDD.n12212 0.0180394
R4059 DVDD.n13542 DVDD.n13541 0.0180394
R4060 DVDD.n13623 DVDD.n13622 0.0180394
R4061 DVDD.n2735 DVDD.n2734 0.0180394
R4062 DVDD.n2776 DVDD.n2775 0.0180394
R4063 DVDD.n2811 DVDD.n2810 0.0180394
R4064 DVDD.n10070 DVDD.n10069 0.0180394
R4065 DVDD.n14825 DVDD.n14824 0.0180394
R4066 DVDD.n14716 DVDD.n14715 0.0180394
R4067 DVDD.n14633 DVDD.n14632 0.0180394
R4068 DVDD.n14579 DVDD.n14578 0.0180394
R4069 DVDD.n14491 DVDD.n14490 0.0180394
R4070 DVDD.n4789 DVDD.n4788 0.0180394
R4071 DVDD.n5209 DVDD.n5208 0.0180394
R4072 DVDD.n5556 DVDD.n5555 0.0180394
R4073 DVDD.n6087 DVDD.n6086 0.0180394
R4074 DVDD.n11615 DVDD.n11614 0.0180394
R4075 DVDD.n12389 DVDD.n12388 0.0180394
R4076 DVDD.n12861 DVDD.n12860 0.0180394
R4077 DVDD.n12719 DVDD.n12718 0.0180394
R4078 DVDD.n773 DVDD.n772 0.0180394
R4079 DVDD.n810 DVDD.n809 0.0180394
R4080 DVDD.n843 DVDD.n842 0.0180394
R4081 DVDD.n10102 DVDD.n10101 0.0180394
R4082 DVDD.n18213 DVDD.n18212 0.0180394
R4083 DVDD.n18069 DVDD.n18068 0.0180394
R4084 DVDD.n17991 DVDD.n17990 0.0180394
R4085 DVDD.n17939 DVDD.n17938 0.0180394
R4086 DVDD.n17858 DVDD.n17857 0.0180394
R4087 DVDD.n6895 DVDD.n6894 0.0180394
R4088 DVDD.n6473 DVDD.n6472 0.0180394
R4089 DVDD.n6240 DVDD.n6239 0.0180394
R4090 DVDD.n4537 DVDD.n4536 0.0180394
R4091 DVDD.n7871 DVDD.n7870 0.0180394
R4092 DVDD.n8410 DVDD.n8409 0.0180394
R4093 DVDD.n8942 DVDD.n8941 0.0180394
R4094 DVDD.n8804 DVDD.n8803 0.0180394
R4095 DVDD.n9891 DVDD.n9890 0.0180105
R4096 DVDD.n13516 DVDD.n13515 0.0178622
R4097 DVDD.n13568 DVDD.n13567 0.0178622
R4098 DVDD.n13596 DVDD.n13595 0.0178622
R4099 DVDD.n13649 DVDD.n13648 0.0178622
R4100 DVDD.n13677 DVDD.n13676 0.0178622
R4101 DVDD.n15415 DVDD.n15414 0.0178622
R4102 DVDD.n15446 DVDD.n15445 0.0178622
R4103 DVDD.n14688 DVDD.n14687 0.0178622
R4104 DVDD.n14605 DVDD.n14604 0.0178622
R4105 DVDD.n14551 DVDD.n14550 0.0178622
R4106 DVDD.n14520 DVDD.n14519 0.0178622
R4107 DVDD.n14463 DVDD.n14462 0.0178622
R4108 DVDD.n14416 DVDD.n14415 0.0178622
R4109 DVDD.n5482 DVDD.n5481 0.0178622
R4110 DVDD.n5605 DVDD.n5604 0.0178622
R4111 DVDD.n6031 DVDD.n6030 0.0178622
R4112 DVDD.n5974 DVDD.n5973 0.0178622
R4113 DVDD.n12981 DVDD.n12980 0.0178622
R4114 DVDD.n12822 DVDD.n12821 0.0178622
R4115 DVDD.n12682 DVDD.n12681 0.0178622
R4116 DVDD.n12637 DVDD.n12636 0.0178622
R4117 DVDD.n18187 DVDD.n18186 0.0178622
R4118 DVDD.n18159 DVDD.n18158 0.0178622
R4119 DVDD.n18043 DVDD.n18042 0.0178622
R4120 DVDD.n17965 DVDD.n17964 0.0178622
R4121 DVDD.n17913 DVDD.n17912 0.0178622
R4122 DVDD.n17885 DVDD.n17884 0.0178622
R4123 DVDD.n17832 DVDD.n17831 0.0178622
R4124 DVDD.n17790 DVDD.n17789 0.0178622
R4125 DVDD.n6277 DVDD.n6276 0.0178622
R4126 DVDD.n6200 DVDD.n6199 0.0178622
R4127 DVDD.n4482 DVDD.n4481 0.0178622
R4128 DVDD.n4437 DVDD.n4436 0.0178622
R4129 DVDD.n9063 DVDD.n9062 0.0178622
R4130 DVDD.n8902 DVDD.n8901 0.0178622
R4131 DVDD.n8768 DVDD.n8767 0.0178622
R4132 DVDD.n8711 DVDD.n8710 0.0178622
R4133 DVDD.n3806 DVDD.n3805 0.017825
R4134 DVDD.n3811 DVDD.n3810 0.017825
R4135 DVDD.n3816 DVDD.n3815 0.017825
R4136 DVDD.n18829 DVDD.n18828 0.017825
R4137 DVDD.n18824 DVDD.n18823 0.017825
R4138 DVDD.n18819 DVDD.n18818 0.017825
R4139 DVDD.n18814 DVDD.n18813 0.017825
R4140 DVDD.n10084 DVDD.n10083 0.017825
R4141 DVDD.n3894 DVDD.n3893 0.017825
R4142 DVDD.n3899 DVDD.n3898 0.017825
R4143 DVDD.n3904 DVDD.n3903 0.017825
R4144 DVDD.n3909 DVDD.n3908 0.017825
R4145 DVDD.n7129 DVDD.n7128 0.017825
R4146 DVDD.n7124 DVDD.n7123 0.017825
R4147 DVDD.n7119 DVDD.n7118 0.017825
R4148 DVDD.n7114 DVDD.n7113 0.017825
R4149 DVDD.n1820 DVDD.n1819 0.017825
R4150 DVDD.n3783 DVDD.n3782 0.017825
R4151 DVDD.n3788 DVDD.n3787 0.017825
R4152 DVDD.n3793 DVDD.n3792 0.017825
R4153 DVDD.n3798 DVDD.n3797 0.017825
R4154 DVDD.n2831 DVDD.n2830 0.017825
R4155 DVDD.n2826 DVDD.n2825 0.017825
R4156 DVDD.n2821 DVDD.n2820 0.017825
R4157 DVDD.n2816 DVDD.n2815 0.017825
R4158 DVDD.n14842 DVDD.n14841 0.017825
R4159 DVDD.n14847 DVDD.n14846 0.017825
R4160 DVDD.n14852 DVDD.n14851 0.017825
R4161 DVDD.n14877 DVDD.n14876 0.017825
R4162 DVDD.n14872 DVDD.n14871 0.017825
R4163 DVDD.n14867 DVDD.n14866 0.017825
R4164 DVDD.n14862 DVDD.n14861 0.017825
R4165 DVDD.n13517 DVDD.n13516 0.017685
R4166 DVDD.n13569 DVDD.n13568 0.017685
R4167 DVDD.n13595 DVDD.n13594 0.017685
R4168 DVDD.n13650 DVDD.n13649 0.017685
R4169 DVDD.n13676 DVDD.n13675 0.017685
R4170 DVDD.n15416 DVDD.n15415 0.017685
R4171 DVDD.n15445 DVDD.n15444 0.017685
R4172 DVDD.n14687 DVDD.n14686 0.017685
R4173 DVDD.n14604 DVDD.n14603 0.017685
R4174 DVDD.n14550 DVDD.n14549 0.017685
R4175 DVDD.n14521 DVDD.n14520 0.017685
R4176 DVDD.n14462 DVDD.n14461 0.017685
R4177 DVDD.n14417 DVDD.n14416 0.017685
R4178 DVDD.n5483 DVDD.n5482 0.017685
R4179 DVDD.n5606 DVDD.n5605 0.017685
R4180 DVDD.n5656 DVDD.n5655 0.017685
R4181 DVDD.n6030 DVDD.n6029 0.017685
R4182 DVDD.n5975 DVDD.n5974 0.017685
R4183 DVDD.n12980 DVDD.n12979 0.017685
R4184 DVDD.n12821 DVDD.n12820 0.017685
R4185 DVDD.n12781 DVDD.n12780 0.017685
R4186 DVDD.n12681 DVDD.n12680 0.017685
R4187 DVDD.n12638 DVDD.n12637 0.017685
R4188 DVDD.n18186 DVDD.n18185 0.017685
R4189 DVDD.n18160 DVDD.n18159 0.017685
R4190 DVDD.n18042 DVDD.n18041 0.017685
R4191 DVDD.n17964 DVDD.n17963 0.017685
R4192 DVDD.n17912 DVDD.n17911 0.017685
R4193 DVDD.n17886 DVDD.n17885 0.017685
R4194 DVDD.n17831 DVDD.n17830 0.017685
R4195 DVDD.n17791 DVDD.n17790 0.017685
R4196 DVDD.n6276 DVDD.n6275 0.017685
R4197 DVDD.n6199 DVDD.n6198 0.017685
R4198 DVDD.n6158 DVDD.n6157 0.017685
R4199 DVDD.n4481 DVDD.n4480 0.017685
R4200 DVDD.n4438 DVDD.n4437 0.017685
R4201 DVDD.n9062 DVDD.n9061 0.017685
R4202 DVDD.n8901 DVDD.n8900 0.017685
R4203 DVDD.n8860 DVDD.n8859 0.017685
R4204 DVDD.n8767 DVDD.n8766 0.017685
R4205 DVDD.n8712 DVDD.n8711 0.017685
R4206 DVDD.n3821 DVDD.n3820 0.0176
R4207 DVDD.n19004 DVDD.n19003 0.0176
R4208 DVDD.n14857 DVDD.n14856 0.0176
R4209 DVDD.n10607 DVDD.n10606 0.0176
R4210 DVDD.n17240 DVDD.n17239 0.0174947
R4211 DVDD.n17407 DVDD.n17406 0.0174947
R4212 DVDD.n17589 DVDD.n17588 0.0174947
R4213 DVDD.n16537 DVDD.n16536 0.0174336
R4214 DVDD.n16832 DVDD.n16831 0.0174336
R4215 DVDD.n16488 DVDD.n16487 0.0174336
R4216 DVDD.n14317 DVDD.n14316 0.0173307
R4217 DVDD.n14234 DVDD.n14164 0.0173307
R4218 DVDD.n14156 DVDD.n14155 0.0173307
R4219 DVDD.n14121 DVDD.n14065 0.0173307
R4220 DVDD.n14057 DVDD.n14056 0.0173307
R4221 DVDD.n14023 DVDD.n13968 0.0173307
R4222 DVDD.n13960 DVDD.n13959 0.0173307
R4223 DVDD.n13926 DVDD.n13883 0.0173307
R4224 DVDD.n17685 DVDD.n17684 0.0173307
R4225 DVDD.n17601 DVDD.n17504 0.0173307
R4226 DVDD.n17496 DVDD.n17495 0.0173307
R4227 DVDD.n17462 DVDD.n17461 0.0173307
R4228 DVDD.n17453 DVDD.n17452 0.0173307
R4229 DVDD.n17419 DVDD.n17345 0.0173307
R4230 DVDD.n17337 DVDD.n17336 0.0173307
R4231 DVDD.n17303 DVDD.n17261 0.0173307
R4232 DVDD.n14090 DVDD.n14089 0.0172553
R4233 DVDD.n14001 DVDD.n14000 0.0172553
R4234 DVDD.n14210 DVDD.n14209 0.0172553
R4235 DVDD.n1564 DVDD.n1563 0.0171535
R4236 DVDD.n16706 DVDD.n16705 0.0170308
R4237 DVDD.n11475 DVDD.n11474 0.0169764
R4238 DVDD.n1662 DVDD.n1661 0.0167992
R4239 DVDD.n19464 DVDD.n18833 0.0167
R4240 DVDD.n19464 DVDD.n19163 0.0167
R4241 DVDD.n7301 DVDD.n7272 0.0167
R4242 DVDD.n14882 DVDD.n14881 0.0167
R4243 DVDD.n15104 DVDD.n15097 0.0167
R4244 DVDD.n10716 DVDD.n10715 0.0167
R4245 DVDD.n10633 DVDD.n10625 0.0167
R4246 DVDD.n7301 DVDD.n7285 0.0167
R4247 DVDD.n5544 DVDD.n5543 0.016622
R4248 DVDD.n12873 DVDD.n12872 0.016622
R4249 DVDD.n6252 DVDD.n6251 0.016622
R4250 DVDD.n8954 DVDD.n8953 0.016622
R4251 DVDD.n18333 DVDD.n3857 0.016475
R4252 DVDD.n7662 DVDD.n7621 0.016475
R4253 DVDD.n18333 DVDD.n3913 0.016475
R4254 DVDD.n7662 DVDD.n7648 0.016475
R4255 DVDD.n20215 DVDD.n142 0.016475
R4256 DVDD.n20215 DVDD.n3802 0.016475
R4257 DVDD.n20338 DVDD.n20289 0.016475
R4258 DVDD.n20338 DVDD.n20336 0.016475
R4259 DVDD.n1159 DVDD.n1158 0.0164449
R4260 DVDD.n10163 DVDD.n10162 0.0162677
R4261 DVDD.n12583 DVDD.n12582 0.0162646
R4262 DVDD.n4351 DVDD.n4350 0.0162646
R4263 DVDD.n8625 DVDD.n8624 0.0162646
R4264 DVDD.n13832 DVDD.n11224 0.016049
R4265 DVDD.n2486 DVDD.n2485 0.016049
R4266 DVDD.n870 DVDD.n869 0.0157362
R4267 DVDD.n12580 DVDD.n12579 0.0155982
R4268 DVDD.n4350 DVDD.n4349 0.0155982
R4269 DVDD.n8624 DVDD.n8623 0.0155982
R4270 DVDD.n19464 DVDD.n3822 0.015575
R4271 DVDD.n19464 DVDD.n19005 0.015575
R4272 DVDD.n7301 DVDD.n7225 0.015575
R4273 DVDD.n18333 DVDD.n10085 0.015575
R4274 DVDD.n7662 DVDD.n7635 0.015575
R4275 DVDD.n18333 DVDD.n7130 0.015575
R4276 DVDD.n7662 DVDD.n7659 0.015575
R4277 DVDD.n20215 DVDD.n1821 0.015575
R4278 DVDD.n20215 DVDD.n2832 0.015575
R4279 DVDD.n20338 DVDD.n20301 0.015575
R4280 DVDD.n20338 DVDD.n20323 0.015575
R4281 DVDD.n14882 DVDD.n14858 0.015575
R4282 DVDD.n15104 DVDD.n15084 0.015575
R4283 DVDD.n10716 DVDD.n10702 0.015575
R4284 DVDD.n10633 DVDD.n10608 0.015575
R4285 DVDD.n7301 DVDD.n7296 0.015575
R4286 DVDD.n18981 DVDD.n18980 0.0153088
R4287 DVDD.n7207 DVDD.n7206 0.0153088
R4288 DVDD.n7208 DVDD.n7207 0.0153088
R4289 DVDD.n7209 DVDD.n7208 0.0153088
R4290 DVDD.n7214 DVDD.n7213 0.0153088
R4291 DVDD.n7213 DVDD.n7212 0.0153088
R4292 DVDD.n7212 DVDD.n7211 0.0153088
R4293 DVDD.n3840 DVDD.n3839 0.0153088
R4294 DVDD.n7601 DVDD.n7600 0.0153088
R4295 DVDD.n7602 DVDD.n7601 0.0153088
R4296 DVDD.n7603 DVDD.n7602 0.0153088
R4297 DVDD.n7608 DVDD.n7607 0.0153088
R4298 DVDD.n7607 DVDD.n7606 0.0153088
R4299 DVDD.n7606 DVDD.n7605 0.0153088
R4300 DVDD.n125 DVDD.n124 0.0153088
R4301 DVDD.n20310 DVDD.n20309 0.0153088
R4302 DVDD.n20311 DVDD.n20310 0.0153088
R4303 DVDD.n20312 DVDD.n20311 0.0153088
R4304 DVDD.n20307 DVDD.n20306 0.0153088
R4305 DVDD.n20306 DVDD.n20305 0.0153088
R4306 DVDD.n20305 DVDD.n20304 0.0153088
R4307 DVDD.n10548 DVDD.n10547 0.0153088
R4308 DVDD.n10657 DVDD.n10656 0.0153088
R4309 DVDD.n10658 DVDD.n10657 0.0153088
R4310 DVDD.n10659 DVDD.n10658 0.0153088
R4311 DVDD.n10664 DVDD.n10663 0.0153088
R4312 DVDD.n10663 DVDD.n10662 0.0153088
R4313 DVDD.n10662 DVDD.n10661 0.0153088
R4314 DVDD.n13919 DVDD.n13918 0.0150946
R4315 DVDD.n14308 DVDD.n14307 0.0150946
R4316 DVDD.n8136 DVDD.n8135 0.0149979
R4317 DVDD.n5666 DVDD.n5665 0.0149
R4318 DVDD.n12419 DVDD.n12418 0.0149
R4319 DVDD.n5573 DVDD.n5572 0.0149
R4320 DVDD.n8439 DVDD.n8438 0.0149
R4321 DVDD.n5590 DVDD.n5589 0.0148504
R4322 DVDD.n12837 DVDD.n12836 0.0148504
R4323 DVDD.n6217 DVDD.n6216 0.0148504
R4324 DVDD.n8919 DVDD.n8918 0.0148504
R4325 DVDD.n17689 DVDD.n17688 0.0147488
R4326 DVDD.n7201 DVDD.n7200 0.0147
R4327 DVDD.n7202 DVDD.n7201 0.0147
R4328 DVDD.n7203 DVDD.n7202 0.0147
R4329 DVDD.n7346 DVDD.n7345 0.0147
R4330 DVDD.n7345 DVDD.n7344 0.0147
R4331 DVDD.n7344 DVDD.n7343 0.0147
R4332 DVDD.n7555 DVDD.n7554 0.0147
R4333 DVDD.n7556 DVDD.n7555 0.0147
R4334 DVDD.n7557 DVDD.n7556 0.0147
R4335 DVDD.n7516 DVDD.n7515 0.0147
R4336 DVDD.n7515 DVDD.n7514 0.0147
R4337 DVDD.n7514 DVDD.n7513 0.0147
R4338 DVDD.n7667 DVDD.n7666 0.0147
R4339 DVDD.n7668 DVDD.n7667 0.0147
R4340 DVDD.n7669 DVDD.n7668 0.0147
R4341 DVDD.n7673 DVDD.n7672 0.0147
R4342 DVDD.n7672 DVDD.n7671 0.0147
R4343 DVDD.n7671 DVDD.n7670 0.0147
R4344 DVDD.n7428 DVDD.n7427 0.0147
R4345 DVDD.n7429 DVDD.n7428 0.0147
R4346 DVDD.n7430 DVDD.n7429 0.0147
R4347 DVDD.n7434 DVDD.n7433 0.0147
R4348 DVDD.n7433 DVDD.n7432 0.0147
R4349 DVDD.n7432 DVDD.n7431 0.0147
R4350 DVDD.n30 DVDD.n29 0.0147
R4351 DVDD.n31 DVDD.n30 0.0147
R4352 DVDD.n32 DVDD.n31 0.0147
R4353 DVDD.n28 DVDD.n27 0.0147
R4354 DVDD.n27 DVDD.n26 0.0147
R4355 DVDD.n26 DVDD.n25 0.0147
R4356 DVDD.n15137 DVDD.n15136 0.0147
R4357 DVDD.n15138 DVDD.n15137 0.0147
R4358 DVDD.n15139 DVDD.n15138 0.0147
R4359 DVDD.n15146 DVDD.n15145 0.0147
R4360 DVDD.n15145 DVDD.n15144 0.0147
R4361 DVDD.n15144 DVDD.n15143 0.0147
R4362 DVDD.n10207 DVDD.n10206 0.0147
R4363 DVDD.n10208 DVDD.n10207 0.0147
R4364 DVDD.n10209 DVDD.n10208 0.0147
R4365 DVDD.n10217 DVDD.n10216 0.0147
R4366 DVDD.n10216 DVDD.n10215 0.0147
R4367 DVDD.n10215 DVDD.n10214 0.0147
R4368 DVDD.n20218 DVDD.n20217 0.0147
R4369 DVDD.n20219 DVDD.n20218 0.0147
R4370 DVDD.n20220 DVDD.n20219 0.0147
R4371 DVDD.n20224 DVDD.n20223 0.0147
R4372 DVDD.n20223 DVDD.n20222 0.0147
R4373 DVDD.n20222 DVDD.n20221 0.0147
R4374 DVDD.n17297 DVDD.n17266 0.0146892
R4375 DVDD.n17676 DVDD.n17644 0.0146892
R4376 DVDD.n3114 DVDD.n3113 0.0145625
R4377 DVDD.n3098 DVDD.n3097 0.0145625
R4378 DVDD.n3091 DVDD.n3090 0.0145625
R4379 DVDD.n3077 DVDD.n3076 0.0145625
R4380 DVDD.n3071 DVDD.n3070 0.0145625
R4381 DVDD.n3062 DVDD.n3061 0.0145625
R4382 DVDD.n3053 DVDD.n3052 0.0145625
R4383 DVDD.n15121 DVDD.n15120 0.0144331
R4384 DVDD.n18975 DVDD.n18974 0.0143702
R4385 DVDD.n18985 DVDD.n18984 0.0143702
R4386 DVDD.n3827 DVDD.n3826 0.0143702
R4387 DVDD.n3834 DVDD.n3833 0.0143702
R4388 DVDD.n112 DVDD.n111 0.0143702
R4389 DVDD.n119 DVDD.n118 0.0143702
R4390 DVDD.n10542 DVDD.n10541 0.0143702
R4391 DVDD.n10552 DVDD.n10551 0.0143702
R4392 DVDD.n18977 DVDD.n18976 0.0142659
R4393 DVDD.n10544 DVDD.n10543 0.0142659
R4394 DVDD.n5107 DVDD.n5106 0.0141977
R4395 DVDD.n5389 DVDD.n5388 0.0141977
R4396 DVDD.n11648 DVDD.n11647 0.0141977
R4397 DVDD.n13072 DVDD.n13071 0.0141977
R4398 DVDD.n6575 DVDD.n6574 0.0141977
R4399 DVDD.n6372 DVDD.n6371 0.0141977
R4400 DVDD.n9543 DVDD.n9542 0.0141977
R4401 DVDD.n9158 DVDD.n9157 0.0141977
R4402 DVDD.n18983 DVDD.n18982 0.0141616
R4403 DVDD.n3836 DVDD.n3835 0.0141616
R4404 DVDD.n121 DVDD.n120 0.0141616
R4405 DVDD.n10550 DVDD.n10549 0.0141616
R4406 DVDD.n2802 DVDD.n2801 0.0141417
R4407 DVDD.n18570 DVDD.n18569 0.0141417
R4408 DVDD.n18672 DVDD.n18671 0.0141417
R4409 DVDD.n18475 DVDD.n18474 0.0141417
R4410 DVDD.n10061 DVDD.n10060 0.0141417
R4411 DVDD.n14810 DVDD.n14809 0.0141417
R4412 DVDD.n3862 DVDD.n3861 0.0141417
R4413 DVDD.n10109 DVDD.n10108 0.0141417
R4414 DVDD.n834 DVDD.n833 0.0141417
R4415 DVDD.n239 DVDD.n238 0.0141417
R4416 DVDD.n151 DVDD.n150 0.0141417
R4417 DVDD.n19171 DVDD.n19170 0.0141417
R4418 DVDD.n10093 DVDD.n10092 0.0141417
R4419 DVDD.n18228 DVDD.n18227 0.0141417
R4420 DVDD.n7083 DVDD.n7082 0.0141417
R4421 DVDD.n7141 DVDD.n7140 0.0141417
R4422 DVDD.n14321 DVDD.n14320 0.0140824
R4423 DVDD.n3825 DVDD.n3824 0.0140574
R4424 DVDD.n110 DVDD.n109 0.0140574
R4425 DVDD.n5170 DVDD.n5169 0.0138437
R4426 DVDD.n12351 DVDD.n12350 0.0138437
R4427 DVDD.n6512 DVDD.n6511 0.0138437
R4428 DVDD.n8371 DVDD.n8370 0.0138437
R4429 DVDD.n3083 DVDD.n3082 0.0137589
R4430 DVDD.n3829 DVDD.n3828 0.0137445
R4431 DVDD.n114 DVDD.n113 0.0137445
R4432 DVDD.n5542 DVDD.n5503 0.0137198
R4433 DVDD.n6254 DVDD.n6253 0.0137198
R4434 DVDD.n12957 DVDD.n12935 0.0137065
R4435 DVDD.n12957 DVDD.n12954 0.0137065
R4436 DVDD.n5522 DVDD.n5519 0.0137065
R4437 DVDD.n5525 DVDD.n5522 0.0137065
R4438 DVDD.n4020 DVDD.n4017 0.0137065
R4439 DVDD.n4023 DVDD.n4020 0.0137065
R4440 DVDD.n8976 DVDD.n8973 0.0137065
R4441 DVDD.n8979 DVDD.n8976 0.0137065
R4442 DVDD.n12899 DVDD.n12896 0.0137065
R4443 DVDD.n12896 DVDD.n12895 0.0137065
R4444 DVDD.n6068 DVDD.n6065 0.0137065
R4445 DVDD.n4518 DVDD.n4515 0.0137065
R4446 DVDD.n9003 DVDD.n9000 0.0137065
R4447 DVDD.n9006 DVDD.n9003 0.0137065
R4448 DVDD.n8266 DVDD.n8265 0.0136799
R4449 DVDD.n8260 DVDD.n8259 0.0136799
R4450 DVDD.n8203 DVDD.n8202 0.0136799
R4451 DVDD.n8197 DVDD.n8196 0.0136799
R4452 DVDD.n8339 DVDD.n8338 0.0136799
R4453 DVDD.n8333 DVDD.n8332 0.0136799
R4454 DVDD.n8303 DVDD.n8302 0.0136799
R4455 DVDD.n7961 DVDD.n7960 0.0136799
R4456 DVDD.n7986 DVDD.n7985 0.0136799
R4457 DVDD.n7995 DVDD.n7994 0.0136799
R4458 DVDD.n8025 DVDD.n8024 0.0136799
R4459 DVDD.n8050 DVDD.n8049 0.0136799
R4460 DVDD.n8059 DVDD.n8058 0.0136799
R4461 DVDD.n18987 DVDD.n18986 0.0136402
R4462 DVDD.n10554 DVDD.n10553 0.0136402
R4463 DVDD.n3105 DVDD.n3104 0.013558
R4464 DVDD.n9441 DVDD.n9440 0.0134916
R4465 DVDD.n9439 DVDD.n9438 0.0134916
R4466 DVDD.n5394 DVDD.n5393 0.0134897
R4467 DVDD.n13084 DVDD.n13083 0.0134897
R4468 DVDD.n13067 DVDD.n13066 0.0134897
R4469 DVDD.n6385 DVDD.n6384 0.0134897
R4470 DVDD.n6367 DVDD.n6366 0.0134897
R4471 DVDD.n9171 DVDD.n9170 0.0134897
R4472 DVDD.n9153 DVDD.n9152 0.0134897
R4473 DVDD.n20000 DVDD.n19999 0.0134331
R4474 DVDD.n1688 DVDD.n1687 0.0134331
R4475 DVDD.n2221 DVDD.n2220 0.0134331
R4476 DVDD.n3561 DVDD.n3560 0.0134331
R4477 DVDD.n17236 DVDD.n17234 0.0134255
R4478 DVDD.n17234 DVDD.n17232 0.0134255
R4479 DVDD.n17232 DVDD.n17230 0.0134255
R4480 DVDD.n17230 DVDD.n17228 0.0134255
R4481 DVDD.n17228 DVDD.n17226 0.0134255
R4482 DVDD.n17226 DVDD.n17224 0.0134255
R4483 DVDD.n17224 DVDD.n17222 0.0134255
R4484 DVDD.n17222 DVDD.n17220 0.0134255
R4485 DVDD.n17216 DVDD.n17214 0.0134255
R4486 DVDD.n17214 DVDD.n17212 0.0134255
R4487 DVDD.n17212 DVDD.n17210 0.0134255
R4488 DVDD.n17210 DVDD.n17208 0.0134255
R4489 DVDD.n17208 DVDD.n17206 0.0134255
R4490 DVDD.n17206 DVDD.n17204 0.0134255
R4491 DVDD.n17204 DVDD.n17202 0.0134255
R4492 DVDD.n17202 DVDD.n17200 0.0134255
R4493 DVDD.n4200 DVDD.n4198 0.0134255
R4494 DVDD.n4206 DVDD.n4200 0.0134255
R4495 DVDD.n4206 DVDD.n4204 0.0134255
R4496 DVDD.n4204 DVDD.n4202 0.0134255
R4497 DVDD.n4287 DVDD.n4281 0.0134255
R4498 DVDD.n4287 DVDD.n4285 0.0134255
R4499 DVDD.n4285 DVDD.n4283 0.0134255
R4500 DVDD.n14072 DVDD.n14070 0.0134255
R4501 DVDD.n14074 DVDD.n14072 0.0134255
R4502 DVDD.n14076 DVDD.n14074 0.0134255
R4503 DVDD.n14078 DVDD.n14076 0.0134255
R4504 DVDD.n14080 DVDD.n14078 0.0134255
R4505 DVDD.n14082 DVDD.n14080 0.0134255
R4506 DVDD.n14084 DVDD.n14082 0.0134255
R4507 DVDD.n14086 DVDD.n14084 0.0134255
R4508 DVDD.n17403 DVDD.n17401 0.0134255
R4509 DVDD.n17401 DVDD.n17399 0.0134255
R4510 DVDD.n17399 DVDD.n17397 0.0134255
R4511 DVDD.n17397 DVDD.n17395 0.0134255
R4512 DVDD.n17395 DVDD.n17393 0.0134255
R4513 DVDD.n17393 DVDD.n17391 0.0134255
R4514 DVDD.n17391 DVDD.n17389 0.0134255
R4515 DVDD.n17389 DVDD.n17387 0.0134255
R4516 DVDD.n17383 DVDD.n17381 0.0134255
R4517 DVDD.n17381 DVDD.n17379 0.0134255
R4518 DVDD.n17379 DVDD.n17377 0.0134255
R4519 DVDD.n17377 DVDD.n17375 0.0134255
R4520 DVDD.n17375 DVDD.n17373 0.0134255
R4521 DVDD.n17373 DVDD.n17371 0.0134255
R4522 DVDD.n17371 DVDD.n17369 0.0134255
R4523 DVDD.n17369 DVDD.n17367 0.0134255
R4524 DVDD.n4212 DVDD.n4210 0.0134255
R4525 DVDD.n4218 DVDD.n4212 0.0134255
R4526 DVDD.n4218 DVDD.n4216 0.0134255
R4527 DVDD.n4216 DVDD.n4214 0.0134255
R4528 DVDD.n4262 DVDD.n4256 0.0134255
R4529 DVDD.n4262 DVDD.n4260 0.0134255
R4530 DVDD.n4260 DVDD.n4258 0.0134255
R4531 DVDD.n13983 DVDD.n13981 0.0134255
R4532 DVDD.n13985 DVDD.n13983 0.0134255
R4533 DVDD.n13987 DVDD.n13985 0.0134255
R4534 DVDD.n13989 DVDD.n13987 0.0134255
R4535 DVDD.n13991 DVDD.n13989 0.0134255
R4536 DVDD.n13993 DVDD.n13991 0.0134255
R4537 DVDD.n13995 DVDD.n13993 0.0134255
R4538 DVDD.n13997 DVDD.n13995 0.0134255
R4539 DVDD.n17583 DVDD.n17582 0.0134255
R4540 DVDD.n17582 DVDD.n17579 0.0134255
R4541 DVDD.n17579 DVDD.n17578 0.0134255
R4542 DVDD.n17578 DVDD.n17575 0.0134255
R4543 DVDD.n17575 DVDD.n17574 0.0134255
R4544 DVDD.n17574 DVDD.n17571 0.0134255
R4545 DVDD.n17571 DVDD.n17570 0.0134255
R4546 DVDD.n17570 DVDD.n17567 0.0134255
R4547 DVDD.n17563 DVDD.n17562 0.0134255
R4548 DVDD.n17562 DVDD.n17559 0.0134255
R4549 DVDD.n17559 DVDD.n17558 0.0134255
R4550 DVDD.n17558 DVDD.n17555 0.0134255
R4551 DVDD.n17555 DVDD.n17554 0.0134255
R4552 DVDD.n17554 DVDD.n17551 0.0134255
R4553 DVDD.n17551 DVDD.n17550 0.0134255
R4554 DVDD.n17550 DVDD.n17547 0.0134255
R4555 DVDD.n4185 DVDD.n4182 0.0134255
R4556 DVDD.n4194 DVDD.n4185 0.0134255
R4557 DVDD.n4194 DVDD.n4193 0.0134255
R4558 DVDD.n4193 DVDD.n4190 0.0134255
R4559 DVDD.n4316 DVDD.n4307 0.0134255
R4560 DVDD.n4316 DVDD.n4315 0.0134255
R4561 DVDD.n4315 DVDD.n4312 0.0134255
R4562 DVDD.n14183 DVDD.n14180 0.0134255
R4563 DVDD.n14186 DVDD.n14183 0.0134255
R4564 DVDD.n14189 DVDD.n14186 0.0134255
R4565 DVDD.n14192 DVDD.n14189 0.0134255
R4566 DVDD.n14195 DVDD.n14192 0.0134255
R4567 DVDD.n14198 DVDD.n14195 0.0134255
R4568 DVDD.n14201 DVDD.n14198 0.0134255
R4569 DVDD.n14204 DVDD.n14201 0.0134255
R4570 DVDD.n3044 DVDD.n3043 0.0133571
R4571 DVDD.n18979 DVDD.n18978 0.0133273
R4572 DVDD.n10546 DVDD.n10545 0.0133273
R4573 DVDD.n3822 DVDD.n3821 0.013325
R4574 DVDD.n19005 DVDD.n19004 0.013325
R4575 DVDD.n10085 DVDD.n10084 0.013325
R4576 DVDD.n7130 DVDD.n7129 0.013325
R4577 DVDD.n1821 DVDD.n1820 0.013325
R4578 DVDD.n2832 DVDD.n2831 0.013325
R4579 DVDD.n14858 DVDD.n14857 0.013325
R4580 DVDD.n10608 DVDD.n10607 0.013325
R4581 DVDD.n5327 DVDD.n5326 0.0133126
R4582 DVDD.n5444 DVDD.n5443 0.0133126
R4583 DVDD.n13132 DVDD.n13131 0.0133126
R4584 DVDD.n13019 DVDD.n13018 0.0133126
R4585 DVDD.n6434 DVDD.n6433 0.0133126
R4586 DVDD.n6317 DVDD.n6316 0.0133126
R4587 DVDD.n9220 DVDD.n9219 0.0133126
R4588 DVDD.n9103 DVDD.n9102 0.0133126
R4589 DVDD.n8081 DVDD.n8080 0.0133033
R4590 DVDD.n15130 DVDD.n15129 0.0132748
R4591 DVDD.n15975 DVDD.n15974 0.0132384
R4592 DVDD.n16067 DVDD.n15951 0.0132384
R4593 DVDD.n15692 DVDD.n15678 0.0132384
R4594 DVDD.n9407 DVDD.n9406 0.0132384
R4595 DVDD.n8123 DVDD.n8122 0.0132384
R4596 DVDD.n3838 DVDD.n3837 0.0132231
R4597 DVDD.n123 DVDD.n122 0.0132231
R4598 DVDD.n11655 DVDD.n11654 0.0131355
R4599 DVDD.n13112 DVDD.n13111 0.0131355
R4600 DVDD.n6583 DVDD.n6582 0.0131355
R4601 DVDD.n6413 DVDD.n6412 0.0131355
R4602 DVDD.n9551 DVDD.n9550 0.0131355
R4603 DVDD.n9199 DVDD.n9198 0.0131355
R4604 DVDD.n8017 DVDD.n8016 0.0131151
R4605 DVDD.n5036 DVDD.n5035 0.0130787
R4606 DVDD.n5638 DVDD.n5637 0.0130787
R4607 DVDD.n11718 DVDD.n11717 0.0130787
R4608 DVDD.n12799 DVDD.n12798 0.0130787
R4609 DVDD.n6648 DVDD.n6647 0.0130787
R4610 DVDD.n6179 DVDD.n6178 0.0130787
R4611 DVDD.n9616 DVDD.n9615 0.0130787
R4612 DVDD.n8881 DVDD.n8880 0.0130787
R4613 DVDD.n15974 DVDD.n15973 0.0129857
R4614 DVDD.n16067 DVDD.n16066 0.0129857
R4615 DVDD.n15692 DVDD.n15691 0.0129857
R4616 DVDD.n9406 DVDD.n9405 0.0129857
R4617 DVDD.n8122 DVDD.n8121 0.0129857
R4618 DVDD.n13039 DVDD.n13038 0.0129585
R4619 DVDD.n6338 DVDD.n6337 0.0129585
R4620 DVDD.n9124 DVDD.n9123 0.0129585
R4621 DVDD.n8288 DVDD.n8287 0.0129268
R4622 DVDD.n7953 DVDD.n7952 0.0129268
R4623 DVDD.n8041 DVDD.n8040 0.0129268
R4624 DVDD.n8100 DVDD.n8099 0.0129044
R4625 DVDD.n1235 DVDD.n1234 0.0129016
R4626 DVDD.n1219 DVDD.n1218 0.0129016
R4627 DVDD.n1212 DVDD.n1211 0.0129016
R4628 DVDD.n1197 DVDD.n1196 0.0129016
R4629 DVDD.n1191 DVDD.n1190 0.0129016
R4630 DVDD.n1183 DVDD.n1182 0.0129016
R4631 DVDD.n1175 DVDD.n1174 0.0129016
R4632 DVDD.n1571 DVDD.n1570 0.0129016
R4633 DVDD.n1578 DVDD.n1577 0.0129016
R4634 DVDD.n1585 DVDD.n1584 0.0129016
R4635 DVDD.n1593 DVDD.n1592 0.0129016
R4636 DVDD.n1601 DVDD.n1600 0.0129016
R4637 DVDD.n1607 DVDD.n1606 0.0129016
R4638 DVDD.n1613 DVDD.n1612 0.0129016
R4639 DVDD.n1620 DVDD.n1619 0.0129016
R4640 DVDD.n1627 DVDD.n1626 0.0129016
R4641 DVDD.n1634 DVDD.n1633 0.0129016
R4642 DVDD.n1655 DVDD.n1654 0.0129016
R4643 DVDD.n1648 DVDD.n1647 0.0129016
R4644 DVDD.n924 DVDD.n923 0.0129016
R4645 DVDD.n917 DVDD.n916 0.0129016
R4646 DVDD.n910 DVDD.n909 0.0129016
R4647 DVDD.n905 DVDD.n904 0.0129016
R4648 DVDD.n900 DVDD.n899 0.0129016
R4649 DVDD.n893 DVDD.n892 0.0129016
R4650 DVDD.n886 DVDD.n885 0.0129016
R4651 DVDD.n879 DVDD.n878 0.0129016
R4652 DVDD.n19284 DVDD.n19283 0.0129016
R4653 DVDD.n19291 DVDD.n19290 0.0129016
R4654 DVDD.n19296 DVDD.n19295 0.0129016
R4655 DVDD.n19308 DVDD.n19307 0.0129016
R4656 DVDD.n19338 DVDD.n19337 0.0129016
R4657 DVDD.n10176 DVDD.n10175 0.0129016
R4658 DVDD.n10181 DVDD.n10180 0.0129016
R4659 DVDD.n11428 DVDD.n11427 0.0129016
R4660 DVDD.n11435 DVDD.n11434 0.0129016
R4661 DVDD.n12016 DVDD.n12015 0.0129016
R4662 DVDD.n12041 DVDD.n12040 0.0129016
R4663 DVDD.n12049 DVDD.n12048 0.0129016
R4664 DVDD.n12082 DVDD.n12081 0.0129016
R4665 DVDD.n12107 DVDD.n12106 0.0129016
R4666 DVDD.n12115 DVDD.n12114 0.0129016
R4667 DVDD.n13326 DVDD.n13325 0.0129016
R4668 DVDD.n13332 DVDD.n13331 0.0129016
R4669 DVDD.n13365 DVDD.n13364 0.0129016
R4670 DVDD.n13405 DVDD.n13404 0.0129016
R4671 DVDD.n13411 DVDD.n13410 0.0129016
R4672 DVDD.n13471 DVDD.n13470 0.0129016
R4673 DVDD.n13477 DVDD.n13476 0.0129016
R4674 DVDD.n19727 DVDD.n19726 0.0128699
R4675 DVDD.n1372 DVDD.n1371 0.0128699
R4676 DVDD.n1391 DVDD.n1390 0.0128699
R4677 DVDD.n1949 DVDD.n1948 0.0128699
R4678 DVDD.n1968 DVDD.n1967 0.0128699
R4679 DVDD.n3231 DVDD.n3230 0.0128699
R4680 DVDD.n3212 DVDD.n3211 0.0128699
R4681 DVDD.n3831 DVDD.n3830 0.0128059
R4682 DVDD.n116 DVDD.n115 0.0128059
R4683 DVDD.n8225 DVDD.n8224 0.0127385
R4684 DVDD.n7977 DVDD.n7976 0.0127385
R4685 DVDD.n12928 DVDD.n12927 0.0127283
R4686 DVDD.n12947 DVDD.n12946 0.0127283
R4687 DVDD.n5512 DVDD.n5511 0.0127283
R4688 DVDD.n5538 DVDD.n5537 0.0127283
R4689 DVDD.n4010 DVDD.n4009 0.0127283
R4690 DVDD.n4033 DVDD.n4032 0.0127283
R4691 DVDD.n8966 DVDD.n8965 0.0127283
R4692 DVDD.n9035 DVDD.n9034 0.0127283
R4693 DVDD.n12907 DVDD.n12904 0.0127283
R4694 DVDD.n12888 DVDD.n12887 0.0127283
R4695 DVDD.n5716 DVDD.n5715 0.0127283
R4696 DVDD.n6058 DVDD.n6057 0.0127283
R4697 DVDD.n4087 DVDD.n4086 0.0127283
R4698 DVDD.n4501 DVDD.n4500 0.0127283
R4699 DVDD.n8993 DVDD.n8992 0.0127283
R4700 DVDD.n9014 DVDD.n9011 0.0127283
R4701 DVDD.n19324 DVDD.n19323 0.0127244
R4702 DVDD.n11442 DVDD.n11441 0.0127244
R4703 DVDD.n12246 DVDD.n12245 0.0127244
R4704 DVDD.n12244 DVDD.n12243 0.0127244
R4705 DVDD.n19852 DVDD.n19851 0.0127244
R4706 DVDD.n1524 DVDD.n1523 0.0127244
R4707 DVDD.n2074 DVDD.n2073 0.0127244
R4708 DVDD.n3473 DVDD.n3472 0.0127244
R4709 DVDD.n18989 DVDD.n18988 0.0127016
R4710 DVDD.n10556 DVDD.n10555 0.0127016
R4711 DVDD.n19893 DVDD.n19892 0.0126928
R4712 DVDD.n1484 DVDD.n1483 0.0126928
R4713 DVDD.n2114 DVDD.n2113 0.0126928
R4714 DVDD.n3513 DVDD.n3512 0.0126928
R4715 DVDD.n4976 DVDD.n4975 0.0126042
R4716 DVDD.n11645 DVDD.n11644 0.0126042
R4717 DVDD.n11777 DVDD.n11776 0.0126042
R4718 DVDD.n6865 DVDD.n6864 0.0126042
R4719 DVDD.n6708 DVDD.n6707 0.0126042
R4720 DVDD.n7901 DVDD.n7900 0.0126042
R4721 DVDD.n9676 DVDD.n9675 0.0126042
R4722 DVDD.n12212 DVDD.n12211 0.0125559
R4723 DVDD.n13544 DVDD.n13543 0.0125559
R4724 DVDD.n13624 DVDD.n13623 0.0125559
R4725 DVDD.n14490 DVDD.n14489 0.0125559
R4726 DVDD.n14577 DVDD.n14576 0.0125559
R4727 DVDD.n14660 DVDD.n14659 0.0125559
R4728 DVDD.n2737 DVDD.n2736 0.0125559
R4729 DVDD.n14715 DVDD.n14714 0.0125559
R4730 DVDD.n15517 DVDD.n14741 0.0125559
R4731 DVDD.n15482 DVDD.n15481 0.0125559
R4732 DVDD.n15388 DVDD.n14825 0.0125559
R4733 DVDD.n2778 DVDD.n2777 0.0125559
R4734 DVDD.n14632 DVDD.n14631 0.0125559
R4735 DVDD.n5558 DVDD.n5557 0.0125559
R4736 DVDD.n6086 DVDD.n6085 0.0125559
R4737 DVDD.n5210 DVDD.n5209 0.0125559
R4738 DVDD.n5042 DVDD.n5041 0.0125559
R4739 DVDD.n5885 DVDD.n5884 0.0125559
R4740 DVDD.n11712 DVDD.n11711 0.0125559
R4741 DVDD.n12390 DVDD.n12389 0.0125559
R4742 DVDD.n12718 DVDD.n12717 0.0125559
R4743 DVDD.n12859 DVDD.n12858 0.0125559
R4744 DVDD.n17736 DVDD.n17695 0.0125559
R4745 DVDD.n17692 DVDD.n17691 0.0125559
R4746 DVDD.n18016 DVDD.n18015 0.0125559
R4747 DVDD.n18068 DVDD.n18067 0.0125559
R4748 DVDD.n18094 DVDD.n18093 0.0125559
R4749 DVDD.n18127 DVDD.n18126 0.0125559
R4750 DVDD.n18212 DVDD.n18211 0.0125559
R4751 DVDD.n812 DVDD.n811 0.0125559
R4752 DVDD.n775 DVDD.n774 0.0125559
R4753 DVDD.n17990 DVDD.n17989 0.0125559
R4754 DVDD.n17937 DVDD.n17936 0.0125559
R4755 DVDD.n17857 DVDD.n17856 0.0125559
R4756 DVDD.n4378 DVDD.n4377 0.0125559
R4757 DVDD.n6472 DVDD.n6471 0.0125559
R4758 DVDD.n6642 DVDD.n6641 0.0125559
R4759 DVDD.n6238 DVDD.n6237 0.0125559
R4760 DVDD.n4536 DVDD.n4535 0.0125559
R4761 DVDD.n4402 DVDD.n4401 0.0125559
R4762 DVDD.n14381 DVDD.n14380 0.0125559
R4763 DVDD.n5943 DVDD.n5942 0.0125559
R4764 DVDD.n12606 DVDD.n12605 0.0125559
R4765 DVDD.n17759 DVDD.n17758 0.0125559
R4766 DVDD.n13728 DVDD.n13707 0.0125559
R4767 DVDD.n8652 DVDD.n8651 0.0125559
R4768 DVDD.n9610 DVDD.n9609 0.0125559
R4769 DVDD.n8940 DVDD.n8939 0.0125559
R4770 DVDD.n8411 DVDD.n8410 0.0125559
R4771 DVDD.n8803 DVDD.n8802 0.0125559
R4772 DVDD.n8676 DVDD.n8675 0.0125559
R4773 DVDD.n8251 DVDD.n8250 0.0125502
R4774 DVDD.n19277 DVDD.n19276 0.0125472
R4775 DVDD.n10171 DVDD.n10170 0.0125472
R4776 DVDD.n12139 DVDD.n12138 0.0125472
R4777 DVDD.n5011 DVDD.n5010 0.0125472
R4778 DVDD.n5699 DVDD.n5698 0.0125472
R4779 DVDD.n11743 DVDD.n11742 0.0125472
R4780 DVDD.n12742 DVDD.n12741 0.0125472
R4781 DVDD.n6673 DVDD.n6672 0.0125472
R4782 DVDD.n6124 DVDD.n6123 0.0125472
R4783 DVDD.n9641 DVDD.n9640 0.0125472
R4784 DVDD.n8826 DVDD.n8825 0.0125472
R4785 DVDD.n14064 DVDD.n14063 0.0124793
R4786 DVDD.n13967 DVDD.n13966 0.0124793
R4787 DVDD.n17460 DVDD.n17459 0.0124793
R4788 DVDD.n17344 DVDD.n17343 0.0124793
R4789 DVDD.n17503 DVDD.n17502 0.0124793
R4790 DVDD.n13528 DVDD.n13527 0.0124644
R4791 DVDD.n13580 DVDD.n13579 0.0124644
R4792 DVDD.n13661 DVDD.n13660 0.0124644
R4793 DVDD.n5641 DVDD.n5640 0.0124644
R4794 DVDD.n12796 DVDD.n12795 0.0124644
R4795 DVDD.n18175 DVDD.n18174 0.0124644
R4796 DVDD.n18031 DVDD.n18030 0.0124644
R4797 DVDD.n17901 DVDD.n17900 0.0124644
R4798 DVDD.n12358 DVDD.n12357 0.0124271
R4799 DVDD.n13139 DVDD.n13138 0.0124271
R4800 DVDD.n6504 DVDD.n6503 0.0124271
R4801 DVDD.n6442 DVDD.n6441 0.0124271
R4802 DVDD.n8379 DVDD.n8378 0.0124271
R4803 DVDD.n9228 DVDD.n9227 0.0124271
R4804 DVDD.n17185 DVDD.n17182 0.0124231
R4805 DVDD.n17817 DVDD.n17811 0.0124231
R4806 DVDD.n17817 DVDD.n17814 0.0124231
R4807 DVDD.n12484 DVDD.n12481 0.0124231
R4808 DVDD.n12661 DVDD.n12658 0.0124231
R4809 DVDD.n12667 DVDD.n12664 0.0124231
R4810 DVDD.n6007 DVDD.n6004 0.0124231
R4811 DVDD.n5998 DVDD.n5995 0.0124231
R4812 DVDD.n6016 DVDD.n6013 0.0124231
R4813 DVDD.n4109 DVDD.n4106 0.0124231
R4814 DVDD.n4461 DVDD.n4458 0.0124231
R4815 DVDD.n4100 DVDD.n4097 0.0124231
R4816 DVDD.n8744 DVDD.n8738 0.0124231
R4817 DVDD.n8744 DVDD.n8741 0.0124231
R4818 DVDD.n8753 DVDD.n8747 0.0124231
R4819 DVDD.n14439 DVDD.n14436 0.0124231
R4820 DVDD.n14448 DVDD.n14442 0.0124231
R4821 DVDD.n14448 DVDD.n14445 0.0124231
R4822 DVDD.n17708 DVDD.n17705 0.0124231
R4823 DVDD.n17711 DVDD.n17708 0.0124231
R4824 DVDD.n17735 DVDD.n17711 0.0124231
R4825 DVDD.n17735 DVDD.n17732 0.0124231
R4826 DVDD.n17732 DVDD.n17729 0.0124231
R4827 DVDD.n17723 DVDD.n17720 0.0124231
R4828 DVDD.n17720 DVDD.n17717 0.0124231
R4829 DVDD.n17717 DVDD.n17714 0.0124231
R4830 DVDD.n5892 DVDD.n5889 0.0124231
R4831 DVDD.n5895 DVDD.n5892 0.0124231
R4832 DVDD.n5919 DVDD.n5916 0.0124231
R4833 DVDD.n5916 DVDD.n5913 0.0124231
R4834 DVDD.n5913 DVDD.n5910 0.0124231
R4835 DVDD.n5910 DVDD.n5907 0.0124231
R4836 DVDD.n5907 DVDD.n5906 0.0124231
R4837 DVDD.n5906 DVDD.n5903 0.0124231
R4838 DVDD.n4361 DVDD.n4358 0.0124231
R4839 DVDD.n4376 DVDD.n4361 0.0124231
R4840 DVDD.n4376 DVDD.n4373 0.0124231
R4841 DVDD.n4373 DVDD.n4370 0.0124231
R4842 DVDD.n4370 DVDD.n4367 0.0124231
R4843 DVDD.n4367 DVDD.n4364 0.0124231
R4844 DVDD.n8635 DVDD.n8632 0.0124231
R4845 DVDD.n8650 DVDD.n8635 0.0124231
R4846 DVDD.n8650 DVDD.n8647 0.0124231
R4847 DVDD.n8647 DVDD.n8644 0.0124231
R4848 DVDD.n8644 DVDD.n8641 0.0124231
R4849 DVDD.n8641 DVDD.n8638 0.0124231
R4850 DVDD.n14355 DVDD.n14352 0.0124231
R4851 DVDD.n14352 DVDD.n14349 0.0124231
R4852 DVDD.n14349 DVDD.n14346 0.0124231
R4853 DVDD.n14346 DVDD.n14343 0.0124231
R4854 DVDD.n14343 DVDD.n14340 0.0124231
R4855 DVDD.n9042 DVDD.n9041 0.0123889
R4856 DVDD.n12073 DVDD.n12072 0.0123701
R4857 DVDD.n19927 DVDD.n19926 0.0123701
R4858 DVDD.n1450 DVDD.n1449 0.0123701
R4859 DVDD.n2148 DVDD.n2147 0.0123701
R4860 DVDD.n3547 DVDD.n3546 0.0123701
R4861 DVDD.n8188 DVDD.n8187 0.0123619
R4862 DVDD.n9453 DVDD.n9452 0.0123619
R4863 DVDD.n8311 DVDD.n8310 0.0123619
R4864 DVDD.n12211 DVDD.n12210 0.0123034
R4865 DVDD.n13625 DVDD.n13624 0.0123034
R4866 DVDD.n13728 DVDD.n13727 0.0123034
R4867 DVDD.n13543 DVDD.n13542 0.0123034
R4868 DVDD.n15389 DVDD.n15388 0.0123034
R4869 DVDD.n14631 DVDD.n14630 0.0123034
R4870 DVDD.n14659 DVDD.n14658 0.0123034
R4871 DVDD.n15517 DVDD.n15516 0.0123034
R4872 DVDD.n2777 DVDD.n2776 0.0123034
R4873 DVDD.n15481 DVDD.n15480 0.0123034
R4874 DVDD.n2736 DVDD.n2735 0.0123034
R4875 DVDD.n14714 DVDD.n14713 0.0123034
R4876 DVDD.n14578 DVDD.n14577 0.0123034
R4877 DVDD.n14489 DVDD.n14488 0.0123034
R4878 DVDD.n5211 DVDD.n5210 0.0123034
R4879 DVDD.n6085 DVDD.n6084 0.0123034
R4880 DVDD.n5942 DVDD.n5941 0.0123034
R4881 DVDD.n5041 DVDD.n5040 0.0123034
R4882 DVDD.n5886 DVDD.n5885 0.0123034
R4883 DVDD.n5557 DVDD.n5556 0.0123034
R4884 DVDD.n12391 DVDD.n12390 0.0123034
R4885 DVDD.n12605 DVDD.n12604 0.0123034
R4886 DVDD.n11713 DVDD.n11712 0.0123034
R4887 DVDD.n12860 DVDD.n12859 0.0123034
R4888 DVDD.n12717 DVDD.n12716 0.0123034
R4889 DVDD.n18211 DVDD.n18210 0.0123034
R4890 DVDD.n17989 DVDD.n17988 0.0123034
R4891 DVDD.n17856 DVDD.n17855 0.0123034
R4892 DVDD.n17758 DVDD.n17757 0.0123034
R4893 DVDD.n17693 DVDD.n17692 0.0123034
R4894 DVDD.n18015 DVDD.n18014 0.0123034
R4895 DVDD.n18067 DVDD.n18066 0.0123034
R4896 DVDD.n18093 DVDD.n18092 0.0123034
R4897 DVDD.n811 DVDD.n810 0.0123034
R4898 DVDD.n18128 DVDD.n18127 0.0123034
R4899 DVDD.n774 DVDD.n773 0.0123034
R4900 DVDD.n17737 DVDD.n17736 0.0123034
R4901 DVDD.n17938 DVDD.n17937 0.0123034
R4902 DVDD.n4535 DVDD.n4534 0.0123034
R4903 DVDD.n6643 DVDD.n6642 0.0123034
R4904 DVDD.n6471 DVDD.n6470 0.0123034
R4905 DVDD.n4377 DVDD.n4352 0.0123034
R4906 DVDD.n6239 DVDD.n6238 0.0123034
R4907 DVDD.n14380 DVDD.n14379 0.0123034
R4908 DVDD.n4401 DVDD.n4400 0.0123034
R4909 DVDD.n8412 DVDD.n8411 0.0123034
R4910 DVDD.n8802 DVDD.n8801 0.0123034
R4911 DVDD.n8675 DVDD.n8674 0.0123034
R4912 DVDD.n9611 DVDD.n9610 0.0123034
R4913 DVDD.n8651 DVDD.n8626 0.0123034
R4914 DVDD.n8941 DVDD.n8940 0.0123034
R4915 DVDD.n3364 DVDD.n3363 0.0122996
R4916 DVDD.n12203 DVDD.n12202 0.0122877
R4917 DVDD.n11750 DVDD.n11749 0.01225
R4918 DVDD.n6680 DVDD.n6679 0.01225
R4919 DVDD.n9648 DVDD.n9647 0.01225
R4920 DVDD.n5360 DVDD.n5359 0.0122499
R4921 DVDD.n5449 DVDD.n5448 0.0122499
R4922 DVDD.n13014 DVDD.n13013 0.0122499
R4923 DVDD.n6312 DVDD.n6311 0.0122499
R4924 DVDD.n9098 DVDD.n9097 0.0122499
R4925 DVDD.n14340 DVDD.n14337 0.0122308
R4926 DVDD.n18342 DVDD.n18341 0.0122
R4927 DVDD.n1203 DVDD.n1202 0.0121929
R4928 DVDD.n12007 DVDD.n12006 0.0121929
R4929 DVDD.n12098 DVDD.n12097 0.0121929
R4930 DVDD.n13381 DVDD.n13380 0.0121929
R4931 DVDD.n13060 DVDD.n13059 0.0120728
R4932 DVDD.n6359 DVDD.n6358 0.0120728
R4933 DVDD.n9145 DVDD.n9144 0.0120728
R4934 DVDD.n17182 DVDD.n17179 0.0120385
R4935 DVDD.n17705 DVDD.n17702 0.0120385
R4936 DVDD.n1226 DVDD.n1225 0.0120157
R4937 DVDD.n12032 DVDD.n12031 0.0120157
R4938 DVDD.n13447 DVDD.n13446 0.0120157
R4939 DVDD.n19760 DVDD.n19759 0.0120157
R4940 DVDD.n1405 DVDD.n1404 0.0120157
R4941 DVDD.n1982 DVDD.n1981 0.0120157
R4942 DVDD.n3198 DVDD.n3197 0.0120157
R4943 DVDD.n9434 DVDD.n9433 0.0119854
R4944 DVDD.n8348 DVDD.n8347 0.0119854
R4945 DVDD.n14059 DVDD.n14058 0.0119755
R4946 DVDD.n17339 DVDD.n17338 0.0119755
R4947 DVDD.n13962 DVDD.n13961 0.0119755
R4948 DVDD.n17498 DVDD.n17497 0.0119755
R4949 DVDD.n12581 DVDD.n12580 0.0119575
R4950 DVDD.n12582 DVDD.n12581 0.0119575
R4951 DVDD.n17694 DVDD.n17693 0.0119575
R4952 DVDD.n17695 DVDD.n17694 0.0119575
R4953 DVDD.n12182 DVDD.n12181 0.0119309
R4954 DVDD.n12181 DVDD.n12180 0.0119309
R4955 DVDD.n14357 DVDD.n14356 0.0119309
R4956 DVDD.n14326 DVDD.n14325 0.0119309
R4957 DVDD.n14324 DVDD.n14323 0.0119309
R4958 DVDD.n14325 DVDD.n14324 0.0119309
R4959 DVDD.n14356 DVDD.n14327 0.0119309
R4960 DVDD.n14327 DVDD.n14326 0.0119309
R4961 DVDD.n5921 DVDD.n5920 0.0119309
R4962 DVDD.n5884 DVDD.n5883 0.0119309
R4963 DVDD.n5883 DVDD.n5882 0.0119309
R4964 DVDD.n5920 DVDD.n5886 0.0119309
R4965 DVDD.n17455 DVDD.n17454 0.0118543
R4966 DVDD.n17597 DVDD.n17513 0.0118514
R4967 DVDD.n17257 DVDD.n17256 0.0118514
R4968 DVDD.n17414 DVDD.n17354 0.0118514
R4969 DVDD.n17298 DVDD.n17297 0.0118514
R4970 DVDD.n14118 DVDD.n14117 0.0118514
R4971 DVDD.n14020 DVDD.n14019 0.0118514
R4972 DVDD.n14019 DVDD.n13977 0.0118514
R4973 DVDD.n13920 DVDD.n13919 0.0118514
R4974 DVDD.n17256 DVDD.n17255 0.0118514
R4975 DVDD.n17415 DVDD.n17414 0.0118514
R4976 DVDD.n14309 DVDD.n14308 0.0118514
R4977 DVDD.n14232 DVDD.n14231 0.0118514
R4978 DVDD.n14231 DVDD.n14174 0.0118514
R4979 DVDD.n14119 DVDD.n14118 0.0118514
R4980 DVDD.n17677 DVDD.n17676 0.0118514
R4981 DVDD.n17598 DVDD.n17597 0.0118514
R4982 DVDD.n1166 DVDD.n1165 0.0118386
R4983 DVDD.n13420 DVDD.n13419 0.0118386
R4984 DVDD.n14449 DVDD.n14433 0.0118386
R4985 DVDD.n5467 DVDD.n5466 0.0118386
R4986 DVDD.n6017 DVDD.n5992 0.0118386
R4987 DVDD.n12996 DVDD.n12995 0.0118386
R4988 DVDD.n12668 DVDD.n12655 0.0118386
R4989 DVDD.n17818 DVDD.n17808 0.0118386
R4990 DVDD.n6294 DVDD.n6293 0.0118386
R4991 DVDD.n4468 DVDD.n4455 0.0118386
R4992 DVDD.n9080 DVDD.n9079 0.0118386
R4993 DVDD.n8754 DVDD.n8729 0.0118386
R4994 DVDD.n17256 DVDD.n17246 0.01175
R4995 DVDD.n17414 DVDD.n17413 0.01175
R4996 DVDD.n17597 DVDD.n17596 0.01175
R4997 DVDD.n12961 DVDD.n12960 0.0117224
R4998 DVDD.n4796 DVDD.n4795 0.0117185
R4999 DVDD.n11622 DVDD.n11621 0.0117185
R5000 DVDD.n6888 DVDD.n6887 0.0117185
R5001 DVDD.n7878 DVDD.n7877 0.0117185
R5002 DVDD.n12258 DVDD.n12257 0.0116614
R5003 DVDD.n13356 DVDD.n13355 0.0116614
R5004 DVDD.n13486 DVDD.n13485 0.0116614
R5005 DVDD.n14421 DVDD.n14420 0.0116614
R5006 DVDD.n20179 DVDD.n20178 0.0116614
R5007 DVDD.n20084 DVDD.n20083 0.0116614
R5008 DVDD.n5979 DVDD.n5978 0.0116614
R5009 DVDD.n257 DVDD.n256 0.0116614
R5010 DVDD.n19182 DVDD.n19181 0.0116614
R5011 DVDD.n12642 DVDD.n12641 0.0116614
R5012 DVDD.n17795 DVDD.n17794 0.0116614
R5013 DVDD.n19564 DVDD.n19563 0.0116614
R5014 DVDD.n19469 DVDD.n19468 0.0116614
R5015 DVDD.n4442 DVDD.n4441 0.0116614
R5016 DVDD.n3743 DVDD.n3742 0.0116614
R5017 DVDD.n18486 DVDD.n18485 0.0116614
R5018 DVDD.n8716 DVDD.n8715 0.0116614
R5019 DVDD.n7789 DVDD.n7788 0.01166
R5020 DVDD.n7788 DVDD.n7787 0.01166
R5021 DVDD.n7787 DVDD.n7786 0.01166
R5022 DVDD.n7786 DVDD.n7785 0.01166
R5023 DVDD.n7785 DVDD.n7784 0.01166
R5024 DVDD.n7784 DVDD.n7783 0.01166
R5025 DVDD.n7783 DVDD.n7782 0.01166
R5026 DVDD.n7782 DVDD.n7781 0.01166
R5027 DVDD.n7781 DVDD.n7780 0.01166
R5028 DVDD.n7780 DVDD.n7779 0.01166
R5029 DVDD.n7779 DVDD.n7778 0.01166
R5030 DVDD.n7778 DVDD.n7777 0.01166
R5031 DVDD.n7777 DVDD.n7776 0.01166
R5032 DVDD.n7776 DVDD.n7775 0.01166
R5033 DVDD.n7775 DVDD.n7774 0.01166
R5034 DVDD.n7774 DVDD.n7773 0.01166
R5035 DVDD.n7773 DVDD.n7772 0.01166
R5036 DVDD.n3006 DVDD.n3005 0.01166
R5037 DVDD.n3007 DVDD.n3006 0.01166
R5038 DVDD.n3008 DVDD.n3007 0.01166
R5039 DVDD.n3009 DVDD.n3008 0.01166
R5040 DVDD.n3010 DVDD.n3009 0.01166
R5041 DVDD.n3011 DVDD.n3010 0.01166
R5042 DVDD.n3012 DVDD.n3011 0.01166
R5043 DVDD.n3013 DVDD.n3012 0.01166
R5044 DVDD.n3014 DVDD.n3013 0.01166
R5045 DVDD.n3015 DVDD.n3014 0.01166
R5046 DVDD.n3016 DVDD.n3015 0.01166
R5047 DVDD.n3017 DVDD.n3016 0.01166
R5048 DVDD.n3018 DVDD.n3017 0.01166
R5049 DVDD.n3019 DVDD.n3018 0.01166
R5050 DVDD.n3020 DVDD.n3019 0.01166
R5051 DVDD.n3021 DVDD.n3020 0.01166
R5052 DVDD.n3022 DVDD.n3021 0.01166
R5053 DVDD.n3023 DVDD.n3022 0.01166
R5054 DVDD.n3024 DVDD.n3023 0.01166
R5055 DVDD.n3025 DVDD.n3024 0.01166
R5056 DVDD.n3026 DVDD.n3025 0.01166
R5057 DVDD.n3027 DVDD.n3026 0.01166
R5058 DVDD.n3447 DVDD.n3027 0.01166
R5059 DVDD.n2911 DVDD.n2910 0.01166
R5060 DVDD.n2910 DVDD.n2909 0.01166
R5061 DVDD.n2909 DVDD.n2908 0.01166
R5062 DVDD.n2908 DVDD.n2907 0.01166
R5063 DVDD.n2907 DVDD.n2906 0.01166
R5064 DVDD.n2906 DVDD.n2905 0.01166
R5065 DVDD.n2871 DVDD.n2870 0.01166
R5066 DVDD.n2870 DVDD.n2869 0.01166
R5067 DVDD.n2869 DVDD.n2868 0.01166
R5068 DVDD.n2868 DVDD.n2867 0.01166
R5069 DVDD.n3579 DVDD.n2867 0.01166
R5070 DVDD.n9931 DVDD.n9930 0.01166
R5071 DVDD.n9932 DVDD.n9931 0.01166
R5072 DVDD.n9933 DVDD.n9932 0.01166
R5073 DVDD.n9934 DVDD.n9933 0.01166
R5074 DVDD.n9935 DVDD.n9934 0.01166
R5075 DVDD.n9936 DVDD.n9935 0.01166
R5076 DVDD.n9937 DVDD.n9936 0.01166
R5077 DVDD.n9938 DVDD.n9937 0.01166
R5078 DVDD.n9939 DVDD.n9938 0.01166
R5079 DVDD.n9940 DVDD.n9939 0.01166
R5080 DVDD.n9941 DVDD.n9940 0.01166
R5081 DVDD.n9942 DVDD.n9941 0.01166
R5082 DVDD.n9943 DVDD.n9942 0.01166
R5083 DVDD.n9944 DVDD.n9943 0.01166
R5084 DVDD.n9945 DVDD.n9944 0.01166
R5085 DVDD.n9946 DVDD.n9945 0.01166
R5086 DVDD.n9947 DVDD.n9946 0.01166
R5087 DVDD.n9948 DVDD.n9947 0.01166
R5088 DVDD.n9949 DVDD.n9948 0.01166
R5089 DVDD.n9950 DVDD.n9949 0.01166
R5090 DVDD.n9951 DVDD.n9950 0.01166
R5091 DVDD.n9952 DVDD.n9951 0.01166
R5092 DVDD.n9953 DVDD.n9952 0.01166
R5093 DVDD.n9822 DVDD.n9821 0.01166
R5094 DVDD.n9821 DVDD.n9820 0.01166
R5095 DVDD.n9820 DVDD.n9819 0.01166
R5096 DVDD.n9493 DVDD.n9492 0.01166
R5097 DVDD.n9494 DVDD.n9493 0.01166
R5098 DVDD.n9495 DVDD.n9494 0.01166
R5099 DVDD.n9496 DVDD.n9495 0.01166
R5100 DVDD.n9497 DVDD.n9496 0.01166
R5101 DVDD.n9498 DVDD.n9497 0.01166
R5102 DVDD.n9499 DVDD.n9498 0.01166
R5103 DVDD.n9500 DVDD.n9499 0.01166
R5104 DVDD.n9501 DVDD.n9500 0.01166
R5105 DVDD.n9502 DVDD.n9501 0.01166
R5106 DVDD.n9503 DVDD.n9502 0.01166
R5107 DVDD.n9504 DVDD.n9503 0.01166
R5108 DVDD.n9505 DVDD.n9504 0.01166
R5109 DVDD.n9506 DVDD.n9505 0.01166
R5110 DVDD.n9507 DVDD.n9506 0.01166
R5111 DVDD.n9508 DVDD.n9507 0.01166
R5112 DVDD.n9509 DVDD.n9508 0.01166
R5113 DVDD.n9510 DVDD.n9509 0.01166
R5114 DVDD.n9511 DVDD.n9510 0.01166
R5115 DVDD.n9512 DVDD.n9511 0.01166
R5116 DVDD.n9513 DVDD.n9512 0.01166
R5117 DVDD.n9514 DVDD.n9513 0.01166
R5118 DVDD.n1084 DVDD.n1083 0.01166
R5119 DVDD.n1083 DVDD.n1082 0.01166
R5120 DVDD.n1082 DVDD.n1081 0.01166
R5121 DVDD.n1081 DVDD.n1080 0.01166
R5122 DVDD.n1080 DVDD.n1079 0.01166
R5123 DVDD.n1079 DVDD.n1078 0.01166
R5124 DVDD.n1078 DVDD.n1077 0.01166
R5125 DVDD.n1077 DVDD.n1076 0.01166
R5126 DVDD.n1076 DVDD.n1075 0.01166
R5127 DVDD.n1075 DVDD.n1074 0.01166
R5128 DVDD.n1074 DVDD.n1073 0.01166
R5129 DVDD.n1073 DVDD.n1072 0.01166
R5130 DVDD.n1072 DVDD.n1071 0.01166
R5131 DVDD.n1071 DVDD.n1070 0.01166
R5132 DVDD.n1070 DVDD.n1069 0.01166
R5133 DVDD.n1069 DVDD.n1068 0.01166
R5134 DVDD.n1068 DVDD.n1067 0.01166
R5135 DVDD.n1067 DVDD.n1066 0.01166
R5136 DVDD.n1066 DVDD.n1065 0.01166
R5137 DVDD.n1065 DVDD.n1064 0.01166
R5138 DVDD.n1064 DVDD.n1063 0.01166
R5139 DVDD.n1063 DVDD.n1062 0.01166
R5140 DVDD.n1549 DVDD.n1062 0.01166
R5141 DVDD.n1017 DVDD.n1016 0.01166
R5142 DVDD.n1018 DVDD.n1017 0.01166
R5143 DVDD.n1019 DVDD.n1018 0.01166
R5144 DVDD.n1020 DVDD.n1019 0.01166
R5145 DVDD.n1021 DVDD.n1020 0.01166
R5146 DVDD.n1022 DVDD.n1021 0.01166
R5147 DVDD.n1057 DVDD.n1056 0.01166
R5148 DVDD.n1058 DVDD.n1057 0.01166
R5149 DVDD.n1059 DVDD.n1058 0.01166
R5150 DVDD.n1060 DVDD.n1059 0.01166
R5151 DVDD.n1670 DVDD.n1060 0.01166
R5152 DVDD.n1754 DVDD.n1753 0.01166
R5153 DVDD.n11515 DVDD.n11514 0.01166
R5154 DVDD.n11516 DVDD.n11515 0.01166
R5155 DVDD.n11517 DVDD.n11516 0.01166
R5156 DVDD.n11518 DVDD.n11517 0.01166
R5157 DVDD.n11519 DVDD.n11518 0.01166
R5158 DVDD.n11520 DVDD.n11519 0.01166
R5159 DVDD.n11521 DVDD.n11520 0.01166
R5160 DVDD.n11522 DVDD.n11521 0.01166
R5161 DVDD.n11523 DVDD.n11522 0.01166
R5162 DVDD.n11524 DVDD.n11523 0.01166
R5163 DVDD.n11525 DVDD.n11524 0.01166
R5164 DVDD.n11526 DVDD.n11525 0.01166
R5165 DVDD.n11527 DVDD.n11526 0.01166
R5166 DVDD.n11528 DVDD.n11527 0.01166
R5167 DVDD.n11529 DVDD.n11528 0.01166
R5168 DVDD.n11530 DVDD.n11529 0.01166
R5169 DVDD.n11531 DVDD.n11530 0.01166
R5170 DVDD.n11532 DVDD.n11531 0.01166
R5171 DVDD.n11533 DVDD.n11532 0.01166
R5172 DVDD.n11534 DVDD.n11533 0.01166
R5173 DVDD.n11535 DVDD.n11534 0.01166
R5174 DVDD.n11536 DVDD.n11535 0.01166
R5175 DVDD.n11537 DVDD.n11536 0.01166
R5176 DVDD.n10145 DVDD.n10144 0.01166
R5177 DVDD.n10144 DVDD.n10143 0.01166
R5178 DVDD.n10143 DVDD.n10142 0.01166
R5179 DVDD.n10142 DVDD.n10141 0.01166
R5180 DVDD.n10141 DVDD.n10140 0.01166
R5181 DVDD.n10140 DVDD.n10139 0.01166
R5182 DVDD.n10139 DVDD.n10138 0.01166
R5183 DVDD.n10138 DVDD.n10137 0.01166
R5184 DVDD.n10137 DVDD.n10136 0.01166
R5185 DVDD.n10136 DVDD.n10135 0.01166
R5186 DVDD.n10135 DVDD.n10134 0.01166
R5187 DVDD.n10134 DVDD.n10133 0.01166
R5188 DVDD.n10133 DVDD.n10132 0.01166
R5189 DVDD.n10132 DVDD.n10131 0.01166
R5190 DVDD.n10131 DVDD.n10130 0.01166
R5191 DVDD.n10130 DVDD.n10129 0.01166
R5192 DVDD.n10129 DVDD.n10128 0.01166
R5193 DVDD.n11923 DVDD.n11922 0.01166
R5194 DVDD.n11922 DVDD.n11921 0.01166
R5195 DVDD.n11921 DVDD.n11920 0.01166
R5196 DVDD.n1274 DVDD.n1273 0.01166
R5197 DVDD.n1275 DVDD.n1274 0.01166
R5198 DVDD.n1276 DVDD.n1275 0.01166
R5199 DVDD.n1277 DVDD.n1276 0.01166
R5200 DVDD.n1278 DVDD.n1277 0.01166
R5201 DVDD.n1279 DVDD.n1278 0.01166
R5202 DVDD.n12298 DVDD.n12297 0.01166
R5203 DVDD.n12299 DVDD.n12298 0.01166
R5204 DVDD.n12300 DVDD.n12299 0.01166
R5205 DVDD.n12301 DVDD.n12300 0.01166
R5206 DVDD.n12302 DVDD.n12301 0.01166
R5207 DVDD.n12303 DVDD.n12302 0.01166
R5208 DVDD.n12304 DVDD.n12303 0.01166
R5209 DVDD.n12305 DVDD.n12304 0.01166
R5210 DVDD.n12306 DVDD.n12305 0.01166
R5211 DVDD.n12307 DVDD.n12306 0.01166
R5212 DVDD.n12308 DVDD.n12307 0.01166
R5213 DVDD.n12309 DVDD.n12308 0.01166
R5214 DVDD.n12310 DVDD.n12309 0.01166
R5215 DVDD.n12311 DVDD.n12310 0.01166
R5216 DVDD.n12312 DVDD.n12311 0.01166
R5217 DVDD.n12313 DVDD.n12312 0.01166
R5218 DVDD.n12314 DVDD.n12313 0.01166
R5219 DVDD.n12315 DVDD.n12314 0.01166
R5220 DVDD.n12316 DVDD.n12315 0.01166
R5221 DVDD.n12317 DVDD.n12316 0.01166
R5222 DVDD.n12318 DVDD.n12317 0.01166
R5223 DVDD.n12319 DVDD.n12318 0.01166
R5224 DVDD.n3124 DVDD.n3123 0.01166
R5225 DVDD.n3123 DVDD.n3122 0.01166
R5226 DVDD.n3122 DVDD.n3121 0.01166
R5227 DVDD.n3030 DVDD.n3029 0.01166
R5228 DVDD.n3324 DVDD.n3030 0.01166
R5229 DVDD.n2690 DVDD.n2689 0.0116222
R5230 DVDD.n8073 DVDD.n8072 0.0116088
R5231 DVDD.n9363 DVDD.n9362 0.01157
R5232 DVDD.n13274 DVDD.n13273 0.01157
R5233 DVDD.n10656 DVDD.n10655 0.0115186
R5234 DVDD.n14118 DVDD.n14096 0.0115106
R5235 DVDD.n14019 DVDD.n14007 0.0115106
R5236 DVDD.n14231 DVDD.n14217 0.0115106
R5237 DVDD.n19691 DVDD.n19690 0.0114843
R5238 DVDD.n19698 DVDD.n19697 0.0114843
R5239 DVDD.n19705 DVDD.n19704 0.0114843
R5240 DVDD.n19740 DVDD.n19739 0.0114843
R5241 DVDD.n19746 DVDD.n19745 0.0114843
R5242 DVDD.n19859 DVDD.n19858 0.0114843
R5243 DVDD.n19866 DVDD.n19865 0.0114843
R5244 DVDD.n19873 DVDD.n19872 0.0114843
R5245 DVDD.n19880 DVDD.n19879 0.0114843
R5246 DVDD.n19906 DVDD.n19905 0.0114843
R5247 DVDD.n19913 DVDD.n19912 0.0114843
R5248 DVDD.n20006 DVDD.n20005 0.0114843
R5249 DVDD.n20053 DVDD.n20052 0.0114843
R5250 DVDD.n20060 DVDD.n20059 0.0114843
R5251 DVDD.n20207 DVDD.n20206 0.0114843
R5252 DVDD.n20200 DVDD.n20199 0.0114843
R5253 DVDD.n20193 DVDD.n20192 0.0114843
R5254 DVDD.n20098 DVDD.n20097 0.0114843
R5255 DVDD.n20105 DVDD.n20104 0.0114843
R5256 DVDD.n20112 DVDD.n20111 0.0114843
R5257 DVDD.n19065 DVDD.n19064 0.0114843
R5258 DVDD.n19058 DVDD.n19057 0.0114843
R5259 DVDD.n19017 DVDD.n19016 0.0114843
R5260 DVDD.n4655 DVDD.n4654 0.0114843
R5261 DVDD.n4662 DVDD.n4661 0.0114843
R5262 DVDD.n4669 DVDD.n4668 0.0114843
R5263 DVDD.n4805 DVDD.n4804 0.0114843
R5264 DVDD.n4812 DVDD.n4811 0.0114843
R5265 DVDD.n4819 DVDD.n4818 0.0114843
R5266 DVDD.n4903 DVDD.n4902 0.0114843
R5267 DVDD.n4910 DVDD.n4909 0.0114843
R5268 DVDD.n4940 DVDD.n4939 0.0114843
R5269 DVDD.n4947 DVDD.n4946 0.0114843
R5270 DVDD.n4960 DVDD.n4959 0.0114843
R5271 DVDD.n4989 DVDD.n4988 0.0114843
R5272 DVDD.n4996 DVDD.n4995 0.0114843
R5273 DVDD.n5004 DVDD.n5003 0.0114843
R5274 DVDD.n5099 DVDD.n5098 0.0114843
R5275 DVDD.n5165 DVDD.n5164 0.0114843
R5276 DVDD.n5178 DVDD.n5177 0.0114843
R5277 DVDD.n5311 DVDD.n5310 0.0114843
R5278 DVDD.n5319 DVDD.n5318 0.0114843
R5279 DVDD.n5340 DVDD.n5339 0.0114843
R5280 DVDD.n5348 DVDD.n5347 0.0114843
R5281 DVDD.n5370 DVDD.n5369 0.0114843
R5282 DVDD.n5376 DVDD.n5375 0.0114843
R5283 DVDD.n5384 DVDD.n5383 0.0114843
R5284 DVDD.n5402 DVDD.n5401 0.0114843
R5285 DVDD.n5409 DVDD.n5408 0.0114843
R5286 DVDD.n5423 DVDD.n5422 0.0114843
R5287 DVDD.n5431 DVDD.n5430 0.0114843
R5288 DVDD.n6050 DVDD.n6049 0.0114843
R5289 DVDD.n1336 DVDD.n1335 0.0114843
R5290 DVDD.n1343 DVDD.n1342 0.0114843
R5291 DVDD.n1350 DVDD.n1349 0.0114843
R5292 DVDD.n1385 DVDD.n1384 0.0114843
R5293 DVDD.n1517 DVDD.n1516 0.0114843
R5294 DVDD.n1510 DVDD.n1509 0.0114843
R5295 DVDD.n1503 DVDD.n1502 0.0114843
R5296 DVDD.n1497 DVDD.n1496 0.0114843
R5297 DVDD.n1471 DVDD.n1470 0.0114843
R5298 DVDD.n1464 DVDD.n1463 0.0114843
R5299 DVDD.n1694 DVDD.n1693 0.0114843
R5300 DVDD.n1720 DVDD.n1719 0.0114843
R5301 DVDD.n1713 DVDD.n1712 0.0114843
R5302 DVDD.n290 DVDD.n289 0.0114843
R5303 DVDD.n285 DVDD.n284 0.0114843
R5304 DVDD.n278 DVDD.n277 0.0114843
R5305 DVDD.n271 DVDD.n270 0.0114843
R5306 DVDD.n19196 DVDD.n19195 0.0114843
R5307 DVDD.n19203 DVDD.n19202 0.0114843
R5308 DVDD.n19210 DVDD.n19209 0.0114843
R5309 DVDD.n19215 DVDD.n19214 0.0114843
R5310 DVDD.n19447 DVDD.n19446 0.0114843
R5311 DVDD.n19440 DVDD.n19439 0.0114843
R5312 DVDD.n19226 DVDD.n19225 0.0114843
R5313 DVDD.n11357 DVDD.n11356 0.0114843
R5314 DVDD.n11362 DVDD.n11361 0.0114843
R5315 DVDD.n11369 DVDD.n11368 0.0114843
R5316 DVDD.n11376 DVDD.n11375 0.0114843
R5317 DVDD.n11631 DVDD.n11630 0.0114843
R5318 DVDD.n11638 DVDD.n11637 0.0114843
R5319 DVDD.n11850 DVDD.n11849 0.0114843
R5320 DVDD.n11843 DVDD.n11842 0.0114843
R5321 DVDD.n11813 DVDD.n11812 0.0114843
R5322 DVDD.n11806 DVDD.n11805 0.0114843
R5323 DVDD.n11793 DVDD.n11792 0.0114843
R5324 DVDD.n11764 DVDD.n11763 0.0114843
R5325 DVDD.n11757 DVDD.n11756 0.0114843
R5326 DVDD.n12346 DVDD.n12345 0.0114843
R5327 DVDD.n13147 DVDD.n13146 0.0114843
R5328 DVDD.n13119 DVDD.n13118 0.0114843
R5329 DVDD.n13090 DVDD.n13089 0.0114843
R5330 DVDD.n13077 DVDD.n13076 0.0114843
R5331 DVDD.n13053 DVDD.n13052 0.0114843
R5332 DVDD.n13032 DVDD.n13031 0.0114843
R5333 DVDD.n12696 DVDD.n12695 0.0114843
R5334 DVDD.n1913 DVDD.n1912 0.0114843
R5335 DVDD.n1920 DVDD.n1919 0.0114843
R5336 DVDD.n1927 DVDD.n1926 0.0114843
R5337 DVDD.n1962 DVDD.n1961 0.0114843
R5338 DVDD.n2081 DVDD.n2080 0.0114843
R5339 DVDD.n2088 DVDD.n2087 0.0114843
R5340 DVDD.n2095 DVDD.n2094 0.0114843
R5341 DVDD.n2101 DVDD.n2100 0.0114843
R5342 DVDD.n2127 DVDD.n2126 0.0114843
R5343 DVDD.n2134 DVDD.n2133 0.0114843
R5344 DVDD.n2227 DVDD.n2226 0.0114843
R5345 DVDD.n2274 DVDD.n2273 0.0114843
R5346 DVDD.n2281 DVDD.n2280 0.0114843
R5347 DVDD.n19592 DVDD.n19591 0.0114843
R5348 DVDD.n19585 DVDD.n19584 0.0114843
R5349 DVDD.n19578 DVDD.n19577 0.0114843
R5350 DVDD.n19483 DVDD.n19482 0.0114843
R5351 DVDD.n19490 DVDD.n19489 0.0114843
R5352 DVDD.n19497 DVDD.n19496 0.0114843
R5353 DVDD.n18957 DVDD.n18956 0.0114843
R5354 DVDD.n18950 DVDD.n18949 0.0114843
R5355 DVDD.n18944 DVDD.n18943 0.0114843
R5356 DVDD.n7029 DVDD.n7028 0.0114843
R5357 DVDD.n7022 DVDD.n7021 0.0114843
R5358 DVDD.n7015 DVDD.n7014 0.0114843
R5359 DVDD.n6879 DVDD.n6878 0.0114843
R5360 DVDD.n6872 DVDD.n6871 0.0114843
R5361 DVDD.n6781 DVDD.n6780 0.0114843
R5362 DVDD.n6774 DVDD.n6773 0.0114843
R5363 DVDD.n6744 DVDD.n6743 0.0114843
R5364 DVDD.n6737 DVDD.n6736 0.0114843
R5365 DVDD.n6724 DVDD.n6723 0.0114843
R5366 DVDD.n6695 DVDD.n6694 0.0114843
R5367 DVDD.n6688 DVDD.n6687 0.0114843
R5368 DVDD.n6517 DVDD.n6516 0.0114843
R5369 DVDD.n6450 DVDD.n6449 0.0114843
R5370 DVDD.n6421 DVDD.n6420 0.0114843
R5371 DVDD.n6391 DVDD.n6390 0.0114843
R5372 DVDD.n6377 DVDD.n6376 0.0114843
R5373 DVDD.n6352 DVDD.n6351 0.0114843
R5374 DVDD.n6330 DVDD.n6329 0.0114843
R5375 DVDD.n4507 DVDD.n4506 0.0114843
R5376 DVDD.n3267 DVDD.n3266 0.0114843
R5377 DVDD.n3260 DVDD.n3259 0.0114843
R5378 DVDD.n3253 DVDD.n3252 0.0114843
R5379 DVDD.n3218 DVDD.n3217 0.0114843
R5380 DVDD.n3480 DVDD.n3479 0.0114843
R5381 DVDD.n3487 DVDD.n3486 0.0114843
R5382 DVDD.n3494 DVDD.n3493 0.0114843
R5383 DVDD.n3500 DVDD.n3499 0.0114843
R5384 DVDD.n3526 DVDD.n3525 0.0114843
R5385 DVDD.n3533 DVDD.n3532 0.0114843
R5386 DVDD.n3555 DVDD.n3554 0.0114843
R5387 DVDD.n3718 DVDD.n3717 0.0114843
R5388 DVDD.n3725 DVDD.n3724 0.0114843
R5389 DVDD.n3776 DVDD.n3775 0.0114843
R5390 DVDD.n3771 DVDD.n3770 0.0114843
R5391 DVDD.n3764 DVDD.n3763 0.0114843
R5392 DVDD.n3757 DVDD.n3756 0.0114843
R5393 DVDD.n18500 DVDD.n18499 0.0114843
R5394 DVDD.n18507 DVDD.n18506 0.0114843
R5395 DVDD.n18514 DVDD.n18513 0.0114843
R5396 DVDD.n18519 DVDD.n18518 0.0114843
R5397 DVDD.n18794 DVDD.n18793 0.0114843
R5398 DVDD.n18787 DVDD.n18786 0.0114843
R5399 DVDD.n18530 DVDD.n18529 0.0114843
R5400 DVDD.n10051 DVDD.n10050 0.0114843
R5401 DVDD.n10046 DVDD.n10045 0.0114843
R5402 DVDD.n10039 DVDD.n10038 0.0114843
R5403 DVDD.n10032 DVDD.n10031 0.0114843
R5404 DVDD.n7887 DVDD.n7886 0.0114843
R5405 DVDD.n7894 DVDD.n7893 0.0114843
R5406 DVDD.n9749 DVDD.n9748 0.0114843
R5407 DVDD.n9742 DVDD.n9741 0.0114843
R5408 DVDD.n9712 DVDD.n9711 0.0114843
R5409 DVDD.n9705 DVDD.n9704 0.0114843
R5410 DVDD.n9692 DVDD.n9691 0.0114843
R5411 DVDD.n9663 DVDD.n9662 0.0114843
R5412 DVDD.n9656 DVDD.n9655 0.0114843
R5413 DVDD.n8366 DVDD.n7903 0.0114843
R5414 DVDD.n9236 DVDD.n9235 0.0114843
R5415 DVDD.n9207 DVDD.n9206 0.0114843
R5416 DVDD.n9177 DVDD.n9176 0.0114843
R5417 DVDD.n9163 DVDD.n9162 0.0114843
R5418 DVDD.n9138 DVDD.n9137 0.0114843
R5419 DVDD.n9116 DVDD.n9115 0.0114843
R5420 DVDD.n8781 DVDD.n8780 0.0114843
R5421 DVDD.n2905 DVDD.n2904 0.01148
R5422 DVDD.n1023 DVDD.n1022 0.01148
R5423 DVDD.n14158 DVDD.n14157 0.011478
R5424 DVDD.n14163 DVDD.n14162 0.011478
R5425 DVDD.n8009 DVDD.n8008 0.0114205
R5426 DVDD.n9364 DVDD.n9363 0.01139
R5427 DVDD.n13275 DVDD.n13274 0.01139
R5428 DVDD.n19301 DVDD.n19300 0.0113071
R5429 DVDD.n12239 DVDD.n12238 0.0113071
R5430 DVDD.n13317 DVDD.n13316 0.0113071
R5431 DVDD.n19732 DVDD.n19731 0.0113071
R5432 DVDD.n5028 DVDD.n5027 0.0113071
R5433 DVDD.n5458 DVDD.n5457 0.0113071
R5434 DVDD.n5684 DVDD.n5683 0.0113071
R5435 DVDD.n1377 DVDD.n1376 0.0113071
R5436 DVDD.n11726 DVDD.n11725 0.0113071
R5437 DVDD.n13005 DVDD.n13004 0.0113071
R5438 DVDD.n12757 DVDD.n12756 0.0113071
R5439 DVDD.n1954 DVDD.n1953 0.0113071
R5440 DVDD.n6656 DVDD.n6655 0.0113071
R5441 DVDD.n6303 DVDD.n6302 0.0113071
R5442 DVDD.n6141 DVDD.n6140 0.0113071
R5443 DVDD.n3226 DVDD.n3225 0.0113071
R5444 DVDD.n9624 DVDD.n9623 0.0113071
R5445 DVDD.n9089 DVDD.n9088 0.0113071
R5446 DVDD.n8843 DVDD.n8842 0.0113071
R5447 DVDD.n3669 DVDD.n2865 0.0113
R5448 DVDD.n1738 DVDD.n1737 0.0113
R5449 DVDD.n3414 DVDD.n3413 0.0113
R5450 DVDD.n3394 DVDD.n3393 0.0113
R5451 DVDD.n3388 DVDD.n3387 0.0113
R5452 DVDD.n19722 DVDD.n19721 0.0112756
R5453 DVDD.n1367 DVDD.n1366 0.0112756
R5454 DVDD.n1944 DVDD.n1943 0.0112756
R5455 DVDD.n3236 DVDD.n3235 0.0112756
R5456 DVDD.n8280 DVDD.n8279 0.0112322
R5457 DVDD.n8109 DVDD.n8108 0.0112322
R5458 DVDD.n7945 DVDD.n7944 0.0112322
R5459 DVDD.n8032 DVDD.n8031 0.0112322
R5460 DVDD.n4923 DVDD.n4922 0.011187
R5461 DVDD.n11830 DVDD.n11829 0.011187
R5462 DVDD.n6761 DVDD.n6760 0.011187
R5463 DVDD.n9729 DVDD.n9728 0.011187
R5464 DVDD.n12958 DVDD.n12873 0.0111514
R5465 DVDD.n9039 DVDD.n8954 0.0111514
R5466 DVDD.n19331 DVDD.n19330 0.0111299
R5467 DVDD.n19713 DVDD.n19712 0.0111299
R5468 DVDD.n3875 DVDD.n3874 0.0111299
R5469 DVDD.n5439 DVDD.n5438 0.0111299
R5470 DVDD.n1358 DVDD.n1357 0.0111299
R5471 DVDD.n10122 DVDD.n10121 0.0111299
R5472 DVDD.n13100 DVDD.n13099 0.0111299
R5473 DVDD.n13024 DVDD.n13023 0.0111299
R5474 DVDD.n1935 DVDD.n1934 0.0111299
R5475 DVDD.n7096 DVDD.n7095 0.0111299
R5476 DVDD.n6401 DVDD.n6400 0.0111299
R5477 DVDD.n6322 DVDD.n6321 0.0111299
R5478 DVDD.n3245 DVDD.n3244 0.0111299
R5479 DVDD.n7154 DVDD.n7153 0.0111299
R5480 DVDD.n9187 DVDD.n9186 0.0111299
R5481 DVDD.n9108 DVDD.n9107 0.0111299
R5482 DVDD.n1273 DVDD.n1272 0.01112
R5483 DVDD.n3125 DVDD.n3124 0.01112
R5484 DVDD.n12737 DVDD.n12735 0.0110796
R5485 DVDD.n6106 DVDD.n6105 0.0110796
R5486 DVDD.n6119 DVDD.n6117 0.0110796
R5487 DVDD.n8821 DVDD.n8819 0.0110796
R5488 DVDD.n12450 DVDD.n12448 0.0110796
R5489 DVDD.n5668 DVDD.n5667 0.0110796
R5490 DVDD.n4557 DVDD.n4058 0.0110796
R5491 DVDD.n8474 DVDD.n8472 0.0110796
R5492 DVDD.n12437 DVDD.n12435 0.0110796
R5493 DVDD.n5622 DVDD.n5620 0.0110796
R5494 DVDD.n4572 DVDD.n4048 0.0110796
R5495 DVDD.n8456 DVDD.n8454 0.0110796
R5496 DVDD.n12417 DVDD.n12416 0.0110796
R5497 DVDD.n5575 DVDD.n5574 0.0110796
R5498 DVDD.n4587 DVDD.n4038 0.0110796
R5499 DVDD.n8437 DVDD.n8436 0.0110796
R5500 DVDD.n14060 DVDD.n14059 0.0110794
R5501 DVDD.n17340 DVDD.n17339 0.0110794
R5502 DVDD.n13963 DVDD.n13962 0.0110794
R5503 DVDD.n17499 DVDD.n17498 0.0110794
R5504 DVDD.n8217 DVDD.n8216 0.0110439
R5505 DVDD.n7968 DVDD.n7967 0.0110439
R5506 DVDD.n9823 DVDD.n9822 0.01103
R5507 DVDD.n11924 DVDD.n11923 0.01103
R5508 DVDD.n5494 DVDD.n5493 0.0109642
R5509 DVDD.n12969 DVDD.n12968 0.0109642
R5510 DVDD.n19270 DVDD.n19269 0.0109528
R5511 DVDD.n12130 DVDD.n12129 0.0109528
R5512 DVDD.n19898 DVDD.n19897 0.0109528
R5513 DVDD.n20075 DVDD.n20074 0.0109528
R5514 DVDD.n19080 DVDD.n19079 0.0109528
R5515 DVDD.n4953 DVDD.n4952 0.0109528
R5516 DVDD.n1479 DVDD.n1478 0.0109528
R5517 DVDD.n1698 DVDD.n1697 0.0109528
R5518 DVDD.n19462 DVDD.n19461 0.0109528
R5519 DVDD.n11800 DVDD.n11799 0.0109528
R5520 DVDD.n2119 DVDD.n2118 0.0109528
R5521 DVDD.n2296 DVDD.n2295 0.0109528
R5522 DVDD.n18972 DVDD.n18971 0.0109528
R5523 DVDD.n6731 DVDD.n6730 0.0109528
R5524 DVDD.n3518 DVDD.n3517 0.0109528
R5525 DVDD.n3740 DVDD.n3739 0.0109528
R5526 DVDD.n18809 DVDD.n18808 0.0109528
R5527 DVDD.n9699 DVDD.n9698 0.0109528
R5528 DVDD.n9492 DVDD.n9491 0.01094
R5529 DVDD.n12297 DVDD.n12296 0.01094
R5530 DVDD.n3417 DVDD.n3416 0.0109
R5531 DVDD.n12959 DVDD.n12958 0.0108992
R5532 DVDD.n9040 DVDD.n9039 0.0108992
R5533 DVDD.n16027 DVDD.n16026 0.0108633
R5534 DVDD.n16028 DVDD.n16027 0.0108633
R5535 DVDD.n15640 DVDD.n15639 0.0108633
R5536 DVDD.n15639 DVDD.n15638 0.0108633
R5537 DVDD.n8242 DVDD.n8241 0.0108556
R5538 DVDD.n9442 DVDD.n9441 0.0108556
R5539 DVDD.n9440 DVDD.n9439 0.0108556
R5540 DVDD.n7939 DVDD.n7938 0.0108556
R5541 DVDD.n3360 DVDD.n3359 0.01085
R5542 DVDD.n13583 DVDD.n13582 0.0107895
R5543 DVDD.n13664 DVDD.n13663 0.0107895
R5544 DVDD.n5644 DVDD.n5643 0.0107895
R5545 DVDD.n12793 DVDD.n12792 0.0107895
R5546 DVDD.n18172 DVDD.n18171 0.0107895
R5547 DVDD.n17898 DVDD.n17897 0.0107895
R5548 DVDD.n12064 DVDD.n12063 0.0107756
R5549 DVDD.n12159 DVDD.n12158 0.0107756
R5550 DVDD.n20067 DVDD.n20066 0.0107756
R5551 DVDD.n5092 DVDD.n5091 0.0107756
R5552 DVDD.n5186 DVDD.n5185 0.0107756
R5553 DVDD.n5332 DVDD.n5331 0.0107756
R5554 DVDD.n5355 DVDD.n5354 0.0107756
R5555 DVDD.n1706 DVDD.n1705 0.0107756
R5556 DVDD.n11662 DVDD.n11661 0.0107756
R5557 DVDD.n12366 DVDD.n12365 0.0107756
R5558 DVDD.n13127 DVDD.n13126 0.0107756
R5559 DVDD.n13105 DVDD.n13104 0.0107756
R5560 DVDD.n2288 DVDD.n2287 0.0107756
R5561 DVDD.n6590 DVDD.n6589 0.0107756
R5562 DVDD.n6496 DVDD.n6495 0.0107756
R5563 DVDD.n6429 DVDD.n6428 0.0107756
R5564 DVDD.n6406 DVDD.n6405 0.0107756
R5565 DVDD.n3732 DVDD.n3731 0.0107756
R5566 DVDD.n9558 DVDD.n9557 0.0107756
R5567 DVDD.n8387 DVDD.n8386 0.0107756
R5568 DVDD.n9215 DVDD.n9214 0.0107756
R5569 DVDD.n9192 DVDD.n9191 0.0107756
R5570 DVDD.n9397 DVDD.n9396 0.0107695
R5571 DVDD.n9396 DVDD.n9395 0.0107695
R5572 DVDD.n18742 DVDD.n18741 0.01076
R5573 DVDD.n1753 DVDD.n1752 0.01076
R5574 DVDD.n13556 DVDD.n13555 0.010701
R5575 DVDD.n13637 DVDD.n13636 0.010701
R5576 DVDD.n13608 DVDD.n13607 0.010701
R5577 DVDD.n13689 DVDD.n13688 0.010701
R5578 DVDD.n5470 DVDD.n5469 0.010701
R5579 DVDD.n5593 DVDD.n5592 0.010701
R5580 DVDD.n5962 DVDD.n5961 0.010701
R5581 DVDD.n5692 DVDD.n5691 0.010701
R5582 DVDD.n12993 DVDD.n12992 0.010701
R5583 DVDD.n12834 DVDD.n12833 0.010701
R5584 DVDD.n12625 DVDD.n12624 0.010701
R5585 DVDD.n12749 DVDD.n12748 0.010701
R5586 DVDD.n787 DVDD.n786 0.010701
R5587 DVDD.n824 DVDD.n823 0.010701
R5588 DVDD.n18199 DVDD.n18198 0.010701
R5589 DVDD.n18055 DVDD.n18054 0.010701
R5590 DVDD.n17977 DVDD.n17976 0.010701
R5591 DVDD.n17925 DVDD.n17924 0.010701
R5592 DVDD.n17844 DVDD.n17843 0.010701
R5593 DVDD.n18147 DVDD.n18146 0.010701
R5594 DVDD.n17873 DVDD.n17872 0.010701
R5595 DVDD.n17778 DVDD.n17777 0.010701
R5596 DVDD.n3385 DVDD.n3384 0.0106747
R5597 DVDD.n9448 DVDD.n9447 0.0106674
R5598 DVDD.n8319 DVDD.n8318 0.0106674
R5599 DVDD.n13696 DVDD.n13695 0.0106125
R5600 DVDD.n5955 DVDD.n5954 0.0106125
R5601 DVDD.n12618 DVDD.n12617 0.0106125
R5602 DVDD.n761 DVDD.n760 0.0106125
R5603 DVDD.n798 DVDD.n797 0.0106125
R5604 DVDD.n18081 DVDD.n18080 0.0106125
R5605 DVDD.n18003 DVDD.n18002 0.0106125
R5606 DVDD.n17771 DVDD.n17770 0.0106125
R5607 DVDD.n18140 DVDD.n18139 0.0106125
R5608 DVDD.n11998 DVDD.n11997 0.0105984
R5609 DVDD.n12089 DVDD.n12088 0.0105984
R5610 DVDD.n12168 DVDD.n12167 0.0105984
R5611 DVDD.n13390 DVDD.n13389 0.0105984
R5612 DVDD.n19920 DVDD.n19919 0.0105984
R5613 DVDD.n19072 DVDD.n19071 0.0105984
R5614 DVDD.n4683 DVDD.n4682 0.0105984
R5615 DVDD.n4932 DVDD.n4931 0.0105984
R5616 DVDD.n5201 DVDD.n5200 0.0105984
R5617 DVDD.n6072 DVDD.n6071 0.0105984
R5618 DVDD.n1457 DVDD.n1456 0.0105984
R5619 DVDD.n19454 DVDD.n19453 0.0105984
R5620 DVDD.n11390 DVDD.n11389 0.0105984
R5621 DVDD.n11821 DVDD.n11820 0.0105984
R5622 DVDD.n12381 DVDD.n12380 0.0105984
R5623 DVDD.n12704 DVDD.n12703 0.0105984
R5624 DVDD.n2141 DVDD.n2140 0.0105984
R5625 DVDD.n18964 DVDD.n18963 0.0105984
R5626 DVDD.n7001 DVDD.n7000 0.0105984
R5627 DVDD.n6752 DVDD.n6751 0.0105984
R5628 DVDD.n6481 DVDD.n6480 0.0105984
R5629 DVDD.n4522 DVDD.n4521 0.0105984
R5630 DVDD.n3540 DVDD.n3539 0.0105984
R5631 DVDD.n18801 DVDD.n18800 0.0105984
R5632 DVDD.n10018 DVDD.n10017 0.0105984
R5633 DVDD.n9720 DVDD.n9719 0.0105984
R5634 DVDD.n8402 DVDD.n8401 0.0105984
R5635 DVDD.n8789 DVDD.n8788 0.0105984
R5636 DVDD.n15124 DVDD.n15123 0.0105854
R5637 DVDD.n15127 DVDD.n15126 0.0105854
R5638 DVDD.n14162 DVDD.n14161 0.0105814
R5639 DVDD.n14159 DVDD.n14158 0.0105814
R5640 DVDD.n17502 DVDD.n17501 0.0105762
R5641 DVDD.n14063 DVDD.n14062 0.0105762
R5642 DVDD.n17459 DVDD.n17458 0.0105762
R5643 DVDD.n13966 DVDD.n13965 0.0105762
R5644 DVDD.n17343 DVDD.n17342 0.0105762
R5645 DVDD.n14160 DVDD.n14159 0.0105466
R5646 DVDD.n14061 DVDD.n14060 0.0105466
R5647 DVDD.n13964 DVDD.n13963 0.0105466
R5648 DVDD.n17500 DVDD.n17499 0.0105466
R5649 DVDD.n17457 DVDD.n17456 0.0105466
R5650 DVDD.n17342 DVDD.n17341 0.0105466
R5651 DVDD.n17341 DVDD.n17340 0.0105466
R5652 DVDD.n13965 DVDD.n13964 0.0105466
R5653 DVDD.n14062 DVDD.n14061 0.0105466
R5654 DVDD.n17458 DVDD.n17457 0.0105466
R5655 DVDD.n14161 DVDD.n14160 0.0105466
R5656 DVDD.n17501 DVDD.n17500 0.0105466
R5657 DVDD.n13504 DVDD.n13503 0.010524
R5658 DVDD.n5055 DVDD.n5054 0.010524
R5659 DVDD.n11699 DVDD.n11698 0.010524
R5660 DVDD.n18114 DVDD.n18113 0.010524
R5661 DVDD.n17745 DVDD.n17744 0.010524
R5662 DVDD.n5929 DVDD.n5928 0.010524
R5663 DVDD.n12592 DVDD.n12591 0.010524
R5664 DVDD.n13715 DVDD.n13714 0.010524
R5665 DVDD.n3411 DVDD.n3410 0.0104984
R5666 DVDD.n9428 DVDD.n9427 0.0104791
R5667 DVDD.n12023 DVDD.n12022 0.0104213
R5668 DVDD.n13456 DVDD.n13455 0.0104213
R5669 DVDD.n4790 DVDD.n4789 0.0104213
R5670 DVDD.n5416 DVDD.n5415 0.0104213
R5671 DVDD.n6040 DVDD.n6034 0.0104213
R5672 DVDD.n11616 DVDD.n11615 0.0104213
R5673 DVDD.n13046 DVDD.n13045 0.0104213
R5674 DVDD.n12686 DVDD.n12685 0.0104213
R5675 DVDD.n6894 DVDD.n6893 0.0104213
R5676 DVDD.n6345 DVDD.n6344 0.0104213
R5677 DVDD.n4491 DVDD.n4485 0.0104213
R5678 DVDD.n7872 DVDD.n7871 0.0104213
R5679 DVDD.n9131 DVDD.n9130 0.0104213
R5680 DVDD.n8772 DVDD.n8771 0.0104213
R5681 DVDD.n12465 DVDD.n12464 0.0104
R5682 DVDD.n12472 DVDD.n12466 0.0104
R5683 DVDD.n5707 DVDD.n5706 0.0104
R5684 DVDD.n4068 DVDD.n4067 0.0104
R5685 DVDD.n4075 DVDD.n4069 0.0104
R5686 DVDD.n8490 DVDD.n8489 0.0104
R5687 DVDD.n8497 DVDD.n8491 0.0104
R5688 DVDD.n12447 DVDD.n12446 0.0104
R5689 DVDD.n12458 DVDD.n12451 0.0104
R5690 DVDD.n5665 DVDD.n5664 0.0104
R5691 DVDD.n4570 DVDD.n4556 0.0104
R5692 DVDD.n4559 DVDD.n4558 0.0104
R5693 DVDD.n4066 DVDD.n4059 0.0104
R5694 DVDD.n8471 DVDD.n8470 0.0104
R5695 DVDD.n8482 DVDD.n8475 0.0104
R5696 DVDD.n12434 DVDD.n12433 0.0104
R5697 DVDD.n12445 DVDD.n12438 0.0104
R5698 DVDD.n5619 DVDD.n5618 0.0104
R5699 DVDD.n4585 DVDD.n4571 0.0104
R5700 DVDD.n4574 DVDD.n4573 0.0104
R5701 DVDD.n4056 DVDD.n4049 0.0104
R5702 DVDD.n8453 DVDD.n8452 0.0104
R5703 DVDD.n8464 DVDD.n8457 0.0104
R5704 DVDD.n12415 DVDD.n12414 0.0104
R5705 DVDD.n12426 DVDD.n12419 0.0104
R5706 DVDD.n5572 DVDD.n5571 0.0104
R5707 DVDD.n4600 DVDD.n4586 0.0104
R5708 DVDD.n4589 DVDD.n4588 0.0104
R5709 DVDD.n4046 DVDD.n4039 0.0104
R5710 DVDD.n8435 DVDD.n8434 0.0104
R5711 DVDD.n8446 DVDD.n8439 0.0104
R5712 DVDD.n3331 DVDD.n3330 0.0104
R5713 DVDD.n3441 DVDD.n3440 0.0104
R5714 DVDD.n3381 DVDD.n3380 0.0104
R5715 DVDD.n3372 DVDD.n3371 0.0104
R5716 DVDD.n3586 DVDD.n3585 0.0104
R5717 DVDD.n3607 DVDD.n3606 0.0104
R5718 DVDD.n3588 DVDD.n3587 0.0104
R5719 DVDD.n18584 DVDD.n18583 0.0104
R5720 DVDD.n18598 DVDD.n18597 0.0104
R5721 DVDD.n18646 DVDD.n18645 0.0104
R5722 DVDD.n9429 DVDD.n9428 0.0102908
R5723 DVDD.n8117 DVDD.n8116 0.0102908
R5724 DVDD.n12927 DVDD.n12924 0.0102826
R5725 DVDD.n12946 DVDD.n12943 0.0102826
R5726 DVDD.n5511 DVDD.n5508 0.0102826
R5727 DVDD.n5537 DVDD.n5534 0.0102826
R5728 DVDD.n4009 DVDD.n4006 0.0102826
R5729 DVDD.n4032 DVDD.n4029 0.0102826
R5730 DVDD.n8965 DVDD.n8962 0.0102826
R5731 DVDD.n9034 DVDD.n9031 0.0102826
R5732 DVDD.n12908 DVDD.n12907 0.0102826
R5733 DVDD.n12887 DVDD.n12884 0.0102826
R5734 DVDD.n5715 DVDD.n5712 0.0102826
R5735 DVDD.n4086 DVDD.n4083 0.0102826
R5736 DVDD.n8992 DVDD.n8989 0.0102826
R5737 DVDD.n9015 DVDD.n9014 0.0102826
R5738 DVDD.n13529 DVDD.n13528 0.010282
R5739 DVDD.n13581 DVDD.n13580 0.010282
R5740 DVDD.n13662 DVDD.n13661 0.010282
R5741 DVDD.n15429 DVDD.n15428 0.010282
R5742 DVDD.n14674 DVDD.n14673 0.010282
R5743 DVDD.n14538 DVDD.n14537 0.010282
R5744 DVDD.n14537 DVDD.n14536 0.010282
R5745 DVDD.n14675 DVDD.n14674 0.010282
R5746 DVDD.n15428 DVDD.n15427 0.010282
R5747 DVDD.n5642 DVDD.n5641 0.010282
R5748 DVDD.n12795 DVDD.n12794 0.010282
R5749 DVDD.n18030 DVDD.n18029 0.010282
R5750 DVDD.n18174 DVDD.n18173 0.010282
R5751 DVDD.n17900 DVDD.n17899 0.010282
R5752 DVDD.n6175 DVDD.n6174 0.010282
R5753 DVDD.n6174 DVDD.n6173 0.010282
R5754 DVDD.n8877 DVDD.n8876 0.010282
R5755 DVDD.n8876 DVDD.n8875 0.010282
R5756 DVDD.n12194 DVDD.n12193 0.0102585
R5757 DVDD.n13716 DVDD.n13715 0.0102585
R5758 DVDD.n5054 DVDD.n5053 0.0102585
R5759 DVDD.n5930 DVDD.n5929 0.0102585
R5760 DVDD.n11700 DVDD.n11699 0.0102585
R5761 DVDD.n12593 DVDD.n12592 0.0102585
R5762 DVDD.n18115 DVDD.n18114 0.0102585
R5763 DVDD.n17746 DVDD.n17745 0.0102585
R5764 DVDD.n11992 DVDD.n11991 0.0102441
R5765 DVDD.n12247 DVDD.n12246 0.0102441
R5766 DVDD.n12245 DVDD.n12244 0.0102441
R5767 DVDD.n13429 DVDD.n13428 0.0102441
R5768 DVDD.n19753 DVDD.n19752 0.0102441
R5769 DVDD.n19889 DVDD.n19888 0.0102441
R5770 DVDD.n1398 DVDD.n1397 0.0102441
R5771 DVDD.n1488 DVDD.n1487 0.0102441
R5772 DVDD.n1975 DVDD.n1974 0.0102441
R5773 DVDD.n2110 DVDD.n2109 0.0102441
R5774 DVDD.n3205 DVDD.n3204 0.0102441
R5775 DVDD.n3509 DVDD.n3508 0.0102441
R5776 DVDD.n7713 DVDD.n7712 0.01022
R5777 DVDD.n7714 DVDD.n7713 0.01022
R5778 DVDD.n7715 DVDD.n7714 0.01022
R5779 DVDD.n7716 DVDD.n7715 0.01022
R5780 DVDD.n7717 DVDD.n7716 0.01022
R5781 DVDD.n7718 DVDD.n7717 0.01022
R5782 DVDD.n7719 DVDD.n7718 0.01022
R5783 DVDD.n7720 DVDD.n7719 0.01022
R5784 DVDD.n7721 DVDD.n7720 0.01022
R5785 DVDD.n7722 DVDD.n7721 0.01022
R5786 DVDD.n7723 DVDD.n7722 0.01022
R5787 DVDD.n7724 DVDD.n7723 0.01022
R5788 DVDD.n7725 DVDD.n7724 0.01022
R5789 DVDD.n7726 DVDD.n7725 0.01022
R5790 DVDD.n7727 DVDD.n7726 0.01022
R5791 DVDD.n7728 DVDD.n7727 0.01022
R5792 DVDD.n7729 DVDD.n7728 0.01022
R5793 DVDD.n7730 DVDD.n7729 0.01022
R5794 DVDD.n7731 DVDD.n7730 0.01022
R5795 DVDD.n7732 DVDD.n7731 0.01022
R5796 DVDD.n3685 DVDD.n3684 0.01022
R5797 DVDD.n3684 DVDD.n3683 0.01022
R5798 DVDD.n2995 DVDD.n2994 0.01022
R5799 DVDD.n2994 DVDD.n2993 0.01022
R5800 DVDD.n2993 DVDD.n2992 0.01022
R5801 DVDD.n2992 DVDD.n2991 0.01022
R5802 DVDD.n2991 DVDD.n2990 0.01022
R5803 DVDD.n2990 DVDD.n2989 0.01022
R5804 DVDD.n2989 DVDD.n2988 0.01022
R5805 DVDD.n2988 DVDD.n2987 0.01022
R5806 DVDD.n2987 DVDD.n2986 0.01022
R5807 DVDD.n2986 DVDD.n2985 0.01022
R5808 DVDD.n2985 DVDD.n2984 0.01022
R5809 DVDD.n2984 DVDD.n2983 0.01022
R5810 DVDD.n2983 DVDD.n2982 0.01022
R5811 DVDD.n2982 DVDD.n2981 0.01022
R5812 DVDD.n2981 DVDD.n2980 0.01022
R5813 DVDD.n2980 DVDD.n2979 0.01022
R5814 DVDD.n2979 DVDD.n2978 0.01022
R5815 DVDD.n2978 DVDD.n2977 0.01022
R5816 DVDD.n2977 DVDD.n2976 0.01022
R5817 DVDD.n2976 DVDD.n2975 0.01022
R5818 DVDD.n2975 DVDD.n2974 0.01022
R5819 DVDD.n2974 DVDD.n2973 0.01022
R5820 DVDD.n2973 DVDD.n2972 0.01022
R5821 DVDD.n2972 DVDD.n2971 0.01022
R5822 DVDD.n2971 DVDD.n2970 0.01022
R5823 DVDD.n3457 DVDD.n2970 0.01022
R5824 DVDD.n2922 DVDD.n2921 0.01022
R5825 DVDD.n2923 DVDD.n2922 0.01022
R5826 DVDD.n2924 DVDD.n2923 0.01022
R5827 DVDD.n2925 DVDD.n2924 0.01022
R5828 DVDD.n2926 DVDD.n2925 0.01022
R5829 DVDD.n2927 DVDD.n2926 0.01022
R5830 DVDD.n2928 DVDD.n2927 0.01022
R5831 DVDD.n2964 DVDD.n2963 0.01022
R5832 DVDD.n2965 DVDD.n2964 0.01022
R5833 DVDD.n2966 DVDD.n2965 0.01022
R5834 DVDD.n2967 DVDD.n2966 0.01022
R5835 DVDD.n2968 DVDD.n2967 0.01022
R5836 DVDD.n3569 DVDD.n2968 0.01022
R5837 DVDD.n9989 DVDD.n9988 0.01022
R5838 DVDD.n9988 DVDD.n9987 0.01022
R5839 DVDD.n9987 DVDD.n9986 0.01022
R5840 DVDD.n9986 DVDD.n9985 0.01022
R5841 DVDD.n9985 DVDD.n9984 0.01022
R5842 DVDD.n9984 DVDD.n9983 0.01022
R5843 DVDD.n9983 DVDD.n9982 0.01022
R5844 DVDD.n9982 DVDD.n9981 0.01022
R5845 DVDD.n9981 DVDD.n9980 0.01022
R5846 DVDD.n9980 DVDD.n9979 0.01022
R5847 DVDD.n9979 DVDD.n9978 0.01022
R5848 DVDD.n9978 DVDD.n9977 0.01022
R5849 DVDD.n9977 DVDD.n9976 0.01022
R5850 DVDD.n9976 DVDD.n9975 0.01022
R5851 DVDD.n9975 DVDD.n9974 0.01022
R5852 DVDD.n9974 DVDD.n9973 0.01022
R5853 DVDD.n9973 DVDD.n9972 0.01022
R5854 DVDD.n9972 DVDD.n9971 0.01022
R5855 DVDD.n9971 DVDD.n9970 0.01022
R5856 DVDD.n9970 DVDD.n9969 0.01022
R5857 DVDD.n9969 DVDD.n9968 0.01022
R5858 DVDD.n9968 DVDD.n9967 0.01022
R5859 DVDD.n9967 DVDD.n9966 0.01022
R5860 DVDD.n9966 DVDD.n9965 0.01022
R5861 DVDD.n9965 DVDD.n9964 0.01022
R5862 DVDD.n9964 DVDD.n9963 0.01022
R5863 DVDD.n9801 DVDD.n9800 0.01022
R5864 DVDD.n9802 DVDD.n9801 0.01022
R5865 DVDD.n7930 DVDD.n7929 0.01022
R5866 DVDD.n7929 DVDD.n7928 0.01022
R5867 DVDD.n7928 DVDD.n7927 0.01022
R5868 DVDD.n7927 DVDD.n7926 0.01022
R5869 DVDD.n7926 DVDD.n7925 0.01022
R5870 DVDD.n7925 DVDD.n7924 0.01022
R5871 DVDD.n7924 DVDD.n7923 0.01022
R5872 DVDD.n7923 DVDD.n7922 0.01022
R5873 DVDD.n7922 DVDD.n7921 0.01022
R5874 DVDD.n7921 DVDD.n7920 0.01022
R5875 DVDD.n7920 DVDD.n7919 0.01022
R5876 DVDD.n7919 DVDD.n7918 0.01022
R5877 DVDD.n7918 DVDD.n7917 0.01022
R5878 DVDD.n7917 DVDD.n7916 0.01022
R5879 DVDD.n7916 DVDD.n7915 0.01022
R5880 DVDD.n7915 DVDD.n7914 0.01022
R5881 DVDD.n7914 DVDD.n7913 0.01022
R5882 DVDD.n9263 DVDD.n9262 0.01022
R5883 DVDD.n9264 DVDD.n9263 0.01022
R5884 DVDD.n2028 DVDD.n2027 0.01022
R5885 DVDD.n2029 DVDD.n2028 0.01022
R5886 DVDD.n2030 DVDD.n2029 0.01022
R5887 DVDD.n2031 DVDD.n2030 0.01022
R5888 DVDD.n2032 DVDD.n2031 0.01022
R5889 DVDD.n2033 DVDD.n2032 0.01022
R5890 DVDD.n2034 DVDD.n2033 0.01022
R5891 DVDD.n2035 DVDD.n2034 0.01022
R5892 DVDD.n2036 DVDD.n2035 0.01022
R5893 DVDD.n2037 DVDD.n2036 0.01022
R5894 DVDD.n2038 DVDD.n2037 0.01022
R5895 DVDD.n2039 DVDD.n2038 0.01022
R5896 DVDD.n2040 DVDD.n2039 0.01022
R5897 DVDD.n2041 DVDD.n2040 0.01022
R5898 DVDD.n2042 DVDD.n2041 0.01022
R5899 DVDD.n2043 DVDD.n2042 0.01022
R5900 DVDD.n2044 DVDD.n2043 0.01022
R5901 DVDD.n2045 DVDD.n2044 0.01022
R5902 DVDD.n2046 DVDD.n2045 0.01022
R5903 DVDD.n2047 DVDD.n2046 0.01022
R5904 DVDD.n2048 DVDD.n2047 0.01022
R5905 DVDD.n2049 DVDD.n2048 0.01022
R5906 DVDD.n2050 DVDD.n2049 0.01022
R5907 DVDD.n2051 DVDD.n2050 0.01022
R5908 DVDD.n2052 DVDD.n2051 0.01022
R5909 DVDD.n2058 DVDD.n2052 0.01022
R5910 DVDD.n2160 DVDD.n2159 0.01022
R5911 DVDD.n2161 DVDD.n2160 0.01022
R5912 DVDD.n2162 DVDD.n2161 0.01022
R5913 DVDD.n2163 DVDD.n2162 0.01022
R5914 DVDD.n2164 DVDD.n2163 0.01022
R5915 DVDD.n2165 DVDD.n2164 0.01022
R5916 DVDD.n2166 DVDD.n2165 0.01022
R5917 DVDD.n2202 DVDD.n2201 0.01022
R5918 DVDD.n2203 DVDD.n2202 0.01022
R5919 DVDD.n2204 DVDD.n2203 0.01022
R5920 DVDD.n2205 DVDD.n2204 0.01022
R5921 DVDD.n2206 DVDD.n2205 0.01022
R5922 DVDD.n2212 DVDD.n2206 0.01022
R5923 DVDD.n2241 DVDD.n2240 0.01022
R5924 DVDD.n2240 DVDD.n2239 0.01022
R5925 DVDD.n7056 DVDD.n7055 0.01022
R5926 DVDD.n7055 DVDD.n7054 0.01022
R5927 DVDD.n7054 DVDD.n7053 0.01022
R5928 DVDD.n7053 DVDD.n7052 0.01022
R5929 DVDD.n7052 DVDD.n7051 0.01022
R5930 DVDD.n7051 DVDD.n7050 0.01022
R5931 DVDD.n7050 DVDD.n7049 0.01022
R5932 DVDD.n7049 DVDD.n7048 0.01022
R5933 DVDD.n7048 DVDD.n7047 0.01022
R5934 DVDD.n7047 DVDD.n7046 0.01022
R5935 DVDD.n7046 DVDD.n7045 0.01022
R5936 DVDD.n7045 DVDD.n7044 0.01022
R5937 DVDD.n7044 DVDD.n7043 0.01022
R5938 DVDD.n7043 DVDD.n7042 0.01022
R5939 DVDD.n7042 DVDD.n7041 0.01022
R5940 DVDD.n7041 DVDD.n7040 0.01022
R5941 DVDD.n7040 DVDD.n7039 0.01022
R5942 DVDD.n7039 DVDD.n7038 0.01022
R5943 DVDD.n7038 DVDD.n7037 0.01022
R5944 DVDD.n7037 DVDD.n7036 0.01022
R5945 DVDD.n6972 DVDD.n6971 0.01022
R5946 DVDD.n6971 DVDD.n6970 0.01022
R5947 DVDD.n6970 DVDD.n6969 0.01022
R5948 DVDD.n6969 DVDD.n6968 0.01022
R5949 DVDD.n6968 DVDD.n6967 0.01022
R5950 DVDD.n6967 DVDD.n6966 0.01022
R5951 DVDD.n6966 DVDD.n6965 0.01022
R5952 DVDD.n6965 DVDD.n6964 0.01022
R5953 DVDD.n6964 DVDD.n6963 0.01022
R5954 DVDD.n6963 DVDD.n6962 0.01022
R5955 DVDD.n6962 DVDD.n6961 0.01022
R5956 DVDD.n6961 DVDD.n6960 0.01022
R5957 DVDD.n6960 DVDD.n6959 0.01022
R5958 DVDD.n6959 DVDD.n6958 0.01022
R5959 DVDD.n6958 DVDD.n6957 0.01022
R5960 DVDD.n6957 DVDD.n6956 0.01022
R5961 DVDD.n6956 DVDD.n6955 0.01022
R5962 DVDD.n6955 DVDD.n6954 0.01022
R5963 DVDD.n6954 DVDD.n6953 0.01022
R5964 DVDD.n6953 DVDD.n6952 0.01022
R5965 DVDD.n6952 DVDD.n6951 0.01022
R5966 DVDD.n6951 DVDD.n6950 0.01022
R5967 DVDD.n6950 DVDD.n6949 0.01022
R5968 DVDD.n6949 DVDD.n6948 0.01022
R5969 DVDD.n6948 DVDD.n6947 0.01022
R5970 DVDD.n6947 DVDD.n6946 0.01022
R5971 DVDD.n6814 DVDD.n6813 0.01022
R5972 DVDD.n6813 DVDD.n6812 0.01022
R5973 DVDD.n6525 DVDD.n6524 0.01022
R5974 DVDD.n6526 DVDD.n6525 0.01022
R5975 DVDD.n6527 DVDD.n6526 0.01022
R5976 DVDD.n6528 DVDD.n6527 0.01022
R5977 DVDD.n6529 DVDD.n6528 0.01022
R5978 DVDD.n6530 DVDD.n6529 0.01022
R5979 DVDD.n6531 DVDD.n6530 0.01022
R5980 DVDD.n6532 DVDD.n6531 0.01022
R5981 DVDD.n6533 DVDD.n6532 0.01022
R5982 DVDD.n6534 DVDD.n6533 0.01022
R5983 DVDD.n6535 DVDD.n6534 0.01022
R5984 DVDD.n6536 DVDD.n6535 0.01022
R5985 DVDD.n6537 DVDD.n6536 0.01022
R5986 DVDD.n6538 DVDD.n6537 0.01022
R5987 DVDD.n6539 DVDD.n6538 0.01022
R5988 DVDD.n6540 DVDD.n6539 0.01022
R5989 DVDD.n6541 DVDD.n6540 0.01022
R5990 DVDD.n1872 DVDD.n1871 0.01022
R5991 DVDD.n1871 DVDD.n1870 0.01022
R5992 DVDD.n1870 DVDD.n1869 0.01022
R5993 DVDD.n1869 DVDD.n1868 0.01022
R5994 DVDD.n1868 DVDD.n1867 0.01022
R5995 DVDD.n1867 DVDD.n1866 0.01022
R5996 DVDD.n1866 DVDD.n1865 0.01022
R5997 DVDD.n3979 DVDD.n3978 0.01022
R5998 DVDD.n3978 DVDD.n3977 0.01022
R5999 DVDD.n19806 DVDD.n19805 0.01022
R6000 DVDD.n19807 DVDD.n19806 0.01022
R6001 DVDD.n19808 DVDD.n19807 0.01022
R6002 DVDD.n19809 DVDD.n19808 0.01022
R6003 DVDD.n19810 DVDD.n19809 0.01022
R6004 DVDD.n19811 DVDD.n19810 0.01022
R6005 DVDD.n19812 DVDD.n19811 0.01022
R6006 DVDD.n19813 DVDD.n19812 0.01022
R6007 DVDD.n19814 DVDD.n19813 0.01022
R6008 DVDD.n19815 DVDD.n19814 0.01022
R6009 DVDD.n19816 DVDD.n19815 0.01022
R6010 DVDD.n19817 DVDD.n19816 0.01022
R6011 DVDD.n19818 DVDD.n19817 0.01022
R6012 DVDD.n19819 DVDD.n19818 0.01022
R6013 DVDD.n19820 DVDD.n19819 0.01022
R6014 DVDD.n19821 DVDD.n19820 0.01022
R6015 DVDD.n19822 DVDD.n19821 0.01022
R6016 DVDD.n19823 DVDD.n19822 0.01022
R6017 DVDD.n19824 DVDD.n19823 0.01022
R6018 DVDD.n19825 DVDD.n19824 0.01022
R6019 DVDD.n19826 DVDD.n19825 0.01022
R6020 DVDD.n19827 DVDD.n19826 0.01022
R6021 DVDD.n19828 DVDD.n19827 0.01022
R6022 DVDD.n19829 DVDD.n19828 0.01022
R6023 DVDD.n19830 DVDD.n19829 0.01022
R6024 DVDD.n19836 DVDD.n19830 0.01022
R6025 DVDD.n19939 DVDD.n19938 0.01022
R6026 DVDD.n19940 DVDD.n19939 0.01022
R6027 DVDD.n19941 DVDD.n19940 0.01022
R6028 DVDD.n19942 DVDD.n19941 0.01022
R6029 DVDD.n19943 DVDD.n19942 0.01022
R6030 DVDD.n19944 DVDD.n19943 0.01022
R6031 DVDD.n19945 DVDD.n19944 0.01022
R6032 DVDD.n19981 DVDD.n19980 0.01022
R6033 DVDD.n19982 DVDD.n19981 0.01022
R6034 DVDD.n19983 DVDD.n19982 0.01022
R6035 DVDD.n19984 DVDD.n19983 0.01022
R6036 DVDD.n19985 DVDD.n19984 0.01022
R6037 DVDD.n19991 DVDD.n19985 0.01022
R6038 DVDD.n20020 DVDD.n20019 0.01022
R6039 DVDD.n20019 DVDD.n20018 0.01022
R6040 DVDD.n4636 DVDD.n4635 0.01022
R6041 DVDD.n4635 DVDD.n4634 0.01022
R6042 DVDD.n4634 DVDD.n4633 0.01022
R6043 DVDD.n4633 DVDD.n4632 0.01022
R6044 DVDD.n4632 DVDD.n4631 0.01022
R6045 DVDD.n4631 DVDD.n4630 0.01022
R6046 DVDD.n4630 DVDD.n4629 0.01022
R6047 DVDD.n4629 DVDD.n4628 0.01022
R6048 DVDD.n4628 DVDD.n4627 0.01022
R6049 DVDD.n4627 DVDD.n4626 0.01022
R6050 DVDD.n4626 DVDD.n4625 0.01022
R6051 DVDD.n4625 DVDD.n4624 0.01022
R6052 DVDD.n4624 DVDD.n4623 0.01022
R6053 DVDD.n4623 DVDD.n4622 0.01022
R6054 DVDD.n4622 DVDD.n4621 0.01022
R6055 DVDD.n4621 DVDD.n4620 0.01022
R6056 DVDD.n4620 DVDD.n4619 0.01022
R6057 DVDD.n4619 DVDD.n4618 0.01022
R6058 DVDD.n4618 DVDD.n4617 0.01022
R6059 DVDD.n4617 DVDD.n4616 0.01022
R6060 DVDD.n4746 DVDD.n4745 0.01022
R6061 DVDD.n4745 DVDD.n4744 0.01022
R6062 DVDD.n4744 DVDD.n4743 0.01022
R6063 DVDD.n4743 DVDD.n4742 0.01022
R6064 DVDD.n4742 DVDD.n4741 0.01022
R6065 DVDD.n4741 DVDD.n4740 0.01022
R6066 DVDD.n4740 DVDD.n4739 0.01022
R6067 DVDD.n4739 DVDD.n4738 0.01022
R6068 DVDD.n4738 DVDD.n4737 0.01022
R6069 DVDD.n4737 DVDD.n4736 0.01022
R6070 DVDD.n4736 DVDD.n4735 0.01022
R6071 DVDD.n4735 DVDD.n4734 0.01022
R6072 DVDD.n4734 DVDD.n4733 0.01022
R6073 DVDD.n4733 DVDD.n4732 0.01022
R6074 DVDD.n4732 DVDD.n4731 0.01022
R6075 DVDD.n4731 DVDD.n4730 0.01022
R6076 DVDD.n4730 DVDD.n4729 0.01022
R6077 DVDD.n4729 DVDD.n4728 0.01022
R6078 DVDD.n4728 DVDD.n4727 0.01022
R6079 DVDD.n4727 DVDD.n4726 0.01022
R6080 DVDD.n4726 DVDD.n4725 0.01022
R6081 DVDD.n4725 DVDD.n4724 0.01022
R6082 DVDD.n4724 DVDD.n4723 0.01022
R6083 DVDD.n4723 DVDD.n4722 0.01022
R6084 DVDD.n4722 DVDD.n4721 0.01022
R6085 DVDD.n4721 DVDD.n4720 0.01022
R6086 DVDD.n4851 DVDD.n4850 0.01022
R6087 DVDD.n4850 DVDD.n4849 0.01022
R6088 DVDD.n5116 DVDD.n5115 0.01022
R6089 DVDD.n5117 DVDD.n5116 0.01022
R6090 DVDD.n5118 DVDD.n5117 0.01022
R6091 DVDD.n5119 DVDD.n5118 0.01022
R6092 DVDD.n5120 DVDD.n5119 0.01022
R6093 DVDD.n5121 DVDD.n5120 0.01022
R6094 DVDD.n5122 DVDD.n5121 0.01022
R6095 DVDD.n5123 DVDD.n5122 0.01022
R6096 DVDD.n5124 DVDD.n5123 0.01022
R6097 DVDD.n5125 DVDD.n5124 0.01022
R6098 DVDD.n5126 DVDD.n5125 0.01022
R6099 DVDD.n5127 DVDD.n5126 0.01022
R6100 DVDD.n5128 DVDD.n5127 0.01022
R6101 DVDD.n5129 DVDD.n5128 0.01022
R6102 DVDD.n5130 DVDD.n5129 0.01022
R6103 DVDD.n5131 DVDD.n5130 0.01022
R6104 DVDD.n5132 DVDD.n5131 0.01022
R6105 DVDD.n19650 DVDD.n19649 0.01022
R6106 DVDD.n19649 DVDD.n19648 0.01022
R6107 DVDD.n19648 DVDD.n19647 0.01022
R6108 DVDD.n19647 DVDD.n19646 0.01022
R6109 DVDD.n19646 DVDD.n19645 0.01022
R6110 DVDD.n19645 DVDD.n19644 0.01022
R6111 DVDD.n19644 DVDD.n19643 0.01022
R6112 DVDD.n5284 DVDD.n5283 0.01022
R6113 DVDD.n5283 DVDD.n5282 0.01022
R6114 DVDD.n1095 DVDD.n1094 0.01022
R6115 DVDD.n1096 DVDD.n1095 0.01022
R6116 DVDD.n1097 DVDD.n1096 0.01022
R6117 DVDD.n1098 DVDD.n1097 0.01022
R6118 DVDD.n1099 DVDD.n1098 0.01022
R6119 DVDD.n1100 DVDD.n1099 0.01022
R6120 DVDD.n1101 DVDD.n1100 0.01022
R6121 DVDD.n1102 DVDD.n1101 0.01022
R6122 DVDD.n1103 DVDD.n1102 0.01022
R6123 DVDD.n1104 DVDD.n1103 0.01022
R6124 DVDD.n1105 DVDD.n1104 0.01022
R6125 DVDD.n1106 DVDD.n1105 0.01022
R6126 DVDD.n1107 DVDD.n1106 0.01022
R6127 DVDD.n1108 DVDD.n1107 0.01022
R6128 DVDD.n1109 DVDD.n1108 0.01022
R6129 DVDD.n1110 DVDD.n1109 0.01022
R6130 DVDD.n1111 DVDD.n1110 0.01022
R6131 DVDD.n1112 DVDD.n1111 0.01022
R6132 DVDD.n1113 DVDD.n1112 0.01022
R6133 DVDD.n1114 DVDD.n1113 0.01022
R6134 DVDD.n1115 DVDD.n1114 0.01022
R6135 DVDD.n1116 DVDD.n1115 0.01022
R6136 DVDD.n1117 DVDD.n1116 0.01022
R6137 DVDD.n1118 DVDD.n1117 0.01022
R6138 DVDD.n1119 DVDD.n1118 0.01022
R6139 DVDD.n1539 DVDD.n1119 0.01022
R6140 DVDD.n1006 DVDD.n1005 0.01022
R6141 DVDD.n1005 DVDD.n1004 0.01022
R6142 DVDD.n1004 DVDD.n1003 0.01022
R6143 DVDD.n1003 DVDD.n1002 0.01022
R6144 DVDD.n1002 DVDD.n1001 0.01022
R6145 DVDD.n1001 DVDD.n1000 0.01022
R6146 DVDD.n1000 DVDD.n999 0.01022
R6147 DVDD.n964 DVDD.n963 0.01022
R6148 DVDD.n963 DVDD.n962 0.01022
R6149 DVDD.n962 DVDD.n961 0.01022
R6150 DVDD.n961 DVDD.n960 0.01022
R6151 DVDD.n960 DVDD.n958 0.01022
R6152 DVDD.n1679 DVDD.n958 0.01022
R6153 DVDD.n928 DVDD.n927 0.01022
R6154 DVDD.n927 DVDD.n926 0.01022
R6155 DVDD.n11572 DVDD.n11571 0.01022
R6156 DVDD.n11571 DVDD.n11570 0.01022
R6157 DVDD.n11570 DVDD.n11569 0.01022
R6158 DVDD.n11569 DVDD.n11568 0.01022
R6159 DVDD.n11568 DVDD.n11567 0.01022
R6160 DVDD.n11567 DVDD.n11566 0.01022
R6161 DVDD.n11566 DVDD.n11565 0.01022
R6162 DVDD.n11565 DVDD.n11564 0.01022
R6163 DVDD.n11564 DVDD.n11563 0.01022
R6164 DVDD.n11563 DVDD.n11562 0.01022
R6165 DVDD.n11562 DVDD.n11561 0.01022
R6166 DVDD.n11561 DVDD.n11560 0.01022
R6167 DVDD.n11560 DVDD.n11559 0.01022
R6168 DVDD.n11559 DVDD.n11558 0.01022
R6169 DVDD.n11558 DVDD.n11557 0.01022
R6170 DVDD.n11557 DVDD.n11556 0.01022
R6171 DVDD.n11556 DVDD.n11555 0.01022
R6172 DVDD.n11555 DVDD.n11554 0.01022
R6173 DVDD.n11554 DVDD.n11553 0.01022
R6174 DVDD.n11553 DVDD.n11552 0.01022
R6175 DVDD.n11552 DVDD.n11551 0.01022
R6176 DVDD.n11551 DVDD.n11550 0.01022
R6177 DVDD.n11550 DVDD.n11549 0.01022
R6178 DVDD.n11549 DVDD.n11548 0.01022
R6179 DVDD.n11548 DVDD.n11547 0.01022
R6180 DVDD.n11547 DVDD.n11546 0.01022
R6181 DVDD.n18312 DVDD.n18311 0.01022
R6182 DVDD.n18311 DVDD.n18310 0.01022
R6183 DVDD.n18310 DVDD.n18309 0.01022
R6184 DVDD.n18309 DVDD.n18308 0.01022
R6185 DVDD.n18308 DVDD.n18307 0.01022
R6186 DVDD.n18307 DVDD.n18306 0.01022
R6187 DVDD.n18306 DVDD.n18305 0.01022
R6188 DVDD.n18305 DVDD.n18304 0.01022
R6189 DVDD.n18304 DVDD.n18303 0.01022
R6190 DVDD.n18303 DVDD.n18302 0.01022
R6191 DVDD.n18302 DVDD.n18301 0.01022
R6192 DVDD.n18301 DVDD.n18300 0.01022
R6193 DVDD.n18300 DVDD.n18299 0.01022
R6194 DVDD.n18299 DVDD.n18298 0.01022
R6195 DVDD.n18298 DVDD.n18297 0.01022
R6196 DVDD.n18297 DVDD.n18296 0.01022
R6197 DVDD.n18296 DVDD.n18295 0.01022
R6198 DVDD.n18295 DVDD.n18294 0.01022
R6199 DVDD.n18294 DVDD.n18293 0.01022
R6200 DVDD.n18293 DVDD.n18292 0.01022
R6201 DVDD.n11902 DVDD.n11901 0.01022
R6202 DVDD.n11903 DVDD.n11902 0.01022
R6203 DVDD.n1295 DVDD.n1294 0.01022
R6204 DVDD.n1294 DVDD.n1293 0.01022
R6205 DVDD.n1293 DVDD.n1292 0.01022
R6206 DVDD.n1292 DVDD.n1291 0.01022
R6207 DVDD.n1291 DVDD.n1290 0.01022
R6208 DVDD.n1290 DVDD.n1289 0.01022
R6209 DVDD.n1289 DVDD.n1288 0.01022
R6210 DVDD.n11332 DVDD.n11331 0.01022
R6211 DVDD.n11331 DVDD.n11330 0.01022
R6212 DVDD.n11330 DVDD.n11329 0.01022
R6213 DVDD.n11329 DVDD.n11328 0.01022
R6214 DVDD.n11328 DVDD.n11327 0.01022
R6215 DVDD.n11327 DVDD.n11326 0.01022
R6216 DVDD.n11326 DVDD.n11325 0.01022
R6217 DVDD.n11325 DVDD.n11324 0.01022
R6218 DVDD.n11324 DVDD.n11323 0.01022
R6219 DVDD.n11323 DVDD.n11322 0.01022
R6220 DVDD.n11322 DVDD.n11321 0.01022
R6221 DVDD.n11321 DVDD.n11320 0.01022
R6222 DVDD.n11320 DVDD.n11319 0.01022
R6223 DVDD.n11319 DVDD.n11318 0.01022
R6224 DVDD.n11318 DVDD.n11317 0.01022
R6225 DVDD.n11317 DVDD.n11316 0.01022
R6226 DVDD.n11316 DVDD.n11315 0.01022
R6227 DVDD.n13174 DVDD.n13173 0.01022
R6228 DVDD.n13175 DVDD.n13174 0.01022
R6229 DVDD.n3308 DVDD.n3307 0.01022
R6230 DVDD.n3309 DVDD.n3308 0.01022
R6231 DVDD.n3310 DVDD.n3309 0.01022
R6232 DVDD.n3311 DVDD.n3310 0.01022
R6233 DVDD.n3312 DVDD.n3311 0.01022
R6234 DVDD.n3313 DVDD.n3312 0.01022
R6235 DVDD.n3314 DVDD.n3313 0.01022
R6236 DVDD.n17456 DVDD.n17455 0.0102034
R6237 DVDD.n12202 DVDD.n12201 0.0101938
R6238 DVDD.n13695 DVDD.n13694 0.01017
R6239 DVDD.n5956 DVDD.n5955 0.01017
R6240 DVDD.n12619 DVDD.n12618 0.01017
R6241 DVDD.n762 DVDD.n761 0.01017
R6242 DVDD.n799 DVDD.n798 0.01017
R6243 DVDD.n18141 DVDD.n18140 0.01017
R6244 DVDD.n17772 DVDD.n17771 0.01017
R6245 DVDD.n18002 DVDD.n18001 0.01017
R6246 DVDD.n18080 DVDD.n18079 0.01017
R6247 DVDD.n9447 DVDD.n9446 0.0101025
R6248 DVDD.n13505 DVDD.n13504 0.0100815
R6249 DVDD.n13607 DVDD.n13606 0.0100815
R6250 DVDD.n13688 DVDD.n13687 0.0100815
R6251 DVDD.n13557 DVDD.n13556 0.0100815
R6252 DVDD.n13638 DVDD.n13637 0.0100815
R6253 DVDD.n5471 DVDD.n5470 0.0100815
R6254 DVDD.n5691 DVDD.n5690 0.0100815
R6255 DVDD.n5963 DVDD.n5962 0.0100815
R6256 DVDD.n5594 DVDD.n5593 0.0100815
R6257 DVDD.n12992 DVDD.n12991 0.0100815
R6258 DVDD.n12750 DVDD.n12749 0.0100815
R6259 DVDD.n12626 DVDD.n12625 0.0100815
R6260 DVDD.n12833 DVDD.n12832 0.0100815
R6261 DVDD.n788 DVDD.n787 0.0100815
R6262 DVDD.n825 DVDD.n824 0.0100815
R6263 DVDD.n18148 DVDD.n18147 0.0100815
R6264 DVDD.n18054 DVDD.n18053 0.0100815
R6265 DVDD.n17976 DVDD.n17975 0.0100815
R6266 DVDD.n17874 DVDD.n17873 0.0100815
R6267 DVDD.n17779 DVDD.n17778 0.0100815
R6268 DVDD.n18198 DVDD.n18197 0.0100815
R6269 DVDD.n17843 DVDD.n17842 0.0100815
R6270 DVDD.n17924 DVDD.n17923 0.0100815
R6271 DVDD.n12253 DVDD.n12252 0.0100669
R6272 DVDD.n13347 DVDD.n13346 0.0100669
R6273 DVDD.n14426 DVDD.n14425 0.0100669
R6274 DVDD.n5984 DVDD.n5983 0.0100669
R6275 DVDD.n12647 DVDD.n12646 0.0100669
R6276 DVDD.n17800 DVDD.n17799 0.0100669
R6277 DVDD.n4447 DVDD.n4446 0.0100669
R6278 DVDD.n8721 DVDD.n8720 0.0100669
R6279 DVDD.n7733 DVDD.n7732 0.01004
R6280 DVDD.n3457 DVDD.n3456 0.01004
R6281 DVDD.n3570 DVDD.n3569 0.01004
R6282 DVDD.n9963 DVDD.n9962 0.01004
R6283 DVDD.n2058 DVDD.n2057 0.01004
R6284 DVDD.n2212 DVDD.n2211 0.01004
R6285 DVDD.n7036 DVDD.n7035 0.01004
R6286 DVDD.n6946 DVDD.n6945 0.01004
R6287 DVDD.n1865 DVDD.n1864 0.01004
R6288 DVDD.n19836 DVDD.n19835 0.01004
R6289 DVDD.n19991 DVDD.n19990 0.01004
R6290 DVDD.n4616 DVDD.n4615 0.01004
R6291 DVDD.n4720 DVDD.n4719 0.01004
R6292 DVDD.n19643 DVDD.n19642 0.01004
R6293 DVDD.n1540 DVDD.n1539 0.01004
R6294 DVDD.n1679 DVDD.n1678 0.01004
R6295 DVDD.n11546 DVDD.n11545 0.01004
R6296 DVDD.n18292 DVDD.n18291 0.01004
R6297 DVDD.n1288 DVDD.n1287 0.01004
R6298 DVDD.n3315 DVDD.n3314 0.01004
R6299 DVDD.n13665 DVDD.n13664 0.00999298
R6300 DVDD.n13584 DVDD.n13583 0.00999298
R6301 DVDD.n5645 DVDD.n5644 0.00999298
R6302 DVDD.n12792 DVDD.n12791 0.00999298
R6303 DVDD.n18171 DVDD.n18170 0.00999298
R6304 DVDD.n17897 DVDD.n17896 0.00999298
R6305 DVDD.n3679 DVDD.n3678 0.00995
R6306 DVDD.n2996 DVDD.n2995 0.00995
R6307 DVDD.n2921 DVDD.n2920 0.00995
R6308 DVDD.n9989 DVDD.n7157 0.00995
R6309 DVDD.n2027 DVDD.n2026 0.00995
R6310 DVDD.n2159 DVDD.n2158 0.00995
R6311 DVDD.n2235 DVDD.n2234 0.00995
R6312 DVDD.n6972 DVDD.n6940 0.00995
R6313 DVDD.n19805 DVDD.n19804 0.00995
R6314 DVDD.n19938 DVDD.n19937 0.00995
R6315 DVDD.n20014 DVDD.n20013 0.00995
R6316 DVDD.n4746 DVDD.n4714 0.00995
R6317 DVDD.n1094 DVDD.n1093 0.00995
R6318 DVDD.n1007 DVDD.n1006 0.00995
R6319 DVDD.n1728 DVDD.n1727 0.00995
R6320 DVDD.n11572 DVDD.n11417 0.00995
R6321 DVDD.n3445 DVDD.n3444 0.00995
R6322 DVDD.n3425 DVDD.n3424 0.00995
R6323 DVDD.n3582 DVDD.n3581 0.00995
R6324 DVDD.n3653 DVDD.n3652 0.00995
R6325 DVDD.n3591 DVDD.n3590 0.00995
R6326 DVDD.n18582 DVDD.n18581 0.00995
R6327 DVDD.n18344 DVDD.n18343 0.00995
R6328 DVDD.n7809 DVDD.n7808 0.00995
R6329 DVDD.n8065 DVDD.n8064 0.00991423
R6330 DVDD.n12233 DVDD.n12232 0.00988976
R6331 DVDD.n20186 DVDD.n20185 0.00988976
R6332 DVDD.n4968 DVDD.n4967 0.00988976
R6333 DVDD.n264 DVDD.n263 0.00988976
R6334 DVDD.n11785 DVDD.n11784 0.00988976
R6335 DVDD.n19571 DVDD.n19570 0.00988976
R6336 DVDD.n6716 DVDD.n6715 0.00988976
R6337 DVDD.n3750 DVDD.n3749 0.00988976
R6338 DVDD.n9684 DVDD.n9683 0.00988976
R6339 DVDD.n7789 DVDD.n7694 0.00986
R6340 DVDD.n10146 DVDD.n10145 0.00986
R6341 DVDD.n17294 DVDD.n17291 0.00982432
R6342 DVDD.n13911 DVDD.n13908 0.00982432
R6343 DVDD.n17673 DVDD.n17670 0.00982432
R6344 DVDD.n14300 DVDD.n14297 0.00982432
R6345 DVDD.n7772 DVDD.n7771 0.00977
R6346 DVDD.n3448 DVDD.n3447 0.00977
R6347 DVDD.n3579 DVDD.n3578 0.00977
R6348 DVDD.n9954 DVDD.n9953 0.00977
R6349 DVDD.n9819 DVDD.n9818 0.00977
R6350 DVDD.n9515 DVDD.n9514 0.00977
R6351 DVDD.n1549 DVDD.n1548 0.00977
R6352 DVDD.n1671 DVDD.n1670 0.00977
R6353 DVDD.n11538 DVDD.n11537 0.00977
R6354 DVDD.n10128 DVDD.n10127 0.00977
R6355 DVDD.n11920 DVDD.n11919 0.00977
R6356 DVDD.n1280 DVDD.n1279 0.00977
R6357 DVDD.n12320 DVDD.n12319 0.00977
R6358 DVDD.n3324 DVDD.n3323 0.00977
R6359 DVDD.n8001 DVDD.n8000 0.00972594
R6360 DVDD.n8089 DVDD.n8088 0.00972594
R6361 DVDD.n12176 DVDD.n12175 0.0097126
R6362 DVDD.n12234 DVDD.n12233 0.0097126
R6363 DVDD.n20091 DVDD.n20090 0.0097126
R6364 DVDD.n5193 DVDD.n5192 0.0097126
R6365 DVDD.n19189 DVDD.n19188 0.0097126
R6366 DVDD.n12373 DVDD.n12372 0.0097126
R6367 DVDD.n19476 DVDD.n19475 0.0097126
R6368 DVDD.n6489 DVDD.n6488 0.0097126
R6369 DVDD.n18493 DVDD.n18492 0.0097126
R6370 DVDD.n8394 DVDD.n8393 0.0097126
R6371 DVDD.n3670 DVDD.n3669 0.00968
R6372 DVDD.n18643 DVDD.n18642 0.00968
R6373 DVDD.n3005 DVDD.n3004 0.00968
R6374 DVDD.n2912 DVDD.n2911 0.00968
R6375 DVDD.n9930 DVDD.n7165 0.00968
R6376 DVDD.n1085 DVDD.n1084 0.00968
R6377 DVDD.n1016 DVDD.n1015 0.00968
R6378 DVDD.n1737 DVDD.n1736 0.00968
R6379 DVDD.n1755 DVDD.n1754 0.00968
R6380 DVDD.n11514 DVDD.n11426 0.00968
R6381 DVDD.n11260 DVDD.n11259 0.00962857
R6382 DVDD.n11259 DVDD.n11258 0.00962857
R6383 DVDD.n11258 DVDD.n11257 0.00962857
R6384 DVDD.n11257 DVDD.n11256 0.00962857
R6385 DVDD.n11256 DVDD.n11255 0.00962857
R6386 DVDD.n11248 DVDD.n11247 0.00962857
R6387 DVDD.n11247 DVDD.n11246 0.00962857
R6388 DVDD.n11246 DVDD.n11245 0.00962857
R6389 DVDD.n11245 DVDD.n11244 0.00962857
R6390 DVDD.n11244 DVDD.n11243 0.00962857
R6391 DVDD.n11243 DVDD.n11242 0.00962857
R6392 DVDD.n11242 DVDD.n11241 0.00962857
R6393 DVDD.n11241 DVDD.n11240 0.00962857
R6394 DVDD.n11240 DVDD.n11239 0.00962857
R6395 DVDD.n11232 DVDD.n11231 0.00962857
R6396 DVDD.n11231 DVDD.n11230 0.00962857
R6397 DVDD.n11230 DVDD.n11229 0.00962857
R6398 DVDD.n11229 DVDD.n11228 0.00962857
R6399 DVDD.n11228 DVDD.n11227 0.00962857
R6400 DVDD.n11227 DVDD.n11226 0.00962857
R6401 DVDD.n11226 DVDD.n11225 0.00962857
R6402 DVDD.n5730 DVDD.n5729 0.00962857
R6403 DVDD.n5736 DVDD.n5735 0.00962857
R6404 DVDD.n5755 DVDD.n5754 0.00962857
R6405 DVDD.n5751 DVDD.n5750 0.00962857
R6406 DVDD.n5750 DVDD.n5749 0.00962857
R6407 DVDD.n4113 DVDD.n4112 0.00962857
R6408 DVDD.n4114 DVDD.n4113 0.00962857
R6409 DVDD.n4118 DVDD.n4117 0.00962857
R6410 DVDD.n4122 DVDD.n4121 0.00962857
R6411 DVDD.n4126 DVDD.n4125 0.00962857
R6412 DVDD.n4153 DVDD.n4152 0.00962857
R6413 DVDD.n4152 DVDD.n4151 0.00962857
R6414 DVDD.n4142 DVDD.n4141 0.00962857
R6415 DVDD.n4138 DVDD.n4137 0.00962857
R6416 DVDD.n8502 DVDD.n8501 0.00962857
R6417 DVDD.n8507 DVDD.n8506 0.00962857
R6418 DVDD.n8508 DVDD.n8507 0.00962857
R6419 DVDD.n8535 DVDD.n8534 0.00962857
R6420 DVDD.n8522 DVDD.n8521 0.00962857
R6421 DVDD.n13867 DVDD.n13866 0.00962857
R6422 DVDD.n298 DVDD.n297 0.00962857
R6423 DVDD.n297 DVDD.n296 0.00962857
R6424 DVDD.n296 DVDD.n295 0.00962857
R6425 DVDD.n295 DVDD.n294 0.00962857
R6426 DVDD.n473 DVDD.n472 0.00962857
R6427 DVDD.n2418 DVDD.n2417 0.00962857
R6428 DVDD.n394 DVDD.n393 0.00962857
R6429 DVDD.n395 DVDD.n394 0.00962857
R6430 DVDD.n396 DVDD.n395 0.00962857
R6431 DVDD.n398 DVDD.n396 0.00962857
R6432 DVDD.n520 DVDD.n518 0.00962857
R6433 DVDD.n518 DVDD.n516 0.00962857
R6434 DVDD.n516 DVDD.n514 0.00962857
R6435 DVDD.n514 DVDD.n512 0.00962857
R6436 DVDD.n512 DVDD.n510 0.00962857
R6437 DVDD.n510 DVDD.n508 0.00962857
R6438 DVDD.n508 DVDD.n506 0.00962857
R6439 DVDD.n506 DVDD.n504 0.00962857
R6440 DVDD.n478 DVDD.n476 0.00962857
R6441 DVDD.n476 DVDD.n474 0.00962857
R6442 DVDD.n474 DVDD.n471 0.00962857
R6443 DVDD.n471 DVDD.n470 0.00962857
R6444 DVDD.n470 DVDD.n468 0.00962857
R6445 DVDD.n468 DVDD.n466 0.00962857
R6446 DVDD.n466 DVDD.n464 0.00962857
R6447 DVDD.n464 DVDD.n462 0.00962857
R6448 DVDD.n462 DVDD.n460 0.00962857
R6449 DVDD.n460 DVDD.n458 0.00962857
R6450 DVDD.n458 DVDD.n456 0.00962857
R6451 DVDD.n456 DVDD.n454 0.00962857
R6452 DVDD.n430 DVDD.n428 0.00962857
R6453 DVDD.n428 DVDD.n426 0.00962857
R6454 DVDD.n426 DVDD.n424 0.00962857
R6455 DVDD.n424 DVDD.n422 0.00962857
R6456 DVDD.n422 DVDD.n420 0.00962857
R6457 DVDD.n420 DVDD.n418 0.00962857
R6458 DVDD.n418 DVDD.n416 0.00962857
R6459 DVDD.n2305 DVDD.n2303 0.00962857
R6460 DVDD.n2307 DVDD.n2305 0.00962857
R6461 DVDD.n2309 DVDD.n2307 0.00962857
R6462 DVDD.n2311 DVDD.n2309 0.00962857
R6463 DVDD.n2313 DVDD.n2311 0.00962857
R6464 DVDD.n2315 DVDD.n2313 0.00962857
R6465 DVDD.n2317 DVDD.n2315 0.00962857
R6466 DVDD.n2350 DVDD.n2348 0.00962857
R6467 DVDD.n2352 DVDD.n2350 0.00962857
R6468 DVDD.n2354 DVDD.n2352 0.00962857
R6469 DVDD.n2356 DVDD.n2354 0.00962857
R6470 DVDD.n2358 DVDD.n2356 0.00962857
R6471 DVDD.n2360 DVDD.n2358 0.00962857
R6472 DVDD.n2362 DVDD.n2360 0.00962857
R6473 DVDD.n2364 DVDD.n2362 0.00962857
R6474 DVDD.n2366 DVDD.n2364 0.00962857
R6475 DVDD.n2368 DVDD.n2366 0.00962857
R6476 DVDD.n2370 DVDD.n2368 0.00962857
R6477 DVDD.n2372 DVDD.n2370 0.00962857
R6478 DVDD.n2405 DVDD.n2403 0.00962857
R6479 DVDD.n2407 DVDD.n2405 0.00962857
R6480 DVDD.n2409 DVDD.n2407 0.00962857
R6481 DVDD.n2411 DVDD.n2409 0.00962857
R6482 DVDD.n2413 DVDD.n2411 0.00962857
R6483 DVDD.n2415 DVDD.n2413 0.00962857
R6484 DVDD.n2416 DVDD.n2415 0.00962857
R6485 DVDD.n2419 DVDD.n2416 0.00962857
R6486 DVDD.n2460 DVDD.n2458 0.00962857
R6487 DVDD.n2462 DVDD.n2460 0.00962857
R6488 DVDD.n2464 DVDD.n2462 0.00962857
R6489 DVDD.n2467 DVDD.n2464 0.00962857
R6490 DVDD.n2484 DVDD.n2482 0.00962857
R6491 DVDD.n529 DVDD.n528 0.00962857
R6492 DVDD.n528 DVDD.n527 0.00962857
R6493 DVDD.n527 DVDD.n526 0.00962857
R6494 DVDD.n526 DVDD.n525 0.00962857
R6495 DVDD.n699 DVDD.n698 0.00962857
R6496 DVDD.n661 DVDD.n660 0.00962857
R6497 DVDD.n2510 DVDD.n2509 0.00962857
R6498 DVDD.n2563 DVDD.n2562 0.00962857
R6499 DVDD.n625 DVDD.n624 0.00962857
R6500 DVDD.n626 DVDD.n625 0.00962857
R6501 DVDD.n627 DVDD.n626 0.00962857
R6502 DVDD.n629 DVDD.n627 0.00962857
R6503 DVDD.n750 DVDD.n748 0.00962857
R6504 DVDD.n748 DVDD.n746 0.00962857
R6505 DVDD.n746 DVDD.n744 0.00962857
R6506 DVDD.n744 DVDD.n742 0.00962857
R6507 DVDD.n742 DVDD.n740 0.00962857
R6508 DVDD.n740 DVDD.n738 0.00962857
R6509 DVDD.n738 DVDD.n736 0.00962857
R6510 DVDD.n736 DVDD.n734 0.00962857
R6511 DVDD.n710 DVDD.n708 0.00962857
R6512 DVDD.n708 DVDD.n706 0.00962857
R6513 DVDD.n706 DVDD.n704 0.00962857
R6514 DVDD.n704 DVDD.n702 0.00962857
R6515 DVDD.n702 DVDD.n700 0.00962857
R6516 DVDD.n700 DVDD.n697 0.00962857
R6517 DVDD.n697 DVDD.n696 0.00962857
R6518 DVDD.n696 DVDD.n694 0.00962857
R6519 DVDD.n694 DVDD.n692 0.00962857
R6520 DVDD.n692 DVDD.n690 0.00962857
R6521 DVDD.n690 DVDD.n688 0.00962857
R6522 DVDD.n688 DVDD.n686 0.00962857
R6523 DVDD.n662 DVDD.n659 0.00962857
R6524 DVDD.n659 DVDD.n658 0.00962857
R6525 DVDD.n658 DVDD.n656 0.00962857
R6526 DVDD.n656 DVDD.n654 0.00962857
R6527 DVDD.n654 DVDD.n652 0.00962857
R6528 DVDD.n652 DVDD.n650 0.00962857
R6529 DVDD.n650 DVDD.n648 0.00962857
R6530 DVDD.n2505 DVDD.n2503 0.00962857
R6531 DVDD.n2507 DVDD.n2505 0.00962857
R6532 DVDD.n2508 DVDD.n2507 0.00962857
R6533 DVDD.n2511 DVDD.n2508 0.00962857
R6534 DVDD.n2513 DVDD.n2511 0.00962857
R6535 DVDD.n2515 DVDD.n2513 0.00962857
R6536 DVDD.n2517 DVDD.n2515 0.00962857
R6537 DVDD.n2548 DVDD.n2546 0.00962857
R6538 DVDD.n2550 DVDD.n2548 0.00962857
R6539 DVDD.n2552 DVDD.n2550 0.00962857
R6540 DVDD.n2554 DVDD.n2552 0.00962857
R6541 DVDD.n2556 DVDD.n2554 0.00962857
R6542 DVDD.n2558 DVDD.n2556 0.00962857
R6543 DVDD.n2560 DVDD.n2558 0.00962857
R6544 DVDD.n2561 DVDD.n2560 0.00962857
R6545 DVDD.n2564 DVDD.n2561 0.00962857
R6546 DVDD.n2566 DVDD.n2564 0.00962857
R6547 DVDD.n2568 DVDD.n2566 0.00962857
R6548 DVDD.n2570 DVDD.n2568 0.00962857
R6549 DVDD.n2601 DVDD.n2599 0.00962857
R6550 DVDD.n2603 DVDD.n2601 0.00962857
R6551 DVDD.n2605 DVDD.n2603 0.00962857
R6552 DVDD.n2607 DVDD.n2605 0.00962857
R6553 DVDD.n2609 DVDD.n2607 0.00962857
R6554 DVDD.n2611 DVDD.n2609 0.00962857
R6555 DVDD.n2613 DVDD.n2611 0.00962857
R6556 DVDD.n2615 DVDD.n2613 0.00962857
R6557 DVDD.n2658 DVDD.n2656 0.00962857
R6558 DVDD.n2660 DVDD.n2658 0.00962857
R6559 DVDD.n2662 DVDD.n2660 0.00962857
R6560 DVDD.n2665 DVDD.n2662 0.00962857
R6561 DVDD.n11291 DVDD.n11290 0.00962857
R6562 DVDD.n11290 DVDD.n11289 0.00962857
R6563 DVDD.n11289 DVDD.n11288 0.00962857
R6564 DVDD.n11288 DVDD.n11287 0.00962857
R6565 DVDD.n11273 DVDD.n11272 0.00962857
R6566 DVDD.n11272 DVDD.n11271 0.00962857
R6567 DVDD.n11271 DVDD.n11270 0.00962857
R6568 DVDD.n11270 DVDD.n11269 0.00962857
R6569 DVDD.n11269 DVDD.n11268 0.00962857
R6570 DVDD.n11268 DVDD.n11267 0.00962857
R6571 DVDD.n12486 DVDD.n12485 0.00962857
R6572 DVDD.n12497 DVDD.n12496 0.00962857
R6573 DVDD.n12496 DVDD.n12495 0.00962857
R6574 DVDD.n12495 DVDD.n12494 0.00962857
R6575 DVDD.n12494 DVDD.n12493 0.00962857
R6576 DVDD.n5725 DVDD.n5724 0.00962857
R6577 DVDD.n5727 DVDD.n5725 0.00962857
R6578 DVDD.n5728 DVDD.n5727 0.00962857
R6579 DVDD.n5731 DVDD.n5728 0.00962857
R6580 DVDD.n5733 DVDD.n5731 0.00962857
R6581 DVDD.n5734 DVDD.n5733 0.00962857
R6582 DVDD.n5737 DVDD.n5734 0.00962857
R6583 DVDD.n5760 DVDD.n5758 0.00962857
R6584 DVDD.n5758 DVDD.n5756 0.00962857
R6585 DVDD.n5756 DVDD.n5753 0.00962857
R6586 DVDD.n5753 DVDD.n5752 0.00962857
R6587 DVDD.n5752 DVDD.n5748 0.00962857
R6588 DVDD.n5748 DVDD.n5747 0.00962857
R6589 DVDD.n4111 DVDD.n4110 0.00962857
R6590 DVDD.n4115 DVDD.n4111 0.00962857
R6591 DVDD.n4116 DVDD.n4115 0.00962857
R6592 DVDD.n4119 DVDD.n4116 0.00962857
R6593 DVDD.n4120 DVDD.n4119 0.00962857
R6594 DVDD.n4123 DVDD.n4120 0.00962857
R6595 DVDD.n4124 DVDD.n4123 0.00962857
R6596 DVDD.n4127 DVDD.n4124 0.00962857
R6597 DVDD.n4146 DVDD.n4145 0.00962857
R6598 DVDD.n4145 DVDD.n4144 0.00962857
R6599 DVDD.n4144 DVDD.n4143 0.00962857
R6600 DVDD.n4143 DVDD.n4140 0.00962857
R6601 DVDD.n4140 DVDD.n4139 0.00962857
R6602 DVDD.n4139 DVDD.n4136 0.00962857
R6603 DVDD.n8500 DVDD.n8499 0.00962857
R6604 DVDD.n8503 DVDD.n8500 0.00962857
R6605 DVDD.n8504 DVDD.n8503 0.00962857
R6606 DVDD.n8505 DVDD.n8504 0.00962857
R6607 DVDD.n8509 DVDD.n8505 0.00962857
R6608 DVDD.n8529 DVDD.n8528 0.00962857
R6609 DVDD.n8528 DVDD.n8527 0.00962857
R6610 DVDD.n8527 DVDD.n8525 0.00962857
R6611 DVDD.n8525 DVDD.n8523 0.00962857
R6612 DVDD.n8523 DVDD.n8520 0.00962857
R6613 DVDD.n8520 DVDD.n8519 0.00962857
R6614 DVDD.n11211 DVDD.n11209 0.00962857
R6615 DVDD.n13861 DVDD.n13860 0.00962857
R6616 DVDD.n13860 DVDD.n13859 0.00962857
R6617 DVDD.n13859 DVDD.n13857 0.00962857
R6618 DVDD.n13857 DVDD.n13855 0.00962857
R6619 DVDD.n3680 DVDD.n3679 0.00959
R6620 DVDD.n2236 DVDD.n2235 0.00959
R6621 DVDD.n20015 DVDD.n20014 0.00959
R6622 DVDD.n1727 DVDD.n1726 0.00959
R6623 DVDD.n8272 DVDD.n8271 0.00953766
R6624 DVDD.n8110 DVDD.n8109 0.00953766
R6625 DVDD.n12252 DVDD.n12251 0.00953543
R6626 DVDD.n14427 DVDD.n14426 0.00953543
R6627 DVDD.n4981 DVDD.n4980 0.00953543
R6628 DVDD.n5058 DVDD.n5057 0.00953543
R6629 DVDD.n5985 DVDD.n5984 0.00953543
R6630 DVDD.n11772 DVDD.n11771 0.00953543
R6631 DVDD.n11696 DVDD.n11695 0.00953543
R6632 DVDD.n12648 DVDD.n12647 0.00953543
R6633 DVDD.n17801 DVDD.n17800 0.00953543
R6634 DVDD.n6703 DVDD.n6702 0.00953543
R6635 DVDD.n6624 DVDD.n6623 0.00953543
R6636 DVDD.n4448 DVDD.n4447 0.00953543
R6637 DVDD.n9671 DVDD.n9670 0.00953543
R6638 DVDD.n9592 DVDD.n9591 0.00953543
R6639 DVDD.n8722 DVDD.n8721 0.00953543
R6640 DVDD.n2872 DVDD.n2871 0.0095
R6641 DVDD.n1056 DVDD.n1055 0.0095
R6642 DVDD.n3368 DVDD.n3367 0.0095
R6643 DVDD.n18626 DVDD.n18625 0.0095
R6644 DVDD.n18641 DVDD.n18640 0.0095
R6645 DVDD.n14747 DVDD.n14746 0.0095
R6646 DVDD.n14752 DVDD.n14751 0.0095
R6647 DVDD.n14770 DVDD.n14769 0.0095
R6648 DVDD.n7693 DVDD.n7692 0.0095
R6649 DVDD.n13847 DVDD.n13846 0.00943572
R6650 DVDD.n2332 DVDD.n2331 0.00943572
R6651 DVDD.n2383 DVDD.n2382 0.00943572
R6652 DVDD.n2430 DVDD.n2429 0.00943572
R6653 DVDD.n2530 DVDD.n2529 0.00943572
R6654 DVDD.n2581 DVDD.n2580 0.00943572
R6655 DVDD.n2626 DVDD.n2625 0.00943572
R6656 DVDD.n11261 DVDD.n11260 0.00937143
R6657 DVDD.n11249 DVDD.n11248 0.00937143
R6658 DVDD.n11233 DVDD.n11232 0.00937143
R6659 DVDD.n299 DVDD.n298 0.00937143
R6660 DVDD.n530 DVDD.n529 0.00937143
R6661 DVDD.n12121 DVDD.n12120 0.00935827
R6662 DVDD.n13882 DVDD.n13881 0.00935592
R6663 DVDD.n17260 DVDD.n17259 0.00935592
R6664 DVDD.n8209 DVDD.n8208 0.00934937
R6665 DVDD.n9481 DVDD.n9480 0.00934937
R6666 DVDD.n7759 DVDD.n7758 0.00932
R6667 DVDD.n7756 DVDD.n7755 0.00932
R6668 DVDD.n7753 DVDD.n7752 0.00932
R6669 DVDD.n7750 DVDD.n7749 0.00932
R6670 DVDD.n7747 DVDD.n7746 0.00932
R6671 DVDD.n2863 DVDD.n2862 0.00932
R6672 DVDD.n2860 DVDD.n2859 0.00932
R6673 DVDD.n2857 DVDD.n2856 0.00932
R6674 DVDD.n2854 DVDD.n2853 0.00932
R6675 DVDD.n2851 DVDD.n2850 0.00932
R6676 DVDD.n2848 DVDD.n2847 0.00932
R6677 DVDD.n2845 DVDD.n2844 0.00932
R6678 DVDD.n2842 DVDD.n2841 0.00932
R6679 DVDD.n2839 DVDD.n2838 0.00932
R6680 DVDD.n2836 DVDD.n2835 0.00932
R6681 DVDD.n18745 DVDD.n18744 0.00932
R6682 DVDD.n18748 DVDD.n18747 0.00932
R6683 DVDD.n18751 DVDD.n18750 0.00932
R6684 DVDD.n18754 DVDD.n18753 0.00932
R6685 DVDD.n18757 DVDD.n18756 0.00932
R6686 DVDD.n18760 DVDD.n18759 0.00932
R6687 DVDD.n18763 DVDD.n18762 0.00932
R6688 DVDD.n18766 DVDD.n18765 0.00932
R6689 DVDD.n18769 DVDD.n18768 0.00932
R6690 DVDD.n2902 DVDD.n2901 0.00932
R6691 DVDD.n2899 DVDD.n2898 0.00932
R6692 DVDD.n2896 DVDD.n2895 0.00932
R6693 DVDD.n2893 DVDD.n2892 0.00932
R6694 DVDD.n2890 DVDD.n2889 0.00932
R6695 DVDD.n2887 DVDD.n2886 0.00932
R6696 DVDD.n2884 DVDD.n2883 0.00932
R6697 DVDD.n2881 DVDD.n2880 0.00932
R6698 DVDD.n2878 DVDD.n2877 0.00932
R6699 DVDD.n2875 DVDD.n2874 0.00932
R6700 DVDD.n9880 DVDD.n9879 0.00932
R6701 DVDD.n9877 DVDD.n9876 0.00932
R6702 DVDD.n9874 DVDD.n9873 0.00932
R6703 DVDD.n9871 DVDD.n9870 0.00932
R6704 DVDD.n9868 DVDD.n9867 0.00932
R6705 DVDD.n9865 DVDD.n9864 0.00932
R6706 DVDD.n9862 DVDD.n9861 0.00932
R6707 DVDD.n9859 DVDD.n9858 0.00932
R6708 DVDD.n9856 DVDD.n9855 0.00932
R6709 DVDD.n9853 DVDD.n9852 0.00932
R6710 DVDD.n9850 DVDD.n9849 0.00932
R6711 DVDD.n9847 DVDD.n9846 0.00932
R6712 DVDD.n9844 DVDD.n9843 0.00932
R6713 DVDD.n9841 DVDD.n9840 0.00932
R6714 DVDD.n9838 DVDD.n9837 0.00932
R6715 DVDD.n9835 DVDD.n9834 0.00932
R6716 DVDD.n9832 DVDD.n9831 0.00932
R6717 DVDD.n9829 DVDD.n9828 0.00932
R6718 DVDD.n9826 DVDD.n9825 0.00932
R6719 DVDD.n9385 DVDD.n9384 0.00932
R6720 DVDD.n9382 DVDD.n9381 0.00932
R6721 DVDD.n9379 DVDD.n9378 0.00932
R6722 DVDD.n9376 DVDD.n9375 0.00932
R6723 DVDD.n9373 DVDD.n9372 0.00932
R6724 DVDD.n9370 DVDD.n9369 0.00932
R6725 DVDD.n9367 DVDD.n9366 0.00932
R6726 DVDD.n9360 DVDD.n9359 0.00932
R6727 DVDD.n9357 DVDD.n9356 0.00932
R6728 DVDD.n9354 DVDD.n9353 0.00932
R6729 DVDD.n9351 DVDD.n9350 0.00932
R6730 DVDD.n9348 DVDD.n9347 0.00932
R6731 DVDD.n9345 DVDD.n9344 0.00932
R6732 DVDD.n9342 DVDD.n9341 0.00932
R6733 DVDD.n9339 DVDD.n9338 0.00932
R6734 DVDD.n9336 DVDD.n9335 0.00932
R6735 DVDD.n9333 DVDD.n9332 0.00932
R6736 DVDD.n9330 DVDD.n9329 0.00932
R6737 DVDD.n9327 DVDD.n9326 0.00932
R6738 DVDD.n9324 DVDD.n9323 0.00932
R6739 DVDD.n9321 DVDD.n9320 0.00932
R6740 DVDD.n1026 DVDD.n1025 0.00932
R6741 DVDD.n1029 DVDD.n1028 0.00932
R6742 DVDD.n1032 DVDD.n1031 0.00932
R6743 DVDD.n1035 DVDD.n1034 0.00932
R6744 DVDD.n1038 DVDD.n1037 0.00932
R6745 DVDD.n1041 DVDD.n1040 0.00932
R6746 DVDD.n1044 DVDD.n1043 0.00932
R6747 DVDD.n1047 DVDD.n1046 0.00932
R6748 DVDD.n1050 DVDD.n1049 0.00932
R6749 DVDD.n1053 DVDD.n1052 0.00932
R6750 DVDD.n1741 DVDD.n1740 0.00932
R6751 DVDD.n1781 DVDD.n1743 0.00932
R6752 DVDD.n1779 DVDD.n1778 0.00932
R6753 DVDD.n1776 DVDD.n1775 0.00932
R6754 DVDD.n1773 DVDD.n1772 0.00932
R6755 DVDD.n1770 DVDD.n1769 0.00932
R6756 DVDD.n1767 DVDD.n1766 0.00932
R6757 DVDD.n1764 DVDD.n1763 0.00932
R6758 DVDD.n1761 DVDD.n1760 0.00932
R6759 DVDD.n1758 DVDD.n1757 0.00932
R6760 DVDD.n1750 DVDD.n1749 0.00932
R6761 DVDD.n1747 DVDD.n1746 0.00932
R6762 DVDD.n19259 DVDD.n19258 0.00932
R6763 DVDD.n19262 DVDD.n19261 0.00932
R6764 DVDD.n19265 DVDD.n19264 0.00932
R6765 DVDD.n19416 DVDD.n19267 0.00932
R6766 DVDD.n19419 DVDD.n19418 0.00932
R6767 DVDD.n19422 DVDD.n19421 0.00932
R6768 DVDD.n18271 DVDD.n18270 0.00932
R6769 DVDD.n18268 DVDD.n18267 0.00932
R6770 DVDD.n10155 DVDD.n10154 0.00932
R6771 DVDD.n10152 DVDD.n10151 0.00932
R6772 DVDD.n10149 DVDD.n10148 0.00932
R6773 DVDD.n11981 DVDD.n11980 0.00932
R6774 DVDD.n11978 DVDD.n11977 0.00932
R6775 DVDD.n11975 DVDD.n11974 0.00932
R6776 DVDD.n11972 DVDD.n11971 0.00932
R6777 DVDD.n11969 DVDD.n11968 0.00932
R6778 DVDD.n11966 DVDD.n11965 0.00932
R6779 DVDD.n11963 DVDD.n11962 0.00932
R6780 DVDD.n11960 DVDD.n11959 0.00932
R6781 DVDD.n11957 DVDD.n11956 0.00932
R6782 DVDD.n11954 DVDD.n11953 0.00932
R6783 DVDD.n11951 DVDD.n11950 0.00932
R6784 DVDD.n11948 DVDD.n11947 0.00932
R6785 DVDD.n11945 DVDD.n11944 0.00932
R6786 DVDD.n11942 DVDD.n11941 0.00932
R6787 DVDD.n11939 DVDD.n11938 0.00932
R6788 DVDD.n11936 DVDD.n11935 0.00932
R6789 DVDD.n11933 DVDD.n11932 0.00932
R6790 DVDD.n11930 DVDD.n11929 0.00932
R6791 DVDD.n11927 DVDD.n11926 0.00932
R6792 DVDD.n1243 DVDD.n1242 0.00932
R6793 DVDD.n1246 DVDD.n1245 0.00932
R6794 DVDD.n1249 DVDD.n1248 0.00932
R6795 DVDD.n1252 DVDD.n1251 0.00932
R6796 DVDD.n1255 DVDD.n1254 0.00932
R6797 DVDD.n1258 DVDD.n1257 0.00932
R6798 DVDD.n1261 DVDD.n1260 0.00932
R6799 DVDD.n1264 DVDD.n1263 0.00932
R6800 DVDD.n1267 DVDD.n1266 0.00932
R6801 DVDD.n1270 DVDD.n1269 0.00932
R6802 DVDD.n13296 DVDD.n13295 0.00932
R6803 DVDD.n13293 DVDD.n13292 0.00932
R6804 DVDD.n13290 DVDD.n13289 0.00932
R6805 DVDD.n13287 DVDD.n13286 0.00932
R6806 DVDD.n13284 DVDD.n13283 0.00932
R6807 DVDD.n13281 DVDD.n13280 0.00932
R6808 DVDD.n13278 DVDD.n13277 0.00932
R6809 DVDD.n13271 DVDD.n13270 0.00932
R6810 DVDD.n13268 DVDD.n13267 0.00932
R6811 DVDD.n13265 DVDD.n13264 0.00932
R6812 DVDD.n13262 DVDD.n13261 0.00932
R6813 DVDD.n13259 DVDD.n13258 0.00932
R6814 DVDD.n13256 DVDD.n13255 0.00932
R6815 DVDD.n13253 DVDD.n13252 0.00932
R6816 DVDD.n13250 DVDD.n13249 0.00932
R6817 DVDD.n13247 DVDD.n13246 0.00932
R6818 DVDD.n13244 DVDD.n13243 0.00932
R6819 DVDD.n13241 DVDD.n13240 0.00932
R6820 DVDD.n13238 DVDD.n13237 0.00932
R6821 DVDD.n13235 DVDD.n13234 0.00932
R6822 DVDD.n13232 DVDD.n13231 0.00932
R6823 DVDD.n3155 DVDD.n3154 0.00932
R6824 DVDD.n3152 DVDD.n3151 0.00932
R6825 DVDD.n3149 DVDD.n3148 0.00932
R6826 DVDD.n3146 DVDD.n3145 0.00932
R6827 DVDD.n3143 DVDD.n3142 0.00932
R6828 DVDD.n3140 DVDD.n3139 0.00932
R6829 DVDD.n3137 DVDD.n3136 0.00932
R6830 DVDD.n3134 DVDD.n3133 0.00932
R6831 DVDD.n3131 DVDD.n3130 0.00932
R6832 DVDD.n3128 DVDD.n3127 0.00932
R6833 DVDD.n2929 DVDD.n2928 0.00923
R6834 DVDD.n2167 DVDD.n2166 0.00923
R6835 DVDD.n19946 DVDD.n19945 0.00923
R6836 DVDD.n999 DVDD.n998 0.00923
R6837 DVDD.n12055 DVDD.n12054 0.0091811
R6838 DVDD.n12148 DVDD.n12147 0.0091811
R6839 DVDD.n4676 DVDD.n4675 0.0091811
R6840 DVDD.n5067 DVDD.n5066 0.0091811
R6841 DVDD.n6091 DVDD.n6090 0.0091811
R6842 DVDD.n6041 DVDD.n6040 0.0091811
R6843 DVDD.n11383 DVDD.n11382 0.0091811
R6844 DVDD.n11687 DVDD.n11686 0.0091811
R6845 DVDD.n12723 DVDD.n12722 0.0091811
R6846 DVDD.n12687 DVDD.n12686 0.0091811
R6847 DVDD.n7008 DVDD.n7007 0.0091811
R6848 DVDD.n6615 DVDD.n6614 0.0091811
R6849 DVDD.n4541 DVDD.n4540 0.0091811
R6850 DVDD.n4492 DVDD.n4491 0.0091811
R6851 DVDD.n10025 DVDD.n10024 0.0091811
R6852 DVDD.n9583 DVDD.n9582 0.0091811
R6853 DVDD.n8808 DVDD.n8807 0.0091811
R6854 DVDD.n8773 DVDD.n8772 0.0091811
R6855 DVDD.n2466 DVDD.n2465 0.00917857
R6856 DVDD.n19532 DVDD.n19531 0.00917
R6857 DVDD.n20147 DVDD.n20146 0.00917
R6858 DVDD.n199 DVDD.n198 0.00917
R6859 DVDD.n18654 DVDD.n18653 0.00917
R6860 DVDD.n8233 DVDD.n8232 0.00916109
R6861 DVDD.n7762 DVDD.n7761 0.00914
R6862 DVDD.n9800 DVDD.n9799 0.00914
R6863 DVDD.n6815 DVDD.n6814 0.00914
R6864 DVDD.n4852 DVDD.n4851 0.00914
R6865 DVDD.n18274 DVDD.n18273 0.00914
R6866 DVDD.n11901 DVDD.n11900 0.00914
R6867 DVDD.n14118 DVDD.n14108 0.00911702
R6868 DVDD.n14019 DVDD.n14018 0.00911702
R6869 DVDD.n14231 DVDD.n14230 0.00911702
R6870 DVDD.n2963 DVDD.n2962 0.00905
R6871 DVDD.n2201 DVDD.n2200 0.00905
R6872 DVDD.n19980 DVDD.n19979 0.00905
R6873 DVDD.n965 DVDD.n964 0.00905
R6874 DVDD.n3421 DVDD.n3420 0.00905
R6875 DVDD.n3660 DVDD.n3659 0.00905
R6876 DVDD.n18596 DVDD.n18595 0.00905
R6877 DVDD.n7132 DVDD.n7131 0.00905
R6878 DVDD.n14749 DVDD.n14748 0.00905
R6879 DVDD.n14754 DVDD.n14753 0.00905
R6880 DVDD.n7168 DVDD.n7167 0.00905
R6881 DVDD.n5503 DVDD.n5502 0.00904661
R6882 DVDD.n5502 DVDD.n5501 0.00904661
R6883 DVDD.n6255 DVDD.n6254 0.00904661
R6884 DVDD.n6256 DVDD.n6255 0.00904661
R6885 DVDD.n12169 DVDD.n12168 0.00900394
R6886 DVDD.n13399 DVDD.n13398 0.00900394
R6887 DVDD.n5014 DVDD.n5013 0.00900394
R6888 DVDD.n11740 DVDD.n11739 0.00900394
R6889 DVDD.n6670 DVDD.n6669 0.00900394
R6890 DVDD.n9638 DVDD.n9637 0.00900394
R6891 DVDD.n9443 DVDD.n9442 0.0089728
R6892 DVDD.n8327 DVDD.n8326 0.0089728
R6893 DVDD.n18861 DVDD.n18860 0.00893
R6894 DVDD.n19110 DVDD.n19109 0.00893
R6895 DVDD.n19385 DVDD.n19384 0.00893
R6896 DVDD.n18381 DVDD.n18380 0.00893
R6897 DVDD.n17256 DVDD.n17198 0.00887766
R6898 DVDD.n17414 DVDD.n17365 0.00887766
R6899 DVDD.n17597 DVDD.n17526 0.00887766
R6900 DVDD.n1873 DVDD.n1872 0.00887
R6901 DVDD.n19651 DVDD.n19650 0.00887
R6902 DVDD.n1296 DVDD.n1295 0.00887
R6903 DVDD.n3307 DVDD.n3306 0.00887
R6904 DVDD.n12286 DVDD.n12285 0.00882677
R6905 DVDD.n13465 DVDD.n13464 0.00882677
R6906 DVDD.n4918 DVDD.n4917 0.00882677
R6907 DVDD.n5580 DVDD.n5579 0.00882677
R6908 DVDD.n11835 DVDD.n11834 0.00882677
R6909 DVDD.n12847 DVDD.n12846 0.00882677
R6910 DVDD.n6766 DVDD.n6765 0.00882677
R6911 DVDD.n6227 DVDD.n6226 0.00882677
R6912 DVDD.n9734 DVDD.n9733 0.00882677
R6913 DVDD.n8929 DVDD.n8928 0.00882677
R6914 DVDD.n9433 DVDD.n9432 0.00878452
R6915 DVDD.n5495 DVDD.n5494 0.0087818
R6916 DVDD.n12968 DVDD.n12967 0.0087818
R6917 DVDD.n6264 DVDD.n6263 0.0087818
R6918 DVDD.n6263 DVDD.n6262 0.0087818
R6919 DVDD.n9049 DVDD.n9048 0.0087818
R6920 DVDD.n9050 DVDD.n9049 0.0087818
R6921 DVDD.n3686 DVDD.n3685 0.00869
R6922 DVDD.n2242 DVDD.n2241 0.00869
R6923 DVDD.n20021 DVDD.n20020 0.00869
R6924 DVDD.n929 DVDD.n928 0.00869
R6925 DVDD.n11255 DVDD.n11254 0.00866429
R6926 DVDD.n11239 DVDD.n11238 0.00866429
R6927 DVDD.n13438 DVDD.n13437 0.00864961
R6928 DVDD.n5185 DVDD.n5184 0.00864961
R6929 DVDD.n12365 DVDD.n12364 0.00864961
R6930 DVDD.n6497 DVDD.n6496 0.00864961
R6931 DVDD.n8386 DVDD.n8385 0.00864961
R6932 DVDD.n12584 DVDD.n12583 0.00863101
R6933 DVDD.n4352 DVDD.n4351 0.00863101
R6934 DVDD.n8626 DVDD.n8625 0.00863101
R6935 DVDD.n7697 DVDD.n7696 0.0086
R6936 DVDD.n7700 DVDD.n7699 0.0086
R6937 DVDD.n7706 DVDD.n7705 0.0086
R6938 DVDD.n7709 DVDD.n7708 0.0086
R6939 DVDD.n3711 DVDD.n3710 0.0086
R6940 DVDD.n3708 DVDD.n3707 0.0086
R6941 DVDD.n3701 DVDD.n3700 0.0086
R6942 DVDD.n3698 DVDD.n3697 0.0086
R6943 DVDD.n3692 DVDD.n3691 0.0086
R6944 DVDD.n3689 DVDD.n3688 0.0086
R6945 DVDD.n18535 DVDD.n18534 0.0086
R6946 DVDD.n18538 DVDD.n18537 0.0086
R6947 DVDD.n18544 DVDD.n18543 0.0086
R6948 DVDD.n18547 DVDD.n18546 0.0086
R6949 DVDD.n18554 DVDD.n18553 0.0086
R6950 DVDD.n18557 DVDD.n18556 0.0086
R6951 DVDD.n2932 DVDD.n2931 0.0086
R6952 DVDD.n2938 DVDD.n2937 0.0086
R6953 DVDD.n2941 DVDD.n2940 0.0086
R6954 DVDD.n2948 DVDD.n2947 0.0086
R6955 DVDD.n2951 DVDD.n2950 0.0086
R6956 DVDD.n2954 DVDD.n2953 0.0086
R6957 DVDD.n2960 DVDD.n2959 0.0086
R6958 DVDD.n7825 DVDD.n7824 0.0086
R6959 DVDD.n7828 DVDD.n7827 0.0086
R6960 DVDD.n9754 DVDD.n9753 0.0086
R6961 DVDD.n9757 DVDD.n9756 0.0086
R6962 DVDD.n9760 DVDD.n9759 0.0086
R6963 DVDD.n9767 DVDD.n9766 0.0086
R6964 DVDD.n9770 DVDD.n9769 0.0086
R6965 DVDD.n9776 DVDD.n9775 0.0086
R6966 DVDD.n9779 DVDD.n9778 0.0086
R6967 DVDD.n9782 DVDD.n9781 0.0086
R6968 DVDD.n9785 DVDD.n9784 0.0086
R6969 DVDD.n9788 DVDD.n9787 0.0086
R6970 DVDD.n9791 DVDD.n9790 0.0086
R6971 DVDD.n9797 DVDD.n9796 0.0086
R6972 DVDD.n9806 DVDD.n9805 0.0086
R6973 DVDD.n9809 DVDD.n9808 0.0086
R6974 DVDD.n7910 DVDD.n7909 0.0086
R6975 DVDD.n7907 DVDD.n7906 0.0086
R6976 DVDD.n9539 DVDD.n7904 0.0086
R6977 DVDD.n9535 DVDD.n9534 0.0086
R6978 DVDD.n9532 DVDD.n9531 0.0086
R6979 DVDD.n9525 DVDD.n9524 0.0086
R6980 DVDD.n9241 DVDD.n9240 0.0086
R6981 DVDD.n9244 DVDD.n9243 0.0086
R6982 DVDD.n9247 DVDD.n9246 0.0086
R6983 DVDD.n9250 DVDD.n9249 0.0086
R6984 DVDD.n9256 DVDD.n9255 0.0086
R6985 DVDD.n9259 DVDD.n9258 0.0086
R6986 DVDD.n9268 DVDD.n9267 0.0086
R6987 DVDD.n9271 DVDD.n9270 0.0086
R6988 DVDD.n9277 DVDD.n9276 0.0086
R6989 DVDD.n9280 DVDD.n9279 0.0086
R6990 DVDD.n9283 DVDD.n9282 0.0086
R6991 DVDD.n9286 DVDD.n9285 0.0086
R6992 DVDD.n9289 DVDD.n9288 0.0086
R6993 DVDD.n9292 DVDD.n9291 0.0086
R6994 DVDD.n9298 DVDD.n9297 0.0086
R6995 DVDD.n9301 DVDD.n9300 0.0086
R6996 DVDD.n9308 DVDD.n9307 0.0086
R6997 DVDD.n2170 DVDD.n2169 0.0086
R6998 DVDD.n2176 DVDD.n2175 0.0086
R6999 DVDD.n2179 DVDD.n2178 0.0086
R7000 DVDD.n2186 DVDD.n2185 0.0086
R7001 DVDD.n2189 DVDD.n2188 0.0086
R7002 DVDD.n2192 DVDD.n2191 0.0086
R7003 DVDD.n2198 DVDD.n2197 0.0086
R7004 DVDD.n2267 DVDD.n2266 0.0086
R7005 DVDD.n2264 DVDD.n2263 0.0086
R7006 DVDD.n2257 DVDD.n2256 0.0086
R7007 DVDD.n2254 DVDD.n2253 0.0086
R7008 DVDD.n2248 DVDD.n2247 0.0086
R7009 DVDD.n2245 DVDD.n2244 0.0086
R7010 DVDD.n18904 DVDD.n18903 0.0086
R7011 DVDD.n18907 DVDD.n18906 0.0086
R7012 DVDD.n18913 DVDD.n18912 0.0086
R7013 DVDD.n18916 DVDD.n18915 0.0086
R7014 DVDD.n18923 DVDD.n18922 0.0086
R7015 DVDD.n18926 DVDD.n18925 0.0086
R7016 DVDD.n7069 DVDD.n7068 0.0086
R7017 DVDD.n7063 DVDD.n7062 0.0086
R7018 DVDD.n7060 DVDD.n7059 0.0086
R7019 DVDD.n6794 DVDD.n6793 0.0086
R7020 DVDD.n6797 DVDD.n6796 0.0086
R7021 DVDD.n6861 DVDD.n6860 0.0086
R7022 DVDD.n6858 DVDD.n6857 0.0086
R7023 DVDD.n6855 DVDD.n6854 0.0086
R7024 DVDD.n6848 DVDD.n6847 0.0086
R7025 DVDD.n6845 DVDD.n6844 0.0086
R7026 DVDD.n6839 DVDD.n6838 0.0086
R7027 DVDD.n6836 DVDD.n6835 0.0086
R7028 DVDD.n6833 DVDD.n6832 0.0086
R7029 DVDD.n6830 DVDD.n6829 0.0086
R7030 DVDD.n6827 DVDD.n6826 0.0086
R7031 DVDD.n6824 DVDD.n6823 0.0086
R7032 DVDD.n6818 DVDD.n6817 0.0086
R7033 DVDD.n6809 DVDD.n6808 0.0086
R7034 DVDD.n6806 DVDD.n6805 0.0086
R7035 DVDD.n6545 DVDD.n6544 0.0086
R7036 DVDD.n6548 DVDD.n6547 0.0086
R7037 DVDD.n6571 DVDD.n6550 0.0086
R7038 DVDD.n6567 DVDD.n6566 0.0086
R7039 DVDD.n6564 DVDD.n6563 0.0086
R7040 DVDD.n6557 DVDD.n6556 0.0086
R7041 DVDD.n1902 DVDD.n1901 0.0086
R7042 DVDD.n1896 DVDD.n1895 0.0086
R7043 DVDD.n1893 DVDD.n1892 0.0086
R7044 DVDD.n1886 DVDD.n1885 0.0086
R7045 DVDD.n1883 DVDD.n1882 0.0086
R7046 DVDD.n1876 DVDD.n1875 0.0086
R7047 DVDD.n4001 DVDD.n4000 0.0086
R7048 DVDD.n3998 DVDD.n3997 0.0086
R7049 DVDD.n3995 DVDD.n3994 0.0086
R7050 DVDD.n3992 DVDD.n3991 0.0086
R7051 DVDD.n3986 DVDD.n3985 0.0086
R7052 DVDD.n3983 DVDD.n3982 0.0086
R7053 DVDD.n3974 DVDD.n3973 0.0086
R7054 DVDD.n3971 DVDD.n3970 0.0086
R7055 DVDD.n3965 DVDD.n3964 0.0086
R7056 DVDD.n3962 DVDD.n3961 0.0086
R7057 DVDD.n3959 DVDD.n3958 0.0086
R7058 DVDD.n3956 DVDD.n3955 0.0086
R7059 DVDD.n3953 DVDD.n3952 0.0086
R7060 DVDD.n3950 DVDD.n3949 0.0086
R7061 DVDD.n3944 DVDD.n3943 0.0086
R7062 DVDD.n3941 DVDD.n3940 0.0086
R7063 DVDD.n3934 DVDD.n3933 0.0086
R7064 DVDD.n19949 DVDD.n19948 0.0086
R7065 DVDD.n19955 DVDD.n19954 0.0086
R7066 DVDD.n19958 DVDD.n19957 0.0086
R7067 DVDD.n19965 DVDD.n19964 0.0086
R7068 DVDD.n19968 DVDD.n19967 0.0086
R7069 DVDD.n19971 DVDD.n19970 0.0086
R7070 DVDD.n19977 DVDD.n19976 0.0086
R7071 DVDD.n20046 DVDD.n20045 0.0086
R7072 DVDD.n20043 DVDD.n20042 0.0086
R7073 DVDD.n20036 DVDD.n20035 0.0086
R7074 DVDD.n20033 DVDD.n20032 0.0086
R7075 DVDD.n20027 DVDD.n20026 0.0086
R7076 DVDD.n20024 DVDD.n20023 0.0086
R7077 DVDD.n19022 DVDD.n19021 0.0086
R7078 DVDD.n19025 DVDD.n19024 0.0086
R7079 DVDD.n19031 DVDD.n19030 0.0086
R7080 DVDD.n19034 DVDD.n19033 0.0086
R7081 DVDD.n19041 DVDD.n19040 0.0086
R7082 DVDD.n19044 DVDD.n19043 0.0086
R7083 DVDD.n4649 DVDD.n4648 0.0086
R7084 DVDD.n4643 DVDD.n4642 0.0086
R7085 DVDD.n4640 DVDD.n4639 0.0086
R7086 DVDD.n4831 DVDD.n4830 0.0086
R7087 DVDD.n4834 DVDD.n4833 0.0086
R7088 DVDD.n4898 DVDD.n4897 0.0086
R7089 DVDD.n4895 DVDD.n4894 0.0086
R7090 DVDD.n4892 DVDD.n4891 0.0086
R7091 DVDD.n4885 DVDD.n4884 0.0086
R7092 DVDD.n4882 DVDD.n4881 0.0086
R7093 DVDD.n4876 DVDD.n4875 0.0086
R7094 DVDD.n4873 DVDD.n4872 0.0086
R7095 DVDD.n4870 DVDD.n4869 0.0086
R7096 DVDD.n4867 DVDD.n4866 0.0086
R7097 DVDD.n4864 DVDD.n4863 0.0086
R7098 DVDD.n4861 DVDD.n4860 0.0086
R7099 DVDD.n4855 DVDD.n4854 0.0086
R7100 DVDD.n4846 DVDD.n4845 0.0086
R7101 DVDD.n4843 DVDD.n4842 0.0086
R7102 DVDD.n5136 DVDD.n5135 0.0086
R7103 DVDD.n5139 DVDD.n5138 0.0086
R7104 DVDD.n5162 DVDD.n5141 0.0086
R7105 DVDD.n5158 DVDD.n5157 0.0086
R7106 DVDD.n5155 DVDD.n5154 0.0086
R7107 DVDD.n5148 DVDD.n5147 0.0086
R7108 DVDD.n19680 DVDD.n19679 0.0086
R7109 DVDD.n19674 DVDD.n19673 0.0086
R7110 DVDD.n19671 DVDD.n19670 0.0086
R7111 DVDD.n19664 DVDD.n19663 0.0086
R7112 DVDD.n19661 DVDD.n19660 0.0086
R7113 DVDD.n19654 DVDD.n19653 0.0086
R7114 DVDD.n5306 DVDD.n5305 0.0086
R7115 DVDD.n5303 DVDD.n5302 0.0086
R7116 DVDD.n5300 DVDD.n5299 0.0086
R7117 DVDD.n5297 DVDD.n5296 0.0086
R7118 DVDD.n5291 DVDD.n5290 0.0086
R7119 DVDD.n5288 DVDD.n5287 0.0086
R7120 DVDD.n5279 DVDD.n5278 0.0086
R7121 DVDD.n5276 DVDD.n5275 0.0086
R7122 DVDD.n5270 DVDD.n5269 0.0086
R7123 DVDD.n5267 DVDD.n5266 0.0086
R7124 DVDD.n5264 DVDD.n5263 0.0086
R7125 DVDD.n5261 DVDD.n5260 0.0086
R7126 DVDD.n5258 DVDD.n5257 0.0086
R7127 DVDD.n5255 DVDD.n5254 0.0086
R7128 DVDD.n5249 DVDD.n5248 0.0086
R7129 DVDD.n5246 DVDD.n5245 0.0086
R7130 DVDD.n5239 DVDD.n5238 0.0086
R7131 DVDD.n996 DVDD.n995 0.0086
R7132 DVDD.n990 DVDD.n989 0.0086
R7133 DVDD.n987 DVDD.n986 0.0086
R7134 DVDD.n980 DVDD.n979 0.0086
R7135 DVDD.n977 DVDD.n976 0.0086
R7136 DVDD.n974 DVDD.n973 0.0086
R7137 DVDD.n968 DVDD.n967 0.0086
R7138 DVDD.n954 DVDD.n953 0.0086
R7139 DVDD.n951 DVDD.n950 0.0086
R7140 DVDD.n944 DVDD.n943 0.0086
R7141 DVDD.n941 DVDD.n940 0.0086
R7142 DVDD.n935 DVDD.n934 0.0086
R7143 DVDD.n932 DVDD.n931 0.0086
R7144 DVDD.n19231 DVDD.n19230 0.0086
R7145 DVDD.n19234 DVDD.n19233 0.0086
R7146 DVDD.n19240 DVDD.n19239 0.0086
R7147 DVDD.n19243 DVDD.n19242 0.0086
R7148 DVDD.n19250 DVDD.n19249 0.0086
R7149 DVDD.n19253 DVDD.n19252 0.0086
R7150 DVDD.n18328 DVDD.n18327 0.0086
R7151 DVDD.n18325 DVDD.n18324 0.0086
R7152 DVDD.n18319 DVDD.n18318 0.0086
R7153 DVDD.n18316 DVDD.n18315 0.0086
R7154 DVDD.n11350 DVDD.n11349 0.0086
R7155 DVDD.n11353 DVDD.n11352 0.0086
R7156 DVDD.n11855 DVDD.n11854 0.0086
R7157 DVDD.n11858 DVDD.n11857 0.0086
R7158 DVDD.n11861 DVDD.n11860 0.0086
R7159 DVDD.n11868 DVDD.n11867 0.0086
R7160 DVDD.n11871 DVDD.n11870 0.0086
R7161 DVDD.n11877 DVDD.n11876 0.0086
R7162 DVDD.n11880 DVDD.n11879 0.0086
R7163 DVDD.n11883 DVDD.n11882 0.0086
R7164 DVDD.n11886 DVDD.n11885 0.0086
R7165 DVDD.n11889 DVDD.n11888 0.0086
R7166 DVDD.n11892 DVDD.n11891 0.0086
R7167 DVDD.n11898 DVDD.n11897 0.0086
R7168 DVDD.n11907 DVDD.n11906 0.0086
R7169 DVDD.n11910 DVDD.n11909 0.0086
R7170 DVDD.n1325 DVDD.n1324 0.0086
R7171 DVDD.n1319 DVDD.n1318 0.0086
R7172 DVDD.n1316 DVDD.n1315 0.0086
R7173 DVDD.n1309 DVDD.n1308 0.0086
R7174 DVDD.n1306 DVDD.n1305 0.0086
R7175 DVDD.n1299 DVDD.n1298 0.0086
R7176 DVDD.n11312 DVDD.n11311 0.0086
R7177 DVDD.n11309 DVDD.n11308 0.0086
R7178 DVDD.n12343 DVDD.n11305 0.0086
R7179 DVDD.n12339 DVDD.n12338 0.0086
R7180 DVDD.n12336 DVDD.n12335 0.0086
R7181 DVDD.n12329 DVDD.n12328 0.0086
R7182 DVDD.n13152 DVDD.n13151 0.0086
R7183 DVDD.n13155 DVDD.n13154 0.0086
R7184 DVDD.n13158 DVDD.n13157 0.0086
R7185 DVDD.n13161 DVDD.n13160 0.0086
R7186 DVDD.n13167 DVDD.n13166 0.0086
R7187 DVDD.n13170 DVDD.n13169 0.0086
R7188 DVDD.n13179 DVDD.n13178 0.0086
R7189 DVDD.n13182 DVDD.n13181 0.0086
R7190 DVDD.n13188 DVDD.n13187 0.0086
R7191 DVDD.n13191 DVDD.n13190 0.0086
R7192 DVDD.n13194 DVDD.n13193 0.0086
R7193 DVDD.n13197 DVDD.n13196 0.0086
R7194 DVDD.n13200 DVDD.n13199 0.0086
R7195 DVDD.n13203 DVDD.n13202 0.0086
R7196 DVDD.n13209 DVDD.n13208 0.0086
R7197 DVDD.n13212 DVDD.n13211 0.0086
R7198 DVDD.n13219 DVDD.n13218 0.0086
R7199 DVDD.n3401 DVDD.n3400 0.0086
R7200 DVDD.n3598 DVDD.n3597 0.0086
R7201 DVDD.n14761 DVDD.n14760 0.0086
R7202 DVDD.n3278 DVDD.n3277 0.0086
R7203 DVDD.n3284 DVDD.n3283 0.0086
R7204 DVDD.n3287 DVDD.n3286 0.0086
R7205 DVDD.n3294 DVDD.n3293 0.0086
R7206 DVDD.n3297 DVDD.n3296 0.0086
R7207 DVDD.n3304 DVDD.n3303 0.0086
R7208 DVDD.n9424 DVDD.n9423 0.00859623
R7209 DVDD.n3714 DVDD.n3682 0.00851
R7210 DVDD.n3714 DVDD.n3713 0.00851
R7211 DVDD.n18782 DVDD.n18559 0.00851
R7212 DVDD.n18782 DVDD.n18781 0.00851
R7213 DVDD.n2944 DVDD.n2943 0.00851
R7214 DVDD.n2182 DVDD.n2181 0.00851
R7215 DVDD.n2270 DVDD.n2238 0.00851
R7216 DVDD.n2270 DVDD.n2269 0.00851
R7217 DVDD.n18935 DVDD.n18928 0.00851
R7218 DVDD.n18935 DVDD.n18934 0.00851
R7219 DVDD.n1880 DVDD.n1879 0.00851
R7220 DVDD.n1879 DVDD.n1878 0.00851
R7221 DVDD.n19961 DVDD.n19960 0.00851
R7222 DVDD.n20049 DVDD.n20017 0.00851
R7223 DVDD.n20049 DVDD.n20048 0.00851
R7224 DVDD.n19053 DVDD.n19046 0.00851
R7225 DVDD.n19053 DVDD.n19052 0.00851
R7226 DVDD.n19658 DVDD.n19657 0.00851
R7227 DVDD.n19657 DVDD.n19656 0.00851
R7228 DVDD.n984 DVDD.n983 0.00851
R7229 DVDD.n1724 DVDD.n1723 0.00851
R7230 DVDD.n1723 DVDD.n956 0.00851
R7231 DVDD.n19435 DVDD.n19255 0.00851
R7232 DVDD.n19435 DVDD.n19434 0.00851
R7233 DVDD.n1303 DVDD.n1302 0.00851
R7234 DVDD.n1302 DVDD.n1301 0.00851
R7235 DVDD.n3300 DVDD.n3299 0.00851
R7236 DVDD.n3301 DVDD.n3300 0.00851
R7237 DVDD DVDD.n15339 0.00850632
R7238 DVDD.n15914 DVDD 0.00850632
R7239 DVDD.n20309 DVDD.n20308 0.0084942
R7240 DVDD.n14906 DVDD.n14905 0.0084875
R7241 DVDD.n14907 DVDD.n14906 0.0084875
R7242 DVDD.n14908 DVDD.n14907 0.0084875
R7243 DVDD.n14909 DVDD.n14908 0.0084875
R7244 DVDD.n14910 DVDD.n14909 0.0084875
R7245 DVDD.n14911 DVDD.n14910 0.0084875
R7246 DVDD.n14934 DVDD.n14933 0.0084875
R7247 DVDD.n14933 DVDD.n14932 0.0084875
R7248 DVDD.n14932 DVDD.n14931 0.0084875
R7249 DVDD.n14834 DVDD.n14833 0.0084875
R7250 DVDD.n14835 DVDD.n14834 0.0084875
R7251 DVDD.n14836 DVDD.n14835 0.0084875
R7252 DVDD.n14837 DVDD.n14836 0.0084875
R7253 DVDD.n14838 DVDD.n14837 0.0084875
R7254 DVDD.n14896 DVDD.n14895 0.0084875
R7255 DVDD.n14897 DVDD.n14896 0.0084875
R7256 DVDD.n14898 DVDD.n14897 0.0084875
R7257 DVDD.n14899 DVDD.n14898 0.0084875
R7258 DVDD.n14900 DVDD.n14899 0.0084875
R7259 DVDD.n14901 DVDD.n14900 0.0084875
R7260 DVDD.n14902 DVDD.n14901 0.0084875
R7261 DVDD.n14903 DVDD.n14902 0.0084875
R7262 DVDD.n15229 DVDD.n15228 0.0084875
R7263 DVDD.n15230 DVDD.n15229 0.0084875
R7264 DVDD.n15231 DVDD.n15230 0.0084875
R7265 DVDD.n15232 DVDD.n15231 0.0084875
R7266 DVDD.n15112 DVDD.n15111 0.0084875
R7267 DVDD.n15113 DVDD.n15112 0.0084875
R7268 DVDD.n15114 DVDD.n15113 0.0084875
R7269 DVDD.n15115 DVDD.n15114 0.0084875
R7270 DVDD.n15116 DVDD.n15115 0.0084875
R7271 DVDD.n15117 DVDD.n15116 0.0084875
R7272 DVDD.n15118 DVDD.n15117 0.0084875
R7273 DVDD.n15119 DVDD.n15118 0.0084875
R7274 DVDD.n15301 DVDD.n15300 0.0084875
R7275 DVDD.n15300 DVDD.n15299 0.0084875
R7276 DVDD.n15299 DVDD.n15298 0.0084875
R7277 DVDD.n15298 DVDD.n15297 0.0084875
R7278 DVDD.n14992 DVDD.n14991 0.0084875
R7279 DVDD.n14993 DVDD.n14992 0.0084875
R7280 DVDD.n14994 DVDD.n14993 0.0084875
R7281 DVDD.n14995 DVDD.n14994 0.0084875
R7282 DVDD.n14996 DVDD.n14995 0.0084875
R7283 DVDD.n14997 DVDD.n14996 0.0084875
R7284 DVDD.n15011 DVDD.n15010 0.0084875
R7285 DVDD.n15010 DVDD.n15009 0.0084875
R7286 DVDD.n15009 DVDD.n15008 0.0084875
R7287 DVDD.n15099 DVDD.n15098 0.0084875
R7288 DVDD.n15100 DVDD.n15099 0.0084875
R7289 DVDD.n15101 DVDD.n15100 0.0084875
R7290 DVDD.n15102 DVDD.n15101 0.0084875
R7291 DVDD.n15103 DVDD.n15102 0.0084875
R7292 DVDD.n10691 DVDD.n10690 0.0084875
R7293 DVDD.n10690 DVDD.n10689 0.0084875
R7294 DVDD.n10689 DVDD.n10688 0.0084875
R7295 DVDD.n10688 DVDD.n10687 0.0084875
R7296 DVDD.n10687 DVDD.n10686 0.0084875
R7297 DVDD.n10686 DVDD.n10685 0.0084875
R7298 DVDD.n10464 DVDD.n10463 0.0084875
R7299 DVDD.n10465 DVDD.n10464 0.0084875
R7300 DVDD.n10466 DVDD.n10465 0.0084875
R7301 DVDD.n10476 DVDD.n10475 0.0084875
R7302 DVDD.n10475 DVDD.n10474 0.0084875
R7303 DVDD.n10474 DVDD.n10473 0.0084875
R7304 DVDD.n10473 DVDD.n10472 0.0084875
R7305 DVDD.n10472 DVDD.n10471 0.0084875
R7306 DVDD.n10471 DVDD.n10470 0.0084875
R7307 DVDD.n10673 DVDD.n10672 0.0084875
R7308 DVDD.n10674 DVDD.n10673 0.0084875
R7309 DVDD.n10675 DVDD.n10674 0.0084875
R7310 DVDD.n10676 DVDD.n10675 0.0084875
R7311 DVDD.n10677 DVDD.n10676 0.0084875
R7312 DVDD.n10729 DVDD.n10728 0.0084875
R7313 DVDD.n10728 DVDD.n10727 0.0084875
R7314 DVDD.n10727 DVDD.n10726 0.0084875
R7315 DVDD.n10726 DVDD.n10725 0.0084875
R7316 DVDD.n10725 DVDD.n10724 0.0084875
R7317 DVDD.n10724 DVDD.n10723 0.0084875
R7318 DVDD.n10723 DVDD.n10722 0.0084875
R7319 DVDD.n10722 DVDD.n10721 0.0084875
R7320 DVDD.n10632 DVDD.n10631 0.0084875
R7321 DVDD.n10631 DVDD.n10630 0.0084875
R7322 DVDD.n10630 DVDD.n10629 0.0084875
R7323 DVDD.n10629 DVDD.n10628 0.0084875
R7324 DVDD.n10628 DVDD.n10627 0.0084875
R7325 DVDD.n10627 DVDD.n10626 0.0084875
R7326 DVDD.n10384 DVDD.n10383 0.0084875
R7327 DVDD.n10385 DVDD.n10384 0.0084875
R7328 DVDD.n10386 DVDD.n10385 0.0084875
R7329 DVDD.n10393 DVDD.n10392 0.0084875
R7330 DVDD.n10392 DVDD.n10391 0.0084875
R7331 DVDD.n10391 DVDD.n10390 0.0084875
R7332 DVDD.n10390 DVDD.n10389 0.0084875
R7333 DVDD.n10389 DVDD.n10388 0.0084875
R7334 DVDD.n10578 DVDD.n10577 0.0084875
R7335 DVDD.n10579 DVDD.n10578 0.0084875
R7336 DVDD.n10580 DVDD.n10579 0.0084875
R7337 DVDD.n10581 DVDD.n10580 0.0084875
R7338 DVDD.n10652 DVDD.n10651 0.0084875
R7339 DVDD.n10651 DVDD.n10650 0.0084875
R7340 DVDD.n10650 DVDD.n10649 0.0084875
R7341 DVDD.n10649 DVDD.n10648 0.0084875
R7342 DVDD.n10648 DVDD.n10647 0.0084875
R7343 DVDD.n10647 DVDD.n10646 0.0084875
R7344 DVDD.n10646 DVDD.n10645 0.0084875
R7345 DVDD.n10645 DVDD.n10644 0.0084875
R7346 DVDD.n12248 DVDD.n12247 0.00847244
R7347 DVDD.n13338 DVDD.n13337 0.00847244
R7348 DVDD.n14431 DVDD.n14430 0.00847244
R7349 DVDD.n5989 DVDD.n5988 0.00847244
R7350 DVDD.n12652 DVDD.n12651 0.00847244
R7351 DVDD.n17805 DVDD.n17804 0.00847244
R7352 DVDD.n4452 DVDD.n4451 0.00847244
R7353 DVDD.n8726 DVDD.n8725 0.00847244
R7354 DVDD.n4154 DVDD.n4153 0.00847143
R7355 DVDD.n8536 DVDD.n8535 0.00847143
R7356 DVDD.n13868 DVDD.n13867 0.00847143
R7357 DVDD.n2347 DVDD.n2346 0.00847143
R7358 DVDD.n2402 DVDD.n2401 0.00847143
R7359 DVDD.n2545 DVDD.n2544 0.00847143
R7360 DVDD.n2598 DVDD.n2597 0.00847143
R7361 DVDD.n3404 DVDD.n3403 0.00847022
R7362 DVDD.n7737 DVDD.n7155 0.00842
R7363 DVDD.n9753 DVDD.n7830 0.00842
R7364 DVDD.n9764 DVDD.n9763 0.00842
R7365 DVDD.n9262 DVDD.n9261 0.00842
R7366 DVDD.n9265 DVDD.n9264 0.00842
R7367 DVDD.n9304 DVDD.n9303 0.00842
R7368 DVDD.n7105 DVDD.n7102 0.00842
R7369 DVDD.n6861 DVDD.n6799 0.00842
R7370 DVDD.n6851 DVDD.n6850 0.00842
R7371 DVDD.n3980 DVDD.n3979 0.00842
R7372 DVDD.n3977 DVDD.n3976 0.00842
R7373 DVDD.n3938 DVDD.n3937 0.00842
R7374 DVDD.n3884 DVDD.n3881 0.00842
R7375 DVDD.n4898 DVDD.n4836 0.00842
R7376 DVDD.n4888 DVDD.n4887 0.00842
R7377 DVDD.n5285 DVDD.n5284 0.00842
R7378 DVDD.n5282 DVDD.n5281 0.00842
R7379 DVDD.n5243 DVDD.n5242 0.00842
R7380 DVDD.n18330 DVDD.n10124 0.00842
R7381 DVDD.n11854 DVDD.n11355 0.00842
R7382 DVDD.n11865 DVDD.n11864 0.00842
R7383 DVDD.n13173 DVDD.n13172 0.00842
R7384 DVDD.n13176 DVDD.n13175 0.00842
R7385 DVDD.n13215 DVDD.n13214 0.00842
R7386 DVDD.n9452 DVDD.n9451 0.00840795
R7387 DVDD.n7712 DVDD.n7711 0.00833
R7388 DVDD.n3704 DVDD.n3703 0.00833
R7389 DVDD.n18550 DVDD.n18549 0.00833
R7390 DVDD.n18772 DVDD.n18771 0.00833
R7391 DVDD.n2260 DVDD.n2259 0.00833
R7392 DVDD.n18919 DVDD.n18918 0.00833
R7393 DVDD.n7057 DVDD.n7056 0.00833
R7394 DVDD.n1890 DVDD.n1889 0.00833
R7395 DVDD.n20039 DVDD.n20038 0.00833
R7396 DVDD.n19037 DVDD.n19036 0.00833
R7397 DVDD.n4637 DVDD.n4636 0.00833
R7398 DVDD.n19668 DVDD.n19667 0.00833
R7399 DVDD.n947 DVDD.n946 0.00833
R7400 DVDD.n19246 DVDD.n19245 0.00833
R7401 DVDD.n19425 DVDD.n19424 0.00833
R7402 DVDD.n18313 DVDD.n18312 0.00833
R7403 DVDD.n1313 DVDD.n1312 0.00833
R7404 DVDD.n3290 DVDD.n3289 0.00833
R7405 DVDD.n12935 DVDD.n12932 0.00832609
R7406 DVDD.n12954 DVDD.n12951 0.00832609
R7407 DVDD.n5519 DVDD.n5516 0.00832609
R7408 DVDD.n5526 DVDD.n5525 0.00832609
R7409 DVDD.n4017 DVDD.n4014 0.00832609
R7410 DVDD.n4024 DVDD.n4023 0.00832609
R7411 DVDD.n8973 DVDD.n8970 0.00832609
R7412 DVDD.n8980 DVDD.n8979 0.00832609
R7413 DVDD.n12900 DVDD.n12899 0.00832609
R7414 DVDD.n12895 DVDD.n12892 0.00832609
R7415 DVDD.n5720 DVDD.n5719 0.00832609
R7416 DVDD.n6065 DVDD.n6062 0.00832609
R7417 DVDD.n4091 DVDD.n4090 0.00832609
R7418 DVDD.n4515 DVDD.n4512 0.00832609
R7419 DVDD.n9000 DVDD.n8997 0.00832609
R7420 DVDD.n9007 DVDD.n9006 0.00832609
R7421 DVDD.n19464 DVDD.n18990 0.00832155
R7422 DVDD.n7301 DVDD.n7214 0.00832155
R7423 DVDD.n18333 DVDD.n3832 0.00832155
R7424 DVDD.n7662 DVDD.n7603 0.00832155
R7425 DVDD.n20215 DVDD.n117 0.00832155
R7426 DVDD.n20338 DVDD.n20312 0.00832155
R7427 DVDD.n10558 DVDD.n10557 0.00832155
R7428 DVDD.n10665 DVDD.n10664 0.00832155
R7429 DVDD.n15308 DVDD.n15307 0.00831875
R7430 DVDD.n15294 DVDD.n15293 0.00831875
R7431 DVDD.n15001 DVDD.n15000 0.00831875
R7432 DVDD.n12579 DVDD.n12578 0.00829908
R7433 DVDD.n4349 DVDD.n4348 0.00829908
R7434 DVDD.n8623 DVDD.n8622 0.00829908
R7435 DVDD.n12238 DVDD.n12237 0.00829528
R7436 DVDD.n19888 DVDD.n19887 0.00829528
R7437 DVDD.n5021 DVDD.n5020 0.00829528
R7438 DVDD.n1489 DVDD.n1488 0.00829528
R7439 DVDD.n11733 DVDD.n11732 0.00829528
R7440 DVDD.n2109 DVDD.n2108 0.00829528
R7441 DVDD.n6663 DVDD.n6662 0.00829528
R7442 DVDD.n3508 DVDD.n3507 0.00829528
R7443 DVDD.n9631 DVDD.n9630 0.00829528
R7444 DVDD.n10477 DVDD.n10476 0.0082625
R7445 DVDD.n10672 DVDD.n10671 0.0082625
R7446 DVDD.n10684 DVDD.n10683 0.0082625
R7447 DVDD.n5877 DVDD.n5876 0.00825207
R7448 DVDD.n5863 DVDD.n5862 0.00825207
R7449 DVDD.n5857 DVDD.n5856 0.00825207
R7450 DVDD.n5846 DVDD.n5845 0.00825207
R7451 DVDD.n5840 DVDD.n5839 0.00825207
R7452 DVDD.n5829 DVDD.n5828 0.00825207
R7453 DVDD.n5823 DVDD.n5822 0.00825207
R7454 DVDD.n5809 DVDD.n5808 0.00825207
R7455 DVDD.n12572 DVDD.n12571 0.00825207
R7456 DVDD.n12561 DVDD.n12560 0.00825207
R7457 DVDD.n12555 DVDD.n12554 0.00825207
R7458 DVDD.n12544 DVDD.n12543 0.00825207
R7459 DVDD.n12538 DVDD.n12537 0.00825207
R7460 DVDD.n12527 DVDD.n12526 0.00825207
R7461 DVDD.n12521 DVDD.n12520 0.00825207
R7462 DVDD.n12510 DVDD.n12509 0.00825207
R7463 DVDD.n5810 DVDD.n5809 0.00825207
R7464 DVDD.n12511 DVDD.n12510 0.00825207
R7465 DVDD.n12545 DVDD.n12544 0.00825207
R7466 DVDD.n5847 DVDD.n5846 0.00825207
R7467 DVDD.n12539 DVDD.n12538 0.00825207
R7468 DVDD.n5841 DVDD.n5840 0.00825207
R7469 DVDD.n12528 DVDD.n12527 0.00825207
R7470 DVDD.n5830 DVDD.n5829 0.00825207
R7471 DVDD.n12522 DVDD.n12521 0.00825207
R7472 DVDD.n5824 DVDD.n5823 0.00825207
R7473 DVDD.n12556 DVDD.n12555 0.00825207
R7474 DVDD.n5858 DVDD.n5857 0.00825207
R7475 DVDD.n5864 DVDD.n5863 0.00825207
R7476 DVDD.n12562 DVDD.n12561 0.00825207
R7477 DVDD.n5876 DVDD.n5873 0.00825207
R7478 DVDD.n12573 DVDD.n12572 0.00825207
R7479 DVDD.n4332 DVDD.n4331 0.00825207
R7480 DVDD.n4321 DVDD.n4320 0.00825207
R7481 DVDD.n4303 DVDD.n4302 0.00825207
R7482 DVDD.n4292 DVDD.n4291 0.00825207
R7483 DVDD.n4278 DVDD.n4277 0.00825207
R7484 DVDD.n4267 DVDD.n4266 0.00825207
R7485 DVDD.n4253 DVDD.n4252 0.00825207
R7486 DVDD.n4238 DVDD.n4237 0.00825207
R7487 DVDD.n4304 DVDD.n4303 0.00825207
R7488 DVDD.n4293 DVDD.n4292 0.00825207
R7489 DVDD.n4279 DVDD.n4278 0.00825207
R7490 DVDD.n4268 DVDD.n4267 0.00825207
R7491 DVDD.n4254 DVDD.n4253 0.00825207
R7492 DVDD.n4333 DVDD.n4332 0.00825207
R7493 DVDD.n4322 DVDD.n4321 0.00825207
R7494 DVDD.n4239 DVDD.n4238 0.00825207
R7495 DVDD.n8617 DVDD.n8616 0.00825207
R7496 DVDD.n8605 DVDD.n8604 0.00825207
R7497 DVDD.n8600 DVDD.n8599 0.00825207
R7498 DVDD.n8588 DVDD.n8587 0.00825207
R7499 DVDD.n8583 DVDD.n8582 0.00825207
R7500 DVDD.n8571 DVDD.n8570 0.00825207
R7501 DVDD.n8566 DVDD.n8565 0.00825207
R7502 DVDD.n8554 DVDD.n8553 0.00825207
R7503 DVDD.n8599 DVDD.n8598 0.00825207
R7504 DVDD.n8589 DVDD.n8588 0.00825207
R7505 DVDD.n8582 DVDD.n8581 0.00825207
R7506 DVDD.n8572 DVDD.n8571 0.00825207
R7507 DVDD.n8565 DVDD.n8564 0.00825207
R7508 DVDD.n8606 DVDD.n8605 0.00825207
R7509 DVDD.n8616 DVDD.n8615 0.00825207
R7510 DVDD.n8555 DVDD.n8554 0.00825207
R7511 DVDD.n7821 DVDD.n7820 0.00824
R7512 DVDD.n7822 DVDD.n7821 0.00824
R7513 DVDD.n9529 DVDD.n9528 0.00824
R7514 DVDD.n9528 DVDD.n9527 0.00824
R7515 DVDD.n6790 DVDD.n6789 0.00824
R7516 DVDD.n6791 DVDD.n6790 0.00824
R7517 DVDD.n6561 DVDD.n6560 0.00824
R7518 DVDD.n6560 DVDD.n6559 0.00824
R7519 DVDD.n4827 DVDD.n4826 0.00824
R7520 DVDD.n4828 DVDD.n4827 0.00824
R7521 DVDD.n5152 DVDD.n5151 0.00824
R7522 DVDD.n5151 DVDD.n5150 0.00824
R7523 DVDD.n11346 DVDD.n11345 0.00824
R7524 DVDD.n11347 DVDD.n11346 0.00824
R7525 DVDD.n12333 DVDD.n12332 0.00824
R7526 DVDD.n12332 DVDD.n12331 0.00824
R7527 DVDD.n15988 DVDD.n15987 0.0082373
R7528 DVDD.n15961 DVDD.n15960 0.0082373
R7529 DVDD.n15960 DVDD.n15959 0.0082373
R7530 DVDD.n15989 DVDD.n15988 0.0082373
R7531 DVDD.n16053 DVDD.n16052 0.0082373
R7532 DVDD.n16024 DVDD.n16023 0.0082373
R7533 DVDD.n15997 DVDD.n15996 0.0082373
R7534 DVDD.n16054 DVDD.n16053 0.0082373
R7535 DVDD.n16023 DVDD.n16022 0.0082373
R7536 DVDD.n15998 DVDD.n15997 0.0082373
R7537 DVDD.n15665 DVDD.n15664 0.0082373
R7538 DVDD.n15636 DVDD.n15635 0.0082373
R7539 DVDD.n15935 DVDD.n15934 0.0082373
R7540 DVDD.n15934 DVDD.n15933 0.0082373
R7541 DVDD.n15666 DVDD.n15665 0.0082373
R7542 DVDD.n15635 DVDD.n15634 0.0082373
R7543 DVDD.n8168 DVDD.n8167 0.0082373
R7544 DVDD.n8169 DVDD.n8168 0.0082373
R7545 DVDD.n7206 DVDD.n7205 0.00823251
R7546 DVDD.n7211 DVDD.n7210 0.00823251
R7547 DVDD.n7600 DVDD.n7599 0.00823251
R7548 DVDD.n7605 DVDD.n7604 0.00823251
R7549 DVDD.n20304 DVDD.n20303 0.00823251
R7550 DVDD.n10661 DVDD.n10660 0.00823251
R7551 DVDD.n9419 DVDD.n9418 0.00821966
R7552 DVDD.n13913 DVDD.n13912 0.0082027
R7553 DVDD.n13917 DVDD.n13916 0.0082027
R7554 DVDD.n14302 DVDD.n14301 0.0082027
R7555 DVDD.n14306 DVDD.n14305 0.0082027
R7556 DVDD.n3705 DVDD.n3704 0.00815
R7557 DVDD.n18551 DVDD.n18550 0.00815
R7558 DVDD.n7931 DVDD.n7930 0.00815
R7559 DVDD.n2261 DVDD.n2260 0.00815
R7560 DVDD.n18920 DVDD.n18919 0.00815
R7561 DVDD.n6524 DVDD.n6523 0.00815
R7562 DVDD.n1889 DVDD.n1888 0.00815
R7563 DVDD.n20040 DVDD.n20039 0.00815
R7564 DVDD.n19038 DVDD.n19037 0.00815
R7565 DVDD.n5115 DVDD.n5114 0.00815
R7566 DVDD.n19667 DVDD.n19666 0.00815
R7567 DVDD.n948 DVDD.n947 0.00815
R7568 DVDD.n19247 DVDD.n19246 0.00815
R7569 DVDD.n1312 DVDD.n1311 0.00815
R7570 DVDD.n11333 DVDD.n11332 0.00815
R7571 DVDD.n3600 DVDD.n3599 0.00815
R7572 DVDD.n18390 DVDD.n18389 0.00815
R7573 DVDD.n14763 DVDD.n14762 0.00815
R7574 DVDD.n3291 DVDD.n3290 0.00815
R7575 DVDD.n12229 DVDD.n12228 0.00811811
R7576 DVDD.n5363 DVDD.n5362 0.00811811
R7577 DVDD.n13097 DVDD.n13096 0.00811811
R7578 DVDD.n6398 DVDD.n6397 0.00811811
R7579 DVDD.n9184 DVDD.n9183 0.00811811
R7580 DVDD.n9763 DVDD.n9762 0.00806
R7581 DVDD.n7913 DVDD.n7912 0.00806
R7582 DVDD.n9489 DVDD.n9488 0.00806
R7583 DVDD.n9305 DVDD.n9304 0.00806
R7584 DVDD.n6852 DVDD.n6851 0.00806
R7585 DVDD.n6542 DVDD.n6541 0.00806
R7586 DVDD.n3937 DVDD.n3936 0.00806
R7587 DVDD.n4889 DVDD.n4888 0.00806
R7588 DVDD.n5133 DVDD.n5132 0.00806
R7589 DVDD.n5242 DVDD.n5241 0.00806
R7590 DVDD.n11864 DVDD.n11863 0.00806
R7591 DVDD.n11315 DVDD.n11314 0.00806
R7592 DVDD.n12294 DVDD.n12293 0.00806
R7593 DVDD.n13216 DVDD.n13215 0.00806
R7594 DVDD.n7475 DVDD.n7346 0.008
R7595 DVDD.n7674 DVDD.n7557 0.008
R7596 DVDD.n7674 DVDD.n7669 0.008
R7597 DVDD.n7475 DVDD.n7434 0.008
R7598 DVDD.n20341 DVDD.n32 0.008
R7599 DVDD.n15147 DVDD.n15146 0.008
R7600 DVDD.n10218 DVDD.n10217 0.008
R7601 DVDD.n20341 DVDD.n20220 0.008
R7602 DVDD.n2945 DVDD.n2944 0.00797
R7603 DVDD.n9803 DVDD.n9802 0.00797
R7604 DVDD.n9883 DVDD.n9882 0.00797
R7605 DVDD.n2183 DVDD.n2182 0.00797
R7606 DVDD.n6812 DVDD.n6811 0.00797
R7607 DVDD.n19962 DVDD.n19961 0.00797
R7608 DVDD.n4849 DVDD.n4848 0.00797
R7609 DVDD.n983 DVDD.n982 0.00797
R7610 DVDD.n11904 DVDD.n11903 0.00797
R7611 DVDD.n11984 DVDD.n11983 0.00797
R7612 DVDD.n13854 DVDD.n13853 0.00795714
R7613 DVDD.n2664 DVDD.n2663 0.00795714
R7614 DVDD.n12257 DVDD.n12256 0.00794094
R7615 DVDD.n14422 DVDD.n14421 0.00794094
R7616 DVDD.n4797 DVDD.n4796 0.00794094
R7617 DVDD.n5980 DVDD.n5979 0.00794094
R7618 DVDD.n11623 DVDD.n11622 0.00794094
R7619 DVDD.n12643 DVDD.n12642 0.00794094
R7620 DVDD.n17796 DVDD.n17795 0.00794094
R7621 DVDD.n6887 DVDD.n6886 0.00794094
R7622 DVDD.n4443 DVDD.n4442 0.00794094
R7623 DVDD.n7879 DVDD.n7878 0.00794094
R7624 DVDD.n8717 DVDD.n8716 0.00794094
R7625 DVDD.n15196 DVDD.n15195 0.00789594
R7626 DVDD.n15201 DVDD.n15200 0.00789594
R7627 DVDD.n15206 DVDD.n15205 0.00789594
R7628 DVDD.n15256 DVDD.n15255 0.00789594
R7629 DVDD.n15261 DVDD.n15260 0.00789594
R7630 DVDD.n15266 DVDD.n15265 0.00789594
R7631 DVDD.n15271 DVDD.n15270 0.00789594
R7632 DVDD.n9784 DVDD.n9783 0.00788
R7633 DVDD.n9243 DVDD.n9242 0.00788
R7634 DVDD.n9285 DVDD.n9284 0.00788
R7635 DVDD.n6831 DVDD.n6830 0.00788
R7636 DVDD.n3999 DVDD.n3998 0.00788
R7637 DVDD.n3957 DVDD.n3956 0.00788
R7638 DVDD.n4868 DVDD.n4867 0.00788
R7639 DVDD.n5304 DVDD.n5303 0.00788
R7640 DVDD.n5262 DVDD.n5261 0.00788
R7641 DVDD.n11885 DVDD.n11884 0.00788
R7642 DVDD.n13154 DVDD.n13153 0.00788
R7643 DVDD.n13196 DVDD.n13195 0.00788
R7644 DVDD.n8105 DVDD.n8104 0.0078431
R7645 DVDD.n2483 DVDD 0.00782857
R7646 DVDD DVDD.n2484 0.00782857
R7647 DVDD.n12195 DVDD.n12194 0.00781054
R7648 DVDD.n2723 DVDD.n2722 0.00781054
R7649 DVDD.n2750 DVDD.n2749 0.00781054
R7650 DVDD.n2764 DVDD.n2763 0.00781054
R7651 DVDD.n2792 DVDD.n2791 0.00781054
R7652 DVDD.n15403 DVDD.n15402 0.00781054
R7653 DVDD.n15433 DVDD.n15432 0.00781054
R7654 DVDD.n15459 DVDD.n15458 0.00781054
R7655 DVDD.n15468 DVDD.n15467 0.00781054
R7656 DVDD.n15496 DVDD.n15495 0.00781054
R7657 DVDD.n14728 DVDD.n14727 0.00781054
R7658 DVDD.n14700 DVDD.n14699 0.00781054
R7659 DVDD.n14645 DVDD.n14644 0.00781054
R7660 DVDD.n14617 DVDD.n14616 0.00781054
R7661 DVDD.n14563 DVDD.n14562 0.00781054
R7662 DVDD.n14534 DVDD.n14533 0.00781054
R7663 DVDD.n14507 DVDD.n14506 0.00781054
R7664 DVDD.n14475 DVDD.n14474 0.00781054
R7665 DVDD.n14403 DVDD.n14402 0.00781054
R7666 DVDD.n14394 DVDD.n14393 0.00781054
R7667 DVDD.n14367 DVDD.n14366 0.00781054
R7668 DVDD.n14646 DVDD.n14645 0.00781054
R7669 DVDD.n2751 DVDD.n2750 0.00781054
R7670 DVDD.n15495 DVDD.n15494 0.00781054
R7671 DVDD.n14729 DVDD.n14728 0.00781054
R7672 DVDD.n15402 DVDD.n15401 0.00781054
R7673 DVDD.n15432 DVDD.n15431 0.00781054
R7674 DVDD.n15458 DVDD.n15457 0.00781054
R7675 DVDD.n15467 DVDD.n15466 0.00781054
R7676 DVDD.n2763 DVDD.n2762 0.00781054
R7677 DVDD.n2791 DVDD.n2790 0.00781054
R7678 DVDD.n2722 DVDD.n2721 0.00781054
R7679 DVDD.n14618 DVDD.n14617 0.00781054
R7680 DVDD.n14476 DVDD.n14475 0.00781054
R7681 DVDD.n14404 DVDD.n14403 0.00781054
R7682 DVDD.n14508 DVDD.n14507 0.00781054
R7683 DVDD.n14564 DVDD.n14563 0.00781054
R7684 DVDD.n14533 DVDD.n14532 0.00781054
R7685 DVDD.n14701 DVDD.n14700 0.00781054
R7686 DVDD.n6629 DVDD.n6628 0.00781054
R7687 DVDD.n6289 DVDD.n6288 0.00781054
R7688 DVDD.n6212 DVDD.n6211 0.00781054
R7689 DVDD.n6171 DVDD.n6170 0.00781054
R7690 DVDD.n6132 DVDD.n6131 0.00781054
R7691 DVDD.n4424 DVDD.n4423 0.00781054
R7692 DVDD.n4415 DVDD.n4414 0.00781054
R7693 DVDD.n4387 DVDD.n4386 0.00781054
R7694 DVDD.n6628 DVDD.n6627 0.00781054
R7695 DVDD.n6290 DVDD.n6289 0.00781054
R7696 DVDD.n4425 DVDD.n4424 0.00781054
R7697 DVDD.n6133 DVDD.n6132 0.00781054
R7698 DVDD.n6213 DVDD.n6212 0.00781054
R7699 DVDD.n6170 DVDD.n6169 0.00781054
R7700 DVDD.n4388 DVDD.n4387 0.00781054
R7701 DVDD.n14366 DVDD.n14365 0.00781054
R7702 DVDD.n4416 DVDD.n4415 0.00781054
R7703 DVDD.n14395 DVDD.n14394 0.00781054
R7704 DVDD.n9597 DVDD.n9596 0.00781054
R7705 DVDD.n9075 DVDD.n9074 0.00781054
R7706 DVDD.n8914 DVDD.n8913 0.00781054
R7707 DVDD.n8873 DVDD.n8872 0.00781054
R7708 DVDD.n8834 DVDD.n8833 0.00781054
R7709 DVDD.n8698 DVDD.n8697 0.00781054
R7710 DVDD.n8689 DVDD.n8688 0.00781054
R7711 DVDD.n8661 DVDD.n8660 0.00781054
R7712 DVDD.n8662 DVDD.n8661 0.00781054
R7713 DVDD.n9596 DVDD.n9595 0.00781054
R7714 DVDD.n9076 DVDD.n9075 0.00781054
R7715 DVDD.n8699 DVDD.n8698 0.00781054
R7716 DVDD.n8835 DVDD.n8834 0.00781054
R7717 DVDD.n8915 DVDD.n8914 0.00781054
R7718 DVDD.n8872 DVDD.n8871 0.00781054
R7719 DVDD.n8690 DVDD.n8689 0.00781054
R7720 DVDD.n15211 DVDD.n15210 0.00779989
R7721 DVDD.n17265 DVDD.n17264 0.0077973
R7722 DVDD.n17296 DVDD.n17295 0.0077973
R7723 DVDD.n17643 DVDD.n17642 0.0077973
R7724 DVDD.n17675 DVDD.n17674 0.0077973
R7725 DVDD.n3397 DVDD.n3396 0.00779377
R7726 DVDD.n3391 DVDD.n3390 0.00779377
R7727 DVDD.n12224 DVDD.n12223 0.00776378
R7728 DVDD.n14450 DVDD.n14449 0.00776378
R7729 DVDD.n6018 DVDD.n6017 0.00776378
R7730 DVDD.n12669 DVDD.n12668 0.00776378
R7731 DVDD.n17819 DVDD.n17818 0.00776378
R7732 DVDD.n4469 DVDD.n4468 0.00776378
R7733 DVDD.n8755 DVDD.n8754 0.00776378
R7734 DVDD.n19464 DVDD.n3823 0.00770384
R7735 DVDD.n7301 DVDD.n7298 0.00770384
R7736 DVDD.n3662 DVDD.n3661 0.0077
R7737 DVDD.n18630 DVDD.n18629 0.0077
R7738 DVDD.n18561 DVDD.n18560 0.0077
R7739 DVDD.n18723 DVDD.n18722 0.0077
R7740 DVDD.n18708 DVDD.n18707 0.0077
R7741 DVDD.n18693 DVDD.n18692 0.0077
R7742 DVDD.n18666 DVDD.n18665 0.0077
R7743 DVDD.n18422 DVDD.n18421 0.0077
R7744 DVDD.n18429 DVDD.n18428 0.0077
R7745 DVDD.n18447 DVDD.n18446 0.0077
R7746 DVDD.n18440 DVDD.n18439 0.0077
R7747 DVDD.n18433 DVDD.n18432 0.0077
R7748 DVDD.n18348 DVDD.n18347 0.0077
R7749 DVDD.n18350 DVDD.n18349 0.0077
R7750 DVDD.n9416 DVDD.n9415 0.00765481
R7751 DVDD.n8104 DVDD.n8103 0.00765481
R7752 DVDD.n9457 DVDD.n9456 0.00764769
R7753 DVDD.n10483 DVDD.n10482 0.00764375
R7754 DVDD.n10678 DVDD.n10677 0.00764375
R7755 DVDD.n10721 DVDD.n10720 0.00764375
R7756 DVDD.n9388 DVDD.n9387 0.00761
R7757 DVDD.n13299 DVDD.n13298 0.00761
R7758 DVDD.n19721 DVDD.n19720 0.00758661
R7759 DVDD.n1366 DVDD.n1365 0.00758661
R7760 DVDD.n1943 DVDD.n1942 0.00758661
R7761 DVDD.n3237 DVDD.n3236 0.00758661
R7762 DVDD.n9318 DVDD.n9317 0.00752
R7763 DVDD.n13229 DVDD.n13228 0.00752
R7764 DVDD.n19464 DVDD.n18981 0.00748725
R7765 DVDD.n7301 DVDD.n7209 0.00748725
R7766 DVDD.n18333 DVDD.n3840 0.00748725
R7767 DVDD.n7662 DVDD.n7608 0.00748725
R7768 DVDD.n20215 DVDD.n125 0.00748725
R7769 DVDD.n20338 DVDD.n20307 0.00748725
R7770 DVDD.n10558 DVDD.n10548 0.00748725
R7771 DVDD.n10665 DVDD.n10659 0.00748725
R7772 DVDD.n15111 DVDD.n15110 0.007475
R7773 DVDD.n15302 DVDD.n15301 0.007475
R7774 DVDD.n15007 DVDD.n15006 0.007475
R7775 DVDD.n12164 DVDD.n12163 0.00740945
R7776 DVDD.n5543 DVDD.n5542 0.00735992
R7777 DVDD.n6253 DVDD.n6252 0.00735992
R7778 DVDD.n11264 DVDD.n11263 0.00725
R7779 DVDD.n11252 DVDD.n11251 0.00725
R7780 DVDD.n11236 DVDD.n11235 0.00725
R7781 DVDD.n302 DVDD.n301 0.00725
R7782 DVDD.n493 DVDD.n492 0.00725
R7783 DVDD.n447 DVDD.n446 0.00725
R7784 DVDD.n2340 DVDD.n2339 0.00725
R7785 DVDD.n2391 DVDD.n2390 0.00725
R7786 DVDD.n533 DVDD.n532 0.00725
R7787 DVDD.n725 DVDD.n724 0.00725
R7788 DVDD.n679 DVDD.n678 0.00725
R7789 DVDD.n2538 DVDD.n2537 0.00725
R7790 DVDD.n2589 DVDD.n2588 0.00725
R7791 DVDD.n10470 DVDD.n10469 0.00725
R7792 DVDD.n10388 DVDD.n10387 0.00725
R7793 DVDD.n3407 DVDD.n3406 0.00725
R7794 DVDD.n3656 DVDD.n3655 0.00725
R7795 DVDD.n18613 DVDD.n18612 0.00725
R7796 DVDD.n18720 DVDD.n18719 0.00725
R7797 DVDD.n18705 DVDD.n18704 0.00725
R7798 DVDD.n18664 DVDD.n18663 0.00725
R7799 DVDD.n18465 DVDD.n18464 0.00725
R7800 DVDD.n18425 DVDD.n18424 0.00725
R7801 DVDD.n18431 DVDD.n18430 0.00725
R7802 DVDD.n18437 DVDD.n18436 0.00725
R7803 DVDD.n18386 DVDD.n18385 0.00725
R7804 DVDD.n18394 DVDD.n18393 0.00725
R7805 DVDD.n12163 DVDD.n12162 0.00723228
R7806 DVDD.n12221 DVDD.n12220 0.00723228
R7807 DVDD.n4924 DVDD.n4923 0.00723228
R7808 DVDD.n5318 DVDD.n5317 0.00723228
R7809 DVDD.n5408 DVDD.n5407 0.00723228
R7810 DVDD.n5450 DVDD.n5449 0.00723228
R7811 DVDD.n11829 DVDD.n11828 0.00723228
R7812 DVDD.n13140 DVDD.n13139 0.00723228
R7813 DVDD.n13054 DVDD.n13053 0.00723228
R7814 DVDD.n13013 DVDD.n13012 0.00723228
R7815 DVDD.n6760 DVDD.n6759 0.00723228
R7816 DVDD.n6443 DVDD.n6442 0.00723228
R7817 DVDD.n6353 DVDD.n6352 0.00723228
R7818 DVDD.n6311 DVDD.n6310 0.00723228
R7819 DVDD.n9728 DVDD.n9727 0.00723228
R7820 DVDD.n9229 DVDD.n9228 0.00723228
R7821 DVDD.n9139 DVDD.n9138 0.00723228
R7822 DVDD.n9097 DVDD.n9096 0.00723228
R7823 DVDD.n7475 DVDD.n7203 0.0072
R7824 DVDD.n7674 DVDD.n7516 0.0072
R7825 DVDD.n7674 DVDD.n7673 0.0072
R7826 DVDD.n7475 DVDD.n7430 0.0072
R7827 DVDD.n20341 DVDD.n28 0.0072
R7828 DVDD.n15147 DVDD.n15139 0.0072
R7829 DVDD.n10218 DVDD.n10209 0.0072
R7830 DVDD.n20341 DVDD.n20224 0.0072
R7831 DVDD.n9438 DVDD.n9437 0.00708996
R7832 DVDD.n2 DVDD.n1 0.00708169
R7833 DVDD.n3 DVDD.n2 0.00708169
R7834 DVDD.n6 DVDD.n5 0.00708169
R7835 DVDD.n5 DVDD.n4 0.00708169
R7836 DVDD.n7348 DVDD.n7347 0.00708169
R7837 DVDD.n7349 DVDD.n7348 0.00708169
R7838 DVDD.n7352 DVDD.n7351 0.00708169
R7839 DVDD.n7351 DVDD.n7350 0.00708169
R7840 DVDD.n7562 DVDD.n7561 0.00708169
R7841 DVDD.n7563 DVDD.n7562 0.00708169
R7842 DVDD.n7560 DVDD.n7559 0.00708169
R7843 DVDD.n7559 DVDD.n7558 0.00708169
R7844 DVDD.n10189 DVDD.n10188 0.00708169
R7845 DVDD.n10190 DVDD.n10189 0.00708169
R7846 DVDD.n10193 DVDD.n10192 0.00708169
R7847 DVDD.n10192 DVDD.n10191 0.00708169
R7848 DVDD.n3431 DVDD.n3430 0.00707472
R7849 DVDD.n5224 DVDD.n5223 0.00705512
R7850 DVDD.n5627 DVDD.n5626 0.00705512
R7851 DVDD.n12404 DVDD.n12403 0.00705512
R7852 DVDD.n12810 DVDD.n12809 0.00705512
R7853 DVDD.n6458 DVDD.n6457 0.00705512
R7854 DVDD.n6189 DVDD.n6188 0.00705512
R7855 DVDD.n8425 DVDD.n8424 0.00705512
R7856 DVDD.n8891 DVDD.n8890 0.00705512
R7857 DVDD.n15297 DVDD.n15296 0.007025
R7858 DVDD.n14998 DVDD.n14997 0.007025
R7859 DVDD.n7663 DVDD.n7662 0.00693543
R7860 DVDD.n15250 DVDD.n15212 0.00693543
R7861 DVDD.n15290 DVDD.n15130 0.00693543
R7862 DVDD.n8179 DVDD.n8178 0.00690167
R7863 DVDD.n9423 DVDD.n9422 0.00690167
R7864 DVDD.n20074 DVDD.n20073 0.00687795
R7865 DVDD.n1699 DVDD.n1698 0.00687795
R7866 DVDD.n2295 DVDD.n2294 0.00687795
R7867 DVDD.n3739 DVDD.n3738 0.00687795
R7868 DVDD.n399 DVDD.n398 0.00686429
R7869 DVDD.n454 DVDD.n452 0.00686429
R7870 DVDD.n630 DVDD.n629 0.00686429
R7871 DVDD.n686 DVDD.n684 0.00686429
R7872 DVDD.n11287 DVDD.n11286 0.00686429
R7873 DVDD.n12487 DVDD.n12486 0.00686429
R7874 DVDD.n5738 DVDD.n5737 0.00686429
R7875 DVDD.n12461 DVDD.n12460 0.0068
R7876 DVDD.n12469 DVDD.n12468 0.0068
R7877 DVDD.n5703 DVDD.n5702 0.0068
R7878 DVDD.n6110 DVDD.n4555 0.0068
R7879 DVDD.n6115 DVDD.n6114 0.0068
R7880 DVDD.n4072 DVDD.n4071 0.0068
R7881 DVDD.n8486 DVDD.n8485 0.0068
R7882 DVDD.n8494 DVDD.n8493 0.0068
R7883 DVDD.n12774 DVDD.n12773 0.0068
R7884 DVDD.n12455 DVDD.n12454 0.0068
R7885 DVDD.n5661 DVDD.n5660 0.0068
R7886 DVDD.n4567 DVDD.n4566 0.0068
R7887 DVDD.n4563 DVDD.n4562 0.0068
R7888 DVDD.n4063 DVDD.n4062 0.0068
R7889 DVDD.n8467 DVDD.n8466 0.0068
R7890 DVDD.n8479 DVDD.n8478 0.0068
R7891 DVDD.n12430 DVDD.n12429 0.0068
R7892 DVDD.n12442 DVDD.n12441 0.0068
R7893 DVDD.n5615 DVDD.n5614 0.0068
R7894 DVDD.n4582 DVDD.n4581 0.0068
R7895 DVDD.n4578 DVDD.n4577 0.0068
R7896 DVDD.n4053 DVDD.n4052 0.0068
R7897 DVDD.n8449 DVDD.n8448 0.0068
R7898 DVDD.n8461 DVDD.n8460 0.0068
R7899 DVDD.n12411 DVDD.n12410 0.0068
R7900 DVDD.n12423 DVDD.n12422 0.0068
R7901 DVDD.n5568 DVDD.n5567 0.0068
R7902 DVDD.n4597 DVDD.n4596 0.0068
R7903 DVDD.n4593 DVDD.n4592 0.0068
R7904 DVDD.n4043 DVDD.n4042 0.0068
R7905 DVDD.n8431 DVDD.n8430 0.0068
R7906 DVDD.n8443 DVDD.n8442 0.0068
R7907 DVDD.n14882 DVDD.n14838 0.0068
R7908 DVDD.n15104 DVDD.n15103 0.0068
R7909 DVDD.n3427 DVDD.n3426 0.0068
R7910 DVDD.n3594 DVDD.n3593 0.0068
R7911 DVDD.n18355 DVDD.n18354 0.0068
R7912 DVDD.n8357 DVDD.n8356 0.00671339
R7913 DVDD.n12243 DVDD.n12242 0.00670079
R7914 DVDD.n19079 DVDD.n19078 0.00670079
R7915 DVDD.n5085 DVDD.n5084 0.00670079
R7916 DVDD.n19461 DVDD.n19460 0.00670079
R7917 DVDD.n11669 DVDD.n11668 0.00670079
R7918 DVDD.n18971 DVDD.n18970 0.00670079
R7919 DVDD.n6597 DVDD.n6596 0.00670079
R7920 DVDD.n18808 DVDD.n18807 0.00670079
R7921 DVDD.n9565 DVDD.n9564 0.00670079
R7922 DVDD.n9041 DVDD.n9040 0.0066935
R7923 DVDD.n17690 DVDD.n17689 0.0066935
R7924 DVDD.n14981 DVDD.n14934 0.0066875
R7925 DVDD.n15013 DVDD.n15011 0.0066875
R7926 DVDD.n13833 DVDD 0.00667143
R7927 DVDD.n2348 DVDD.n2345 0.00667143
R7928 DVDD.n2458 DVDD.n2456 0.00667143
R7929 DVDD DVDD.n2697 0.00667143
R7930 DVDD.n2546 DVDD.n2543 0.00667143
R7931 DVDD.n2656 DVDD.n2654 0.00667143
R7932 DVDD.n4147 DVDD.n4146 0.00667143
R7933 DVDD.n8530 DVDD.n8529 0.00667143
R7934 DVDD.n13862 DVDD.n13861 0.00667143
R7935 DVDD.n3378 DVDD.n3377 0.00662472
R7936 DVDD.n3810 DVDD.n3809 0.006575
R7937 DVDD.n18995 DVDD.n18994 0.006575
R7938 DVDD.n7218 DVDD.n7217 0.006575
R7939 DVDD.n7115 DVDD.n7114 0.006575
R7940 DVDD.n2817 DVDD.n2816 0.006575
R7941 DVDD.n14846 DVDD.n14845 0.006575
R7942 DVDD.n15077 DVDD.n15076 0.006575
R7943 DVDD.n10695 DVDD.n10694 0.006575
R7944 DVDD.n10598 DVDD.n10597 0.006575
R7945 DVDD.n7289 DVDD.n7288 0.006575
R7946 DVDD.n15704 DVDD 0.0065675
R7947 DVDD.n15133 DVDD.n15132 0.0065619
R7948 DVDD.n15134 DVDD.n15133 0.0065619
R7949 DVDD.n15135 DVDD.n15134 0.0065619
R7950 DVDD.n15287 DVDD.n15286 0.0065619
R7951 DVDD.n15286 DVDD.n15282 0.0065619
R7952 DVDD.n15282 DVDD.n15278 0.0065619
R7953 DVDD.n504 DVDD.n502 0.00654286
R7954 DVDD.n734 DVDD.n732 0.00654286
R7955 DVDD.n12228 DVDD.n12227 0.00652362
R7956 DVDD.n13495 DVDD.n13494 0.00652362
R7957 DVDD.n17155 DVDD.n17154 0.0065
R7958 DVDD.n16970 DVDD.n16969 0.0065
R7959 DVDD.n16816 DVDD.n16694 0.0065
R7960 DVDD.n17043 DVDD.n16816 0.0065
R7961 DVDD.n16966 DVDD.n16921 0.0065
R7962 DVDD.n17152 DVDD.n17043 0.0065
R7963 DVDD.n16312 DVDD.n15535 0.0065
R7964 DVDD.n16312 DVDD.n16118 0.0065
R7965 DVDD.n16233 DVDD.n16232 0.0065
R7966 DVDD.n16118 DVDD.n16117 0.0065
R7967 DVDD.n17154 DVDD.n17153 0.0065
R7968 DVDD.n11112 DVDD.n11111 0.0065
R7969 DVDD.n11121 DVDD.n11120 0.0065
R7970 DVDD.n11120 DVDD.n11112 0.0065
R7971 DVDD.n17156 DVDD.n17155 0.0065
R7972 DVDD.n15108 DVDD.n15107 0.00640625
R7973 DVDD.n15305 DVDD.n15304 0.00640625
R7974 DVDD.n15004 DVDD.n15003 0.00640625
R7975 DVDD.n10480 DVDD.n10479 0.00640625
R7976 DVDD.n10669 DVDD.n10668 0.00640625
R7977 DVDD.n10681 DVDD.n10680 0.00640625
R7978 DVDD.n10718 DVDD.n10717 0.00640625
R7979 DVDD.n14322 DVDD.n14321 0.00636121
R7980 DVDD.n12960 DVDD.n12959 0.00636121
R7981 DVDD.n3807 DVDD.n3806 0.00635
R7982 DVDD.n18815 DVDD.n18814 0.00635
R7983 DVDD.n19149 DVDD.n19148 0.00635
R7984 DVDD.n7262 DVDD.n7261 0.00635
R7985 DVDD.n10075 DVDD.n10074 0.00635
R7986 DVDD.n7628 DVDD.n7627 0.00635
R7987 DVDD.n3898 DVDD.n3897 0.00635
R7988 DVDD.n7118 DVDD.n7117 0.00635
R7989 DVDD.n7652 DVDD.n7651 0.00635
R7990 DVDD.n1811 DVDD.n1810 0.00635
R7991 DVDD.n3787 DVDD.n3786 0.00635
R7992 DVDD.n2820 DVDD.n2819 0.00635
R7993 DVDD.n20294 DVDD.n20293 0.00635
R7994 DVDD.n20316 DVDD.n20315 0.00635
R7995 DVDD.n14843 DVDD.n14842 0.00635
R7996 DVDD.n14863 DVDD.n14862 0.00635
R7997 DVDD.n15087 DVDD.n15086 0.00635
R7998 DVDD.n10705 DVDD.n10704 0.00635
R7999 DVDD.n10611 DVDD.n10610 0.00635
R8000 DVDD.n3379 DVDD.n3378 0.00635
R8001 DVDD.n3374 DVDD.n3373 0.00635
R8002 DVDD.n18737 DVDD.n18736 0.00635
R8003 DVDD.n18695 DVDD.n18691 0.00635
R8004 DVDD.n18667 DVDD.n18664 0.00635
R8005 DVDD.n18466 DVDD.n18465 0.00635
R8006 DVDD.n18448 DVDD.n18431 0.00635
R8007 DVDD.n18443 DVDD.n18442 0.00635
R8008 DVDD.n7275 DVDD.n7274 0.00635
R8009 DVDD.n12262 DVDD.n12261 0.00634646
R8010 DVDD.n13308 DVDD.n13307 0.00634646
R8011 DVDD.n3327 DVDD.n3326 0.00633333
R8012 DVDD.n15251 DVDD 0.00626307
R8013 DVDD DVDD.n15289 0.00626307
R8014 DVDD.n10484 DVDD.n10483 0.0062375
R8015 DVDD.n10451 DVDD.n10409 0.0062375
R8016 DVDD.n2403 DVDD.n2400 0.00622143
R8017 DVDD.n2599 DVDD.n2596 0.00622143
R8018 DVDD.n14432 DVDD.n14431 0.00616929
R8019 DVDD.n5990 DVDD.n5989 0.00616929
R8020 DVDD.n12653 DVDD.n12652 0.00616929
R8021 DVDD.n17806 DVDD.n17805 0.00616929
R8022 DVDD.n4453 DVDD.n4452 0.00616929
R8023 DVDD.n8727 DVDD.n8726 0.00616929
R8024 DVDD.n3398 DVDD.n3397 0.00616906
R8025 DVDD.n3392 DVDD.n3391 0.00616906
R8026 DVDD.n2373 DVDD.n2372 0.00615714
R8027 DVDD.n2420 DVDD.n2419 0.00615714
R8028 DVDD.n2571 DVDD.n2570 0.00615714
R8029 DVDD.n2616 DVDD.n2615 0.00615714
R8030 DVDD.n4128 DVDD.n4127 0.00615714
R8031 DVDD.n8510 DVDD.n8509 0.00615714
R8032 DVDD.n11212 DVDD.n11211 0.00615714
R8033 DVDD.n13855 DVDD.n13852 0.00615714
R8034 DVDD.n18832 DVDD.n18831 0.006125
R8035 DVDD.n18818 DVDD.n18817 0.006125
R8036 DVDD.n19162 DVDD.n19161 0.006125
R8037 DVDD.n7271 DVDD.n7270 0.006125
R8038 DVDD.n3843 DVDD.n3842 0.006125
R8039 DVDD.n3855 DVDD.n3854 0.006125
R8040 DVDD.n7611 DVDD.n7610 0.006125
R8041 DVDD.n3895 DVDD.n3894 0.006125
R8042 DVDD.n3911 DVDD.n3910 0.006125
R8043 DVDD.n7638 DVDD.n7637 0.006125
R8044 DVDD.n128 DVDD.n127 0.006125
R8045 DVDD.n140 DVDD.n139 0.006125
R8046 DVDD.n3784 DVDD.n3783 0.006125
R8047 DVDD.n3800 DVDD.n3799 0.006125
R8048 DVDD.n20279 DVDD.n20278 0.006125
R8049 DVDD.n20326 DVDD.n20325 0.006125
R8050 DVDD.n14880 DVDD.n14879 0.006125
R8051 DVDD.n14866 DVDD.n14865 0.006125
R8052 DVDD.n15096 DVDD.n15095 0.006125
R8053 DVDD.n10714 DVDD.n10713 0.006125
R8054 DVDD.n10624 DVDD.n10623 0.006125
R8055 DVDD.n7284 DVDD.n7283 0.006125
R8056 DVDD.n7703 DVDD.n7702 0.00608
R8057 DVDD.n3695 DVDD.n3694 0.00608
R8058 DVDD.n18541 DVDD.n18540 0.00608
R8059 DVDD.n2935 DVDD.n2934 0.00608
R8060 DVDD.n2957 DVDD.n2956 0.00608
R8061 DVDD.n9773 DVDD.n9772 0.00608
R8062 DVDD.n9794 DVDD.n9793 0.00608
R8063 DVDD.n9538 DVDD.n9537 0.00608
R8064 DVDD.n9253 DVDD.n9252 0.00608
R8065 DVDD.n9274 DVDD.n9273 0.00608
R8066 DVDD.n9295 DVDD.n9294 0.00608
R8067 DVDD.n2173 DVDD.n2172 0.00608
R8068 DVDD.n2195 DVDD.n2194 0.00608
R8069 DVDD.n2251 DVDD.n2250 0.00608
R8070 DVDD.n18910 DVDD.n18909 0.00608
R8071 DVDD.n7066 DVDD.n7065 0.00608
R8072 DVDD.n6842 DVDD.n6841 0.00608
R8073 DVDD.n6821 DVDD.n6820 0.00608
R8074 DVDD.n6570 DVDD.n6569 0.00608
R8075 DVDD.n1899 DVDD.n1898 0.00608
R8076 DVDD.n3989 DVDD.n3988 0.00608
R8077 DVDD.n3968 DVDD.n3967 0.00608
R8078 DVDD.n3947 DVDD.n3946 0.00608
R8079 DVDD.n19952 DVDD.n19951 0.00608
R8080 DVDD.n19974 DVDD.n19973 0.00608
R8081 DVDD.n20030 DVDD.n20029 0.00608
R8082 DVDD.n19028 DVDD.n19027 0.00608
R8083 DVDD.n4646 DVDD.n4645 0.00608
R8084 DVDD.n4879 DVDD.n4878 0.00608
R8085 DVDD.n4858 DVDD.n4857 0.00608
R8086 DVDD.n5161 DVDD.n5160 0.00608
R8087 DVDD.n19677 DVDD.n19676 0.00608
R8088 DVDD.n5294 DVDD.n5293 0.00608
R8089 DVDD.n5273 DVDD.n5272 0.00608
R8090 DVDD.n5252 DVDD.n5251 0.00608
R8091 DVDD.n993 DVDD.n992 0.00608
R8092 DVDD.n971 DVDD.n970 0.00608
R8093 DVDD.n938 DVDD.n937 0.00608
R8094 DVDD.n19237 DVDD.n19236 0.00608
R8095 DVDD.n18322 DVDD.n18321 0.00608
R8096 DVDD.n11874 DVDD.n11873 0.00608
R8097 DVDD.n11895 DVDD.n11894 0.00608
R8098 DVDD.n1322 DVDD.n1321 0.00608
R8099 DVDD.n12342 DVDD.n12341 0.00608
R8100 DVDD.n13164 DVDD.n13163 0.00608
R8101 DVDD.n13185 DVDD.n13184 0.00608
R8102 DVDD.n13206 DVDD.n13205 0.00608
R8103 DVDD.n3281 DVDD.n3280 0.00608
R8104 DVDD.n10409 DVDD.n10408 0.00606875
R8105 DVDD.n10582 DVDD.n10581 0.00606875
R8106 DVDD.n11141 DVDD.n11140 0.0060223
R8107 DVDD.n17244 DVDD.n17241 0.00600532
R8108 DVDD.n14094 DVDD.n14091 0.00600532
R8109 DVDD.n17411 DVDD.n17408 0.00600532
R8110 DVDD.n14005 DVDD.n14002 0.00600532
R8111 DVDD.n17594 DVDD.n17590 0.00600532
R8112 DVDD.n14215 DVDD.n14211 0.00600532
R8113 DVDD.n15212 DVDD.n15211 0.00597492
R8114 DVDD.n521 DVDD.n520 0.00596429
R8115 DVDD.n479 DVDD.n478 0.00596429
R8116 DVDD.n751 DVDD.n750 0.00596429
R8117 DVDD.n711 DVDD.n710 0.00596429
R8118 DVDD.n11292 DVDD.n11291 0.00596429
R8119 DVDD.n11274 DVDD.n11273 0.00596429
R8120 DVDD.n12498 DVDD.n12497 0.00596429
R8121 DVDD.n5761 DVDD.n5760 0.00596429
R8122 DVDD.n8294 DVDD.n8293 0.00592158
R8123 DVDD.n18831 DVDD.n18830 0.0059
R8124 DVDD.n12468 DVDD.n12467 0.0059
R8125 DVDD.n5702 DVDD.n5701 0.0059
R8126 DVDD.n6111 DVDD.n6110 0.0059
R8127 DVDD.n6116 DVDD.n6115 0.0059
R8128 DVDD.n4071 DVDD.n4070 0.0059
R8129 DVDD.n8485 DVDD.n8484 0.0059
R8130 DVDD.n12454 DVDD.n12453 0.0059
R8131 DVDD.n5660 DVDD.n5659 0.0059
R8132 DVDD.n4566 DVDD.n4565 0.0059
R8133 DVDD.n4564 DVDD.n4563 0.0059
R8134 DVDD.n4062 DVDD.n4061 0.0059
R8135 DVDD.n8466 DVDD.n8465 0.0059
R8136 DVDD.n12441 DVDD.n12440 0.0059
R8137 DVDD.n5614 DVDD.n5613 0.0059
R8138 DVDD.n4581 DVDD.n4580 0.0059
R8139 DVDD.n4579 DVDD.n4578 0.0059
R8140 DVDD.n4052 DVDD.n4051 0.0059
R8141 DVDD.n8448 DVDD.n8447 0.0059
R8142 DVDD.n12422 DVDD.n12421 0.0059
R8143 DVDD.n5567 DVDD.n5566 0.0059
R8144 DVDD.n4596 DVDD.n4595 0.0059
R8145 DVDD.n4594 DVDD.n4593 0.0059
R8146 DVDD.n4042 DVDD.n4041 0.0059
R8147 DVDD.n8430 DVDD.n8429 0.0059
R8148 DVDD.n19161 DVDD.n19160 0.0059
R8149 DVDD.n3856 DVDD.n3855 0.0059
R8150 DVDD.n7620 DVDD.n7619 0.0059
R8151 DVDD.n3912 DVDD.n3911 0.0059
R8152 DVDD.n7647 DVDD.n7646 0.0059
R8153 DVDD.n141 DVDD.n140 0.0059
R8154 DVDD.n3801 DVDD.n3800 0.0059
R8155 DVDD.n20288 DVDD.n20287 0.0059
R8156 DVDD.n20335 DVDD.n20334 0.0059
R8157 DVDD.n14930 DVDD.n14929 0.0059
R8158 DVDD.n15228 DVDD.n15227 0.0059
R8159 DVDD.n14879 DVDD.n14878 0.0059
R8160 DVDD.n10623 DVDD.n10622 0.0059
R8161 DVDD.n3432 DVDD.n3431 0.0059
R8162 DVDD.n3604 DVDD.n3603 0.0059
R8163 DVDD.n18347 DVDD.n18346 0.0059
R8164 DVDD.n14757 DVDD.n14756 0.0059
R8165 DVDD.n12932 DVDD.n12931 0.00588043
R8166 DVDD.n12951 DVDD.n12950 0.00588043
R8167 DVDD.n5516 DVDD.n5515 0.00588043
R8168 DVDD.n5541 DVDD.n5526 0.00588043
R8169 DVDD.n4014 DVDD.n4013 0.00588043
R8170 DVDD.n4036 DVDD.n4024 0.00588043
R8171 DVDD.n8970 DVDD.n8969 0.00588043
R8172 DVDD.n9038 DVDD.n8980 0.00588043
R8173 DVDD.n12903 DVDD.n12900 0.00588043
R8174 DVDD.n12892 DVDD.n12891 0.00588043
R8175 DVDD.n5723 DVDD.n5720 0.00588043
R8176 DVDD.n6062 DVDD.n6061 0.00588043
R8177 DVDD.n4094 DVDD.n4091 0.00588043
R8178 DVDD.n8997 DVDD.n8996 0.00588043
R8179 DVDD.n9010 DVDD.n9007 0.00588043
R8180 DVDD DVDD.n3823 0.00587887
R8181 DVDD.n7298 DVDD 0.00587887
R8182 DVDD.n7813 DVDD.n7812 0.00585135
R8183 DVDD.n6096 DVDD.n6095 0.00581496
R8184 DVDD.n12728 DVDD.n12727 0.00581496
R8185 DVDD.n4546 DVDD.n4545 0.00581496
R8186 DVDD.n8813 DVDD.n8812 0.00581496
R8187 DVDD.n10730 DVDD.n10729 0.0057875
R8188 DVDD.n10644 DVDD.n10643 0.0057875
R8189 DVDD.n4974 DVDD.n4973 0.00569488
R8190 DVDD.n11802 DVDD.n11801 0.00569487
R8191 DVDD.n6733 DVDD.n6732 0.00569487
R8192 DVDD.n9701 DVDD.n9700 0.00569487
R8193 DVDD.n15311 DVDD.n15310 0.005675
R8194 DVDD.n9905 DVDD.n9904 0.00560811
R8195 DVDD.n16039 DVDD.n16038 0.00558368
R8196 DVDD.n16012 DVDD.n16011 0.00558368
R8197 DVDD.n15651 DVDD.n15650 0.00558368
R8198 DVDD.n8154 DVDD.n8153 0.00558368
R8199 DVDD.n8114 DVDD.n8113 0.00558368
R8200 DVDD.n14895 DVDD.n14894 0.00550625
R8201 DVDD.n3405 DVDD.n3404 0.0054955
R8202 DVDD.n14433 DVDD.n14432 0.00546063
R8203 DVDD.n19890 DVDD.n19889 0.00546063
R8204 DVDD.n4975 DVDD.n4974 0.00546063
R8205 DVDD.n5657 DVDD.n5656 0.00546063
R8206 DVDD.n1487 DVDD.n1486 0.00546063
R8207 DVDD.n11778 DVDD.n11777 0.00546063
R8208 DVDD.n12780 DVDD.n12779 0.00546063
R8209 DVDD.n2111 DVDD.n2110 0.00546063
R8210 DVDD.n6709 DVDD.n6708 0.00546063
R8211 DVDD.n6157 DVDD.n6156 0.00546063
R8212 DVDD.n3510 DVDD.n3509 0.00546063
R8213 DVDD.n9677 DVDD.n9676 0.00546063
R8214 DVDD.n8859 DVDD.n8858 0.00546063
R8215 DVDD.n18820 DVDD.n18819 0.00545
R8216 DVDD.n407 DVDD.n406 0.00545
R8217 DVDD.n490 DVDD.n489 0.00545
R8218 DVDD.n444 DVDD.n443 0.00545
R8219 DVDD.n2338 DVDD.n2337 0.00545
R8220 DVDD.n2389 DVDD.n2388 0.00545
R8221 DVDD.n2500 DVDD.n2499 0.00545
R8222 DVDD.n3849 DVDD.n3848 0.00545
R8223 DVDD.n7615 DVDD.n7614 0.00545
R8224 DVDD.n3903 DVDD.n3902 0.00545
R8225 DVDD.n7642 DVDD.n7641 0.00545
R8226 DVDD.n134 DVDD.n133 0.00545
R8227 DVDD.n3792 DVDD.n3791 0.00545
R8228 DVDD.n20283 DVDD.n20282 0.00545
R8229 DVDD.n20330 DVDD.n20329 0.00545
R8230 DVDD.n638 DVDD.n637 0.00545
R8231 DVDD.n722 DVDD.n721 0.00545
R8232 DVDD.n676 DVDD.n675 0.00545
R8233 DVDD.n2536 DVDD.n2535 0.00545
R8234 DVDD.n2587 DVDD.n2586 0.00545
R8235 DVDD.n2712 DVDD.n2711 0.00545
R8236 DVDD.n14868 DVDD.n14867 0.00545
R8237 DVDD.n13731 DVDD.n13730 0.00545
R8238 DVDD.n11282 DVDD.n11281 0.00545
R8239 DVDD.n12492 DVDD.n12491 0.00545
R8240 DVDD.n5746 DVDD.n5745 0.00545
R8241 DVDD.n4158 DVDD.n4157 0.00545
R8242 DVDD.n8540 DVDD.n8539 0.00545
R8243 DVDD.n13872 DVDD.n13871 0.00545
R8244 DVDD.n13837 DVDD.n13836 0.00545
R8245 DVDD.n3375 DVDD.n3374 0.00545
R8246 DVDD.n3666 DVDD.n3665 0.00545
R8247 DVDD.n18610 DVDD.n18609 0.00545
R8248 DVDD.n18719 DVDD.n18718 0.00545
R8249 DVDD.n18724 DVDD.n18721 0.00545
R8250 DVDD.n18706 DVDD.n18705 0.00545
R8251 DVDD.n18393 DVDD.n18392 0.00545
R8252 DVDD.n18391 DVDD.n18390 0.00545
R8253 DVDD.n8299 DVDD.n8298 0.00543509
R8254 DVDD.n16042 DVDD.n16041 0.0053954
R8255 DVDD.n16009 DVDD.n16008 0.0053954
R8256 DVDD.n15654 DVDD.n15653 0.0053954
R8257 DVDD.n15923 DVDD.n15922 0.0053954
R8258 DVDD.n8269 DVDD.n8268 0.0053954
R8259 DVDD.n8263 DVDD.n8262 0.0053954
R8260 DVDD.n8206 DVDD.n8205 0.0053954
R8261 DVDD.n8200 DVDD.n8199 0.0053954
R8262 DVDD.n8157 DVDD.n8156 0.0053954
R8263 DVDD.n9393 DVDD.n9392 0.0053954
R8264 DVDD.n8336 DVDD.n8335 0.0053954
R8265 DVDD.n8330 DVDD.n8329 0.0053954
R8266 DVDD.n8300 DVDD.n8299 0.0053954
R8267 DVDD.n4925 DVDD.n4924 0.00534051
R8268 DVDD.n1459 DVDD.n1458 0.00534051
R8269 DVDD.n2139 DVDD.n2138 0.00534051
R8270 DVDD.n3538 DVDD.n3537 0.00534051
R8271 DVDD.n12173 DVDD.n12172 0.00528346
R8272 DVDD.n13518 DVDD.n13517 0.00528346
R8273 DVDD.n13570 DVDD.n13569 0.00528346
R8274 DVDD.n13594 DVDD.n13593 0.00528346
R8275 DVDD.n13651 DVDD.n13650 0.00528346
R8276 DVDD.n13675 DVDD.n13674 0.00528346
R8277 DVDD.n18571 DVDD.n18570 0.00528346
R8278 DVDD.n14809 DVDD.n14808 0.00528346
R8279 DVDD.n15417 DVDD.n15416 0.00528346
R8280 DVDD.n15444 DVDD.n15443 0.00528346
R8281 DVDD.n14686 DVDD.n14685 0.00528346
R8282 DVDD.n14603 DVDD.n14602 0.00528346
R8283 DVDD.n14549 DVDD.n14548 0.00528346
R8284 DVDD.n14522 DVDD.n14521 0.00528346
R8285 DVDD.n14461 DVDD.n14460 0.00528346
R8286 DVDD.n14418 DVDD.n14417 0.00528346
R8287 DVDD.n5484 DVDD.n5483 0.00528346
R8288 DVDD.n5655 DVDD.n5654 0.00528346
R8289 DVDD.n6029 DVDD.n6028 0.00528346
R8290 DVDD.n5976 DVDD.n5975 0.00528346
R8291 DVDD.n12979 DVDD.n12978 0.00528346
R8292 DVDD.n12782 DVDD.n12781 0.00528346
R8293 DVDD.n12680 DVDD.n12679 0.00528346
R8294 DVDD.n12639 DVDD.n12638 0.00528346
R8295 DVDD.n240 DVDD.n239 0.00528346
R8296 DVDD.n18229 DVDD.n18228 0.00528346
R8297 DVDD.n18185 DVDD.n18184 0.00528346
R8298 DVDD.n18161 DVDD.n18160 0.00528346
R8299 DVDD.n18041 DVDD.n18040 0.00528346
R8300 DVDD.n17963 DVDD.n17962 0.00528346
R8301 DVDD.n17911 DVDD.n17910 0.00528346
R8302 DVDD.n17887 DVDD.n17886 0.00528346
R8303 DVDD.n17830 DVDD.n17829 0.00528346
R8304 DVDD.n17792 DVDD.n17791 0.00528346
R8305 DVDD.n6275 DVDD.n6274 0.00528346
R8306 DVDD.n6159 DVDD.n6158 0.00528346
R8307 DVDD.n4480 DVDD.n4479 0.00528346
R8308 DVDD.n4439 DVDD.n4438 0.00528346
R8309 DVDD.n9061 DVDD.n9060 0.00528346
R8310 DVDD.n8861 DVDD.n8860 0.00528346
R8311 DVDD.n8766 DVDD.n8765 0.00528346
R8312 DVDD.n8713 DVDD.n8712 0.00528346
R8313 DVDD.n10653 DVDD.n10652 0.00528125
R8314 DVDD.n2482 DVDD.n2480 0.00525714
R8315 DVDD.n3805 DVDD.n3804 0.005225
R8316 DVDD.n18823 DVDD.n18822 0.005225
R8317 DVDD.n19155 DVDD.n19154 0.005225
R8318 DVDD.n7266 DVDD.n7265 0.005225
R8319 DVDD.n3900 DVDD.n3899 0.005225
R8320 DVDD.n3789 DVDD.n3788 0.005225
R8321 DVDD.n14841 DVDD.n14840 0.005225
R8322 DVDD.n14871 DVDD.n14870 0.005225
R8323 DVDD.n15091 DVDD.n15090 0.005225
R8324 DVDD.n10709 DVDD.n10708 0.005225
R8325 DVDD.n10617 DVDD.n10616 0.005225
R8326 DVDD.n7279 DVDD.n7278 0.005225
R8327 DVDD.n15950 DVDD.n15949 0.00520711
R8328 DVDD.n15690 DVDD.n15689 0.00520711
R8329 DVDD.n8286 DVDD.n8285 0.00520711
R8330 DVDD.n8278 DVDD.n8277 0.00520711
R8331 DVDD.n8270 DVDD.n8269 0.00520711
R8332 DVDD.n8264 DVDD.n8263 0.00520711
R8333 DVDD.n8258 DVDD.n8257 0.00520711
R8334 DVDD.n8249 DVDD.n8248 0.00520711
R8335 DVDD.n8240 DVDD.n8239 0.00520711
R8336 DVDD.n8231 DVDD.n8230 0.00520711
R8337 DVDD.n8223 DVDD.n8222 0.00520711
R8338 DVDD.n8215 DVDD.n8214 0.00520711
R8339 DVDD.n8207 DVDD.n8206 0.00520711
R8340 DVDD.n8201 DVDD.n8200 0.00520711
R8341 DVDD.n8195 DVDD.n8194 0.00520711
R8342 DVDD.n8186 DVDD.n8185 0.00520711
R8343 DVDD.n8175 DVDD.n8174 0.00520711
R8344 DVDD.n9409 DVDD.n9408 0.00520711
R8345 DVDD.n8326 DVDD.n8325 0.00520711
R8346 DVDD.n8322 DVDD.n8321 0.00520711
R8347 DVDD.n9892 DVDD.n9891 0.00520711
R8348 DVDD.n1396 DVDD.n1395 0.0051633
R8349 DVDD.n1973 DVDD.n1972 0.0051633
R8350 DVDD.n3207 DVDD.n3206 0.0051633
R8351 DVDD.n2318 DVDD.n2317 0.00512857
R8352 DVDD.n2518 DVDD.n2517 0.00512857
R8353 DVDD.n19311 DVDD.n19310 0.0051063
R8354 DVDD.n13303 DVDD.n11298 0.0051063
R8355 DVDD.n13329 DVDD.n13328 0.0051063
R8356 DVDD.n13335 DVDD.n13334 0.0051063
R8357 DVDD.n13368 DVDD.n13367 0.0051063
R8358 DVDD.n13402 DVDD.n13401 0.0051063
R8359 DVDD.n13408 DVDD.n13407 0.0051063
R8360 DVDD.n13468 DVDD.n13467 0.0051063
R8361 DVDD.n13474 DVDD.n13473 0.0051063
R8362 DVDD.n13515 DVDD.n13514 0.0051063
R8363 DVDD.n13567 DVDD.n13566 0.0051063
R8364 DVDD.n13597 DVDD.n13596 0.0051063
R8365 DVDD.n13648 DVDD.n13647 0.0051063
R8366 DVDD.n13678 DVDD.n13677 0.0051063
R8367 DVDD.n2801 DVDD.n2800 0.0051063
R8368 DVDD.n18673 DVDD.n18672 0.0051063
R8369 DVDD.n10060 DVDD.n10059 0.0051063
R8370 DVDD.n15414 DVDD.n15413 0.0051063
R8371 DVDD.n15447 DVDD.n15446 0.0051063
R8372 DVDD.n14689 DVDD.n14688 0.0051063
R8373 DVDD.n14606 DVDD.n14605 0.0051063
R8374 DVDD.n14552 DVDD.n14551 0.0051063
R8375 DVDD.n14519 DVDD.n14518 0.0051063
R8376 DVDD.n14464 DVDD.n14463 0.0051063
R8377 DVDD.n14415 DVDD.n14414 0.0051063
R8378 DVDD.n19724 DVDD.n19723 0.0051063
R8379 DVDD.n3861 DVDD.n3860 0.0051063
R8380 DVDD.n4969 DVDD.n4968 0.0051063
R8381 DVDD.n4970 DVDD.n4969 0.0051063
R8382 DVDD.n5164 DVDD.n5163 0.0051063
R8383 DVDD.n5312 DVDD.n5311 0.0051063
R8384 DVDD.n5403 DVDD.n5402 0.0051063
R8385 DVDD.n5481 DVDD.n5480 0.0051063
R8386 DVDD.n5604 DVDD.n5603 0.0051063
R8387 DVDD.n6032 DVDD.n6031 0.0051063
R8388 DVDD.n5973 DVDD.n5972 0.0051063
R8389 DVDD.n1369 DVDD.n1368 0.0051063
R8390 DVDD.n10108 DVDD.n10107 0.0051063
R8391 DVDD.n11784 DVDD.n11783 0.0051063
R8392 DVDD.n11783 DVDD.n11782 0.0051063
R8393 DVDD.n11779 DVDD.n11778 0.0051063
R8394 DVDD.n12345 DVDD.n12344 0.0051063
R8395 DVDD.n13146 DVDD.n13145 0.0051063
R8396 DVDD.n13059 DVDD.n13058 0.0051063
R8397 DVDD.n12982 DVDD.n12981 0.0051063
R8398 DVDD.n12823 DVDD.n12822 0.0051063
R8399 DVDD.n12683 DVDD.n12682 0.0051063
R8400 DVDD.n12636 DVDD.n12635 0.0051063
R8401 DVDD.n833 DVDD.n832 0.0051063
R8402 DVDD.n152 DVDD.n151 0.0051063
R8403 DVDD.n10092 DVDD.n10091 0.0051063
R8404 DVDD.n18188 DVDD.n18187 0.0051063
R8405 DVDD.n18158 DVDD.n18157 0.0051063
R8406 DVDD.n18044 DVDD.n18043 0.0051063
R8407 DVDD.n17966 DVDD.n17965 0.0051063
R8408 DVDD.n17914 DVDD.n17913 0.0051063
R8409 DVDD.n17884 DVDD.n17883 0.0051063
R8410 DVDD.n17833 DVDD.n17832 0.0051063
R8411 DVDD.n17789 DVDD.n17788 0.0051063
R8412 DVDD.n1946 DVDD.n1945 0.0051063
R8413 DVDD.n7082 DVDD.n7081 0.0051063
R8414 DVDD.n6715 DVDD.n6714 0.0051063
R8415 DVDD.n6714 DVDD.n6713 0.0051063
R8416 DVDD.n6710 DVDD.n6709 0.0051063
R8417 DVDD.n6572 DVDD.n6517 0.0051063
R8418 DVDD.n6449 DVDD.n6448 0.0051063
R8419 DVDD.n6358 DVDD.n6357 0.0051063
R8420 DVDD.n6278 DVDD.n6277 0.0051063
R8421 DVDD.n6201 DVDD.n6200 0.0051063
R8422 DVDD.n4483 DVDD.n4482 0.0051063
R8423 DVDD.n4436 DVDD.n4435 0.0051063
R8424 DVDD.n3234 DVDD.n3233 0.0051063
R8425 DVDD.n7140 DVDD.n7139 0.0051063
R8426 DVDD.n9683 DVDD.n9682 0.0051063
R8427 DVDD.n9682 DVDD.n9681 0.0051063
R8428 DVDD.n9678 DVDD.n9677 0.0051063
R8429 DVDD.n9540 DVDD.n7903 0.0051063
R8430 DVDD.n9235 DVDD.n9234 0.0051063
R8431 DVDD.n9144 DVDD.n9143 0.0051063
R8432 DVDD.n9064 DVDD.n9063 0.0051063
R8433 DVDD.n8903 DVDD.n8902 0.0051063
R8434 DVDD.n8769 DVDD.n8768 0.0051063
R8435 DVDD.n8710 DVDD.n8709 0.0051063
R8436 DVDD.n379 DVDD.n378 0.00506429
R8437 DVDD.n524 DVDD.n414 0.00506429
R8438 DVDD.n483 DVDD.n482 0.00506429
R8439 DVDD.n437 DVDD.n436 0.00506429
R8440 DVDD.n610 DVDD.n609 0.00506429
R8441 DVDD.n753 DVDD.n645 0.00506429
R8442 DVDD.n715 DVDD.n714 0.00506429
R8443 DVDD.n669 DVDD.n668 0.00506429
R8444 DVDD.n11295 DVDD.n11294 0.00506429
R8445 DVDD.n11277 DVDD.n11276 0.00506429
R8446 DVDD.n12501 DVDD.n12500 0.00506429
R8447 DVDD.n5765 DVDD.n5764 0.00506429
R8448 DVDD.n14096 DVDD.n14095 0.00504787
R8449 DVDD.n14007 DVDD.n14006 0.00504787
R8450 DVDD.n14217 DVDD.n14216 0.00504787
R8451 DVDD.n15972 DVDD.n15971 0.00501883
R8452 DVDD.n8239 DVDD.n8238 0.00501883
R8453 DVDD.n9444 DVDD.n9443 0.00501883
R8454 DVDD.n8125 DVDD.n8124 0.00501883
R8455 DVDD.n3818 DVDD.n3817 0.005
R8456 DVDD.n2330 DVDD.n2329 0.005
R8457 DVDD.n2381 DVDD.n2380 0.005
R8458 DVDD.n2428 DVDD.n2427 0.005
R8459 DVDD.n19001 DVDD.n19000 0.005
R8460 DVDD.n10082 DVDD.n10081 0.005
R8461 DVDD.n7633 DVDD.n7632 0.005
R8462 DVDD.n7127 DVDD.n7126 0.005
R8463 DVDD.n7113 DVDD.n7112 0.005
R8464 DVDD.n7657 DVDD.n7656 0.005
R8465 DVDD.n1818 DVDD.n1817 0.005
R8466 DVDD.n2829 DVDD.n2828 0.005
R8467 DVDD.n2815 DVDD.n2814 0.005
R8468 DVDD.n20299 DVDD.n20298 0.005
R8469 DVDD.n20321 DVDD.n20320 0.005
R8470 DVDD.n2528 DVDD.n2527 0.005
R8471 DVDD.n2579 DVDD.n2578 0.005
R8472 DVDD.n2624 DVDD.n2623 0.005
R8473 DVDD.n2666 DVDD.n2665 0.005
R8474 DVDD.n2688 DVDD.n2687 0.005
R8475 DVDD.n14854 DVDD.n14853 0.005
R8476 DVDD.n10604 DVDD.n10603 0.005
R8477 DVDD.n4166 DVDD.n4165 0.005
R8478 DVDD.n8548 DVDD.n8547 0.005
R8479 DVDD.n13880 DVDD.n13879 0.005
R8480 DVDD.n13844 DVDD.n13843 0.005
R8481 DVDD.n3428 DVDD.n3427 0.005
R8482 DVDD.n3667 DVDD.n3666 0.005
R8483 DVDD.n18611 DVDD.n18610 0.005
R8484 DVDD.n18724 DVDD.n18723 0.005
R8485 DVDD.n18709 DVDD.n18708 0.005
R8486 DVDD.n18667 DVDD.n18666 0.005
R8487 DVDD.n18428 DVDD.n18427 0.005
R8488 DVDD.n18448 DVDD.n18447 0.005
R8489 DVDD.n18438 DVDD.n18437 0.005
R8490 DVDD.n18435 DVDD.n18434 0.005
R8491 DVDD.n18434 DVDD.n18433 0.005
R8492 DVDD.n18388 DVDD.n18387 0.005
R8493 DVDD.n18354 DVDD.n18353 0.005
R8494 DVDD.n14767 DVDD.n14766 0.005
R8495 DVDD.n2329 DVDD.n2328 0.00493571
R8496 DVDD.n2380 DVDD.n2379 0.00493571
R8497 DVDD.n2427 DVDD.n2426 0.00493571
R8498 DVDD.n2527 DVDD.n2526 0.00493571
R8499 DVDD.n2578 DVDD.n2577 0.00493571
R8500 DVDD.n2623 DVDD.n2622 0.00493571
R8501 DVDD.n4166 DVDD.n4135 0.00493571
R8502 DVDD.n8548 DVDD.n8517 0.00493571
R8503 DVDD.n13880 DVDD.n11219 0.00493571
R8504 DVDD.n13845 DVDD.n13844 0.00493571
R8505 DVDD.n11476 DVDD.n11475 0.00492913
R8506 DVDD.n12214 DVDD.n12213 0.00492913
R8507 DVDD.n13339 DVDD.n13338 0.00492913
R8508 DVDD.n13344 DVDD.n13343 0.00492913
R8509 DVDD.n13374 DVDD.n13373 0.00492913
R8510 DVDD.n13383 DVDD.n13382 0.00492913
R8511 DVDD.n13392 DVDD.n13391 0.00492913
R8512 DVDD.n13401 DVDD.n13400 0.00492913
R8513 DVDD.n13407 DVDD.n13406 0.00492913
R8514 DVDD.n13413 DVDD.n13412 0.00492913
R8515 DVDD.n13422 DVDD.n13421 0.00492913
R8516 DVDD.n13431 DVDD.n13430 0.00492913
R8517 DVDD.n13440 DVDD.n13439 0.00492913
R8518 DVDD.n13449 DVDD.n13448 0.00492913
R8519 DVDD.n13458 DVDD.n13457 0.00492913
R8520 DVDD.n13467 DVDD.n13466 0.00492913
R8521 DVDD.n13473 DVDD.n13472 0.00492913
R8522 DVDD.n13479 DVDD.n13478 0.00492913
R8523 DVDD.n13488 DVDD.n13487 0.00492913
R8524 DVDD.n13499 DVDD.n13498 0.00492913
R8525 DVDD.n13541 DVDD.n13540 0.00492913
R8526 DVDD.n13622 DVDD.n13621 0.00492913
R8527 DVDD.n2734 DVDD.n2733 0.00492913
R8528 DVDD.n2775 DVDD.n2774 0.00492913
R8529 DVDD.n2810 DVDD.n2809 0.00492913
R8530 DVDD.n18474 DVDD.n18473 0.00492913
R8531 DVDD.n10069 DVDD.n10068 0.00492913
R8532 DVDD.n14824 DVDD.n14823 0.00492913
R8533 DVDD.n14717 DVDD.n14716 0.00492913
R8534 DVDD.n14634 DVDD.n14633 0.00492913
R8535 DVDD.n14580 DVDD.n14579 0.00492913
R8536 DVDD.n14492 DVDD.n14491 0.00492913
R8537 DVDD.n19891 DVDD.n19890 0.00492913
R8538 DVDD.n20051 DVDD.n20050 0.00492913
R8539 DVDD.n19056 DVDD.n19055 0.00492913
R8540 DVDD.n19018 DVDD.n19017 0.00492913
R8541 DVDD.n3870 DVDD.n3869 0.00492913
R8542 DVDD.n4788 DVDD.n4787 0.00492913
R8543 DVDD.n4921 DVDD.n4920 0.00492913
R8544 DVDD.n5019 DVDD.n5018 0.00492913
R8545 DVDD.n5189 DVDD.n5188 0.00492913
R8546 DVDD.n5208 DVDD.n5207 0.00492913
R8547 DVDD.n5555 DVDD.n5554 0.00492913
R8548 DVDD.n5607 DVDD.n5606 0.00492913
R8549 DVDD.n5611 DVDD.n5610 0.00492913
R8550 DVDD.n5673 DVDD.n5672 0.00492913
R8551 DVDD.n6088 DVDD.n6087 0.00492913
R8552 DVDD.n1486 DVDD.n1485 0.00492913
R8553 DVDD.n1722 DVDD.n1721 0.00492913
R8554 DVDD.n19438 DVDD.n19437 0.00492913
R8555 DVDD.n19227 DVDD.n19226 0.00492913
R8556 DVDD.n10117 DVDD.n10116 0.00492913
R8557 DVDD.n11614 DVDD.n11613 0.00492913
R8558 DVDD.n11832 DVDD.n11831 0.00492913
R8559 DVDD.n11735 DVDD.n11734 0.00492913
R8560 DVDD.n12369 DVDD.n12368 0.00492913
R8561 DVDD.n12388 DVDD.n12387 0.00492913
R8562 DVDD.n12862 DVDD.n12861 0.00492913
R8563 DVDD.n12820 DVDD.n12819 0.00492913
R8564 DVDD.n12816 DVDD.n12815 0.00492913
R8565 DVDD.n12768 DVDD.n12767 0.00492913
R8566 DVDD.n12720 DVDD.n12719 0.00492913
R8567 DVDD.n772 DVDD.n771 0.00492913
R8568 DVDD.n809 DVDD.n808 0.00492913
R8569 DVDD.n842 DVDD.n841 0.00492913
R8570 DVDD.n19170 DVDD.n19169 0.00492913
R8571 DVDD.n10101 DVDD.n10100 0.00492913
R8572 DVDD.n18214 DVDD.n18213 0.00492913
R8573 DVDD.n18070 DVDD.n18069 0.00492913
R8574 DVDD.n17992 DVDD.n17991 0.00492913
R8575 DVDD.n17940 DVDD.n17939 0.00492913
R8576 DVDD.n17859 DVDD.n17858 0.00492913
R8577 DVDD.n2112 DVDD.n2111 0.00492913
R8578 DVDD.n2272 DVDD.n2271 0.00492913
R8579 DVDD.n18948 DVDD.n18947 0.00492913
R8580 DVDD.n18945 DVDD.n18944 0.00492913
R8581 DVDD.n7091 DVDD.n7090 0.00492913
R8582 DVDD.n6896 DVDD.n6895 0.00492913
R8583 DVDD.n6763 DVDD.n6762 0.00492913
R8584 DVDD.n6665 DVDD.n6664 0.00492913
R8585 DVDD.n6493 DVDD.n6492 0.00492913
R8586 DVDD.n6474 DVDD.n6473 0.00492913
R8587 DVDD.n6241 DVDD.n6240 0.00492913
R8588 DVDD.n6198 DVDD.n6197 0.00492913
R8589 DVDD.n6195 DVDD.n6194 0.00492913
R8590 DVDD.n6151 DVDD.n6150 0.00492913
R8591 DVDD.n4538 DVDD.n4537 0.00492913
R8592 DVDD.n3511 DVDD.n3510 0.00492913
R8593 DVDD.n3716 DVDD.n3715 0.00492913
R8594 DVDD.n18785 DVDD.n18784 0.00492913
R8595 DVDD.n18531 DVDD.n18530 0.00492913
R8596 DVDD.n7149 DVDD.n7148 0.00492913
R8597 DVDD.n7870 DVDD.n7869 0.00492913
R8598 DVDD.n9731 DVDD.n9730 0.00492913
R8599 DVDD.n9633 DVDD.n9632 0.00492913
R8600 DVDD.n8390 DVDD.n8389 0.00492913
R8601 DVDD.n8409 DVDD.n8408 0.00492913
R8602 DVDD.n8943 DVDD.n8942 0.00492913
R8603 DVDD.n8900 DVDD.n8899 0.00492913
R8604 DVDD.n8897 DVDD.n8896 0.00492913
R8605 DVDD.n8853 DVDD.n8852 0.00492913
R8606 DVDD.n8805 DVDD.n8804 0.00492913
R8607 DVDD.n7372 DVDD.n7368 0.0049
R8608 DVDD.n74 DVDD.n70 0.0049
R8609 DVDD.n7245 DVDD.n7241 0.0049
R8610 DVDD.n20264 DVDD.n20260 0.0049
R8611 DVDD.n19720 DVDD.n19719 0.00489758
R8612 DVDD.n5022 DVDD.n5021 0.00489753
R8613 DVDD.n2692 DVDD 0.00487143
R8614 DVDD DVDD.n11223 0.00487143
R8615 DVDD.n14925 DVDD.n14924 0.00483125
R8616 DVDD.n14888 DVDD.n14887 0.00483125
R8617 DVDD.n15223 DVDD.n15222 0.00483125
R8618 DVDD.n15291 DVDD.n15290 0.00483125
R8619 DVDD.n10404 DVDD.n10403 0.00483125
R8620 DVDD.n10587 DVDD.n10586 0.00483125
R8621 DVDD.n10637 DVDD.n10636 0.00483125
R8622 DVDD.n8214 DVDD.n8213 0.00483054
R8623 DVDD.n8210 DVDD.n8209 0.00483054
R8624 DVDD.n8350 DVDD.n8349 0.00483054
R8625 DVDD.n8341 DVDD.n8340 0.00483054
R8626 DVDD.n8335 DVDD.n8334 0.00483054
R8627 DVDD.n8329 DVDD.n8328 0.00483054
R8628 DVDD.n8321 DVDD.n8320 0.00483054
R8629 DVDD.n8313 DVDD.n8312 0.00483054
R8630 DVDD.n8305 DVDD.n8304 0.00483054
R8631 DVDD.n5086 DVDD.n5085 0.00480905
R8632 DVDD.n8477 DVDD.n8476 0.00480864
R8633 DVDD.n8459 DVDD.n8458 0.00480864
R8634 DVDD.n8441 DVDD.n8440 0.00480864
R8635 DVDD.n17246 DVDD.n17245 0.00480851
R8636 DVDD.n17413 DVDD.n17412 0.00480851
R8637 DVDD.n17596 DVDD.n17595 0.00480851
R8638 DVDD.n12770 DVDD.n12769 0.00480845
R8639 DVDD.n12428 DVDD.n12427 0.00480845
R8640 DVDD.n12409 DVDD.n12408 0.00480845
R8641 DVDD.n524 DVDD.n523 0.00480714
R8642 DVDD.n482 DVDD.n481 0.00480714
R8643 DVDD.n436 DVDD.n435 0.00480714
R8644 DVDD.n431 DVDD.n430 0.00480714
R8645 DVDD.n753 DVDD.n752 0.00480714
R8646 DVDD.n714 DVDD.n713 0.00480714
R8647 DVDD.n668 DVDD.n667 0.00480714
R8648 DVDD.n663 DVDD.n662 0.00480714
R8649 DVDD.n11294 DVDD.n11293 0.00480714
R8650 DVDD.n11276 DVDD.n11275 0.00480714
R8651 DVDD.n12500 DVDD.n12499 0.00480714
R8652 DVDD.n5764 DVDD.n5763 0.00480714
R8653 DVDD.n3819 DVDD.n3818 0.004775
R8654 DVDD.n19002 DVDD.n19001 0.004775
R8655 DVDD.n7223 DVDD.n7222 0.004775
R8656 DVDD.n10081 DVDD.n10080 0.004775
R8657 DVDD.n7126 DVDD.n7125 0.004775
R8658 DVDD.n1817 DVDD.n1816 0.004775
R8659 DVDD.n2828 DVDD.n2827 0.004775
R8660 DVDD.n14855 DVDD.n14854 0.004775
R8661 DVDD.n15082 DVDD.n15081 0.004775
R8662 DVDD.n10700 DVDD.n10699 0.004775
R8663 DVDD.n10605 DVDD.n10604 0.004775
R8664 DVDD.n7294 DVDD.n7293 0.004775
R8665 DVDD.n10495 DVDD.n10494 0.00476
R8666 DVDD.n10494 DVDD.n10493 0.00476
R8667 DVDD.n10493 DVDD.n10492 0.00476
R8668 DVDD.n10492 DVDD.n10491 0.00476
R8669 DVDD.n10491 DVDD.n10490 0.00476
R8670 DVDD.n10490 DVDD.n10489 0.00476
R8671 DVDD.n10489 DVDD.n10488 0.00476
R8672 DVDD.n10488 DVDD.n10487 0.00476
R8673 DVDD.n10487 DVDD.n10486 0.00476
R8674 DVDD.n10486 DVDD.n10485 0.00476
R8675 DVDD.n10424 DVDD.n10423 0.00476
R8676 DVDD.n10423 DVDD.n10422 0.00476
R8677 DVDD.n10422 DVDD.n10421 0.00476
R8678 DVDD.n10421 DVDD.n10420 0.00476
R8679 DVDD.n10420 DVDD.n10419 0.00476
R8680 DVDD.n10419 DVDD.n10418 0.00476
R8681 DVDD.n10418 DVDD.n10417 0.00476
R8682 DVDD.n14944 DVDD.n14943 0.00476
R8683 DVDD.n14945 DVDD.n14944 0.00476
R8684 DVDD.n14946 DVDD.n14945 0.00476
R8685 DVDD.n14947 DVDD.n14946 0.00476
R8686 DVDD.n14948 DVDD.n14947 0.00476
R8687 DVDD.n14949 DVDD.n14948 0.00476
R8688 DVDD.n15015 DVDD.n15014 0.00476
R8689 DVDD.n15016 DVDD.n15015 0.00476
R8690 DVDD.n15017 DVDD.n15016 0.00476
R8691 DVDD.n15018 DVDD.n15017 0.00476
R8692 DVDD.n15019 DVDD.n15018 0.00476
R8693 DVDD.n15020 DVDD.n15019 0.00476
R8694 DVDD.n15021 DVDD.n15020 0.00476
R8695 DVDD.n15022 DVDD.n15021 0.00476
R8696 DVDD.n15023 DVDD.n15022 0.00476
R8697 DVDD.n10360 DVDD.n10358 0.00476
R8698 DVDD.n10362 DVDD.n10360 0.00476
R8699 DVDD.n10364 DVDD.n10362 0.00476
R8700 DVDD.n10366 DVDD.n10364 0.00476
R8701 DVDD.n10539 DVDD.n10537 0.00476
R8702 DVDD.n10537 DVDD.n10535 0.00476
R8703 DVDD.n10535 DVDD.n10533 0.00476
R8704 DVDD.n10533 DVDD.n10531 0.00476
R8705 DVDD.n10531 DVDD.n10529 0.00476
R8706 DVDD.n10529 DVDD.n10527 0.00476
R8707 DVDD.n10527 DVDD.n10525 0.00476
R8708 DVDD.n10525 DVDD.n10523 0.00476
R8709 DVDD.n10498 DVDD.n10496 0.00476
R8710 DVDD.n10496 DVDD.n10461 0.00476
R8711 DVDD.n10461 DVDD.n10460 0.00476
R8712 DVDD.n10460 DVDD.n10459 0.00476
R8713 DVDD.n10459 DVDD.n10458 0.00476
R8714 DVDD.n10458 DVDD.n10457 0.00476
R8715 DVDD.n10457 DVDD.n10456 0.00476
R8716 DVDD.n10456 DVDD.n10455 0.00476
R8717 DVDD.n10455 DVDD.n10454 0.00476
R8718 DVDD.n10454 DVDD.n10453 0.00476
R8719 DVDD.n10453 DVDD.n10452 0.00476
R8720 DVDD.n10425 DVDD.n10416 0.00476
R8721 DVDD.n10416 DVDD.n10415 0.00476
R8722 DVDD.n10415 DVDD.n10414 0.00476
R8723 DVDD.n10414 DVDD.n10413 0.00476
R8724 DVDD.n10413 DVDD.n10412 0.00476
R8725 DVDD.n10412 DVDD.n10411 0.00476
R8726 DVDD.n10411 DVDD.n10410 0.00476
R8727 DVDD.n14937 DVDD.n14936 0.00476
R8728 DVDD.n14938 DVDD.n14937 0.00476
R8729 DVDD.n14939 DVDD.n14938 0.00476
R8730 DVDD.n14940 DVDD.n14939 0.00476
R8731 DVDD.n14941 DVDD.n14940 0.00476
R8732 DVDD.n14942 DVDD.n14941 0.00476
R8733 DVDD.n14950 DVDD.n14942 0.00476
R8734 DVDD.n14983 DVDD.n14982 0.00476
R8735 DVDD.n14984 DVDD.n14983 0.00476
R8736 DVDD.n14985 DVDD.n14984 0.00476
R8737 DVDD.n14986 DVDD.n14985 0.00476
R8738 DVDD.n14987 DVDD.n14986 0.00476
R8739 DVDD.n14988 DVDD.n14987 0.00476
R8740 DVDD.n14989 DVDD.n14988 0.00476
R8741 DVDD.n14990 DVDD.n14989 0.00476
R8742 DVDD.n15024 DVDD.n14990 0.00476
R8743 DVDD.n15026 DVDD.n15024 0.00476
R8744 DVDD.n15028 DVDD.n15026 0.00476
R8745 DVDD.n15061 DVDD.n15059 0.00476
R8746 DVDD.n15063 DVDD.n15061 0.00476
R8747 DVDD.n15065 DVDD.n15063 0.00476
R8748 DVDD.n15067 DVDD.n15065 0.00476
R8749 DVDD.n15069 DVDD.n15067 0.00476
R8750 DVDD.n15071 DVDD.n15069 0.00476
R8751 DVDD.n15073 DVDD.n15071 0.00476
R8752 DVDD.n15313 DVDD.n15073 0.00476
R8753 DVDD.n15376 DVDD.n15374 0.00476
R8754 DVDD.n15374 DVDD.n15372 0.00476
R8755 DVDD.n15372 DVDD.n15370 0.00476
R8756 DVDD.n15370 DVDD.n15368 0.00476
R8757 DVDD.n16512 DVDD.n16511 0.00476
R8758 DVDD.n16513 DVDD.n16512 0.00476
R8759 DVDD.n16514 DVDD.n16513 0.00476
R8760 DVDD.n16516 DVDD.n16514 0.00476
R8761 DVDD.n17150 DVDD.n17148 0.00476
R8762 DVDD.n17148 DVDD.n17146 0.00476
R8763 DVDD.n17146 DVDD.n17144 0.00476
R8764 DVDD.n17144 DVDD.n17142 0.00476
R8765 DVDD.n17142 DVDD.n17139 0.00476
R8766 DVDD.n17139 DVDD.n17138 0.00476
R8767 DVDD.n17138 DVDD.n17135 0.00476
R8768 DVDD.n17135 DVDD.n17134 0.00476
R8769 DVDD.n17109 DVDD.n17107 0.00476
R8770 DVDD.n17107 DVDD.n17104 0.00476
R8771 DVDD.n17104 DVDD.n17103 0.00476
R8772 DVDD.n17103 DVDD.n17101 0.00476
R8773 DVDD.n17101 DVDD.n17098 0.00476
R8774 DVDD.n17098 DVDD.n17097 0.00476
R8775 DVDD.n17097 DVDD.n17095 0.00476
R8776 DVDD.n17095 DVDD.n17093 0.00476
R8777 DVDD.n17093 DVDD.n17090 0.00476
R8778 DVDD.n17090 DVDD.n17089 0.00476
R8779 DVDD.n17089 DVDD.n17087 0.00476
R8780 DVDD.n17057 DVDD.n17055 0.00476
R8781 DVDD.n17055 DVDD.n17053 0.00476
R8782 DVDD.n17053 DVDD.n17051 0.00476
R8783 DVDD.n17051 DVDD.n17048 0.00476
R8784 DVDD.n17048 DVDD.n17047 0.00476
R8785 DVDD.n17047 DVDD.n17045 0.00476
R8786 DVDD.n10993 DVDD.n10992 0.00476
R8787 DVDD.n10996 DVDD.n10993 0.00476
R8788 DVDD.n10998 DVDD.n10996 0.00476
R8789 DVDD.n11000 DVDD.n10998 0.00476
R8790 DVDD.n11002 DVDD.n11000 0.00476
R8791 DVDD.n11004 DVDD.n11002 0.00476
R8792 DVDD.n11006 DVDD.n11004 0.00476
R8793 DVDD.n11008 DVDD.n11006 0.00476
R8794 DVDD.n11045 DVDD.n11041 0.00476
R8795 DVDD.n11047 DVDD.n11045 0.00476
R8796 DVDD.n11049 DVDD.n11047 0.00476
R8797 DVDD.n11051 DVDD.n11049 0.00476
R8798 DVDD.n11053 DVDD.n11051 0.00476
R8799 DVDD.n11055 DVDD.n11053 0.00476
R8800 DVDD.n11057 DVDD.n11055 0.00476
R8801 DVDD.n11059 DVDD.n11057 0.00476
R8802 DVDD.n11061 DVDD.n11059 0.00476
R8803 DVDD.n11063 DVDD.n11061 0.00476
R8804 DVDD.n11065 DVDD.n11063 0.00476
R8805 DVDD.n11098 DVDD.n11096 0.00476
R8806 DVDD.n11100 DVDD.n11098 0.00476
R8807 DVDD.n11102 DVDD.n11100 0.00476
R8808 DVDD.n11104 DVDD.n11102 0.00476
R8809 DVDD.n11106 DVDD.n11104 0.00476
R8810 DVDD.n11108 DVDD.n11106 0.00476
R8811 DVDD.n11110 DVDD.n11108 0.00476
R8812 DVDD.n11123 DVDD.n11110 0.00476
R8813 DVDD.n11185 DVDD.n11183 0.00476
R8814 DVDD.n11183 DVDD.n11181 0.00476
R8815 DVDD.n11181 DVDD.n11179 0.00476
R8816 DVDD.n11179 DVDD.n11177 0.00476
R8817 DVDD.n16854 DVDD.n16853 0.00476
R8818 DVDD.n16855 DVDD.n16854 0.00476
R8819 DVDD.n16856 DVDD.n16855 0.00476
R8820 DVDD.n16858 DVDD.n16856 0.00476
R8821 DVDD.n17041 DVDD.n17039 0.00476
R8822 DVDD.n17039 DVDD.n17036 0.00476
R8823 DVDD.n17036 DVDD.n17035 0.00476
R8824 DVDD.n17035 DVDD.n17033 0.00476
R8825 DVDD.n17033 DVDD.n17031 0.00476
R8826 DVDD.n17031 DVDD.n17027 0.00476
R8827 DVDD.n17027 DVDD.n17026 0.00476
R8828 DVDD.n17026 DVDD.n17025 0.00476
R8829 DVDD.n16993 DVDD.n16991 0.00476
R8830 DVDD.n16991 DVDD.n16989 0.00476
R8831 DVDD.n16989 DVDD.n16987 0.00476
R8832 DVDD.n16987 DVDD.n16985 0.00476
R8833 DVDD.n16985 DVDD.n16983 0.00476
R8834 DVDD.n16983 DVDD.n16981 0.00476
R8835 DVDD.n16981 DVDD.n16979 0.00476
R8836 DVDD.n16979 DVDD.n16977 0.00476
R8837 DVDD.n16977 DVDD.n16975 0.00476
R8838 DVDD.n16975 DVDD.n16973 0.00476
R8839 DVDD.n16973 DVDD.n16967 0.00476
R8840 DVDD.n16933 DVDD.n16931 0.00476
R8841 DVDD.n16931 DVDD.n16929 0.00476
R8842 DVDD.n16929 DVDD.n16926 0.00476
R8843 DVDD.n16926 DVDD.n16925 0.00476
R8844 DVDD.n16925 DVDD.n16922 0.00476
R8845 DVDD.n16121 DVDD.n16120 0.00476
R8846 DVDD.n16122 DVDD.n16121 0.00476
R8847 DVDD.n16126 DVDD.n16122 0.00476
R8848 DVDD.n16128 DVDD.n16126 0.00476
R8849 DVDD.n16130 DVDD.n16128 0.00476
R8850 DVDD.n16131 DVDD.n16130 0.00476
R8851 DVDD.n16134 DVDD.n16131 0.00476
R8852 DVDD.n16136 DVDD.n16134 0.00476
R8853 DVDD.n16138 DVDD.n16136 0.00476
R8854 DVDD.n16238 DVDD.n16236 0.00476
R8855 DVDD.n16240 DVDD.n16238 0.00476
R8856 DVDD.n16241 DVDD.n16240 0.00476
R8857 DVDD.n16244 DVDD.n16241 0.00476
R8858 DVDD.n16246 DVDD.n16244 0.00476
R8859 DVDD.n16248 DVDD.n16246 0.00476
R8860 DVDD.n16250 DVDD.n16248 0.00476
R8861 DVDD.n16252 DVDD.n16250 0.00476
R8862 DVDD.n16254 DVDD.n16252 0.00476
R8863 DVDD.n16256 DVDD.n16254 0.00476
R8864 DVDD.n16258 DVDD.n16256 0.00476
R8865 DVDD.n16296 DVDD.n16295 0.00476
R8866 DVDD.n16299 DVDD.n16296 0.00476
R8867 DVDD.n16301 DVDD.n16299 0.00476
R8868 DVDD.n16303 DVDD.n16301 0.00476
R8869 DVDD.n16305 DVDD.n16303 0.00476
R8870 DVDD.n16307 DVDD.n16305 0.00476
R8871 DVDD.n16309 DVDD.n16307 0.00476
R8872 DVDD.n16311 DVDD.n16309 0.00476
R8873 DVDD.n16337 DVDD.n16335 0.00476
R8874 DVDD.n16340 DVDD.n16337 0.00476
R8875 DVDD.n16341 DVDD.n16340 0.00476
R8876 DVDD.n16376 DVDD.n16341 0.00476
R8877 DVDD.n16721 DVDD.n16720 0.00476
R8878 DVDD.n16722 DVDD.n16721 0.00476
R8879 DVDD.n16723 DVDD.n16722 0.00476
R8880 DVDD.n16725 DVDD.n16723 0.00476
R8881 DVDD.n16814 DVDD.n16812 0.00476
R8882 DVDD.n16812 DVDD.n16810 0.00476
R8883 DVDD.n16810 DVDD.n16808 0.00476
R8884 DVDD.n16808 DVDD.n16806 0.00476
R8885 DVDD.n16806 DVDD.n16800 0.00476
R8886 DVDD.n16800 DVDD.n16799 0.00476
R8887 DVDD.n16799 DVDD.n16798 0.00476
R8888 DVDD.n16798 DVDD.n16797 0.00476
R8889 DVDD.n16768 DVDD.n16766 0.00476
R8890 DVDD.n16766 DVDD.n16764 0.00476
R8891 DVDD.n16764 DVDD.n16762 0.00476
R8892 DVDD.n16762 DVDD.n16760 0.00476
R8893 DVDD.n16760 DVDD.n16758 0.00476
R8894 DVDD.n16758 DVDD.n16756 0.00476
R8895 DVDD.n16756 DVDD.n16754 0.00476
R8896 DVDD.n16754 DVDD.n16752 0.00476
R8897 DVDD.n16752 DVDD.n16749 0.00476
R8898 DVDD.n16749 DVDD.n16748 0.00476
R8899 DVDD.n16748 DVDD.n16745 0.00476
R8900 DVDD.n16891 DVDD.n16888 0.00476
R8901 DVDD.n16888 DVDD.n16887 0.00476
R8902 DVDD.n16887 DVDD.n16883 0.00476
R8903 DVDD.n16883 DVDD.n16882 0.00476
R8904 DVDD.n16882 DVDD.n16881 0.00476
R8905 DVDD.n16179 DVDD.n16177 0.00476
R8906 DVDD.n16180 DVDD.n16179 0.00476
R8907 DVDD.n16181 DVDD.n16180 0.00476
R8908 DVDD.n16182 DVDD.n16181 0.00476
R8909 DVDD.n16187 DVDD.n16182 0.00476
R8910 DVDD.n16189 DVDD.n16187 0.00476
R8911 DVDD.n16191 DVDD.n16189 0.00476
R8912 DVDD.n16193 DVDD.n16191 0.00476
R8913 DVDD.n16195 DVDD.n16193 0.00476
R8914 DVDD.n15539 DVDD.n15538 0.00476
R8915 DVDD.n15540 DVDD.n15539 0.00476
R8916 DVDD.n15544 DVDD.n15540 0.00476
R8917 DVDD.n15546 DVDD.n15544 0.00476
R8918 DVDD.n15548 DVDD.n15546 0.00476
R8919 DVDD.n15550 DVDD.n15548 0.00476
R8920 DVDD.n15552 DVDD.n15550 0.00476
R8921 DVDD.n15553 DVDD.n15552 0.00476
R8922 DVDD.n15556 DVDD.n15553 0.00476
R8923 DVDD.n15558 DVDD.n15556 0.00476
R8924 DVDD.n15560 DVDD.n15558 0.00476
R8925 DVDD.n15598 DVDD.n15596 0.00476
R8926 DVDD.n15599 DVDD.n15598 0.00476
R8927 DVDD.n15602 DVDD.n15599 0.00476
R8928 DVDD.n15604 DVDD.n15602 0.00476
R8929 DVDD.n15606 DVDD.n15604 0.00476
R8930 DVDD.n15608 DVDD.n15606 0.00476
R8931 DVDD.n15610 DVDD.n15608 0.00476
R8932 DVDD.n15612 DVDD.n15610 0.00476
R8933 DVDD.n15729 DVDD.n15727 0.00476
R8934 DVDD.n15727 DVDD.n15725 0.00476
R8935 DVDD.n15725 DVDD.n15723 0.00476
R8936 DVDD.n15723 DVDD.n15720 0.00476
R8937 DVDD.n16552 DVDD.n16551 0.00476
R8938 DVDD.n16553 DVDD.n16552 0.00476
R8939 DVDD.n16554 DVDD.n16553 0.00476
R8940 DVDD.n16556 DVDD.n16554 0.00476
R8941 DVDD.n16692 DVDD.n16688 0.00476
R8942 DVDD.n16688 DVDD.n16687 0.00476
R8943 DVDD.n16687 DVDD.n16686 0.00476
R8944 DVDD.n16686 DVDD.n16684 0.00476
R8945 DVDD.n16684 DVDD.n16682 0.00476
R8946 DVDD.n16682 DVDD.n16679 0.00476
R8947 DVDD.n16679 DVDD.n16678 0.00476
R8948 DVDD.n16678 DVDD.n16676 0.00476
R8949 DVDD.n16645 DVDD.n16643 0.00476
R8950 DVDD.n16643 DVDD.n16641 0.00476
R8951 DVDD.n16641 DVDD.n16638 0.00476
R8952 DVDD.n16638 DVDD.n16637 0.00476
R8953 DVDD.n16637 DVDD.n16635 0.00476
R8954 DVDD.n16635 DVDD.n16632 0.00476
R8955 DVDD.n16632 DVDD.n16631 0.00476
R8956 DVDD.n16631 DVDD.n16629 0.00476
R8957 DVDD.n16629 DVDD.n16626 0.00476
R8958 DVDD.n16626 DVDD.n16625 0.00476
R8959 DVDD.n16625 DVDD.n16623 0.00476
R8960 DVDD.n16588 DVDD.n16586 0.00476
R8961 DVDD.n16586 DVDD.n16584 0.00476
R8962 DVDD.n16584 DVDD.n16582 0.00476
R8963 DVDD.n16582 DVDD.n16580 0.00476
R8964 DVDD.n16580 DVDD.n16578 0.00476
R8965 DVDD.n15758 DVDD.n15757 0.00476
R8966 DVDD.n15761 DVDD.n15758 0.00476
R8967 DVDD.n15763 DVDD.n15761 0.00476
R8968 DVDD.n15764 DVDD.n15763 0.00476
R8969 DVDD.n15765 DVDD.n15764 0.00476
R8970 DVDD.n15769 DVDD.n15765 0.00476
R8971 DVDD.n15771 DVDD.n15769 0.00476
R8972 DVDD.n15773 DVDD.n15771 0.00476
R8973 DVDD.n15775 DVDD.n15773 0.00476
R8974 DVDD.n15817 DVDD.n15816 0.00476
R8975 DVDD.n15820 DVDD.n15817 0.00476
R8976 DVDD.n15822 DVDD.n15820 0.00476
R8977 DVDD.n15824 DVDD.n15822 0.00476
R8978 DVDD.n15826 DVDD.n15824 0.00476
R8979 DVDD.n15828 DVDD.n15826 0.00476
R8980 DVDD.n15829 DVDD.n15828 0.00476
R8981 DVDD.n15832 DVDD.n15829 0.00476
R8982 DVDD.n15834 DVDD.n15832 0.00476
R8983 DVDD.n15836 DVDD.n15834 0.00476
R8984 DVDD.n15838 DVDD.n15836 0.00476
R8985 DVDD.n15877 DVDD.n15875 0.00476
R8986 DVDD.n15879 DVDD.n15877 0.00476
R8987 DVDD.n15880 DVDD.n15879 0.00476
R8988 DVDD.n15881 DVDD.n15880 0.00476
R8989 DVDD.n15885 DVDD.n15881 0.00476
R8990 DVDD.n15887 DVDD.n15885 0.00476
R8991 DVDD.n15889 DVDD.n15887 0.00476
R8992 DVDD.n15891 DVDD.n15889 0.00476
R8993 DVDD.n16088 DVDD.n16086 0.00476
R8994 DVDD.n16086 DVDD.n16084 0.00476
R8995 DVDD.n16084 DVDD.n16082 0.00476
R8996 DVDD.n16082 DVDD.n16079 0.00476
R8997 DVDD.n16530 DVDD.n16529 0.00476
R8998 DVDD.n16529 DVDD.n16528 0.00476
R8999 DVDD.n16528 DVDD.n16527 0.00476
R9000 DVDD.n16527 DVDD.n16526 0.00476
R9001 DVDD.n16691 DVDD.n16690 0.00476
R9002 DVDD.n16690 DVDD.n16689 0.00476
R9003 DVDD.n16681 DVDD.n16680 0.00476
R9004 DVDD.n16640 DVDD.n16639 0.00476
R9005 DVDD.n16634 DVDD.n16633 0.00476
R9006 DVDD.n16628 DVDD.n16627 0.00476
R9007 DVDD.n15760 DVDD.n15759 0.00476
R9008 DVDD.n15767 DVDD.n15766 0.00476
R9009 DVDD.n15768 DVDD.n15767 0.00476
R9010 DVDD.n15819 DVDD.n15818 0.00476
R9011 DVDD.n15831 DVDD.n15830 0.00476
R9012 DVDD.n15883 DVDD.n15882 0.00476
R9013 DVDD.n15884 DVDD.n15883 0.00476
R9014 DVDD.n16081 DVDD.n16080 0.00476
R9015 DVDD.n16699 DVDD.n16698 0.00476
R9016 DVDD.n16698 DVDD.n16697 0.00476
R9017 DVDD.n16697 DVDD.n16696 0.00476
R9018 DVDD.n16696 DVDD.n16695 0.00476
R9019 DVDD.n16805 DVDD.n16804 0.00476
R9020 DVDD.n16804 DVDD.n16803 0.00476
R9021 DVDD.n16803 DVDD.n16802 0.00476
R9022 DVDD.n16802 DVDD.n16801 0.00476
R9023 DVDD.n16751 DVDD.n16750 0.00476
R9024 DVDD.n16747 DVDD.n16746 0.00476
R9025 DVDD.n16890 DVDD.n16889 0.00476
R9026 DVDD.n16886 DVDD.n16885 0.00476
R9027 DVDD.n16885 DVDD.n16884 0.00476
R9028 DVDD.n16184 DVDD.n16183 0.00476
R9029 DVDD.n16185 DVDD.n16184 0.00476
R9030 DVDD.n16186 DVDD.n16185 0.00476
R9031 DVDD.n15542 DVDD.n15541 0.00476
R9032 DVDD.n15543 DVDD.n15542 0.00476
R9033 DVDD.n15555 DVDD.n15554 0.00476
R9034 DVDD.n15601 DVDD.n15600 0.00476
R9035 DVDD.n15722 DVDD.n15721 0.00476
R9036 DVDD.n16825 DVDD.n16824 0.00476
R9037 DVDD.n16824 DVDD.n16823 0.00476
R9038 DVDD.n16823 DVDD.n16822 0.00476
R9039 DVDD.n16822 DVDD.n16821 0.00476
R9040 DVDD.n17038 DVDD.n17037 0.00476
R9041 DVDD.n17030 DVDD.n17029 0.00476
R9042 DVDD.n17029 DVDD.n17028 0.00476
R9043 DVDD.n16972 DVDD.n16971 0.00476
R9044 DVDD.n16928 DVDD.n16927 0.00476
R9045 DVDD.n16924 DVDD.n16923 0.00476
R9046 DVDD.n16124 DVDD.n16123 0.00476
R9047 DVDD.n16125 DVDD.n16124 0.00476
R9048 DVDD.n16133 DVDD.n16132 0.00476
R9049 DVDD.n16243 DVDD.n16242 0.00476
R9050 DVDD.n16298 DVDD.n16297 0.00476
R9051 DVDD.n16339 DVDD.n16338 0.00476
R9052 DVDD.n16481 DVDD.n16480 0.00476
R9053 DVDD.n16480 DVDD.n16479 0.00476
R9054 DVDD.n16479 DVDD.n16478 0.00476
R9055 DVDD.n16478 DVDD.n16477 0.00476
R9056 DVDD.n17141 DVDD.n17140 0.00476
R9057 DVDD.n17137 DVDD.n17136 0.00476
R9058 DVDD.n17106 DVDD.n17105 0.00476
R9059 DVDD.n17100 DVDD.n17099 0.00476
R9060 DVDD.n17092 DVDD.n17091 0.00476
R9061 DVDD.n17050 DVDD.n17049 0.00476
R9062 DVDD.n10995 DVDD.n10994 0.00476
R9063 DVDD.n11044 DVDD.n11043 0.00476
R9064 DVDD.n1584 DVDD.n1583 0.00475197
R9065 DVDD.n1606 DVDD.n1605 0.00475197
R9066 DVDD.n1612 DVDD.n1611 0.00475197
R9067 DVDD.n12184 DVDD.n12183 0.00475197
R9068 DVDD.n12249 DVDD.n12248 0.00475197
R9069 DVDD.n13432 DVDD.n13431 0.00475197
R9070 DVDD.n13726 DVDD.n13725 0.00475197
R9071 DVDD.n18483 DVDD.n18482 0.00475197
R9072 DVDD.n15484 DVDD.n15483 0.00475197
R9073 DVDD.n15515 DVDD.n15514 0.00475197
R9074 DVDD.n14662 DVDD.n14661 0.00475197
R9075 DVDD.n14378 DVDD.n14377 0.00475197
R9076 DVDD.n19770 DVDD.n19769 0.00475197
R9077 DVDD.n19840 DVDD.n19839 0.00475197
R9078 DVDD.n19995 DVDD.n19994 0.00475197
R9079 DVDD.n20007 DVDD.n20006 0.00475197
R9080 DVDD.n20079 DVDD.n20078 0.00475197
R9081 DVDD.n3873 DVDD.n3872 0.00475197
R9082 DVDD.n4706 DVDD.n4705 0.00475197
R9083 DVDD.n4776 DVDD.n4775 0.00475197
R9084 DVDD.n4920 DVDD.n4919 0.00475197
R9085 DVDD.n4948 DVDD.n4947 0.00475197
R9086 DVDD.n5044 DVDD.n5043 0.00475197
R9087 DVDD.n5090 DVDD.n5089 0.00475197
R9088 DVDD.n5339 DVDD.n5338 0.00475197
R9089 DVDD.n5385 DVDD.n5384 0.00475197
R9090 DVDD.n5456 DVDD.n5455 0.00475197
R9091 DVDD.n5940 DVDD.n5939 0.00475197
R9092 DVDD.n1415 DVDD.n1414 0.00475197
R9093 DVDD.n1536 DVDD.n1535 0.00475197
R9094 DVDD.n1683 DVDD.n1682 0.00475197
R9095 DVDD.n1695 DVDD.n1694 0.00475197
R9096 DVDD.n293 DVDD.n292 0.00475197
R9097 DVDD.n10120 DVDD.n10119 0.00475197
R9098 DVDD.n11413 DVDD.n11412 0.00475197
R9099 DVDD.n11602 DVDD.n11601 0.00475197
R9100 DVDD.n11833 DVDD.n11832 0.00475197
R9101 DVDD.n11805 DVDD.n11804 0.00475197
R9102 DVDD.n11710 DVDD.n11709 0.00475197
R9103 DVDD.n11664 DVDD.n11663 0.00475197
R9104 DVDD.n13120 DVDD.n13119 0.00475197
R9105 DVDD.n13076 DVDD.n13075 0.00475197
R9106 DVDD.n13007 DVDD.n13006 0.00475197
R9107 DVDD.n12603 DVDD.n12602 0.00475197
R9108 DVDD.n19179 DVDD.n19178 0.00475197
R9109 DVDD.n18125 DVDD.n18124 0.00475197
R9110 DVDD.n18096 DVDD.n18095 0.00475197
R9111 DVDD.n18018 DVDD.n18017 0.00475197
R9112 DVDD.n17756 DVDD.n17755 0.00475197
R9113 DVDD.n1992 DVDD.n1991 0.00475197
R9114 DVDD.n2062 DVDD.n2061 0.00475197
R9115 DVDD.n2216 DVDD.n2215 0.00475197
R9116 DVDD.n2228 DVDD.n2227 0.00475197
R9117 DVDD.n2300 DVDD.n2299 0.00475197
R9118 DVDD.n7094 DVDD.n7093 0.00475197
R9119 DVDD.n6978 DVDD.n6977 0.00475197
R9120 DVDD.n6908 DVDD.n6907 0.00475197
R9121 DVDD.n6764 DVDD.n6763 0.00475197
R9122 DVDD.n6736 DVDD.n6735 0.00475197
R9123 DVDD.n6640 DVDD.n6639 0.00475197
R9124 DVDD.n6592 DVDD.n6591 0.00475197
R9125 DVDD.n6422 DVDD.n6421 0.00475197
R9126 DVDD.n6376 DVDD.n6375 0.00475197
R9127 DVDD.n6305 DVDD.n6304 0.00475197
R9128 DVDD.n4399 DVDD.n4398 0.00475197
R9129 DVDD.n3188 DVDD.n3187 0.00475197
R9130 DVDD.n3461 DVDD.n3460 0.00475197
R9131 DVDD.n3566 DVDD.n3565 0.00475197
R9132 DVDD.n3554 DVDD.n3553 0.00475197
R9133 DVDD.n3779 DVDD.n3778 0.00475197
R9134 DVDD.n7152 DVDD.n7151 0.00475197
R9135 DVDD.n9995 DVDD.n9994 0.00475197
R9136 DVDD.n7858 DVDD.n7857 0.00475197
R9137 DVDD.n9732 DVDD.n9731 0.00475197
R9138 DVDD.n9704 DVDD.n9703 0.00475197
R9139 DVDD.n9608 DVDD.n9607 0.00475197
R9140 DVDD.n9560 DVDD.n9559 0.00475197
R9141 DVDD.n9208 DVDD.n9207 0.00475197
R9142 DVDD.n9162 DVDD.n9161 0.00475197
R9143 DVDD.n9091 DVDD.n9090 0.00475197
R9144 DVDD.n8673 DVDD.n8672 0.00475197
R9145 DVDD.n393 DVDD.n392 0.00474286
R9146 DVDD.n624 DVDD.n623 0.00474286
R9147 DVDD.n19887 DVDD.n19886 0.00472036
R9148 DVDD.n7410 DVDD.n7406 0.00468667
R9149 DVDD.n7458 DVDD.n7454 0.00468667
R9150 DVDD.n7499 DVDD.n7495 0.00468667
R9151 DVDD.n7326 DVDD.n7322 0.00468667
R9152 DVDD.n14963 DVDD.n14962 0.00467
R9153 DVDD.n15040 DVDD.n15039 0.00467
R9154 DVDD.n14831 DVDD.n14830 0.00467
R9155 DVDD.n16110 DVDD.n16109 0.00467
R9156 DVDD.n16072 DVDD.n16071 0.00467
R9157 DVDD.n15750 DVDD.n15749 0.00467
R9158 DVDD.n15714 DVDD.n15713 0.00467
R9159 DVDD.n11117 DVDD.n11116 0.00467
R9160 DVDD.n11021 DVDD.n11020 0.00467
R9161 DVDD.n11077 DVDD.n11076 0.00467
R9162 DVDD.n15521 DVDD.n15520 0.00467
R9163 DVDD.n8277 DVDD.n8276 0.00464226
R9164 DVDD.n8273 DVDD.n8272 0.00464226
R9165 DVDD.n9888 DVDD.n9887 0.00464226
R9166 DVDD.n7942 DVDD.n7941 0.00464226
R9167 DVDD.n7964 DVDD.n7963 0.00464226
R9168 DVDD.n7991 DVDD.n7990 0.00464226
R9169 DVDD.n7998 DVDD.n7997 0.00464226
R9170 DVDD.n8028 DVDD.n8027 0.00464226
R9171 DVDD.n8055 DVDD.n8054 0.00464226
R9172 DVDD.n8062 DVDD.n8061 0.00464226
R9173 DVDD.n10434 DVDD.n10433 0.00464
R9174 DVDD.n16531 DVDD.n16530 0.00464
R9175 DVDD.n16575 DVDD.n16574 0.00464
R9176 DVDD.n16700 DVDD.n16699 0.00464
R9177 DVDD.n16743 DVDD.n16742 0.00464
R9178 DVDD.n16826 DVDD.n16825 0.00464
R9179 DVDD.n16878 DVDD.n16877 0.00464
R9180 DVDD.n16482 DVDD.n16481 0.00464
R9181 DVDD.n5680 DVDD.n5679 0.0046318
R9182 DVDD.n12761 DVDD.n12760 0.0046318
R9183 DVDD.n6145 DVDD.n6144 0.0046318
R9184 DVDD.n8847 DVDD.n8846 0.0046318
R9185 DVDD.n4917 DVDD.n4916 0.00463168
R9186 DVDD.n4317 DVDD.n4304 0.00461744
R9187 DVDD.n4288 DVDD.n4279 0.00461744
R9188 DVDD.n4263 DVDD.n4254 0.00461744
R9189 DVDD.n1641 DVDD.n1640 0.0045748
R9190 DVDD.n13315 DVDD.n13314 0.0045748
R9191 DVDD.n13324 DVDD.n13323 0.0045748
R9192 DVDD.n13330 DVDD.n13329 0.0045748
R9193 DVDD.n13336 DVDD.n13335 0.0045748
R9194 DVDD.n13345 DVDD.n13344 0.0045748
R9195 DVDD.n13354 DVDD.n13353 0.0045748
R9196 DVDD.n13363 DVDD.n13362 0.0045748
R9197 DVDD.n13369 DVDD.n13368 0.0045748
R9198 DVDD.n13459 DVDD.n13458 0.0045748
R9199 DVDD.n13464 DVDD.n13463 0.0045748
R9200 DVDD.n19725 DVDD.n19724 0.0045748
R9201 DVDD.n19772 DVDD.n19771 0.0045748
R9202 DVDD.n19842 DVDD.n19841 0.0045748
R9203 DVDD.n19997 DVDD.n19996 0.0045748
R9204 DVDD.n20069 DVDD.n20068 0.0045748
R9205 DVDD.n19074 DVDD.n19073 0.0045748
R9206 DVDD.n4708 DVDD.n4707 0.0045748
R9207 DVDD.n4794 DVDD.n4793 0.0045748
R9208 DVDD.n1370 DVDD.n1369 0.0045748
R9209 DVDD.n1417 DVDD.n1416 0.0045748
R9210 DVDD.n1534 DVDD.n1533 0.0045748
R9211 DVDD.n1685 DVDD.n1684 0.0045748
R9212 DVDD.n1704 DVDD.n1703 0.0045748
R9213 DVDD.n19456 DVDD.n19455 0.0045748
R9214 DVDD.n11415 DVDD.n11414 0.0045748
R9215 DVDD.n11620 DVDD.n11619 0.0045748
R9216 DVDD.n13125 DVDD.n13124 0.0045748
R9217 DVDD.n13026 DVDD.n13025 0.0045748
R9218 DVDD.n1947 DVDD.n1946 0.0045748
R9219 DVDD.n1994 DVDD.n1993 0.0045748
R9220 DVDD.n2064 DVDD.n2063 0.0045748
R9221 DVDD.n2218 DVDD.n2217 0.0045748
R9222 DVDD.n2290 DVDD.n2289 0.0045748
R9223 DVDD.n18966 DVDD.n18965 0.0045748
R9224 DVDD.n6976 DVDD.n6975 0.0045748
R9225 DVDD.n6890 DVDD.n6889 0.0045748
R9226 DVDD.n6427 DVDD.n6426 0.0045748
R9227 DVDD.n6324 DVDD.n6323 0.0045748
R9228 DVDD.n3233 DVDD.n3232 0.0045748
R9229 DVDD.n3186 DVDD.n3185 0.0045748
R9230 DVDD.n3463 DVDD.n3462 0.0045748
R9231 DVDD.n3564 DVDD.n3563 0.0045748
R9232 DVDD.n3734 DVDD.n3733 0.0045748
R9233 DVDD.n18803 DVDD.n18802 0.0045748
R9234 DVDD.n9993 DVDD.n9992 0.0045748
R9235 DVDD.n7876 DVDD.n7875 0.0045748
R9236 DVDD.n9213 DVDD.n9212 0.0045748
R9237 DVDD.n9110 DVDD.n9109 0.0045748
R9238 DVDD.n13738 DVDD.n13737 0.00455714
R9239 DVDD.n13739 DVDD.n13738 0.00455714
R9240 DVDD.n13740 DVDD.n13739 0.00455714
R9241 DVDD.n13741 DVDD.n13740 0.00455714
R9242 DVDD.n13742 DVDD.n13741 0.00455714
R9243 DVDD.n13743 DVDD.n13742 0.00455714
R9244 DVDD.n13744 DVDD.n13743 0.00455714
R9245 DVDD.n13745 DVDD.n13744 0.00455714
R9246 DVDD.n13746 DVDD.n13745 0.00455714
R9247 DVDD.n13747 DVDD.n13746 0.00455714
R9248 DVDD.n13748 DVDD.n13747 0.00455714
R9249 DVDD.n13749 DVDD.n13748 0.00455714
R9250 DVDD.n13750 DVDD.n13749 0.00455714
R9251 DVDD.n13751 DVDD.n13750 0.00455714
R9252 DVDD.n13752 DVDD.n13751 0.00455714
R9253 DVDD.n13753 DVDD.n13752 0.00455714
R9254 DVDD.n13754 DVDD.n13753 0.00455714
R9255 DVDD.n13755 DVDD.n13754 0.00455714
R9256 DVDD.n13756 DVDD.n13755 0.00455714
R9257 DVDD.n13757 DVDD.n13756 0.00455714
R9258 DVDD.n13758 DVDD.n13757 0.00455714
R9259 DVDD.n13759 DVDD.n13758 0.00455714
R9260 DVDD.n13760 DVDD.n13759 0.00455714
R9261 DVDD.n13761 DVDD.n13760 0.00455714
R9262 DVDD.n13762 DVDD.n13761 0.00455714
R9263 DVDD.n13763 DVDD.n13762 0.00455714
R9264 DVDD.n13764 DVDD.n13763 0.00455714
R9265 DVDD.n13765 DVDD.n13764 0.00455714
R9266 DVDD.n13766 DVDD.n13765 0.00455714
R9267 DVDD.n13767 DVDD.n13766 0.00455714
R9268 DVDD.n13768 DVDD.n13767 0.00455714
R9269 DVDD.n13769 DVDD.n13768 0.00455714
R9270 DVDD.n13770 DVDD.n13769 0.00455714
R9271 DVDD.n13771 DVDD.n13770 0.00455714
R9272 DVDD.n13772 DVDD.n13771 0.00455714
R9273 DVDD.n13773 DVDD.n13772 0.00455714
R9274 DVDD.n13774 DVDD.n13773 0.00455714
R9275 DVDD.n13775 DVDD.n13774 0.00455714
R9276 DVDD.n13776 DVDD.n13775 0.00455714
R9277 DVDD.n13777 DVDD.n13776 0.00455714
R9278 DVDD.n13778 DVDD.n13777 0.00455714
R9279 DVDD.n13779 DVDD.n13778 0.00455714
R9280 DVDD.n13780 DVDD.n13779 0.00455714
R9281 DVDD.n13781 DVDD.n13780 0.00455714
R9282 DVDD.n13782 DVDD.n13781 0.00455714
R9283 DVDD.n13783 DVDD.n13782 0.00455714
R9284 DVDD.n13784 DVDD.n13783 0.00455714
R9285 DVDD.n13785 DVDD.n13784 0.00455714
R9286 DVDD.n13786 DVDD.n13785 0.00455714
R9287 DVDD.n13787 DVDD.n13786 0.00455714
R9288 DVDD.n13788 DVDD.n13787 0.00455714
R9289 DVDD.n13789 DVDD.n13788 0.00455714
R9290 DVDD.n13790 DVDD.n13789 0.00455714
R9291 DVDD.n13791 DVDD.n13790 0.00455714
R9292 DVDD.n13792 DVDD.n13791 0.00455714
R9293 DVDD.n13793 DVDD.n13792 0.00455714
R9294 DVDD.n13794 DVDD.n13793 0.00455714
R9295 DVDD.n13795 DVDD.n13794 0.00455714
R9296 DVDD.n13796 DVDD.n13795 0.00455714
R9297 DVDD.n13797 DVDD.n13796 0.00455714
R9298 DVDD.n13798 DVDD.n13797 0.00455714
R9299 DVDD.n13799 DVDD.n13798 0.00455714
R9300 DVDD.n13800 DVDD.n13799 0.00455714
R9301 DVDD.n13801 DVDD.n13800 0.00455714
R9302 DVDD.n13802 DVDD.n13801 0.00455714
R9303 DVDD.n13803 DVDD.n13802 0.00455714
R9304 DVDD.n13804 DVDD.n13803 0.00455714
R9305 DVDD.n13805 DVDD.n13804 0.00455714
R9306 DVDD.n13806 DVDD.n13805 0.00455714
R9307 DVDD.n13807 DVDD.n13806 0.00455714
R9308 DVDD.n13808 DVDD.n13807 0.00455714
R9309 DVDD.n13809 DVDD.n13808 0.00455714
R9310 DVDD.n13810 DVDD.n13809 0.00455714
R9311 DVDD.n13811 DVDD.n13810 0.00455714
R9312 DVDD.n13812 DVDD.n13811 0.00455714
R9313 DVDD.n13813 DVDD.n13812 0.00455714
R9314 DVDD.n13814 DVDD.n13813 0.00455714
R9315 DVDD.n13815 DVDD.n13814 0.00455714
R9316 DVDD.n13816 DVDD.n13815 0.00455714
R9317 DVDD.n13817 DVDD.n13816 0.00455714
R9318 DVDD.n13818 DVDD.n13817 0.00455714
R9319 DVDD.n13819 DVDD.n13818 0.00455714
R9320 DVDD.n13820 DVDD.n13819 0.00455714
R9321 DVDD.n13821 DVDD.n13820 0.00455714
R9322 DVDD.n13822 DVDD.n13821 0.00455714
R9323 DVDD.n13823 DVDD.n13822 0.00455714
R9324 DVDD.n13824 DVDD.n13823 0.00455714
R9325 DVDD.n13825 DVDD.n13824 0.00455714
R9326 DVDD.n13826 DVDD.n13825 0.00455714
R9327 DVDD.n13827 DVDD.n13826 0.00455714
R9328 DVDD.n13828 DVDD.n13827 0.00455714
R9329 DVDD.n13829 DVDD.n13828 0.00455714
R9330 DVDD.n13830 DVDD.n13829 0.00455714
R9331 DVDD.n13831 DVDD.n13830 0.00455714
R9332 DVDD.n372 DVDD.n371 0.00455714
R9333 DVDD.n371 DVDD.n370 0.00455714
R9334 DVDD.n370 DVDD.n369 0.00455714
R9335 DVDD.n369 DVDD.n368 0.00455714
R9336 DVDD.n368 DVDD.n367 0.00455714
R9337 DVDD.n367 DVDD.n366 0.00455714
R9338 DVDD.n366 DVDD.n365 0.00455714
R9339 DVDD.n365 DVDD.n364 0.00455714
R9340 DVDD.n364 DVDD.n363 0.00455714
R9341 DVDD.n363 DVDD.n362 0.00455714
R9342 DVDD.n362 DVDD.n361 0.00455714
R9343 DVDD.n361 DVDD.n360 0.00455714
R9344 DVDD.n360 DVDD.n359 0.00455714
R9345 DVDD.n359 DVDD.n358 0.00455714
R9346 DVDD.n358 DVDD.n357 0.00455714
R9347 DVDD.n357 DVDD.n356 0.00455714
R9348 DVDD.n356 DVDD.n355 0.00455714
R9349 DVDD.n355 DVDD.n354 0.00455714
R9350 DVDD.n354 DVDD.n353 0.00455714
R9351 DVDD.n353 DVDD.n352 0.00455714
R9352 DVDD.n352 DVDD.n351 0.00455714
R9353 DVDD.n351 DVDD.n350 0.00455714
R9354 DVDD.n350 DVDD.n349 0.00455714
R9355 DVDD.n349 DVDD.n348 0.00455714
R9356 DVDD.n348 DVDD.n347 0.00455714
R9357 DVDD.n347 DVDD.n346 0.00455714
R9358 DVDD.n346 DVDD.n345 0.00455714
R9359 DVDD.n345 DVDD.n344 0.00455714
R9360 DVDD.n344 DVDD.n343 0.00455714
R9361 DVDD.n343 DVDD.n342 0.00455714
R9362 DVDD.n342 DVDD.n341 0.00455714
R9363 DVDD.n341 DVDD.n340 0.00455714
R9364 DVDD.n340 DVDD.n339 0.00455714
R9365 DVDD.n339 DVDD.n338 0.00455714
R9366 DVDD.n338 DVDD.n337 0.00455714
R9367 DVDD.n337 DVDD.n336 0.00455714
R9368 DVDD.n336 DVDD.n335 0.00455714
R9369 DVDD.n335 DVDD.n334 0.00455714
R9370 DVDD.n334 DVDD.n333 0.00455714
R9371 DVDD.n333 DVDD.n332 0.00455714
R9372 DVDD.n332 DVDD.n331 0.00455714
R9373 DVDD.n331 DVDD.n330 0.00455714
R9374 DVDD.n330 DVDD.n329 0.00455714
R9375 DVDD.n329 DVDD.n328 0.00455714
R9376 DVDD.n328 DVDD.n327 0.00455714
R9377 DVDD.n327 DVDD.n326 0.00455714
R9378 DVDD.n326 DVDD.n325 0.00455714
R9379 DVDD.n325 DVDD.n324 0.00455714
R9380 DVDD.n324 DVDD.n323 0.00455714
R9381 DVDD.n323 DVDD.n322 0.00455714
R9382 DVDD.n322 DVDD.n321 0.00455714
R9383 DVDD.n321 DVDD.n320 0.00455714
R9384 DVDD.n320 DVDD.n319 0.00455714
R9385 DVDD.n319 DVDD.n318 0.00455714
R9386 DVDD.n318 DVDD.n317 0.00455714
R9387 DVDD.n317 DVDD.n316 0.00455714
R9388 DVDD.n316 DVDD.n315 0.00455714
R9389 DVDD.n315 DVDD.n314 0.00455714
R9390 DVDD.n314 DVDD.n313 0.00455714
R9391 DVDD.n313 DVDD.n312 0.00455714
R9392 DVDD.n312 DVDD.n311 0.00455714
R9393 DVDD.n311 DVDD.n310 0.00455714
R9394 DVDD.n310 DVDD.n309 0.00455714
R9395 DVDD.n309 DVDD.n308 0.00455714
R9396 DVDD.n308 DVDD.n307 0.00455714
R9397 DVDD.n307 DVDD.n306 0.00455714
R9398 DVDD.n306 DVDD.n305 0.00455714
R9399 DVDD.n2432 DVDD.n2431 0.00455714
R9400 DVDD.n2433 DVDD.n2432 0.00455714
R9401 DVDD.n2434 DVDD.n2433 0.00455714
R9402 DVDD.n2435 DVDD.n2434 0.00455714
R9403 DVDD.n2436 DVDD.n2435 0.00455714
R9404 DVDD.n2437 DVDD.n2436 0.00455714
R9405 DVDD.n2438 DVDD.n2437 0.00455714
R9406 DVDD.n2439 DVDD.n2438 0.00455714
R9407 DVDD.n2440 DVDD.n2439 0.00455714
R9408 DVDD.n2441 DVDD.n2440 0.00455714
R9409 DVDD.n2442 DVDD.n2441 0.00455714
R9410 DVDD.n2443 DVDD.n2442 0.00455714
R9411 DVDD.n2444 DVDD.n2443 0.00455714
R9412 DVDD.n2445 DVDD.n2444 0.00455714
R9413 DVDD.n2446 DVDD.n2445 0.00455714
R9414 DVDD.n2447 DVDD.n2446 0.00455714
R9415 DVDD.n2496 DVDD.n2495 0.00455714
R9416 DVDD.n2495 DVDD.n2494 0.00455714
R9417 DVDD.n2494 DVDD.n2493 0.00455714
R9418 DVDD.n2493 DVDD.n2492 0.00455714
R9419 DVDD.n2492 DVDD.n2491 0.00455714
R9420 DVDD.n2491 DVDD.n2490 0.00455714
R9421 DVDD.n2490 DVDD.n2489 0.00455714
R9422 DVDD.n2489 DVDD.n2488 0.00455714
R9423 DVDD.n2488 DVDD.n2487 0.00455714
R9424 DVDD.n603 DVDD.n602 0.00455714
R9425 DVDD.n602 DVDD.n601 0.00455714
R9426 DVDD.n601 DVDD.n600 0.00455714
R9427 DVDD.n600 DVDD.n599 0.00455714
R9428 DVDD.n599 DVDD.n598 0.00455714
R9429 DVDD.n598 DVDD.n597 0.00455714
R9430 DVDD.n597 DVDD.n596 0.00455714
R9431 DVDD.n596 DVDD.n595 0.00455714
R9432 DVDD.n595 DVDD.n594 0.00455714
R9433 DVDD.n594 DVDD.n593 0.00455714
R9434 DVDD.n593 DVDD.n592 0.00455714
R9435 DVDD.n592 DVDD.n591 0.00455714
R9436 DVDD.n591 DVDD.n590 0.00455714
R9437 DVDD.n590 DVDD.n589 0.00455714
R9438 DVDD.n589 DVDD.n588 0.00455714
R9439 DVDD.n588 DVDD.n587 0.00455714
R9440 DVDD.n587 DVDD.n586 0.00455714
R9441 DVDD.n586 DVDD.n585 0.00455714
R9442 DVDD.n585 DVDD.n584 0.00455714
R9443 DVDD.n584 DVDD.n583 0.00455714
R9444 DVDD.n583 DVDD.n582 0.00455714
R9445 DVDD.n582 DVDD.n581 0.00455714
R9446 DVDD.n581 DVDD.n580 0.00455714
R9447 DVDD.n580 DVDD.n579 0.00455714
R9448 DVDD.n579 DVDD.n578 0.00455714
R9449 DVDD.n578 DVDD.n577 0.00455714
R9450 DVDD.n577 DVDD.n576 0.00455714
R9451 DVDD.n576 DVDD.n575 0.00455714
R9452 DVDD.n575 DVDD.n574 0.00455714
R9453 DVDD.n574 DVDD.n573 0.00455714
R9454 DVDD.n573 DVDD.n572 0.00455714
R9455 DVDD.n572 DVDD.n571 0.00455714
R9456 DVDD.n571 DVDD.n570 0.00455714
R9457 DVDD.n570 DVDD.n569 0.00455714
R9458 DVDD.n569 DVDD.n568 0.00455714
R9459 DVDD.n568 DVDD.n567 0.00455714
R9460 DVDD.n567 DVDD.n566 0.00455714
R9461 DVDD.n566 DVDD.n565 0.00455714
R9462 DVDD.n565 DVDD.n564 0.00455714
R9463 DVDD.n564 DVDD.n563 0.00455714
R9464 DVDD.n563 DVDD.n562 0.00455714
R9465 DVDD.n562 DVDD.n561 0.00455714
R9466 DVDD.n561 DVDD.n560 0.00455714
R9467 DVDD.n560 DVDD.n559 0.00455714
R9468 DVDD.n559 DVDD.n558 0.00455714
R9469 DVDD.n558 DVDD.n557 0.00455714
R9470 DVDD.n557 DVDD.n556 0.00455714
R9471 DVDD.n556 DVDD.n555 0.00455714
R9472 DVDD.n555 DVDD.n554 0.00455714
R9473 DVDD.n554 DVDD.n553 0.00455714
R9474 DVDD.n553 DVDD.n552 0.00455714
R9475 DVDD.n552 DVDD.n551 0.00455714
R9476 DVDD.n551 DVDD.n550 0.00455714
R9477 DVDD.n550 DVDD.n549 0.00455714
R9478 DVDD.n549 DVDD.n548 0.00455714
R9479 DVDD.n548 DVDD.n547 0.00455714
R9480 DVDD.n547 DVDD.n546 0.00455714
R9481 DVDD.n546 DVDD.n545 0.00455714
R9482 DVDD.n545 DVDD.n544 0.00455714
R9483 DVDD.n544 DVDD.n543 0.00455714
R9484 DVDD.n543 DVDD.n542 0.00455714
R9485 DVDD.n542 DVDD.n541 0.00455714
R9486 DVDD.n541 DVDD.n540 0.00455714
R9487 DVDD.n540 DVDD.n539 0.00455714
R9488 DVDD.n539 DVDD.n538 0.00455714
R9489 DVDD.n538 DVDD.n537 0.00455714
R9490 DVDD.n537 DVDD.n536 0.00455714
R9491 DVDD.n2629 DVDD.n2628 0.00455714
R9492 DVDD.n2630 DVDD.n2629 0.00455714
R9493 DVDD.n2631 DVDD.n2630 0.00455714
R9494 DVDD.n2632 DVDD.n2631 0.00455714
R9495 DVDD.n2633 DVDD.n2632 0.00455714
R9496 DVDD.n2634 DVDD.n2633 0.00455714
R9497 DVDD.n2635 DVDD.n2634 0.00455714
R9498 DVDD.n2636 DVDD.n2635 0.00455714
R9499 DVDD.n2637 DVDD.n2636 0.00455714
R9500 DVDD.n2638 DVDD.n2637 0.00455714
R9501 DVDD.n2639 DVDD.n2638 0.00455714
R9502 DVDD.n2640 DVDD.n2639 0.00455714
R9503 DVDD.n2641 DVDD.n2640 0.00455714
R9504 DVDD.n2642 DVDD.n2641 0.00455714
R9505 DVDD.n2643 DVDD.n2642 0.00455714
R9506 DVDD.n2644 DVDD.n2643 0.00455714
R9507 DVDD.n2708 DVDD.n2707 0.00455714
R9508 DVDD.n2707 DVDD.n2706 0.00455714
R9509 DVDD.n2706 DVDD.n2705 0.00455714
R9510 DVDD.n2705 DVDD.n2704 0.00455714
R9511 DVDD.n2704 DVDD.n2703 0.00455714
R9512 DVDD.n2703 DVDD.n2702 0.00455714
R9513 DVDD.n2702 DVDD.n2701 0.00455714
R9514 DVDD.n2701 DVDD.n2700 0.00455714
R9515 DVDD.n2700 DVDD.n2699 0.00455714
R9516 DVDD.n2699 DVDD.n2651 0.00455714
R9517 DVDD.n3815 DVDD.n3814 0.00455
R9518 DVDD.n18999 DVDD.n18998 0.00455
R9519 DVDD.n7221 DVDD.n7220 0.00455
R9520 DVDD.n7120 DVDD.n7119 0.00455
R9521 DVDD.n2822 DVDD.n2821 0.00455
R9522 DVDD.n14912 DVDD.n14911 0.00455
R9523 DVDD.n14851 DVDD.n14850 0.00455
R9524 DVDD.n15080 DVDD.n15079 0.00455
R9525 DVDD.n10698 DVDD.n10697 0.00455
R9526 DVDD.n10602 DVDD.n10601 0.00455
R9527 DVDD.n3408 DVDD.n3407 0.00455
R9528 DVDD.n3605 DVDD.n3604 0.00455
R9529 DVDD.n18424 DVDD.n18423 0.00455
R9530 DVDD.n18427 DVDD.n18426 0.00455
R9531 DVDD.n18445 DVDD.n18444 0.00455
R9532 DVDD.n18442 DVDD.n18441 0.00455
R9533 DVDD.n18356 DVDD.n18351 0.00455
R9534 DVDD.n7133 DVDD.n7132 0.00455
R9535 DVDD.n14750 DVDD.n14749 0.00455
R9536 DVDD.n14771 DVDD.n14754 0.00455
R9537 DVDD.n14768 DVDD.n14767 0.00455
R9538 DVDD.n14766 DVDD.n14765 0.00455
R9539 DVDD.n14759 DVDD.n14758 0.00455
R9540 DVDD.n7292 DVDD.n7291 0.00455
R9541 DVDD.n3113 DVDD.n3112 0.00451786
R9542 DVDD.n3097 DVDD.n3096 0.00451786
R9543 DVDD.n3090 DVDD.n3089 0.00451786
R9544 DVDD.n3082 DVDD.n3081 0.00451786
R9545 DVDD.n3076 DVDD.n3075 0.00451786
R9546 DVDD.n3061 DVDD.n3060 0.00451786
R9547 DVDD.n3052 DVDD.n3051 0.00451786
R9548 DVDD.n4320 DVDD.n4319 0.00449949
R9549 DVDD.n4291 DVDD.n4290 0.00449949
R9550 DVDD.n4266 DVDD.n4265 0.00449949
R9551 DVDD.n10399 DVDD.n10398 0.00449375
R9552 DVDD.n10563 DVDD.n10562 0.00449375
R9553 DVDD.n10592 DVDD.n10591 0.00449375
R9554 DVDD.n386 DVDD.n385 0.00448571
R9555 DVDD.n617 DVDD.n616 0.00448571
R9556 DVDD.n5364 DVDD.n5363 0.00445468
R9557 DVDD.n9418 DVDD.n9417 0.00445398
R9558 DVDD.n8115 DVDD.n8114 0.00445398
R9559 DVDD.n8002 DVDD.n8001 0.00445398
R9560 DVDD.n8006 DVDD.n8005 0.00445398
R9561 DVDD.n8095 DVDD.n8094 0.00445398
R9562 DVDD DVDD.n20290 0.0044381
R9563 DVDD.n14920 DVDD.n14919 0.0044375
R9564 DVDD.n15218 DVDD.n15217 0.0044375
R9565 DVDD.n15233 DVDD.n15232 0.0044375
R9566 DVDD.n2678 DVDD.n2677 0.00442143
R9567 DVDD.n1147 DVDD.n1146 0.00439764
R9568 DVDD.n1556 DVDD.n1555 0.00439764
R9569 DVDD.n1619 DVDD.n1618 0.00439764
R9570 DVDD.n1628 DVDD.n1627 0.00439764
R9571 DVDD.n1664 DVDD.n1663 0.00439764
R9572 DVDD.n925 DVDD.n924 0.00439764
R9573 DVDD.n906 DVDD.n905 0.00439764
R9574 DVDD.n901 DVDD.n900 0.00439764
R9575 DVDD.n894 DVDD.n893 0.00439764
R9576 DVDD.n873 DVDD.n872 0.00439764
R9577 DVDD.n11472 DVDD.n11471 0.00439764
R9578 DVDD.n11988 DVDD.n11339 0.00439764
R9579 DVDD.n11995 DVDD.n11994 0.00439764
R9580 DVDD.n12019 DVDD.n12018 0.00439764
R9581 DVDD.n12045 DVDD.n12044 0.00439764
R9582 DVDD.n12052 DVDD.n12051 0.00439764
R9583 DVDD.n12085 DVDD.n12084 0.00439764
R9584 DVDD.n12111 DVDD.n12110 0.00439764
R9585 DVDD.n12118 DVDD.n12117 0.00439764
R9586 DVDD.n13393 DVDD.n13392 0.00439764
R9587 DVDD.n13398 DVDD.n13397 0.00439764
R9588 DVDD.n18476 DVDD.n18475 0.00439764
R9589 DVDD.n19692 DVDD.n19691 0.00439764
R9590 DVDD.n19081 DVDD.n19008 0.00439764
R9591 DVDD.n19078 DVDD.n19077 0.00439764
R9592 DVDD.n19075 DVDD.n19074 0.00439764
R9593 DVDD.n4803 DVDD.n4802 0.00439764
R9594 DVDD.n4929 DVDD.n4928 0.00439764
R9595 DVDD.n4997 DVDD.n4996 0.00439764
R9596 DVDD.n5180 DVDD.n5179 0.00439764
R9597 DVDD.n5432 DVDD.n5431 0.00439764
R9598 DVDD.n1337 DVDD.n1336 0.00439764
R9599 DVDD.n19463 DVDD.n19217 0.00439764
R9600 DVDD.n19460 DVDD.n19459 0.00439764
R9601 DVDD.n19457 DVDD.n19456 0.00439764
R9602 DVDD.n11629 DVDD.n11628 0.00439764
R9603 DVDD.n11828 DVDD.n11827 0.00439764
R9604 DVDD.n11824 DVDD.n11823 0.00439764
R9605 DVDD.n11756 DVDD.n11755 0.00439764
R9606 DVDD.n12360 DVDD.n12359 0.00439764
R9607 DVDD.n13031 DVDD.n13030 0.00439764
R9608 DVDD.n19172 DVDD.n19171 0.00439764
R9609 DVDD.n1914 DVDD.n1913 0.00439764
R9610 DVDD.n18973 DVDD.n18900 0.00439764
R9611 DVDD.n18970 DVDD.n18969 0.00439764
R9612 DVDD.n18967 DVDD.n18966 0.00439764
R9613 DVDD.n6881 DVDD.n6880 0.00439764
R9614 DVDD.n6759 DVDD.n6758 0.00439764
R9615 DVDD.n6755 DVDD.n6754 0.00439764
R9616 DVDD.n6687 DVDD.n6686 0.00439764
R9617 DVDD.n6502 DVDD.n6501 0.00439764
R9618 DVDD.n6329 DVDD.n6328 0.00439764
R9619 DVDD.n3266 DVDD.n3265 0.00439764
R9620 DVDD.n18810 DVDD.n18521 0.00439764
R9621 DVDD.n18807 DVDD.n18806 0.00439764
R9622 DVDD.n18804 DVDD.n18803 0.00439764
R9623 DVDD.n7885 DVDD.n7884 0.00439764
R9624 DVDD.n9727 DVDD.n9726 0.00439764
R9625 DVDD.n9723 DVDD.n9722 0.00439764
R9626 DVDD.n9655 DVDD.n9654 0.00439764
R9627 DVDD.n8381 DVDD.n8380 0.00439764
R9628 DVDD.n9115 DVDD.n9114 0.00439764
R9629 DVDD.n14919 DVDD.n14918 0.00438125
R9630 DVDD.n15217 DVDD.n15216 0.00438125
R9631 DVDD.n3812 DVDD.n3811 0.004325
R9632 DVDD.n10079 DVDD.n10078 0.004325
R9633 DVDD.n7631 DVDD.n7630 0.004325
R9634 DVDD.n3893 DVDD.n3892 0.004325
R9635 DVDD.n7123 DVDD.n7122 0.004325
R9636 DVDD.n7655 DVDD.n7654 0.004325
R9637 DVDD.n1815 DVDD.n1814 0.004325
R9638 DVDD.n3782 DVDD.n3781 0.004325
R9639 DVDD.n2825 DVDD.n2824 0.004325
R9640 DVDD.n20297 DVDD.n20296 0.004325
R9641 DVDD.n20319 DVDD.n20318 0.004325
R9642 DVDD.n14848 DVDD.n14847 0.004325
R9643 DVDD.n17024 DVDD.n17023 0.00431
R9644 DVDD.n16964 DVDD.n16963 0.00431
R9645 DVDD.n17133 DVDD.n17132 0.00431
R9646 DVDD.n17084 DVDD.n17083 0.00431
R9647 DVDD.n5451 DVDD.n5450 0.00427756
R9648 DVDD.n5634 DVDD.n5633 0.00427747
R9649 DVDD.n12803 DVDD.n12802 0.00427747
R9650 DVDD.n6183 DVDD.n6182 0.00427747
R9651 DVDD.n8885 DVDD.n8884 0.00427747
R9652 DVDD.n4982 DVDD.n4981 0.00427717
R9653 DVDD.n10398 DVDD.n10397 0.00426875
R9654 DVDD.n10394 DVDD.n10393 0.00426875
R9655 DVDD.n10593 DVDD.n10592 0.00426875
R9656 DVDD.n15977 DVDD.n15976 0.00426569
R9657 DVDD.n8256 DVDD.n8255 0.00426569
R9658 DVDD.n8178 DVDD.n8177 0.00426569
R9659 DVDD.n8176 DVDD.n8175 0.00426569
R9660 DVDD.n9437 DVDD.n9436 0.00426569
R9661 DVDD.n8120 DVDD.n8119 0.00426569
R9662 DVDD.n8066 DVDD.n8065 0.00426569
R9663 DVDD.n8070 DVDD.n8069 0.00426569
R9664 DVDD.n8096 DVDD.n8095 0.00424228
R9665 DVDD.n1151 DVDD.n1150 0.00422047
R9666 DVDD.n1552 DVDD.n1551 0.00422047
R9667 DVDD.n1572 DVDD.n1571 0.00422047
R9668 DVDD.n1668 DVDD.n1667 0.00422047
R9669 DVDD.n1647 DVDD.n864 0.00422047
R9670 DVDD.n909 DVDD.n908 0.00422047
R9671 DVDD.n904 DVDD.n903 0.00422047
R9672 DVDD.n10158 DVDD.n10157 0.00422047
R9673 DVDD.n11468 DVDD.n11467 0.00422047
R9674 DVDD.n11489 DVDD.n11488 0.00422047
R9675 DVDD.n12056 DVDD.n12055 0.00422047
R9676 DVDD.n12061 DVDD.n12060 0.00422047
R9677 DVDD.n12154 DVDD.n12153 0.00422047
R9678 DVDD.n12174 DVDD.n12173 0.00422047
R9679 DVDD.n12223 DVDD.n12222 0.00422047
R9680 DVDD.n2803 DVDD.n2802 0.00422047
R9681 DVDD.n18671 DVDD.n18670 0.00422047
R9682 DVDD.n10062 DVDD.n10061 0.00422047
R9683 DVDD.n19696 DVDD.n19695 0.00422047
R9684 DVDD.n19715 DVDD.n19714 0.00422047
R9685 DVDD.n19914 DVDD.n19913 0.00422047
R9686 DVDD.n20070 DVDD.n20069 0.00422047
R9687 DVDD.n20073 DVDD.n20072 0.00422047
R9688 DVDD.n20078 DVDD.n20077 0.00422047
R9689 DVDD.n20201 DVDD.n20200 0.00422047
R9690 DVDD.n20106 DVDD.n20105 0.00422047
R9691 DVDD.n19008 DVDD.n19007 0.00422047
R9692 DVDD.n3863 DVDD.n3862 0.00422047
R9693 DVDD.n4661 DVDD.n4660 0.00422047
R9694 DVDD.n4663 DVDD.n4662 0.00422047
R9695 DVDD.n4678 DVDD.n4677 0.00422047
R9696 DVDD.n4978 DVDD.n4977 0.00422047
R9697 DVDD.n5089 DVDD.n5088 0.00422047
R9698 DVDD.n5191 DVDD.n5190 0.00422047
R9699 DVDD.n5323 DVDD.n5322 0.00422047
R9700 DVDD.n5358 DVDD.n5357 0.00422047
R9701 DVDD.n5412 DVDD.n5411 0.00422047
R9702 DVDD.n5447 DVDD.n5446 0.00422047
R9703 DVDD.n1341 DVDD.n1340 0.00422047
R9704 DVDD.n1360 DVDD.n1359 0.00422047
R9705 DVDD.n1463 DVDD.n1462 0.00422047
R9706 DVDD.n1703 DVDD.n1702 0.00422047
R9707 DVDD.n1700 DVDD.n1699 0.00422047
R9708 DVDD.n292 DVDD.n291 0.00422047
R9709 DVDD.n279 DVDD.n278 0.00422047
R9710 DVDD.n19204 DVDD.n19203 0.00422047
R9711 DVDD.n19217 DVDD.n19216 0.00422047
R9712 DVDD.n10110 DVDD.n10109 0.00422047
R9713 DVDD.n11368 DVDD.n11367 0.00422047
R9714 DVDD.n11370 DVDD.n11369 0.00422047
R9715 DVDD.n11385 DVDD.n11384 0.00422047
R9716 DVDD.n11775 DVDD.n11774 0.00422047
R9717 DVDD.n11665 DVDD.n11664 0.00422047
R9718 DVDD.n12371 DVDD.n12370 0.00422047
R9719 DVDD.n13136 DVDD.n13135 0.00422047
R9720 DVDD.n13102 DVDD.n13101 0.00422047
R9721 DVDD.n13050 DVDD.n13049 0.00422047
R9722 DVDD.n13016 DVDD.n13015 0.00422047
R9723 DVDD.n835 DVDD.n834 0.00422047
R9724 DVDD.n150 DVDD.n149 0.00422047
R9725 DVDD.n10094 DVDD.n10093 0.00422047
R9726 DVDD.n1918 DVDD.n1917 0.00422047
R9727 DVDD.n1937 DVDD.n1936 0.00422047
R9728 DVDD.n2135 DVDD.n2134 0.00422047
R9729 DVDD.n2291 DVDD.n2290 0.00422047
R9730 DVDD.n2294 DVDD.n2293 0.00422047
R9731 DVDD.n2299 DVDD.n2298 0.00422047
R9732 DVDD.n19586 DVDD.n19585 0.00422047
R9733 DVDD.n19491 DVDD.n19490 0.00422047
R9734 DVDD.n18900 DVDD.n18899 0.00422047
R9735 DVDD.n7084 DVDD.n7083 0.00422047
R9736 DVDD.n7023 DVDD.n7022 0.00422047
R9737 DVDD.n7021 DVDD.n7020 0.00422047
R9738 DVDD.n7006 DVDD.n7005 0.00422047
R9739 DVDD.n6706 DVDD.n6705 0.00422047
R9740 DVDD.n6593 DVDD.n6592 0.00422047
R9741 DVDD.n6491 DVDD.n6490 0.00422047
R9742 DVDD.n6438 DVDD.n6437 0.00422047
R9743 DVDD.n6403 DVDD.n6402 0.00422047
R9744 DVDD.n6349 DVDD.n6348 0.00422047
R9745 DVDD.n6314 DVDD.n6313 0.00422047
R9746 DVDD.n3262 DVDD.n3261 0.00422047
R9747 DVDD.n3243 DVDD.n3242 0.00422047
R9748 DVDD.n3534 DVDD.n3533 0.00422047
R9749 DVDD.n3735 DVDD.n3734 0.00422047
R9750 DVDD.n3738 DVDD.n3737 0.00422047
R9751 DVDD.n3778 DVDD.n3777 0.00422047
R9752 DVDD.n3765 DVDD.n3764 0.00422047
R9753 DVDD.n18508 DVDD.n18507 0.00422047
R9754 DVDD.n18521 DVDD.n18520 0.00422047
R9755 DVDD.n7142 DVDD.n7141 0.00422047
R9756 DVDD.n10040 DVDD.n10039 0.00422047
R9757 DVDD.n10038 DVDD.n10037 0.00422047
R9758 DVDD.n10023 DVDD.n10022 0.00422047
R9759 DVDD.n9674 DVDD.n9673 0.00422047
R9760 DVDD.n9561 DVDD.n9560 0.00422047
R9761 DVDD.n8392 DVDD.n8391 0.00422047
R9762 DVDD.n9224 DVDD.n9223 0.00422047
R9763 DVDD.n9189 DVDD.n9188 0.00422047
R9764 DVDD.n9135 DVDD.n9134 0.00422047
R9765 DVDD.n9100 DVDD.n9099 0.00422047
R9766 DVDD.n16174 DVDD.n16173 0.00422
R9767 DVDD.n16294 DVDD.n16293 0.00422
R9768 DVDD.n11038 DVDD.n11037 0.00422
R9769 DVDD.n11095 DVDD.n11094 0.00422
R9770 DVDD.n10577 DVDD.n10576 0.0042125
R9771 DVDD.n13044 DVDD.n13043 0.00418891
R9772 DVDD.n6343 DVDD.n6342 0.00418891
R9773 DVDD.n9129 DVDD.n9128 0.00418891
R9774 DVDD.n523 DVDD.n521 0.00416429
R9775 DVDD.n481 DVDD.n479 0.00416429
R9776 DVDD.n752 DVDD.n751 0.00416429
R9777 DVDD.n713 DVDD.n711 0.00416429
R9778 DVDD.n11293 DVDD.n11292 0.00416429
R9779 DVDD.n11275 DVDD.n11274 0.00416429
R9780 DVDD.n12499 DVDD.n12498 0.00416429
R9781 DVDD.n5763 DVDD.n5761 0.00416429
R9782 DVDD.n4798 DVDD.n4797 0.00410038
R9783 DVDD.n18827 DVDD.n18826 0.0041
R9784 DVDD.n18813 DVDD.n18812 0.0041
R9785 DVDD.n19158 DVDD.n19157 0.0041
R9786 DVDD.n7268 DVDD.n7267 0.0041
R9787 DVDD.n3851 DVDD.n3850 0.0041
R9788 DVDD.n3906 DVDD.n3905 0.0041
R9789 DVDD.n136 DVDD.n135 0.0041
R9790 DVDD.n3795 DVDD.n3794 0.0041
R9791 DVDD.n15314 DVDD.n14904 0.0041
R9792 DVDD.n14875 DVDD.n14874 0.0041
R9793 DVDD.n14861 DVDD.n14860 0.0041
R9794 DVDD.n15093 DVDD.n15092 0.0041
R9795 DVDD.n10711 DVDD.n10710 0.0041
R9796 DVDD.n10620 DVDD.n10619 0.0041
R9797 DVDD.n3593 DVDD.n3592 0.0041
R9798 DVDD.n18739 DVDD.n18738 0.0041
R9799 DVDD.n18736 DVDD.n18562 0.0041
R9800 DVDD.n18691 DVDD.n18690 0.0041
R9801 DVDD.n14756 DVDD.n14755 0.0041
R9802 DVDD.n7169 DVDD.n7168 0.0041
R9803 DVDD.n7281 DVDD.n7280 0.0041
R9804 DVDD.n16065 DVDD.n16064 0.00407741
R9805 DVDD.n15677 DVDD.n15676 0.00407741
R9806 DVDD.n8193 DVDD.n8192 0.00407741
R9807 DVDD.n9404 DVDD.n9403 0.00407741
R9808 DVDD.n8358 DVDD.n8357 0.00407741
R9809 DVDD.n7943 DVDD.n7942 0.00407741
R9810 DVDD.n7951 DVDD.n7950 0.00407741
R9811 DVDD.n7959 DVDD.n7958 0.00407741
R9812 DVDD.n7975 DVDD.n7974 0.00407741
R9813 DVDD.n7984 DVDD.n7983 0.00407741
R9814 DVDD.n7999 DVDD.n7998 0.00407741
R9815 DVDD.n8007 DVDD.n8006 0.00407741
R9816 DVDD.n8015 DVDD.n8014 0.00407741
R9817 DVDD.n8023 DVDD.n8022 0.00407741
R9818 DVDD.n8039 DVDD.n8038 0.00407741
R9819 DVDD.n8048 DVDD.n8047 0.00407741
R9820 DVDD.n8063 DVDD.n8062 0.00407741
R9821 DVDD.n8071 DVDD.n8070 0.00407741
R9822 DVDD.n8079 DVDD.n8078 0.00407741
R9823 DVDD.n8087 DVDD.n8086 0.00407741
R9824 DVDD.n15149 DVDD.n15148 0.00405
R9825 DVDD.n15150 DVDD.n15149 0.00405
R9826 DVDD.n15151 DVDD.n15150 0.00405
R9827 DVDD.n15152 DVDD.n15151 0.00405
R9828 DVDD.n15153 DVDD.n15152 0.00405
R9829 DVDD.n15154 DVDD.n15153 0.00405
R9830 DVDD.n15155 DVDD.n15154 0.00405
R9831 DVDD.n15156 DVDD.n15155 0.00405
R9832 DVDD.n15157 DVDD.n15156 0.00405
R9833 DVDD.n15158 DVDD.n15157 0.00405
R9834 DVDD.n15183 DVDD.n15182 0.00405
R9835 DVDD.n15184 DVDD.n15183 0.00405
R9836 DVDD.n15185 DVDD.n15184 0.00405
R9837 DVDD.n15186 DVDD.n15185 0.00405
R9838 DVDD.n15187 DVDD.n15186 0.00405
R9839 DVDD.n15188 DVDD.n15187 0.00405
R9840 DVDD.n15189 DVDD.n15188 0.00405
R9841 DVDD.n15190 DVDD.n15189 0.00405
R9842 DVDD.n15191 DVDD.n15190 0.00405
R9843 DVDD.n10196 DVDD.n10195 0.00405
R9844 DVDD.n10197 DVDD.n10196 0.00405
R9845 DVDD.n10198 DVDD.n10197 0.00405
R9846 DVDD.n10199 DVDD.n10198 0.00405
R9847 DVDD.n10200 DVDD.n10199 0.00405
R9848 DVDD.n10201 DVDD.n10200 0.00405
R9849 DVDD.n10202 DVDD.n10201 0.00405
R9850 DVDD.n10203 DVDD.n10202 0.00405
R9851 DVDD.n10204 DVDD.n10203 0.00405
R9852 DVDD.n10205 DVDD.n10204 0.00405
R9853 DVDD.n10228 DVDD.n10227 0.00405
R9854 DVDD.n10227 DVDD.n10226 0.00405
R9855 DVDD.n10226 DVDD.n10225 0.00405
R9856 DVDD.n10225 DVDD.n10224 0.00405
R9857 DVDD.n10224 DVDD.n10223 0.00405
R9858 DVDD.n10223 DVDD.n10222 0.00405
R9859 DVDD.n10222 DVDD.n10221 0.00405
R9860 DVDD.n10221 DVDD.n10220 0.00405
R9861 DVDD.n10220 DVDD.n10219 0.00405
R9862 DVDD.n10280 DVDD.n10279 0.00405
R9863 DVDD.n10279 DVDD.n10278 0.00405
R9864 DVDD.n10278 DVDD.n10277 0.00405
R9865 DVDD.n10232 DVDD.n10231 0.00405
R9866 DVDD.n10233 DVDD.n10232 0.00405
R9867 DVDD.n10234 DVDD.n10233 0.00405
R9868 DVDD.n10235 DVDD.n10234 0.00405
R9869 DVDD.n10236 DVDD.n10235 0.00405
R9870 DVDD.n10237 DVDD.n10236 0.00405
R9871 DVDD.n10244 DVDD.n10243 0.00405
R9872 DVDD.n10243 DVDD.n10242 0.00405
R9873 DVDD.n10242 DVDD.n10241 0.00405
R9874 DVDD.n10241 DVDD.n10240 0.00405
R9875 DVDD.n10240 DVDD.n10239 0.00405
R9876 DVDD.n10239 DVDD.n10238 0.00405
R9877 DVDD.n15141 DVDD.n15140 0.00405
R9878 DVDD.n15142 DVDD.n15141 0.00405
R9879 DVDD.n10213 DVDD.n10212 0.00405
R9880 DVDD.n10212 DVDD.n10211 0.00405
R9881 DVDD.n10211 DVDD.n10210 0.00405
R9882 DVDD.n10271 DVDD.n10270 0.00405
R9883 DVDD.n10272 DVDD.n10271 0.00405
R9884 DVDD.n10273 DVDD.n10272 0.00405
R9885 DVDD.n10274 DVDD.n10273 0.00405
R9886 DVDD.n10275 DVDD.n10274 0.00405
R9887 DVDD.n10276 DVDD.n10275 0.00405
R9888 DVDD.n10291 DVDD.n10290 0.00405
R9889 DVDD.n10290 DVDD.n10289 0.00405
R9890 DVDD.n10289 DVDD.n10288 0.00405
R9891 DVDD.n10288 DVDD.n10287 0.00405
R9892 DVDD.n10287 DVDD.n10286 0.00405
R9893 DVDD.n10286 DVDD.n10285 0.00405
R9894 DVDD.n10285 DVDD.n10284 0.00405
R9895 DVDD.n10284 DVDD.n10283 0.00405
R9896 DVDD.n10283 DVDD.n10282 0.00405
R9897 DVDD.n1234 DVDD.n1233 0.00404331
R9898 DVDD.n1218 DVDD.n1217 0.00404331
R9899 DVDD.n1211 DVDD.n1210 0.00404331
R9900 DVDD.n1202 DVDD.n1201 0.00404331
R9901 DVDD.n1196 DVDD.n1195 0.00404331
R9902 DVDD.n1182 DVDD.n1181 0.00404331
R9903 DVDD.n1174 DVDD.n1173 0.00404331
R9904 DVDD.n1632 DVDD.n1631 0.00404331
R9905 DVDD.n885 DVDD.n884 0.00404331
R9906 DVDD.n877 DVDD.n876 0.00404331
R9907 DVDD.n10175 DVDD.n10174 0.00404331
R9908 DVDD.n10180 DVDD.n10179 0.00404331
R9909 DVDD.n11427 DVDD.n10183 0.00404331
R9910 DVDD.n11448 DVDD.n11447 0.00404331
R9911 DVDD.n12122 DVDD.n12121 0.00404331
R9912 DVDD.n12127 DVDD.n12126 0.00404331
R9913 DVDD.n12179 DVDD.n12178 0.00404331
R9914 DVDD.n12242 DVDD.n12241 0.00404331
R9915 DVDD.n13415 DVDD.n13414 0.00404331
R9916 DVDD.n13496 DVDD.n13495 0.00404331
R9917 DVDD.n13498 DVDD.n13497 0.00404331
R9918 DVDD.n13706 DVDD.n13705 0.00404331
R9919 DVDD.n18569 DVDD.n18568 0.00404331
R9920 DVDD.n18680 DVDD.n18679 0.00404331
R9921 DVDD.n14811 DVDD.n14810 0.00404331
R9922 DVDD.n15479 DVDD.n15478 0.00404331
R9923 DVDD.n14740 DVDD.n14739 0.00404331
R9924 DVDD.n14657 DVDD.n14656 0.00404331
R9925 DVDD.n14383 DVDD.n14382 0.00404331
R9926 DVDD.n19860 DVDD.n19859 0.00404331
R9927 DVDD.n19895 DVDD.n19894 0.00404331
R9928 DVDD.n20087 DVDD.n20086 0.00404331
R9929 DVDD.n20110 DVDD.n20109 0.00404331
R9930 DVDD.n3888 DVDD.n3887 0.00404331
R9931 DVDD.n4680 DVDD.n4679 0.00404331
R9932 DVDD.n4930 DVDD.n4929 0.00404331
R9933 DVDD.n4995 DVDD.n4994 0.00404331
R9934 DVDD.n5039 DVDD.n5038 0.00404331
R9935 DVDD.n5059 DVDD.n5058 0.00404331
R9936 DVDD.n5061 DVDD.n5060 0.00404331
R9937 DVDD.n5166 DVDD.n5165 0.00404331
R9938 DVDD.n5357 DVDD.n5356 0.00404331
R9939 DVDD.n5368 DVDD.n5367 0.00404331
R9940 DVDD.n5446 DVDD.n5445 0.00404331
R9941 DVDD.n6047 DVDD.n6046 0.00404331
R9942 DVDD.n5945 DVDD.n5944 0.00404331
R9943 DVDD.n1516 DVDD.n1515 0.00404331
R9944 DVDD.n1482 DVDD.n1481 0.00404331
R9945 DVDD.n19185 DVDD.n19184 0.00404331
R9946 DVDD.n19208 DVDD.n19207 0.00404331
R9947 DVDD.n18332 DVDD.n18331 0.00404331
R9948 DVDD.n11387 DVDD.n11386 0.00404331
R9949 DVDD.n11823 DVDD.n11822 0.00404331
R9950 DVDD.n11758 DVDD.n11757 0.00404331
R9951 DVDD.n11715 DVDD.n11714 0.00404331
R9952 DVDD.n11695 DVDD.n11694 0.00404331
R9953 DVDD.n11693 DVDD.n11692 0.00404331
R9954 DVDD.n12347 DVDD.n12346 0.00404331
R9955 DVDD.n13103 DVDD.n13102 0.00404331
R9956 DVDD.n13092 DVDD.n13091 0.00404331
R9957 DVDD.n13017 DVDD.n13016 0.00404331
R9958 DVDD.n12693 DVDD.n12692 0.00404331
R9959 DVDD.n12608 DVDD.n12607 0.00404331
R9960 DVDD.n238 DVDD.n237 0.00404331
R9961 DVDD.n159 DVDD.n158 0.00404331
R9962 DVDD.n18227 DVDD.n18226 0.00404331
R9963 DVDD.n18130 DVDD.n18129 0.00404331
R9964 DVDD.n18091 DVDD.n18090 0.00404331
R9965 DVDD.n18013 DVDD.n18012 0.00404331
R9966 DVDD.n17761 DVDD.n17760 0.00404331
R9967 DVDD.n2082 DVDD.n2081 0.00404331
R9968 DVDD.n2116 DVDD.n2115 0.00404331
R9969 DVDD.n19472 DVDD.n19471 0.00404331
R9970 DVDD.n19495 DVDD.n19494 0.00404331
R9971 DVDD.n7109 DVDD.n7108 0.00404331
R9972 DVDD.n7004 DVDD.n7003 0.00404331
R9973 DVDD.n6754 DVDD.n6753 0.00404331
R9974 DVDD.n6689 DVDD.n6688 0.00404331
R9975 DVDD.n6645 DVDD.n6644 0.00404331
R9976 DVDD.n6623 DVDD.n6622 0.00404331
R9977 DVDD.n6621 DVDD.n6620 0.00404331
R9978 DVDD.n6516 DVDD.n6515 0.00404331
R9979 DVDD.n6404 DVDD.n6403 0.00404331
R9980 DVDD.n6393 DVDD.n6392 0.00404331
R9981 DVDD.n6315 DVDD.n6314 0.00404331
R9982 DVDD.n4497 DVDD.n4496 0.00404331
R9983 DVDD.n4404 DVDD.n4403 0.00404331
R9984 DVDD.n3481 DVDD.n3480 0.00404331
R9985 DVDD.n3515 DVDD.n3514 0.00404331
R9986 DVDD.n18489 DVDD.n18488 0.00404331
R9987 DVDD.n18512 DVDD.n18511 0.00404331
R9988 DVDD.n10054 DVDD.n10053 0.00404331
R9989 DVDD.n10021 DVDD.n10020 0.00404331
R9990 DVDD.n9722 DVDD.n9721 0.00404331
R9991 DVDD.n9657 DVDD.n9656 0.00404331
R9992 DVDD.n9613 DVDD.n9612 0.00404331
R9993 DVDD.n9591 DVDD.n9590 0.00404331
R9994 DVDD.n9589 DVDD.n9588 0.00404331
R9995 DVDD.n8367 DVDD.n8366 0.00404331
R9996 DVDD.n9190 DVDD.n9189 0.00404331
R9997 DVDD.n9179 DVDD.n9178 0.00404331
R9998 DVDD.n9101 DVDD.n9100 0.00404331
R9999 DVDD.n8778 DVDD.n8777 0.00404331
R10000 DVDD.n8678 DVDD.n8677 0.00404331
R10001 DVDD.n2487 DVDD 0.00401429
R10002 DVDD.n13107 DVDD.n13106 0.00401178
R10003 DVDD.n6408 DVDD.n6407 0.00401178
R10004 DVDD.n9194 DVDD.n9193 0.00401178
R10005 DVDD.n11731 DVDD.n11730 0.00401125
R10006 DVDD.n6661 DVDD.n6660 0.00401125
R10007 DVDD.n9629 DVDD.n9628 0.00401125
R10008 DVDD.n19752 DVDD.n19751 0.00401111
R10009 DVDD.n10570 DVDD.n10569 0.0039875
R10010 DVDD.n16380 DVDD.n16379 0.00398
R10011 DVDD.n11176 DVDD.n11175 0.00398
R10012 DVDD.n20341 DVDD.n3 0.00397625
R10013 DVDD.n7475 DVDD.n7352 0.00397625
R10014 DVDD.n7674 DVDD.n7563 0.00397625
R10015 DVDD.n10194 DVDD.n10193 0.00397625
R10016 DVDD.n8084 DVDD.n8083 0.00394684
R10017 DVDD.n9474 DVDD.n9473 0.00394408
R10018 DVDD.n15243 DVDD.n15242 0.00393125
R10019 DVDD.n12924 DVDD.n12923 0.00392391
R10020 DVDD.n12943 DVDD.n12942 0.00392391
R10021 DVDD.n5508 DVDD.n5507 0.00392391
R10022 DVDD.n5534 DVDD.n5533 0.00392391
R10023 DVDD.n4006 DVDD.n4005 0.00392391
R10024 DVDD.n4029 DVDD.n4028 0.00392391
R10025 DVDD.n8962 DVDD.n8961 0.00392391
R10026 DVDD.n9031 DVDD.n9030 0.00392391
R10027 DVDD.n12911 DVDD.n12908 0.00392391
R10028 DVDD.n12884 DVDD.n12883 0.00392391
R10029 DVDD.n5712 DVDD.n5711 0.00392391
R10030 DVDD.n6039 DVDD.n6035 0.00392391
R10031 DVDD.n4083 DVDD.n4082 0.00392391
R10032 DVDD.n4490 DVDD.n4486 0.00392391
R10033 DVDD.n8989 DVDD.n8988 0.00392391
R10034 DVDD.n9018 DVDD.n9015 0.00392391
R10035 DVDD.n5317 DVDD.n5316 0.00392323
R10036 DVDD.n5407 DVDD.n5406 0.00392323
R10037 DVDD.n11724 DVDD.n11723 0.00392323
R10038 DVDD.n6654 DVDD.n6653 0.00392323
R10039 DVDD.n9622 DVDD.n9621 0.00392323
R10040 DVDD.n3086 DVDD.n3085 0.00390971
R10041 DVDD.n16035 DVDD.n16034 0.00388912
R10042 DVDD.n16016 DVDD.n16015 0.00388912
R10043 DVDD.n15647 DVDD.n15646 0.00388912
R10044 DVDD.n15628 DVDD.n15627 0.00388912
R10045 DVDD.n8150 DVDD.n8149 0.00388912
R10046 DVDD.n8360 DVDD.n8359 0.00388912
R10047 DVDD.n8351 DVDD.n8350 0.00388912
R10048 DVDD.n9484 DVDD.n8141 0.00388912
R10049 DVDD.n8046 DVDD.n8045 0.00388912
R10050 DVDD.n18826 DVDD.n18825 0.003875
R10051 DVDD.n19157 DVDD.n19156 0.003875
R10052 DVDD.n3852 DVDD.n3851 0.003875
R10053 DVDD.n7617 DVDD.n7616 0.003875
R10054 DVDD.n3907 DVDD.n3906 0.003875
R10055 DVDD.n7644 DVDD.n7643 0.003875
R10056 DVDD.n137 DVDD.n136 0.003875
R10057 DVDD.n3796 DVDD.n3795 0.003875
R10058 DVDD.n20285 DVDD.n20284 0.003875
R10059 DVDD.n20332 DVDD.n20331 0.003875
R10060 DVDD.n14874 DVDD.n14873 0.003875
R10061 DVDD.n10619 DVDD.n10618 0.003875
R10062 DVDD.n1576 DVDD.n1575 0.00386614
R10063 DVDD.n1615 DVDD.n1614 0.00386614
R10064 DVDD.n1654 DVDD.n1653 0.00386614
R10065 DVDD.n898 DVDD.n897 0.00386614
R10066 DVDD.n10172 DVDD.n10171 0.00386614
R10067 DVDD.n10177 DVDD.n10176 0.00386614
R10068 DVDD.n10182 DVDD.n10181 0.00386614
R10069 DVDD.n11444 DVDD.n11443 0.00386614
R10070 DVDD.n11996 DVDD.n11995 0.00386614
R10071 DVDD.n12005 DVDD.n12004 0.00386614
R10072 DVDD.n12014 DVDD.n12013 0.00386614
R10073 DVDD.n12030 DVDD.n12029 0.00386614
R10074 DVDD.n12039 DVDD.n12038 0.00386614
R10075 DVDD.n12053 DVDD.n12052 0.00386614
R10076 DVDD.n12062 DVDD.n12061 0.00386614
R10077 DVDD.n12071 DVDD.n12070 0.00386614
R10078 DVDD.n12080 DVDD.n12079 0.00386614
R10079 DVDD.n12096 DVDD.n12095 0.00386614
R10080 DVDD.n12105 DVDD.n12104 0.00386614
R10081 DVDD.n12119 DVDD.n12118 0.00386614
R10082 DVDD.n12128 DVDD.n12127 0.00386614
R10083 DVDD.n12137 DVDD.n12136 0.00386614
R10084 DVDD.n12146 DVDD.n12145 0.00386614
R10085 DVDD.n12155 DVDD.n12154 0.00386614
R10086 DVDD.n12209 DVDD.n12208 0.00386614
R10087 DVDD.n13307 DVDD.n13306 0.00386614
R10088 DVDD.n13481 DVDD.n13480 0.00386614
R10089 DVDD.n13546 DVDD.n13545 0.00386614
R10090 DVDD.n13627 DVDD.n13626 0.00386614
R10091 DVDD.n2739 DVDD.n2738 0.00386614
R10092 DVDD.n2780 DVDD.n2779 0.00386614
R10093 DVDD.n18578 DVDD.n18577 0.00386614
R10094 DVDD.n14802 DVDD.n14801 0.00386614
R10095 DVDD.n15391 DVDD.n15390 0.00386614
R10096 DVDD.n14712 DVDD.n14711 0.00386614
R10097 DVDD.n14629 DVDD.n14628 0.00386614
R10098 DVDD.n14575 DVDD.n14574 0.00386614
R10099 DVDD.n14487 DVDD.n14486 0.00386614
R10100 DVDD.n19716 DVDD.n19715 0.00386614
R10101 DVDD.n19739 DVDD.n19738 0.00386614
R10102 DVDD.n19747 DVDD.n19746 0.00386614
R10103 DVDD.n19882 DVDD.n19881 0.00386614
R10104 DVDD.n20005 DVDD.n20004 0.00386614
R10105 DVDD.n20205 DVDD.n20204 0.00386614
R10106 DVDD.n20104 DVDD.n20103 0.00386614
R10107 DVDD.n4657 DVDD.n4656 0.00386614
R10108 DVDD.n4791 DVDD.n4790 0.00386614
R10109 DVDD.n4793 DVDD.n4792 0.00386614
R10110 DVDD.n4899 DVDD.n4820 0.00386614
R10111 DVDD.n4902 DVDD.n4901 0.00386614
R10112 DVDD.n5034 DVDD.n5033 0.00386614
R10113 DVDD.n5213 DVDD.n5212 0.00386614
R10114 DVDD.n5308 DVDD.n5307 0.00386614
R10115 DVDD.n5398 DVDD.n5397 0.00386614
R10116 DVDD.n5658 DVDD.n5657 0.00386614
R10117 DVDD.n6083 DVDD.n6082 0.00386614
R10118 DVDD.n1361 DVDD.n1360 0.00386614
R10119 DVDD.n1365 DVDD.n1364 0.00386614
R10120 DVDD.n1384 DVDD.n1383 0.00386614
R10121 DVDD.n1392 DVDD.n1391 0.00386614
R10122 DVDD.n1495 DVDD.n1494 0.00386614
R10123 DVDD.n1693 DVDD.n1692 0.00386614
R10124 DVDD.n283 DVDD.n282 0.00386614
R10125 DVDD.n19202 DVDD.n19201 0.00386614
R10126 DVDD.n11364 DVDD.n11363 0.00386614
R10127 DVDD.n11617 DVDD.n11616 0.00386614
R10128 DVDD.n11619 DVDD.n11618 0.00386614
R10129 DVDD.n11853 DVDD.n11646 0.00386614
R10130 DVDD.n11851 DVDD.n11850 0.00386614
R10131 DVDD.n11720 DVDD.n11719 0.00386614
R10132 DVDD.n12393 DVDD.n12392 0.00386614
R10133 DVDD.n13150 DVDD.n13149 0.00386614
R10134 DVDD.n13063 DVDD.n13062 0.00386614
R10135 DVDD.n12779 DVDD.n12778 0.00386614
R10136 DVDD.n12715 DVDD.n12714 0.00386614
R10137 DVDD.n777 DVDD.n776 0.00386614
R10138 DVDD.n814 DVDD.n813 0.00386614
R10139 DVDD.n247 DVDD.n246 0.00386614
R10140 DVDD.n18236 DVDD.n18235 0.00386614
R10141 DVDD.n18209 DVDD.n18208 0.00386614
R10142 DVDD.n18065 DVDD.n18064 0.00386614
R10143 DVDD.n17987 DVDD.n17986 0.00386614
R10144 DVDD.n17935 DVDD.n17934 0.00386614
R10145 DVDD.n17854 DVDD.n17853 0.00386614
R10146 DVDD.n1938 DVDD.n1937 0.00386614
R10147 DVDD.n1942 DVDD.n1941 0.00386614
R10148 DVDD.n1961 DVDD.n1960 0.00386614
R10149 DVDD.n1969 DVDD.n1968 0.00386614
R10150 DVDD.n2103 DVDD.n2102 0.00386614
R10151 DVDD.n2226 DVDD.n2225 0.00386614
R10152 DVDD.n19590 DVDD.n19589 0.00386614
R10153 DVDD.n19489 DVDD.n19488 0.00386614
R10154 DVDD.n7027 DVDD.n7026 0.00386614
R10155 DVDD.n6893 DVDD.n6892 0.00386614
R10156 DVDD.n6891 DVDD.n6890 0.00386614
R10157 DVDD.n6863 DVDD.n6862 0.00386614
R10158 DVDD.n6782 DVDD.n6781 0.00386614
R10159 DVDD.n6650 DVDD.n6649 0.00386614
R10160 DVDD.n6469 DVDD.n6468 0.00386614
R10161 DVDD.n6453 DVDD.n6452 0.00386614
R10162 DVDD.n6363 DVDD.n6362 0.00386614
R10163 DVDD.n6156 DVDD.n6155 0.00386614
R10164 DVDD.n4533 DVDD.n4532 0.00386614
R10165 DVDD.n3242 DVDD.n3241 0.00386614
R10166 DVDD.n3238 DVDD.n3237 0.00386614
R10167 DVDD.n3219 DVDD.n3218 0.00386614
R10168 DVDD.n3211 DVDD.n3210 0.00386614
R10169 DVDD.n3502 DVDD.n3501 0.00386614
R10170 DVDD.n3556 DVDD.n3555 0.00386614
R10171 DVDD.n3769 DVDD.n3768 0.00386614
R10172 DVDD.n18506 DVDD.n18505 0.00386614
R10173 DVDD.n10044 DVDD.n10043 0.00386614
R10174 DVDD.n7873 DVDD.n7872 0.00386614
R10175 DVDD.n7875 DVDD.n7874 0.00386614
R10176 DVDD.n9752 DVDD.n7902 0.00386614
R10177 DVDD.n9750 DVDD.n9749 0.00386614
R10178 DVDD.n9618 DVDD.n9617 0.00386614
R10179 DVDD.n8414 DVDD.n8413 0.00386614
R10180 DVDD.n9239 DVDD.n9238 0.00386614
R10181 DVDD.n9149 DVDD.n9148 0.00386614
R10182 DVDD.n8858 DVDD.n8857 0.00386614
R10183 DVDD.n8800 DVDD.n8799 0.00386614
R10184 DVDD.n8020 DVDD.n8019 0.00385277
R10185 DVDD.n12375 DVDD.n12374 0.00383447
R10186 DVDD.n6487 DVDD.n6486 0.00383447
R10187 DVDD.n8396 DVDD.n8395 0.00383447
R10188 DVDD.n19919 DVDD.n19918 0.0038338
R10189 DVDD.n15014 DVDD.n15013 0.0038
R10190 DVDD.n14982 DVDD.n14981 0.0038
R10191 DVDD.n11041 DVDD.n11040 0.0038
R10192 DVDD.n16236 DVDD.n16233 0.0038
R10193 DVDD.n15816 DVDD.n15814 0.0038
R10194 DVDD.n15537 DVDD.n15536 0.0038
R10195 DVDD.n16235 DVDD.n16234 0.0038
R10196 DVDD.n11043 DVDD.n11042 0.0038
R10197 DVDD.n18333 DVDD 0.00376574
R10198 DVDD.n7662 DVDD 0.00376574
R10199 DVDD.n20215 DVDD 0.00376574
R10200 DVDD.n20338 DVDD 0.00376574
R10201 DVDD.n7956 DVDD.n7955 0.00375871
R10202 DVDD.n8291 DVDD.n8290 0.00375845
R10203 DVDD.n5194 DVDD.n5193 0.00374585
R10204 DVDD.n5333 DVDD.n5332 0.00374514
R10205 DVDD.n4952 DVDD.n4951 0.00374497
R10206 DVDD.n17266 DVDD.n17265 0.00374324
R10207 DVDD.n17295 DVDD.n17294 0.00374324
R10208 DVDD.n17644 DVDD.n17643 0.00374324
R10209 DVDD.n17674 DVDD.n17673 0.00374324
R10210 DVDD.n2675 DVDD.n2674 0.00371429
R10211 DVDD.n3093 DVDD.n3092 0.00371429
R10212 DVDD.n15287 DVDD.n15192 0.00370171
R10213 DVDD.n20342 DVDD.n20341 0.00370171
R10214 DVDD.n7475 DVDD.n7204 0.00370171
R10215 DVDD.n16046 DVDD.n16045 0.00370084
R10216 DVDD.n16005 DVDD.n16004 0.00370084
R10217 DVDD.n15658 DVDD.n15657 0.00370084
R10218 DVDD.n15927 DVDD.n15926 0.00370084
R10219 DVDD.n8161 DVDD.n8160 0.00370084
R10220 DVDD.n8343 DVDD.n8342 0.00370084
R10221 DVDD.n7982 DVDD.n7981 0.00370084
R10222 DVDD.n10219 DVDD.n10218 0.0037
R10223 DVDD.n1599 DVDD.n1598 0.00368898
R10224 DVDD.n916 DVDD.n915 0.00368898
R10225 DVDD.n11436 DVDD.n11435 0.00368898
R10226 DVDD.n12103 DVDD.n12102 0.00368898
R10227 DVDD.n12196 DVDD.n12195 0.00368898
R10228 DVDD.n12289 DVDD.n12199 0.00368898
R10229 DVDD.n12279 DVDD.n12278 0.00368898
R10230 DVDD.n13305 DVDD.n13304 0.00368898
R10231 DVDD.n13314 DVDD.n13313 0.00368898
R10232 DVDD.n13522 DVDD.n13521 0.00368898
R10233 DVDD.n13574 DVDD.n13573 0.00368898
R10234 DVDD.n13590 DVDD.n13589 0.00368898
R10235 DVDD.n13655 DVDD.n13654 0.00368898
R10236 DVDD.n13671 DVDD.n13670 0.00368898
R10237 DVDD.n18574 DVDD.n18573 0.00368898
R10238 DVDD.n14806 DVDD.n14805 0.00368898
R10239 DVDD.n15421 DVDD.n15420 0.00368898
R10240 DVDD.n15440 DVDD.n15439 0.00368898
R10241 DVDD.n14682 DVDD.n14681 0.00368898
R10242 DVDD.n14599 DVDD.n14598 0.00368898
R10243 DVDD.n14545 DVDD.n14544 0.00368898
R10244 DVDD.n14526 DVDD.n14525 0.00368898
R10245 DVDD.n14457 DVDD.n14456 0.00368898
R10246 DVDD.n14423 DVDD.n14422 0.00368898
R10247 DVDD.n19729 DVDD.n19728 0.00368898
R10248 DVDD.n20199 DVDD.n20198 0.00368898
R10249 DVDD.n20195 DVDD.n20194 0.00368898
R10250 DVDD.n20188 DVDD.n20187 0.00368898
R10251 DVDD.n20182 DVDD.n20181 0.00368898
R10252 DVDD.n4667 DVDD.n4666 0.00368898
R10253 DVDD.n4813 DVDD.n4812 0.00368898
R10254 DVDD.n4904 DVDD.n4903 0.00368898
R10255 DVDD.n4962 DVDD.n4961 0.00368898
R10256 DVDD.n4979 DVDD.n4978 0.00368898
R10257 DVDD.n5025 DVDD.n5024 0.00368898
R10258 DVDD.n5455 DVDD.n5454 0.00368898
R10259 DVDD.n5488 DVDD.n5487 0.00368898
R10260 DVDD.n5651 DVDD.n5650 0.00368898
R10261 DVDD.n5674 DVDD.n5673 0.00368898
R10262 DVDD.n6025 DVDD.n6024 0.00368898
R10263 DVDD.n5981 DVDD.n5980 0.00368898
R10264 DVDD.n1374 DVDD.n1373 0.00368898
R10265 DVDD.n1379 DVDD.n1378 0.00368898
R10266 DVDD.n277 DVDD.n276 0.00368898
R10267 DVDD.n273 DVDD.n272 0.00368898
R10268 DVDD.n266 DVDD.n265 0.00368898
R10269 DVDD.n260 DVDD.n259 0.00368898
R10270 DVDD.n11374 DVDD.n11373 0.00368898
R10271 DVDD.n11639 DVDD.n11638 0.00368898
R10272 DVDD.n11849 DVDD.n11848 0.00368898
R10273 DVDD.n11791 DVDD.n11790 0.00368898
R10274 DVDD.n11774 DVDD.n11773 0.00368898
R10275 DVDD.n11729 DVDD.n11728 0.00368898
R10276 DVDD.n13012 DVDD.n13011 0.00368898
R10277 DVDD.n13008 DVDD.n13007 0.00368898
R10278 DVDD.n12975 DVDD.n12974 0.00368898
R10279 DVDD.n12786 DVDD.n12785 0.00368898
R10280 DVDD.n12767 DVDD.n12766 0.00368898
R10281 DVDD.n12676 DVDD.n12675 0.00368898
R10282 DVDD.n12644 DVDD.n12643 0.00368898
R10283 DVDD.n243 DVDD.n242 0.00368898
R10284 DVDD.n18232 DVDD.n18231 0.00368898
R10285 DVDD.n18181 DVDD.n18180 0.00368898
R10286 DVDD.n18165 DVDD.n18164 0.00368898
R10287 DVDD.n18037 DVDD.n18036 0.00368898
R10288 DVDD.n17959 DVDD.n17958 0.00368898
R10289 DVDD.n17907 DVDD.n17906 0.00368898
R10290 DVDD.n17891 DVDD.n17890 0.00368898
R10291 DVDD.n17826 DVDD.n17825 0.00368898
R10292 DVDD.n17797 DVDD.n17796 0.00368898
R10293 DVDD.n1951 DVDD.n1950 0.00368898
R10294 DVDD.n1956 DVDD.n1955 0.00368898
R10295 DVDD.n19584 DVDD.n19583 0.00368898
R10296 DVDD.n19580 DVDD.n19579 0.00368898
R10297 DVDD.n19573 DVDD.n19572 0.00368898
R10298 DVDD.n19567 DVDD.n19566 0.00368898
R10299 DVDD.n7017 DVDD.n7016 0.00368898
R10300 DVDD.n6871 DVDD.n6870 0.00368898
R10301 DVDD.n6780 DVDD.n6779 0.00368898
R10302 DVDD.n6722 DVDD.n6721 0.00368898
R10303 DVDD.n6705 DVDD.n6704 0.00368898
R10304 DVDD.n6659 DVDD.n6658 0.00368898
R10305 DVDD.n6310 DVDD.n6309 0.00368898
R10306 DVDD.n6306 DVDD.n6305 0.00368898
R10307 DVDD.n6271 DVDD.n6270 0.00368898
R10308 DVDD.n6163 DVDD.n6162 0.00368898
R10309 DVDD.n6150 DVDD.n6149 0.00368898
R10310 DVDD.n4476 DVDD.n4475 0.00368898
R10311 DVDD.n4444 DVDD.n4443 0.00368898
R10312 DVDD.n3229 DVDD.n3228 0.00368898
R10313 DVDD.n3224 DVDD.n3223 0.00368898
R10314 DVDD.n3763 DVDD.n3762 0.00368898
R10315 DVDD.n3759 DVDD.n3758 0.00368898
R10316 DVDD.n3752 DVDD.n3751 0.00368898
R10317 DVDD.n3746 DVDD.n3745 0.00368898
R10318 DVDD.n10034 DVDD.n10033 0.00368898
R10319 DVDD.n7895 DVDD.n7894 0.00368898
R10320 DVDD.n9748 DVDD.n9747 0.00368898
R10321 DVDD.n9690 DVDD.n9689 0.00368898
R10322 DVDD.n9673 DVDD.n9672 0.00368898
R10323 DVDD.n9627 DVDD.n9626 0.00368898
R10324 DVDD.n9096 DVDD.n9095 0.00368898
R10325 DVDD.n9092 DVDD.n9091 0.00368898
R10326 DVDD.n9057 DVDD.n9056 0.00368898
R10327 DVDD.n8865 DVDD.n8864 0.00368898
R10328 DVDD.n8852 DVDD.n8851 0.00368898
R10329 DVDD.n8762 DVDD.n8761 0.00368898
R10330 DVDD.n8718 DVDD.n8717 0.00368898
R10331 DVDD.n8228 DVDD.n8227 0.0036644
R10332 DVDD.n4549 DVDD.n4548 0.00365742
R10333 DVDD.n8816 DVDD.n8815 0.00365742
R10334 DVDD.n6186 DVDD.n6185 0.00365731
R10335 DVDD.n8888 DVDD.n8887 0.00365731
R10336 DVDD.n6108 DVDD.n6107 0.00365678
R10337 DVDD.n12739 DVDD.n12738 0.00365678
R10338 DVDD.n6121 DVDD.n6120 0.00365678
R10339 DVDD.n8823 DVDD.n8822 0.00365678
R10340 DVDD.n2472 DVDD.n2471 0.00365
R10341 DVDD.n16534 DVDD.n16533 0.00365
R10342 DVDD.n16703 DVDD.n16702 0.00365
R10343 DVDD.n16829 DVDD.n16828 0.00365
R10344 DVDD.n16875 DVDD.n16874 0.00365
R10345 DVDD.n11114 DVDD.n11113 0.00365
R10346 DVDD.n16485 DVDD.n16484 0.00365
R10347 DVDD.n17130 DVDD.n17129 0.00365
R10348 DVDD.n17081 DVDD.n17080 0.00365
R10349 DVDD.n11092 DVDD.n11091 0.00365
R10350 DVDD.n3665 DVDD.n3664 0.00365
R10351 DVDD.n3658 DVDD.n3657 0.00365
R10352 DVDD.n3655 DVDD.n3654 0.00365
R10353 DVDD.n3652 DVDD.n3651 0.00365
R10354 DVDD.n3603 DVDD.n3602 0.00365
R10355 DVDD.n3596 DVDD.n3595 0.00365
R10356 DVDD.n3590 DVDD.n3589 0.00365
R10357 DVDD.n18585 DVDD.n18582 0.00365
R10358 DVDD.n18600 DVDD.n18596 0.00365
R10359 DVDD.n18615 DVDD.n18611 0.00365
R10360 DVDD.n18614 DVDD.n18613 0.00365
R10361 DVDD.n18631 DVDD.n18627 0.00365
R10362 DVDD.n18648 DVDD.n18641 0.00365
R10363 DVDD.n18738 DVDD.n18737 0.00365
R10364 DVDD.n18690 DVDD.n18689 0.00365
R10365 DVDD.n18695 DVDD.n18694 0.00365
R10366 DVDD.n18345 DVDD.n18344 0.00365
R10367 DVDD.n16025 DVDD.n16024 0.00363444
R10368 DVDD.n16026 DVDD.n16025 0.00363444
R10369 DVDD.n15637 DVDD.n15636 0.00363444
R10370 DVDD.n15638 DVDD.n15637 0.00363444
R10371 DVDD DVDD.n20342 0.00361633
R10372 DVDD.n20341 DVDD.n6 0.00360545
R10373 DVDD.n7475 DVDD.n7349 0.00360545
R10374 DVDD.n7674 DVDD.n7560 0.00360545
R10375 DVDD.n10194 DVDD.n10190 0.00360545
R10376 DVDD.n14883 DVDD.n14882 0.00359375
R10377 DVDD.n15105 DVDD.n15104 0.00359375
R10378 DVDD.n389 DVDD.n388 0.00358571
R10379 DVDD.n390 DVDD.n389 0.00358571
R10380 DVDD.n620 DVDD.n619 0.00358571
R10381 DVDD.n621 DVDD.n620 0.00358571
R10382 DVDD.n12460 DVDD.n12459 0.00358566
R10383 DVDD.n12774 DVDD.n12770 0.00358566
R10384 DVDD.n12429 DVDD.n12428 0.00358566
R10385 DVDD.n12410 DVDD.n12409 0.00358566
R10386 DVDD.n8493 DVDD.n8492 0.00358546
R10387 DVDD.n8478 DVDD.n8477 0.00358546
R10388 DVDD.n8460 DVDD.n8459 0.00358546
R10389 DVDD.n8442 DVDD.n8441 0.00358546
R10390 DVDD.n5184 DVDD.n5183 0.00356885
R10391 DVDD.n5586 DVDD.n5585 0.00356881
R10392 DVDD.n12841 DVDD.n12840 0.00356881
R10393 DVDD.n6221 DVDD.n6220 0.00356881
R10394 DVDD.n8923 DVDD.n8922 0.00356881
R10395 DVDD.n10484 DVDD.n10462 0.00356
R10396 DVDD.n10451 DVDD.n10450 0.00356
R10397 DVDD.n17079 DVDD.n17078 0.00356
R10398 DVDD.n16966 DVDD.n16965 0.00356
R10399 DVDD.n16921 DVDD.n16920 0.00356
R10400 DVDD.n16620 DVDD.n16619 0.00356
R10401 DVDD.n16969 DVDD.n16968 0.00356
R10402 DVDD.n17085 DVDD.n17084 0.00356
R10403 DVDD.n16055 DVDD.n16054 0.00354041
R10404 DVDD.n15996 DVDD.n15995 0.00354041
R10405 DVDD.n15995 DVDD.n15994 0.00354041
R10406 DVDD.n16056 DVDD.n16055 0.00354041
R10407 DVDD.n15667 DVDD.n15666 0.00354041
R10408 DVDD.n15937 DVDD.n15936 0.00354041
R10409 DVDD.n15668 DVDD.n15667 0.00354041
R10410 DVDD.n15936 DVDD.n15935 0.00354041
R10411 DVDD.n1587 DVDD.n1586 0.00353694
R10412 DVDD.n13038 DVDD.n13037 0.00353694
R10413 DVDD.n13113 DVDD.n13112 0.00353693
R10414 DVDD.n1636 DVDD.n1635 0.00353669
R10415 DVDD.n1595 DVDD.n1594 0.00353669
R10416 DVDD.n11751 DVDD.n11750 0.00353669
R10417 DVDD.n1580 DVDD.n1579 0.00353663
R10418 DVDD.n435 DVDD.n433 0.00352143
R10419 DVDD.n667 DVDD.n665 0.00352143
R10420 DVDD.n15946 DVDD.n15945 0.00351255
R10421 DVDD.n15686 DVDD.n15685 0.00351255
R10422 DVDD.n8185 DVDD.n8184 0.00351255
R10423 DVDD.n9413 DVDD.n9412 0.00351255
R10424 DVDD.n8318 DVDD.n8317 0.00351255
R10425 DVDD.n8314 DVDD.n8313 0.00351255
R10426 DVDD.n9896 DVDD.n9895 0.00351255
R10427 DVDD.n918 DVDD.n917 0.00351181
R10428 DVDD.n19314 DVDD.n19313 0.00351181
R10429 DVDD.n11434 DVDD.n11433 0.00351181
R10430 DVDD.n12037 DVDD.n12036 0.00351181
R10431 DVDD.n13322 DVDD.n13321 0.00351181
R10432 DVDD.n13511 DVDD.n13510 0.00351181
R10433 DVDD.n13563 DVDD.n13562 0.00351181
R10434 DVDD.n13601 DVDD.n13600 0.00351181
R10435 DVDD.n13644 DVDD.n13643 0.00351181
R10436 DVDD.n13682 DVDD.n13681 0.00351181
R10437 DVDD.n2798 DVDD.n2797 0.00351181
R10438 DVDD.n18676 DVDD.n18675 0.00351181
R10439 DVDD.n10057 DVDD.n10056 0.00351181
R10440 DVDD.n15410 DVDD.n15409 0.00351181
R10441 DVDD.n15451 DVDD.n15450 0.00351181
R10442 DVDD.n14693 DVDD.n14692 0.00351181
R10443 DVDD.n14610 DVDD.n14609 0.00351181
R10444 DVDD.n14556 DVDD.n14555 0.00351181
R10445 DVDD.n14515 DVDD.n14514 0.00351181
R10446 DVDD.n14468 DVDD.n14467 0.00351181
R10447 DVDD.n14411 DVDD.n14410 0.00351181
R10448 DVDD.n19690 DVDD.n19689 0.00351181
R10449 DVDD.n19744 DVDD.n19743 0.00351181
R10450 DVDD.n19864 DVDD.n19863 0.00351181
R10451 DVDD.n19872 DVDD.n19871 0.00351181
R10452 DVDD.n19883 DVDD.n19882 0.00351181
R10453 DVDD.n19896 DVDD.n19895 0.00351181
R10454 DVDD.n19905 DVDD.n19904 0.00351181
R10455 DVDD.n20192 DVDD.n20191 0.00351181
R10456 DVDD.n20097 DVDD.n20096 0.00351181
R10457 DVDD.n20100 DVDD.n20099 0.00351181
R10458 DVDD.n19016 DVDD.n19015 0.00351181
R10459 DVDD.n3887 DVDD.n3886 0.00351181
R10460 DVDD.n4654 DVDD.n4653 0.00351181
R10461 DVDD.n4808 DVDD.n4807 0.00351181
R10462 DVDD.n4908 DVDD.n4907 0.00351181
R10463 DVDD.n4991 DVDD.n4990 0.00351181
R10464 DVDD.n5026 DVDD.n5025 0.00351181
R10465 DVDD.n5367 DVDD.n5366 0.00351181
R10466 DVDD.n5377 DVDD.n5376 0.00351181
R10467 DVDD.n5396 DVDD.n5395 0.00351181
R10468 DVDD.n5477 DVDD.n5476 0.00351181
R10469 DVDD.n5600 DVDD.n5599 0.00351181
R10470 DVDD.n5612 DVDD.n5611 0.00351181
R10471 DVDD.n5685 DVDD.n5684 0.00351181
R10472 DVDD.n5969 DVDD.n5968 0.00351181
R10473 DVDD.n1335 DVDD.n1334 0.00351181
R10474 DVDD.n1389 DVDD.n1388 0.00351181
R10475 DVDD.n1512 DVDD.n1511 0.00351181
R10476 DVDD.n1504 DVDD.n1503 0.00351181
R10477 DVDD.n1494 DVDD.n1493 0.00351181
R10478 DVDD.n1490 DVDD.n1489 0.00351181
R10479 DVDD.n1481 DVDD.n1480 0.00351181
R10480 DVDD.n1472 DVDD.n1471 0.00351181
R10481 DVDD.n270 DVDD.n269 0.00351181
R10482 DVDD.n19195 DVDD.n19194 0.00351181
R10483 DVDD.n19198 DVDD.n19197 0.00351181
R10484 DVDD.n19225 DVDD.n19224 0.00351181
R10485 DVDD.n10105 DVDD.n10104 0.00351181
R10486 DVDD.n18331 DVDD.n10123 0.00351181
R10487 DVDD.n11361 DVDD.n11360 0.00351181
R10488 DVDD.n11634 DVDD.n11633 0.00351181
R10489 DVDD.n11845 DVDD.n11844 0.00351181
R10490 DVDD.n11762 DVDD.n11761 0.00351181
R10491 DVDD.n11728 DVDD.n11727 0.00351181
R10492 DVDD.n13093 DVDD.n13092 0.00351181
R10493 DVDD.n13065 DVDD.n13064 0.00351181
R10494 DVDD.n12986 DVDD.n12985 0.00351181
R10495 DVDD.n12827 DVDD.n12826 0.00351181
R10496 DVDD.n12815 DVDD.n12814 0.00351181
R10497 DVDD.n12756 DVDD.n12755 0.00351181
R10498 DVDD.n12632 DVDD.n12631 0.00351181
R10499 DVDD.n830 DVDD.n829 0.00351181
R10500 DVDD.n155 DVDD.n154 0.00351181
R10501 DVDD.n10089 DVDD.n10088 0.00351181
R10502 DVDD.n18192 DVDD.n18191 0.00351181
R10503 DVDD.n18154 DVDD.n18153 0.00351181
R10504 DVDD.n18048 DVDD.n18047 0.00351181
R10505 DVDD.n17970 DVDD.n17969 0.00351181
R10506 DVDD.n17918 DVDD.n17917 0.00351181
R10507 DVDD.n17880 DVDD.n17879 0.00351181
R10508 DVDD.n17837 DVDD.n17836 0.00351181
R10509 DVDD.n17785 DVDD.n17784 0.00351181
R10510 DVDD.n1912 DVDD.n1911 0.00351181
R10511 DVDD.n1966 DVDD.n1965 0.00351181
R10512 DVDD.n2086 DVDD.n2085 0.00351181
R10513 DVDD.n2094 DVDD.n2093 0.00351181
R10514 DVDD.n2104 DVDD.n2103 0.00351181
R10515 DVDD.n2108 DVDD.n2107 0.00351181
R10516 DVDD.n2117 DVDD.n2116 0.00351181
R10517 DVDD.n2126 DVDD.n2125 0.00351181
R10518 DVDD.n19577 DVDD.n19576 0.00351181
R10519 DVDD.n19482 DVDD.n19481 0.00351181
R10520 DVDD.n19485 DVDD.n19484 0.00351181
R10521 DVDD.n18943 DVDD.n18942 0.00351181
R10522 DVDD.n7079 DVDD.n7078 0.00351181
R10523 DVDD.n7108 DVDD.n7107 0.00351181
R10524 DVDD.n7030 DVDD.n7029 0.00351181
R10525 DVDD.n6876 DVDD.n6875 0.00351181
R10526 DVDD.n6776 DVDD.n6775 0.00351181
R10527 DVDD.n6693 DVDD.n6692 0.00351181
R10528 DVDD.n6658 DVDD.n6657 0.00351181
R10529 DVDD.n6394 DVDD.n6393 0.00351181
R10530 DVDD.n6365 DVDD.n6364 0.00351181
R10531 DVDD.n6282 DVDD.n6281 0.00351181
R10532 DVDD.n6205 DVDD.n6204 0.00351181
R10533 DVDD.n6194 DVDD.n6193 0.00351181
R10534 DVDD.n6140 DVDD.n6139 0.00351181
R10535 DVDD.n4432 DVDD.n4431 0.00351181
R10536 DVDD.n3268 DVDD.n3267 0.00351181
R10537 DVDD.n3214 DVDD.n3213 0.00351181
R10538 DVDD.n3485 DVDD.n3484 0.00351181
R10539 DVDD.n3493 DVDD.n3492 0.00351181
R10540 DVDD.n3503 DVDD.n3502 0.00351181
R10541 DVDD.n3507 DVDD.n3506 0.00351181
R10542 DVDD.n3516 DVDD.n3515 0.00351181
R10543 DVDD.n3525 DVDD.n3524 0.00351181
R10544 DVDD.n3756 DVDD.n3755 0.00351181
R10545 DVDD.n18499 DVDD.n18498 0.00351181
R10546 DVDD.n18502 DVDD.n18501 0.00351181
R10547 DVDD.n18529 DVDD.n18528 0.00351181
R10548 DVDD.n7137 DVDD.n7136 0.00351181
R10549 DVDD.n10053 DVDD.n10052 0.00351181
R10550 DVDD.n10047 DVDD.n10046 0.00351181
R10551 DVDD.n7890 DVDD.n7889 0.00351181
R10552 DVDD.n9744 DVDD.n9743 0.00351181
R10553 DVDD.n9661 DVDD.n9660 0.00351181
R10554 DVDD.n9626 DVDD.n9625 0.00351181
R10555 DVDD.n9180 DVDD.n9179 0.00351181
R10556 DVDD.n9151 DVDD.n9150 0.00351181
R10557 DVDD.n9068 DVDD.n9067 0.00351181
R10558 DVDD.n8907 DVDD.n8906 0.00351181
R10559 DVDD.n8896 DVDD.n8895 0.00351181
R10560 DVDD.n8842 DVDD.n8841 0.00351181
R10561 DVDD.n8706 DVDD.n8705 0.00351181
R10562 DVDD.n10282 DVDD.n10281 0.0035
R10563 DVDD.n4495 DVDD.n4494 0.00348025
R10564 DVDD.n8776 DVDD.n8775 0.00348025
R10565 DVDD.n13582 DVDD.n13581 0.00347895
R10566 DVDD.n13663 DVDD.n13662 0.00347895
R10567 DVDD.n15431 DVDD.n15430 0.00347895
R10568 DVDD.n14535 DVDD.n14534 0.00347895
R10569 DVDD.n14536 DVDD.n14535 0.00347895
R10570 DVDD.n15430 DVDD.n15429 0.00347895
R10571 DVDD.n5991 DVDD.n5990 0.00347895
R10572 DVDD.n5643 DVDD.n5642 0.00347895
R10573 DVDD.n5992 DVDD.n5991 0.00347895
R10574 DVDD.n12654 DVDD.n12653 0.00347895
R10575 DVDD.n12655 DVDD.n12654 0.00347895
R10576 DVDD.n12794 DVDD.n12793 0.00347895
R10577 DVDD.n17807 DVDD.n17806 0.00347895
R10578 DVDD.n17808 DVDD.n17807 0.00347895
R10579 DVDD.n18173 DVDD.n18172 0.00347895
R10580 DVDD.n17899 DVDD.n17898 0.00347895
R10581 DVDD.n6172 DVDD.n6171 0.00347895
R10582 DVDD.n4455 DVDD.n4454 0.00347895
R10583 DVDD.n6173 DVDD.n6172 0.00347895
R10584 DVDD.n4454 DVDD.n4453 0.00347895
R10585 DVDD.n8874 DVDD.n8873 0.00347895
R10586 DVDD.n8728 DVDD.n8727 0.00347895
R10587 DVDD.n8875 DVDD.n8874 0.00347895
R10588 DVDD.n8729 DVDD.n8728 0.00347895
R10589 DVDD.n8308 DVDD.n8307 0.00347627
R10590 DVDD.n3412 DVDD.n3411 0.00347364
R10591 DVDD.n10367 DVDD.n10366 0.00347
R10592 DVDD.n10450 DVDD.n10449 0.00347
R10593 DVDD.n16517 DVDD.n16516 0.00347
R10594 DVDD.n17078 DVDD.n17077 0.00347
R10595 DVDD.n16859 DVDD.n16858 0.00347
R10596 DVDD.n16726 DVDD.n16725 0.00347
R10597 DVDD.n16557 DVDD.n16556 0.00347
R10598 DVDD.n15182 DVDD.n15181 0.00345
R10599 DVDD.n15986 DVDD.n15985 0.00344637
R10600 DVDD.n15987 DVDD.n15986 0.00344637
R10601 DVDD.n9425 DVDD.n9424 0.00344637
R10602 DVDD.n9426 DVDD.n9425 0.00344637
R10603 DVDD.n8107 DVDD.n8106 0.00344637
R10604 DVDD.n8106 DVDD.n8105 0.00344637
R10605 DVDD.n12923 DVDD.n12920 0.00343478
R10606 DVDD.n12942 DVDD.n12941 0.00343478
R10607 DVDD.n5507 DVDD.n5504 0.00343478
R10608 DVDD.n5533 DVDD.n5530 0.00343478
R10609 DVDD.n4005 DVDD.n4002 0.00343478
R10610 DVDD.n4028 DVDD.n4025 0.00343478
R10611 DVDD.n8961 DVDD.n8958 0.00343478
R10612 DVDD.n9030 DVDD.n9027 0.00343478
R10613 DVDD.n12912 DVDD.n12911 0.00343478
R10614 DVDD.n12883 DVDD.n12882 0.00343478
R10615 DVDD.n5711 DVDD.n5708 0.00343478
R10616 DVDD.n6039 DVDD.n6036 0.00343478
R10617 DVDD.n4082 DVDD.n4079 0.00343478
R10618 DVDD.n4490 DVDD.n4489 0.00343478
R10619 DVDD.n8988 DVDD.n8985 0.00343478
R10620 DVDD.n9019 DVDD.n9018 0.00343478
R10621 DVDD.n18825 DVDD.n18824 0.003425
R10622 DVDD.n3853 DVDD.n3852 0.003425
R10623 DVDD.n7618 DVDD.n7617 0.003425
R10624 DVDD.n3908 DVDD.n3907 0.003425
R10625 DVDD.n7645 DVDD.n7644 0.003425
R10626 DVDD.n138 DVDD.n137 0.003425
R10627 DVDD.n3797 DVDD.n3796 0.003425
R10628 DVDD.n20286 DVDD.n20285 0.003425
R10629 DVDD.n20333 DVDD.n20332 0.003425
R10630 DVDD.n14873 DVDD.n14872 0.003425
R10631 DVDD.n11205 DVDD.n11204 0.00340256
R10632 DVDD.n11206 DVDD.n11205 0.00340256
R10633 DVDD.n14332 DVDD.n14331 0.00340256
R10634 DVDD.n14333 DVDD.n14332 0.00340256
R10635 DVDD.n4967 DVDD.n4966 0.00339159
R10636 DVDD.n5417 DVDD.n5416 0.00339134
R10637 DVDD.n13095 DVDD.n13094 0.00339123
R10638 DVDD.n6396 DVDD.n6395 0.00339123
R10639 DVDD.n9182 DVDD.n9181 0.00339123
R10640 DVDD.n5438 DVDD.n5437 0.00339081
R10641 DVDD.n13609 DVDD.n13608 0.00339046
R10642 DVDD.n13690 DVDD.n13689 0.00339046
R10643 DVDD.n13555 DVDD.n13554 0.00339046
R10644 DVDD.n13636 DVDD.n13635 0.00339046
R10645 DVDD.n2749 DVDD.n2748 0.00339046
R10646 DVDD.n2790 DVDD.n2789 0.00339046
R10647 DVDD.n15401 DVDD.n15400 0.00339046
R10648 DVDD.n15461 DVDD.n15460 0.00339046
R10649 DVDD.n14702 DVDD.n14701 0.00339046
R10650 DVDD.n14619 DVDD.n14618 0.00339046
R10651 DVDD.n14565 DVDD.n14564 0.00339046
R10652 DVDD.n14505 DVDD.n14504 0.00339046
R10653 DVDD.n14477 DVDD.n14476 0.00339046
R10654 DVDD.n14402 DVDD.n14401 0.00339046
R10655 DVDD.n14401 DVDD.n14400 0.00339046
R10656 DVDD.n14478 DVDD.n14477 0.00339046
R10657 DVDD.n14566 DVDD.n14565 0.00339046
R10658 DVDD.n14620 DVDD.n14619 0.00339046
R10659 DVDD.n15400 DVDD.n15399 0.00339046
R10660 DVDD.n2789 DVDD.n2788 0.00339046
R10661 DVDD.n15460 DVDD.n15459 0.00339046
R10662 DVDD.n2748 DVDD.n2747 0.00339046
R10663 DVDD.n14506 DVDD.n14505 0.00339046
R10664 DVDD.n14703 DVDD.n14702 0.00339046
R10665 DVDD.n5223 DVDD.n5222 0.00339046
R10666 DVDD.n5693 DVDD.n5692 0.00339046
R10667 DVDD.n6073 DVDD.n6072 0.00339046
R10668 DVDD.n5592 DVDD.n5591 0.00339046
R10669 DVDD.n6074 DVDD.n6073 0.00339046
R10670 DVDD.n5961 DVDD.n5960 0.00339046
R10671 DVDD.n5469 DVDD.n5468 0.00339046
R10672 DVDD.n5222 DVDD.n5221 0.00339046
R10673 DVDD.n12403 DVDD.n12402 0.00339046
R10674 DVDD.n12748 DVDD.n12747 0.00339046
R10675 DVDD.n12705 DVDD.n12704 0.00339046
R10676 DVDD.n12994 DVDD.n12993 0.00339046
R10677 DVDD.n12706 DVDD.n12705 0.00339046
R10678 DVDD.n12835 DVDD.n12834 0.00339046
R10679 DVDD.n12624 DVDD.n12623 0.00339046
R10680 DVDD.n12402 DVDD.n12401 0.00339046
R10681 DVDD.n18146 DVDD.n18145 0.00339046
R10682 DVDD.n17872 DVDD.n17871 0.00339046
R10683 DVDD.n17777 DVDD.n17776 0.00339046
R10684 DVDD.n17978 DVDD.n17977 0.00339046
R10685 DVDD.n18200 DVDD.n18199 0.00339046
R10686 DVDD.n823 DVDD.n822 0.00339046
R10687 DVDD.n786 DVDD.n785 0.00339046
R10688 DVDD.n17926 DVDD.n17925 0.00339046
R10689 DVDD.n17845 DVDD.n17844 0.00339046
R10690 DVDD.n18056 DVDD.n18055 0.00339046
R10691 DVDD.n6459 DVDD.n6458 0.00339046
R10692 DVDD.n6291 DVDD.n6290 0.00339046
R10693 DVDD.n6214 DVDD.n6213 0.00339046
R10694 DVDD.n6130 DVDD.n6129 0.00339046
R10695 DVDD.n4523 DVDD.n4522 0.00339046
R10696 DVDD.n4422 DVDD.n4421 0.00339046
R10697 DVDD.n6292 DVDD.n6291 0.00339046
R10698 DVDD.n6215 DVDD.n6214 0.00339046
R10699 DVDD.n4524 DVDD.n4523 0.00339046
R10700 DVDD.n6131 DVDD.n6130 0.00339046
R10701 DVDD.n4423 DVDD.n4422 0.00339046
R10702 DVDD.n6460 DVDD.n6459 0.00339046
R10703 DVDD.n8423 DVDD.n8422 0.00339046
R10704 DVDD.n9077 DVDD.n9076 0.00339046
R10705 DVDD.n8916 DVDD.n8915 0.00339046
R10706 DVDD.n8832 DVDD.n8831 0.00339046
R10707 DVDD.n8790 DVDD.n8789 0.00339046
R10708 DVDD.n8697 DVDD.n8696 0.00339046
R10709 DVDD.n9078 DVDD.n9077 0.00339046
R10710 DVDD.n8917 DVDD.n8916 0.00339046
R10711 DVDD.n8791 DVDD.n8790 0.00339046
R10712 DVDD.n8696 DVDD.n8695 0.00339046
R10713 DVDD.n8833 DVDD.n8832 0.00339046
R10714 DVDD.n8424 DVDD.n8423 0.00339046
R10715 DVDD.n15340 DVDD 0.00338
R10716 DVDD.n14980 DVDD.n14979 0.00338
R10717 DVDD.n15377 DVDD.n15376 0.00338
R10718 DVDD.n11039 DVDD.n11034 0.00338
R10719 DVDD.n11186 DVDD.n11185 0.00338
R10720 DVDD.n16335 DVDD.n16333 0.00338
R10721 DVDD.n15730 DVDD.n15729 0.00338
R10722 DVDD.n16089 DVDD.n16088 0.00338
R10723 DVDD DVDD.n15913 0.00338
R10724 DVDD.n15697 DVDD 0.00338
R10725 DVDD.n16350 DVDD 0.00338
R10726 DVDD.n11145 DVDD 0.00338
R10727 DVDD.n7674 DVDD.n7665 0.00336019
R10728 DVDD.n1185 DVDD.n1184 0.00335984
R10729 DVDD.n1237 DVDD.n1236 0.0033597
R10730 DVDD.n13083 DVDD.n13082 0.0033597
R10731 DVDD.n1177 DVDD.n1176 0.00335966
R10732 DVDD.n15958 DVDD.n15957 0.00335233
R10733 DVDD.n15959 DVDD.n15958 0.00335233
R10734 DVDD.n8171 DVDD.n8170 0.00335233
R10735 DVDD.n8170 DVDD.n8169 0.00335233
R10736 DVDD.n16965 DVDD.n16960 0.00335
R10737 DVDD.n16797 DVDD.n16796 0.00335
R10738 DVDD.n16920 DVDD.n16919 0.00335
R10739 DVDD.n16676 DVDD.n16674 0.00335
R10740 DVDD.n16619 DVDD.n16617 0.00335
R10741 DVDD.n13912 DVDD.n13911 0.00333784
R10742 DVDD.n13918 DVDD.n13917 0.00333784
R10743 DVDD.n14301 DVDD.n14300 0.00333784
R10744 DVDD.n14307 DVDD.n14306 0.00333784
R10745 DVDD.n1214 DVDD.n1213 0.00333465
R10746 DVDD.n1656 DVDD.n1655 0.00333465
R10747 DVDD.n881 DVDD.n880 0.00333465
R10748 DVDD.n19269 DVDD.n19268 0.00333465
R10749 DVDD.n19276 DVDD.n19275 0.00333465
R10750 DVDD.n19283 DVDD.n19282 0.00333465
R10751 DVDD.n19290 DVDD.n19289 0.00333465
R10752 DVDD.n19295 DVDD.n19294 0.00333465
R10753 DVDD.n19300 DVDD.n19299 0.00333465
R10754 DVDD.n19307 DVDD.n19306 0.00333465
R10755 DVDD.n19339 DVDD.n19338 0.00333465
R10756 DVDD.n19332 DVDD.n19331 0.00333465
R10757 DVDD.n19325 DVDD.n19324 0.00333465
R10758 DVDD.n10162 DVDD.n10161 0.00333465
R10759 DVDD.n10164 DVDD.n10163 0.00333465
R10760 DVDD.n11480 DVDD.n11479 0.00333465
R10761 DVDD.n12218 DVDD.n12217 0.00333465
R10762 DVDD.n13348 DVDD.n13347 0.00333465
R10763 DVDD.n13353 DVDD.n13352 0.00333465
R10764 DVDD.n13489 DVDD.n13488 0.00333465
R10765 DVDD.n13537 DVDD.n13536 0.00333465
R10766 DVDD.n13618 DVDD.n13617 0.00333465
R10767 DVDD.n2730 DVDD.n2729 0.00333465
R10768 DVDD.n2771 DVDD.n2770 0.00333465
R10769 DVDD.n2807 DVDD.n2806 0.00333465
R10770 DVDD.n18471 DVDD.n18470 0.00333465
R10771 DVDD.n10066 DVDD.n10065 0.00333465
R10772 DVDD.n14820 DVDD.n14819 0.00333465
R10773 DVDD.n14721 DVDD.n14720 0.00333465
R10774 DVDD.n14638 DVDD.n14637 0.00333465
R10775 DVDD.n14584 DVDD.n14583 0.00333465
R10776 DVDD.n14496 DVDD.n14495 0.00333465
R10777 DVDD.n19741 DVDD.n19740 0.00333465
R10778 DVDD.n19757 DVDD.n19756 0.00333465
R10779 DVDD.n20210 DVDD.n20209 0.00333465
R10780 DVDD.n20089 DVDD.n20088 0.00333465
R10781 DVDD.n20093 DVDD.n20092 0.00333465
R10782 DVDD.n3867 DVDD.n3866 0.00333465
R10783 DVDD.n4610 DVDD.n4601 0.00333465
R10784 DVDD.n4784 DVDD.n4783 0.00333465
R10785 DVDD.n4802 DVDD.n4801 0.00333465
R10786 DVDD.n4912 DVDD.n4911 0.00333465
R10787 DVDD.n4954 DVDD.n4953 0.00333465
R10788 DVDD.n4988 DVDD.n4987 0.00333465
R10789 DVDD.n5097 DVDD.n5096 0.00333465
R10790 DVDD.n5204 DVDD.n5203 0.00333465
R10791 DVDD.n5313 DVDD.n5312 0.00333465
R10792 DVDD.n5331 DVDD.n5330 0.00333465
R10793 DVDD.n5390 DVDD.n5389 0.00333465
R10794 DVDD.n5404 DVDD.n5403 0.00333465
R10795 DVDD.n5422 DVDD.n5421 0.00333465
R10796 DVDD.n5551 DVDD.n5550 0.00333465
R10797 DVDD.n5678 DVDD.n5677 0.00333465
R10798 DVDD.n1386 DVDD.n1385 0.00333465
R10799 DVDD.n1402 DVDD.n1401 0.00333465
R10800 DVDD.n1498 DVDD.n1497 0.00333465
R10801 DVDD.n1477 DVDD.n1476 0.00333465
R10802 DVDD.n288 DVDD.n287 0.00333465
R10803 DVDD.n19187 DVDD.n19186 0.00333465
R10804 DVDD.n19191 DVDD.n19190 0.00333465
R10805 DVDD.n10114 DVDD.n10113 0.00333465
R10806 DVDD.n11358 DVDD.n11357 0.00333465
R10807 DVDD.n11610 DVDD.n11609 0.00333465
R10808 DVDD.n11624 DVDD.n11623 0.00333465
R10809 DVDD.n11628 DVDD.n11627 0.00333465
R10810 DVDD.n11841 DVDD.n11840 0.00333465
R10811 DVDD.n11799 DVDD.n11798 0.00333465
R10812 DVDD.n11765 DVDD.n11764 0.00333465
R10813 DVDD.n11657 DVDD.n11656 0.00333465
R10814 DVDD.n12384 DVDD.n12383 0.00333465
R10815 DVDD.n13145 DVDD.n13144 0.00333465
R10816 DVDD.n13141 DVDD.n13140 0.00333465
R10817 DVDD.n13128 DVDD.n13127 0.00333465
R10818 DVDD.n13071 DVDD.n13070 0.00333465
R10819 DVDD.n13058 DVDD.n13057 0.00333465
R10820 DVDD.n13040 DVDD.n13039 0.00333465
R10821 DVDD.n12866 DVDD.n12865 0.00333465
R10822 DVDD.n12763 DVDD.n12762 0.00333465
R10823 DVDD.n768 DVDD.n767 0.00333465
R10824 DVDD.n805 DVDD.n804 0.00333465
R10825 DVDD.n839 DVDD.n838 0.00333465
R10826 DVDD.n19167 DVDD.n19166 0.00333465
R10827 DVDD.n10098 DVDD.n10097 0.00333465
R10828 DVDD.n18218 DVDD.n18217 0.00333465
R10829 DVDD.n18074 DVDD.n18073 0.00333465
R10830 DVDD.n17996 DVDD.n17995 0.00333465
R10831 DVDD.n17944 DVDD.n17943 0.00333465
R10832 DVDD.n17863 DVDD.n17862 0.00333465
R10833 DVDD.n1963 DVDD.n1962 0.00333465
R10834 DVDD.n1979 DVDD.n1978 0.00333465
R10835 DVDD.n2100 DVDD.n2099 0.00333465
R10836 DVDD.n2121 DVDD.n2120 0.00333465
R10837 DVDD.n19595 DVDD.n19594 0.00333465
R10838 DVDD.n19474 DVDD.n19473 0.00333465
R10839 DVDD.n19478 DVDD.n19477 0.00333465
R10840 DVDD.n7088 DVDD.n7087 0.00333465
R10841 DVDD.n7073 DVDD.n3922 0.00333465
R10842 DVDD.n6900 DVDD.n6899 0.00333465
R10843 DVDD.n6886 DVDD.n6885 0.00333465
R10844 DVDD.n6882 DVDD.n6881 0.00333465
R10845 DVDD.n6772 DVDD.n6771 0.00333465
R10846 DVDD.n6730 DVDD.n6729 0.00333465
R10847 DVDD.n6696 DVDD.n6695 0.00333465
R10848 DVDD.n6585 DVDD.n6584 0.00333465
R10849 DVDD.n6478 DVDD.n6477 0.00333465
R10850 DVDD.n6448 DVDD.n6447 0.00333465
R10851 DVDD.n6444 DVDD.n6443 0.00333465
R10852 DVDD.n6430 DVDD.n6429 0.00333465
R10853 DVDD.n6371 DVDD.n6370 0.00333465
R10854 DVDD.n6357 DVDD.n6356 0.00333465
R10855 DVDD.n6339 DVDD.n6338 0.00333465
R10856 DVDD.n6245 DVDD.n6244 0.00333465
R10857 DVDD.n6147 DVDD.n6146 0.00333465
R10858 DVDD.n3217 DVDD.n3216 0.00333465
R10859 DVDD.n3201 DVDD.n3200 0.00333465
R10860 DVDD.n3499 DVDD.n3498 0.00333465
R10861 DVDD.n3520 DVDD.n3519 0.00333465
R10862 DVDD.n3774 DVDD.n3773 0.00333465
R10863 DVDD.n18491 DVDD.n18490 0.00333465
R10864 DVDD.n18495 DVDD.n18494 0.00333465
R10865 DVDD.n7146 DVDD.n7145 0.00333465
R10866 DVDD.n10050 DVDD.n10049 0.00333465
R10867 DVDD.n7866 DVDD.n7865 0.00333465
R10868 DVDD.n7880 DVDD.n7879 0.00333465
R10869 DVDD.n7884 DVDD.n7883 0.00333465
R10870 DVDD.n9740 DVDD.n9739 0.00333465
R10871 DVDD.n9698 DVDD.n9697 0.00333465
R10872 DVDD.n9664 DVDD.n9663 0.00333465
R10873 DVDD.n9553 DVDD.n9552 0.00333465
R10874 DVDD.n8405 DVDD.n8404 0.00333465
R10875 DVDD.n9234 DVDD.n9233 0.00333465
R10876 DVDD.n9230 DVDD.n9229 0.00333465
R10877 DVDD.n9216 DVDD.n9215 0.00333465
R10878 DVDD.n9157 DVDD.n9156 0.00333465
R10879 DVDD.n9143 DVDD.n9142 0.00333465
R10880 DVDD.n9125 DVDD.n9124 0.00333465
R10881 DVDD.n8947 DVDD.n8946 0.00333465
R10882 DVDD.n8849 DVDD.n8848 0.00333465
R10883 DVDD.n15968 DVDD.n15967 0.00332427
R10884 DVDD.n8248 DVDD.n8247 0.00332427
R10885 DVDD.n9449 DVDD.n9448 0.00332427
R10886 DVDD.n8129 DVDD.n8128 0.00332427
R10887 DVDD.n9887 DVDD.n7814 0.00332427
R10888 DVDD.n7938 DVDD.n7937 0.00332427
R10889 DVDD.n7993 DVDD.n7992 0.00332427
R10890 DVDD.n10523 DVDD.n10521 0.00332
R10891 DVDD.n17134 DVDD.n17128 0.00332
R10892 DVDD.n17025 DVDD.n17020 0.00332
R10893 DVDD.n15240 DVDD.n15239 0.0033125
R10894 DVDD.n3099 DVDD.n3098 0.0033125
R10895 DVDD.n3070 DVDD.n3069 0.0033125
R10896 DVDD.n17175 DVDD.n17174 0.00330651
R10897 DVDD.n17698 DVDD.n17697 0.00330651
R10898 DVDD.n17174 DVDD.n17173 0.00330651
R10899 DVDD.n17697 DVDD.n17696 0.00330651
R10900 DVDD.n12166 DVDD.n12165 0.00330197
R10901 DVDD.n12230 DVDD.n12229 0.00330197
R10902 DVDD.n13697 DVDD.n13696 0.00330197
R10903 DVDD.n12165 DVDD.n12164 0.00330197
R10904 DVDD.n12231 DVDD.n12230 0.00330197
R10905 DVDD.n2720 DVDD.n2719 0.00330197
R10906 DVDD.n2762 DVDD.n2761 0.00330197
R10907 DVDD.n15470 DVDD.n15469 0.00330197
R10908 DVDD.n14730 DVDD.n14729 0.00330197
R10909 DVDD.n14647 DVDD.n14646 0.00330197
R10910 DVDD.n14392 DVDD.n14391 0.00330197
R10911 DVDD.n14648 DVDD.n14647 0.00330197
R10912 DVDD.n14731 DVDD.n14730 0.00330197
R10913 DVDD.n2761 DVDD.n2760 0.00330197
R10914 DVDD.n15469 DVDD.n15468 0.00330197
R10915 DVDD.n2721 DVDD.n2720 0.00330197
R10916 DVDD.n5954 DVDD.n5953 0.00330197
R10917 DVDD.n12617 DVDD.n12616 0.00330197
R10918 DVDD.n18139 DVDD.n18138 0.00330197
R10919 DVDD.n17770 DVDD.n17769 0.00330197
R10920 DVDD.n18004 DVDD.n18003 0.00330197
R10921 DVDD.n18082 DVDD.n18081 0.00330197
R10922 DVDD.n797 DVDD.n796 0.00330197
R10923 DVDD.n760 DVDD.n759 0.00330197
R10924 DVDD.n4413 DVDD.n4412 0.00330197
R10925 DVDD.n14393 DVDD.n14392 0.00330197
R10926 DVDD.n4414 DVDD.n4413 0.00330197
R10927 DVDD.n8687 DVDD.n8686 0.00330197
R10928 DVDD.n8688 DVDD.n8687 0.00330197
R10929 DVDD.n15147 DVDD.n15142 0.0033
R10930 DVDD.n14105 DVDD.n14104 0.00327279
R10931 DVDD.n14106 DVDD.n14105 0.00327279
R10932 DVDD.n14015 DVDD.n14014 0.00327279
R10933 DVDD.n14016 DVDD.n14015 0.00327279
R10934 DVDD.n14227 DVDD.n14226 0.00327279
R10935 DVDD.n14228 DVDD.n14227 0.00327279
R10936 DVDD.n11120 DVDD.n11119 0.00326
R10937 DVDD.n8235 DVDD.n8234 0.00325828
R10938 DVDD.n8234 DVDD.n8233 0.00325828
R10939 DVDD.n10245 DVDD.n10244 0.00325
R10940 DVDD.n16175 DVDD.n16170 0.00323
R10941 DVDD.n16231 DVDD.n16229 0.00323
R10942 DVDD.n15596 DVDD.n15594 0.00323
R10943 DVDD.n15813 DVDD.n15810 0.00323
R10944 DVDD.n15875 DVDD.n15873 0.00323
R10945 DVDD.n13503 DVDD.n13502 0.00321348
R10946 DVDD.n13714 DVDD.n13713 0.00321348
R10947 DVDD.n15498 DVDD.n15497 0.00321348
R10948 DVDD.n14364 DVDD.n14363 0.00321348
R10949 DVDD.n15497 DVDD.n15496 0.00321348
R10950 DVDD.n5056 DVDD.n5055 0.00321348
R10951 DVDD.n5859 DVDD.n5858 0.00321348
R10952 DVDD.n5853 DVDD.n5852 0.00321348
R10953 DVDD.n5842 DVDD.n5841 0.00321348
R10954 DVDD.n5836 DVDD.n5835 0.00321348
R10955 DVDD.n5825 DVDD.n5824 0.00321348
R10956 DVDD.n5819 DVDD.n5818 0.00321348
R10957 DVDD.n5388 DVDD.n5387 0.00321348
R10958 DVDD.n4951 DVDD.n4950 0.00321348
R10959 DVDD.n5108 DVDD.n5107 0.00321348
R10960 DVDD.n11698 DVDD.n11697 0.00321348
R10961 DVDD.n12557 DVDD.n12556 0.00321348
R10962 DVDD.n12551 DVDD.n12550 0.00321348
R10963 DVDD.n12540 DVDD.n12539 0.00321348
R10964 DVDD.n12534 DVDD.n12533 0.00321348
R10965 DVDD.n12523 DVDD.n12522 0.00321348
R10966 DVDD.n12517 DVDD.n12516 0.00321348
R10967 DVDD.n13073 DVDD.n13072 0.00321348
R10968 DVDD.n11647 DVDD.n11304 0.00321348
R10969 DVDD.n18113 DVDD.n18112 0.00321348
R10970 DVDD.n17744 DVDD.n17743 0.00321348
R10971 DVDD.n5837 DVDD.n5836 0.00321348
R10972 DVDD.n12535 DVDD.n12534 0.00321348
R10973 DVDD.n5820 DVDD.n5819 0.00321348
R10974 DVDD.n12518 DVDD.n12517 0.00321348
R10975 DVDD.n12524 DVDD.n12523 0.00321348
R10976 DVDD.n5826 DVDD.n5825 0.00321348
R10977 DVDD.n12541 DVDD.n12540 0.00321348
R10978 DVDD.n5843 DVDD.n5842 0.00321348
R10979 DVDD.n12558 DVDD.n12557 0.00321348
R10980 DVDD.n5860 DVDD.n5859 0.00321348
R10981 DVDD.n5854 DVDD.n5853 0.00321348
R10982 DVDD.n12552 DVDD.n12551 0.00321348
R10983 DVDD.n6626 DVDD.n6625 0.00321348
R10984 DVDD.n4385 DVDD.n4384 0.00321348
R10985 DVDD.n4299 DVDD.n4298 0.00321348
R10986 DVDD.n4274 DVDD.n4273 0.00321348
R10987 DVDD.n4249 DVDD.n4248 0.00321348
R10988 DVDD.n4250 DVDD.n4249 0.00321348
R10989 DVDD.n4275 DVDD.n4274 0.00321348
R10990 DVDD.n4300 DVDD.n4299 0.00321348
R10991 DVDD.n6373 DVDD.n6372 0.00321348
R10992 DVDD.n6627 DVDD.n6626 0.00321348
R10993 DVDD.n6574 DVDD.n6573 0.00321348
R10994 DVDD.n14365 DVDD.n14364 0.00321348
R10995 DVDD.n4386 DVDD.n4385 0.00321348
R10996 DVDD.n12591 DVDD.n12590 0.00321348
R10997 DVDD.n5928 DVDD.n5927 0.00321348
R10998 DVDD.n9594 DVDD.n9593 0.00321348
R10999 DVDD.n8659 DVDD.n8658 0.00321348
R11000 DVDD.n8601 DVDD.n8600 0.00321348
R11001 DVDD.n8595 DVDD.n8594 0.00321348
R11002 DVDD.n8584 DVDD.n8583 0.00321348
R11003 DVDD.n8578 DVDD.n8577 0.00321348
R11004 DVDD.n8567 DVDD.n8566 0.00321348
R11005 DVDD.n8561 DVDD.n8560 0.00321348
R11006 DVDD.n8596 DVDD.n8595 0.00321348
R11007 DVDD.n8585 DVDD.n8584 0.00321348
R11008 DVDD.n8579 DVDD.n8578 0.00321348
R11009 DVDD.n8568 DVDD.n8567 0.00321348
R11010 DVDD.n8562 DVDD.n8561 0.00321348
R11011 DVDD.n8602 DVDD.n8601 0.00321348
R11012 DVDD.n8660 DVDD.n8659 0.00321348
R11013 DVDD.n9159 DVDD.n9158 0.00321348
R11014 DVDD.n9595 DVDD.n9594 0.00321348
R11015 DVDD.n9542 DVDD.n9541 0.00321348
R11016 DVDD.n18828 DVDD.n18827 0.0032
R11017 DVDD.n18812 DVDD.n18811 0.0032
R11018 DVDD.n19159 DVDD.n19158 0.0032
R11019 DVDD.n7269 DVDD.n7268 0.0032
R11020 DVDD.n3905 DVDD.n3904 0.0032
R11021 DVDD.n3794 DVDD.n3793 0.0032
R11022 DVDD.n14876 DVDD.n14875 0.0032
R11023 DVDD.n14860 DVDD.n14859 0.0032
R11024 DVDD.n15094 DVDD.n15093 0.0032
R11025 DVDD.n10730 DVDD.n10684 0.0032
R11026 DVDD.n10712 DVDD.n10711 0.0032
R11027 DVDD.n10621 DVDD.n10620 0.0032
R11028 DVDD.n10573 DVDD.n10572 0.0032
R11029 DVDD.n10574 DVDD.n10573 0.0032
R11030 DVDD.n10654 DVDD.n10593 0.0032
R11031 DVDD.n3400 DVDD.n3399 0.0032
R11032 DVDD.n3663 DVDD.n3662 0.0032
R11033 DVDD.n18629 DVDD.n18628 0.0032
R11034 DVDD.n18444 DVDD.n18443 0.0032
R11035 DVDD.n14751 DVDD.n14750 0.0032
R11036 DVDD.n14771 DVDD.n14770 0.0032
R11037 DVDD.n14765 DVDD.n14764 0.0032
R11038 DVDD.n14758 DVDD.n14757 0.0032
R11039 DVDD.n7692 DVDD.n7691 0.0032
R11040 DVDD.n7282 DVDD.n7281 0.0032
R11041 DVDD.n15059 DVDD.n15057 0.00317
R11042 DVDD.n11096 DVDD.n11090 0.00317
R11043 DVDD.n16295 DVDD.n16290 0.00317
R11044 DVDD.n10805 DVDD.n10769 0.00316667
R11045 DVDD.n10887 DVDD.n10862 0.00316667
R11046 DVDD.n10837 DVDD.n10805 0.00316667
R11047 DVDD.n10912 DVDD.n10887 0.00316667
R11048 DVDD.n16415 DVDD.n10987 0.00316667
R11049 DVDD.n16440 DVDD.n10912 0.00316667
R11050 DVDD.n16465 DVDD.n10837 0.00316667
R11051 DVDD.n16390 DVDD.n16389 0.00316667
R11052 DVDD.n16389 DVDD.n10989 0.00316667
R11053 DVDD.n10987 DVDD.n10986 0.00316667
R11054 DVDD.n10986 DVDD.n10961 0.00316667
R11055 DVDD.n15894 DVDD.n10989 0.00316667
R11056 DVDD.n1592 DVDD.n1591 0.00315748
R11057 DVDD.n1650 DVDD.n1649 0.00315748
R11058 DVDD.n887 DVDD.n886 0.00315748
R11059 DVDD.n19272 DVDD.n19271 0.00315748
R11060 DVDD.n19279 DVDD.n19278 0.00315748
R11061 DVDD.n19292 DVDD.n19291 0.00315748
R11062 DVDD.n19297 DVDD.n19296 0.00315748
R11063 DVDD.n19303 DVDD.n19302 0.00315748
R11064 DVDD.n19309 DVDD.n19308 0.00315748
R11065 DVDD.n19329 DVDD.n19328 0.00315748
R11066 DVDD.n19322 DVDD.n19321 0.00315748
R11067 DVDD.n19318 DVDD.n19317 0.00315748
R11068 DVDD.n11989 DVDD.n11988 0.00315748
R11069 DVDD.n11991 DVDD.n11990 0.00315748
R11070 DVDD.n12047 DVDD.n12046 0.00315748
R11071 DVDD.n12188 DVDD.n12187 0.00315748
R11072 DVDD.n12254 DVDD.n12253 0.00315748
R11073 DVDD.n13423 DVDD.n13422 0.00315748
R11074 DVDD.n13722 DVDD.n13721 0.00315748
R11075 DVDD.n18480 DVDD.n18479 0.00315748
R11076 DVDD.n15488 DVDD.n15487 0.00315748
R11077 DVDD.n15511 DVDD.n15510 0.00315748
R11078 DVDD.n14666 DVDD.n14665 0.00315748
R11079 DVDD.n14374 DVDD.n14373 0.00315748
R11080 DVDD.n19704 DVDD.n19703 0.00315748
R11081 DVDD.n19730 DVDD.n19729 0.00315748
R11082 DVDD.n19858 DVDD.n19857 0.00315748
R11083 DVDD.n19874 DVDD.n19873 0.00315748
R11084 DVDD.n20062 DVDD.n20061 0.00315748
R11085 DVDD.n20184 DVDD.n20183 0.00315748
R11086 DVDD.n19067 DVDD.n19066 0.00315748
R11087 DVDD.n4913 DVDD.n4912 0.00315748
R11088 DVDD.n5048 DVDD.n5047 0.00315748
R11089 DVDD.n5095 DVDD.n5094 0.00315748
R11090 DVDD.n5174 DVDD.n5173 0.00315748
R11091 DVDD.n5225 DVDD.n5224 0.00315748
R11092 DVDD.n5373 DVDD.n5372 0.00315748
R11093 DVDD.n5430 DVDD.n5429 0.00315748
R11094 DVDD.n5560 DVDD.n5559 0.00315748
R11095 DVDD.n5564 DVDD.n5563 0.00315748
R11096 DVDD.n5565 DVDD.n5564 0.00315748
R11097 DVDD.n5936 DVDD.n5935 0.00315748
R11098 DVDD.n1349 DVDD.n1348 0.00315748
R11099 DVDD.n1375 DVDD.n1374 0.00315748
R11100 DVDD.n1518 DVDD.n1517 0.00315748
R11101 DVDD.n1502 DVDD.n1501 0.00315748
R11102 DVDD.n1711 DVDD.n1710 0.00315748
R11103 DVDD.n262 DVDD.n261 0.00315748
R11104 DVDD.n19449 DVDD.n19448 0.00315748
R11105 DVDD.n11840 DVDD.n11839 0.00315748
R11106 DVDD.n11836 DVDD.n11835 0.00315748
R11107 DVDD.n11770 DVDD.n11769 0.00315748
R11108 DVDD.n11706 DVDD.n11705 0.00315748
R11109 DVDD.n11659 DVDD.n11658 0.00315748
R11110 DVDD.n12355 DVDD.n12354 0.00315748
R11111 DVDD.n12405 DVDD.n12404 0.00315748
R11112 DVDD.n13087 DVDD.n13086 0.00315748
R11113 DVDD.n13033 DVDD.n13032 0.00315748
R11114 DVDD.n12857 DVDD.n12856 0.00315748
R11115 DVDD.n12853 DVDD.n12852 0.00315748
R11116 DVDD.n12852 DVDD.n12851 0.00315748
R11117 DVDD.n12599 DVDD.n12598 0.00315748
R11118 DVDD.n19176 DVDD.n19175 0.00315748
R11119 DVDD.n18121 DVDD.n18120 0.00315748
R11120 DVDD.n18100 DVDD.n18099 0.00315748
R11121 DVDD.n18022 DVDD.n18021 0.00315748
R11122 DVDD.n17752 DVDD.n17751 0.00315748
R11123 DVDD.n1926 DVDD.n1925 0.00315748
R11124 DVDD.n1952 DVDD.n1951 0.00315748
R11125 DVDD.n2080 DVDD.n2079 0.00315748
R11126 DVDD.n2096 DVDD.n2095 0.00315748
R11127 DVDD.n2283 DVDD.n2282 0.00315748
R11128 DVDD.n19569 DVDD.n19568 0.00315748
R11129 DVDD.n18959 DVDD.n18958 0.00315748
R11130 DVDD.n6771 DVDD.n6770 0.00315748
R11131 DVDD.n6767 DVDD.n6766 0.00315748
R11132 DVDD.n6701 DVDD.n6700 0.00315748
R11133 DVDD.n6636 DVDD.n6635 0.00315748
R11134 DVDD.n6587 DVDD.n6586 0.00315748
R11135 DVDD.n6508 DVDD.n6507 0.00315748
R11136 DVDD.n6457 DVDD.n6456 0.00315748
R11137 DVDD.n6388 DVDD.n6387 0.00315748
R11138 DVDD.n6331 DVDD.n6330 0.00315748
R11139 DVDD.n6236 DVDD.n6235 0.00315748
R11140 DVDD.n6233 DVDD.n6232 0.00315748
R11141 DVDD.n6232 DVDD.n6231 0.00315748
R11142 DVDD.n4395 DVDD.n4394 0.00315748
R11143 DVDD.n3254 DVDD.n3253 0.00315748
R11144 DVDD.n3228 DVDD.n3227 0.00315748
R11145 DVDD.n3479 DVDD.n3478 0.00315748
R11146 DVDD.n3495 DVDD.n3494 0.00315748
R11147 DVDD.n3727 DVDD.n3726 0.00315748
R11148 DVDD.n3748 DVDD.n3747 0.00315748
R11149 DVDD.n18796 DVDD.n18795 0.00315748
R11150 DVDD.n9739 DVDD.n9738 0.00315748
R11151 DVDD.n9735 DVDD.n9734 0.00315748
R11152 DVDD.n9669 DVDD.n9668 0.00315748
R11153 DVDD.n9604 DVDD.n9603 0.00315748
R11154 DVDD.n9555 DVDD.n9554 0.00315748
R11155 DVDD.n8375 DVDD.n8374 0.00315748
R11156 DVDD.n8426 DVDD.n8425 0.00315748
R11157 DVDD.n9174 DVDD.n9173 0.00315748
R11158 DVDD.n9117 DVDD.n9116 0.00315748
R11159 DVDD.n8938 DVDD.n8937 0.00315748
R11160 DVDD.n8935 DVDD.n8934 0.00315748
R11161 DVDD.n8934 DVDD.n8933 0.00315748
R11162 DVDD.n8669 DVDD.n8668 0.00315748
R11163 DVDD.n17195 DVDD.n17194 0.00315322
R11164 DVDD.n17196 DVDD.n17195 0.00315322
R11165 DVDD.n17363 DVDD.n17362 0.00315322
R11166 DVDD.n17362 DVDD.n17361 0.00315322
R11167 DVDD.n17523 DVDD.n17522 0.00315322
R11168 DVDD.n17524 DVDD.n17523 0.00315322
R11169 DVDD.n10397 DVDD.n10396 0.00314375
R11170 DVDD.n15029 DVDD.n15028 0.00314
R11171 DVDD.n11066 DVDD.n11065 0.00314
R11172 DVDD.n15720 DVDD.n15719 0.00314
R11173 DVDD.n16079 DVDD.n16078 0.00314
R11174 DVDD.n8222 DVDD.n8221 0.00313598
R11175 DVDD.n8218 DVDD.n8217 0.00313598
R11176 DVDD.n9484 DVDD.n9483 0.00313598
R11177 DVDD.n9482 DVDD.n9481 0.00313598
R11178 DVDD.n7966 DVDD.n7965 0.00313598
R11179 DVDD.n7974 DVDD.n7973 0.00313598
R11180 DVDD.n8057 DVDD.n8056 0.00313598
R11181 DVDD.n13436 DVDD.n13435 0.00312498
R11182 DVDD.n13437 DVDD.n13436 0.00312498
R11183 DVDD.n5867 DVDD.n5866 0.00312498
R11184 DVDD.n5861 DVDD.n5860 0.00312498
R11185 DVDD.n5850 DVDD.n5849 0.00312498
R11186 DVDD.n5844 DVDD.n5843 0.00312498
R11187 DVDD.n5833 DVDD.n5832 0.00312498
R11188 DVDD.n5827 DVDD.n5826 0.00312498
R11189 DVDD.n12565 DVDD.n12564 0.00312498
R11190 DVDD.n12559 DVDD.n12558 0.00312498
R11191 DVDD.n12548 DVDD.n12547 0.00312498
R11192 DVDD.n12542 DVDD.n12541 0.00312498
R11193 DVDD.n12531 DVDD.n12530 0.00312498
R11194 DVDD.n12525 DVDD.n12524 0.00312498
R11195 DVDD.n5845 DVDD.n5844 0.00312498
R11196 DVDD.n12543 DVDD.n12542 0.00312498
R11197 DVDD.n5828 DVDD.n5827 0.00312498
R11198 DVDD.n12526 DVDD.n12525 0.00312498
R11199 DVDD.n12532 DVDD.n12531 0.00312498
R11200 DVDD.n5834 DVDD.n5833 0.00312498
R11201 DVDD.n12549 DVDD.n12548 0.00312498
R11202 DVDD.n5851 DVDD.n5850 0.00312498
R11203 DVDD.n5862 DVDD.n5861 0.00312498
R11204 DVDD.n12560 DVDD.n12559 0.00312498
R11205 DVDD.n5868 DVDD.n5867 0.00312498
R11206 DVDD.n12566 DVDD.n12565 0.00312498
R11207 DVDD.n4325 DVDD.n4324 0.00312498
R11208 DVDD.n4296 DVDD.n4295 0.00312498
R11209 DVDD.n4271 DVDD.n4270 0.00312498
R11210 DVDD.n4272 DVDD.n4271 0.00312498
R11211 DVDD.n4297 DVDD.n4296 0.00312498
R11212 DVDD.n4326 DVDD.n4325 0.00312498
R11213 DVDD.n8609 DVDD.n8608 0.00312498
R11214 DVDD.n8603 DVDD.n8602 0.00312498
R11215 DVDD.n8592 DVDD.n8591 0.00312498
R11216 DVDD.n8586 DVDD.n8585 0.00312498
R11217 DVDD.n8575 DVDD.n8574 0.00312498
R11218 DVDD.n8569 DVDD.n8568 0.00312498
R11219 DVDD.n8604 DVDD.n8603 0.00312498
R11220 DVDD.n8587 DVDD.n8586 0.00312498
R11221 DVDD.n8570 DVDD.n8569 0.00312498
R11222 DVDD.n8576 DVDD.n8575 0.00312498
R11223 DVDD.n8593 DVDD.n8592 0.00312498
R11224 DVDD.n8610 DVDD.n8609 0.00312498
R11225 DVDD.n3043 DVDD.n3042 0.00311161
R11226 DVDD.n3038 DVDD.n3037 0.00311161
R11227 DVDD.n3108 DVDD.n3107 0.00310839
R11228 DVDD.n3085 DVDD.n3084 0.00310839
R11229 DVDD.n3078 DVDD.n3077 0.00310839
R11230 DVDD.n3072 DVDD.n3071 0.00310839
R11231 DVDD.n3047 DVDD.n3046 0.00310839
R11232 DVDD.n3073 DVDD.n3072 0.00310839
R11233 DVDD.n3079 DVDD.n3078 0.00310839
R11234 DVDD.n3109 DVDD.n3108 0.00310839
R11235 DVDD.n3048 DVDD.n3047 0.00310839
R11236 DVDD.n18990 DVDD.n18989 0.00310718
R11237 DVDD.n10557 DVDD.n10556 0.00310718
R11238 DVDD.n8076 DVDD.n8075 0.00310011
R11239 DVDD.n15192 DVDD.n15191 0.0031
R11240 DVDD.n15200 DVDD.n15199 0.00309338
R11241 DVDD.n15123 DVDD.n15122 0.00309338
R11242 DVDD.n15962 DVDD.n15961 0.00307018
R11243 DVDD.n15963 DVDD.n15962 0.00307018
R11244 DVDD.n8292 DVDD.n8291 0.00307018
R11245 DVDD.n9455 DVDD.n9454 0.00307018
R11246 DVDD.n9456 DVDD.n9455 0.00307018
R11247 DVDD.n8135 DVDD.n8134 0.00307018
R11248 DVDD.n8134 DVDD.n8133 0.00307018
R11249 DVDD.n10292 DVDD.n10291 0.00305
R11250 DVDD.n10540 DVDD.n10539 0.00305
R11251 DVDD.n10499 DVDD.n10498 0.00305
R11252 DVDD.n17151 DVDD.n17150 0.00305
R11253 DVDD.n17110 DVDD.n17109 0.00305
R11254 DVDD.n17042 DVDD.n17041 0.00305
R11255 DVDD.n16720 DVDD.n16719 0.00305
R11256 DVDD.n16815 DVDD.n16814 0.00305
R11257 DVDD.n16551 DVDD.n16550 0.00305
R11258 DVDD.n16693 DVDD.n16692 0.00305
R11259 DVDD.n4933 DVDD.n4932 0.00303711
R11260 DVDD.n5354 DVDD.n5353 0.00303701
R11261 DVDD.n11667 DVDD.n11666 0.00303663
R11262 DVDD.n6595 DVDD.n6594 0.00303663
R11263 DVDD.n9563 DVDD.n9562 0.00303663
R11264 DVDD.n5334 DVDD.n5333 0.00303648
R11265 DVDD.n5437 DVDD.n5436 0.00303648
R11266 DVDD.n1603 DVDD.n1602 0.00303648
R11267 DVDD.n1609 DVDD.n1608 0.00303648
R11268 DVDD.n1602 DVDD.n1601 0.00303648
R11269 DVDD.n1608 DVDD.n1607 0.00303648
R11270 DVDD.n3424 DVDD.n3423 0.00302472
R11271 DVDD.n8012 DVDD.n8011 0.00300601
R11272 DVDD.n11654 DVDD.n11653 0.00300558
R11273 DVDD.n3832 DVDD.n3831 0.0030029
R11274 DVDD.n117 DVDD.n116 0.0030029
R11275 DVDD.n15197 DVDD.n15196 0.00299733
R11276 DVDD.n15270 DVDD.n15269 0.00299733
R11277 DVDD.n15277 DVDD.n15276 0.00299733
R11278 DVDD.n1220 DVDD.n1219 0.00298032
R11279 DVDD.n1190 DVDD.n1189 0.00298032
R11280 DVDD.n1570 DVDD.n1569 0.00298032
R11281 DVDD.n912 DVDD.n911 0.00298032
R11282 DVDD.n10168 DVDD.n10167 0.00298032
R11283 DVDD.n12021 DVDD.n12020 0.00298032
R11284 DVDD.n12029 DVDD.n12028 0.00298032
R11285 DVDD.n12113 DVDD.n12112 0.00298032
R11286 DVDD.n12289 DVDD.n12288 0.00298032
R11287 DVDD.n12287 DVDD.n12286 0.00298032
R11288 DVDD.n13450 DVDD.n13449 0.00298032
R11289 DVDD.n13455 DVDD.n13454 0.00298032
R11290 DVDD.n19855 DVDD.n19854 0.00298032
R11291 DVDD.n19868 DVDD.n19867 0.00298032
R11292 DVDD.n19907 DVDD.n19906 0.00298032
R11293 DVDD.n19924 DVDD.n19923 0.00298032
R11294 DVDD.n20116 DVDD.n20114 0.00298032
R11295 DVDD.n20116 DVDD.n20115 0.00298032
R11296 DVDD.n19059 DVDD.n19058 0.00298032
R11297 DVDD.n4674 DVDD.n4673 0.00298032
R11298 DVDD.n4939 DVDD.n4938 0.00298032
R11299 DVDD.n4946 DVDD.n4945 0.00298032
R11300 DVDD.n5010 DVDD.n5009 0.00298032
R11301 DVDD.n5199 DVDD.n5198 0.00298032
R11302 DVDD.n5227 DVDD.n5226 0.00298032
R11303 DVDD.n5349 DVDD.n5348 0.00298032
R11304 DVDD.n5375 DVDD.n5374 0.00298032
R11305 DVDD.n5440 DVDD.n5439 0.00298032
R11306 DVDD.n5464 DVDD.n5463 0.00298032
R11307 DVDD.n5466 DVDD.n5465 0.00298032
R11308 DVDD.n6053 DVDD.n6052 0.00298032
R11309 DVDD.n1356 DVDD.n1355 0.00298032
R11310 DVDD.n1521 DVDD.n1520 0.00298032
R11311 DVDD.n1508 DVDD.n1507 0.00298032
R11312 DVDD.n1470 DVDD.n1469 0.00298032
R11313 DVDD.n1453 DVDD.n1452 0.00298032
R11314 DVDD.n19213 DVDD.n19212 0.00298032
R11315 DVDD.n19214 DVDD.n19213 0.00298032
R11316 DVDD.n19441 DVDD.n19440 0.00298032
R11317 DVDD.n11381 DVDD.n11380 0.00298032
R11318 DVDD.n11814 DVDD.n11813 0.00298032
R11319 DVDD.n11807 DVDD.n11806 0.00298032
R11320 DVDD.n11744 DVDD.n11743 0.00298032
R11321 DVDD.n12379 DVDD.n12378 0.00298032
R11322 DVDD.n12407 DVDD.n12406 0.00298032
R11323 DVDD.n13111 DVDD.n13110 0.00298032
R11324 DVDD.n13085 DVDD.n13084 0.00298032
R11325 DVDD.n13023 DVDD.n13022 0.00298032
R11326 DVDD.n12999 DVDD.n12998 0.00298032
R11327 DVDD.n12997 DVDD.n12996 0.00298032
R11328 DVDD.n12699 DVDD.n12698 0.00298032
R11329 DVDD.n1933 DVDD.n1932 0.00298032
R11330 DVDD.n2077 DVDD.n2076 0.00298032
R11331 DVDD.n2090 DVDD.n2089 0.00298032
R11332 DVDD.n2128 DVDD.n2127 0.00298032
R11333 DVDD.n2145 DVDD.n2144 0.00298032
R11334 DVDD.n19501 DVDD.n19499 0.00298032
R11335 DVDD.n19501 DVDD.n19500 0.00298032
R11336 DVDD.n18951 DVDD.n18950 0.00298032
R11337 DVDD.n7010 DVDD.n7009 0.00298032
R11338 DVDD.n6745 DVDD.n6744 0.00298032
R11339 DVDD.n6738 DVDD.n6737 0.00298032
R11340 DVDD.n6674 DVDD.n6673 0.00298032
R11341 DVDD.n6483 DVDD.n6482 0.00298032
R11342 DVDD.n6455 DVDD.n6454 0.00298032
R11343 DVDD.n6412 DVDD.n6411 0.00298032
R11344 DVDD.n6386 DVDD.n6385 0.00298032
R11345 DVDD.n6321 DVDD.n6320 0.00298032
R11346 DVDD.n6297 DVDD.n6296 0.00298032
R11347 DVDD.n6295 DVDD.n6294 0.00298032
R11348 DVDD.n4510 DVDD.n4509 0.00298032
R11349 DVDD.n3247 DVDD.n3246 0.00298032
R11350 DVDD.n3476 DVDD.n3475 0.00298032
R11351 DVDD.n3489 DVDD.n3488 0.00298032
R11352 DVDD.n3527 DVDD.n3526 0.00298032
R11353 DVDD.n3544 DVDD.n3543 0.00298032
R11354 DVDD.n18517 DVDD.n18516 0.00298032
R11355 DVDD.n18518 DVDD.n18517 0.00298032
R11356 DVDD.n18788 DVDD.n18787 0.00298032
R11357 DVDD.n10027 DVDD.n10026 0.00298032
R11358 DVDD.n9713 DVDD.n9712 0.00298032
R11359 DVDD.n9706 DVDD.n9705 0.00298032
R11360 DVDD.n9642 DVDD.n9641 0.00298032
R11361 DVDD.n8400 DVDD.n8399 0.00298032
R11362 DVDD.n8428 DVDD.n8427 0.00298032
R11363 DVDD.n9198 DVDD.n9197 0.00298032
R11364 DVDD.n9172 DVDD.n9171 0.00298032
R11365 DVDD.n9107 DVDD.n9106 0.00298032
R11366 DVDD.n9083 DVDD.n9082 0.00298032
R11367 DVDD.n9081 DVDD.n9080 0.00298032
R11368 DVDD.n8784 DVDD.n8783 0.00298032
R11369 DVDD.n15990 DVDD.n15989 0.00297612
R11370 DVDD.n15991 DVDD.n15990 0.00297612
R11371 DVDD.n15941 DVDD.n15940 0.00297612
R11372 DVDD.n15940 DVDD.n15939 0.00297612
R11373 DVDD.n15681 DVDD.n15680 0.00297612
R11374 DVDD.n15680 DVDD.n15679 0.00297612
R11375 DVDD.n8229 DVDD.n8228 0.00297612
R11376 DVDD.n9421 DVDD.n9420 0.00297612
R11377 DVDD.n9422 DVDD.n9421 0.00297612
R11378 DVDD.n8103 DVDD.n8102 0.00297612
R11379 DVDD.n8102 DVDD.n8101 0.00297612
R11380 DVDD.n9901 DVDD.n9900 0.00297612
R11381 DVDD.n8091 DVDD.n8090 0.00297612
R11382 DVDD.n8090 DVDD.n8089 0.00297612
R11383 DVDD.n9902 DVDD.n9901 0.00297612
R11384 DVDD.n7475 DVDD 0.00297599
R11385 DVDD.n3813 DVDD.n3812 0.002975
R11386 DVDD.n18997 DVDD.n18996 0.002975
R11387 DVDD.n10078 DVDD.n10077 0.002975
R11388 DVDD.n7630 DVDD.n7629 0.002975
R11389 DVDD.n3892 DVDD.n3891 0.002975
R11390 DVDD.n7122 DVDD.n7121 0.002975
R11391 DVDD.n7654 DVDD.n7653 0.002975
R11392 DVDD.n1814 DVDD.n1813 0.002975
R11393 DVDD.n3781 DVDD.n3780 0.002975
R11394 DVDD.n2824 DVDD.n2823 0.002975
R11395 DVDD.n20296 DVDD.n20295 0.002975
R11396 DVDD.n20318 DVDD.n20317 0.002975
R11397 DVDD.n14849 DVDD.n14848 0.002975
R11398 DVDD.n10600 DVDD.n10599 0.002975
R11399 DVDD.n11660 DVDD.n11659 0.00294879
R11400 DVDD.n6588 DVDD.n6587 0.00294879
R11401 DVDD.n6234 DVDD.n6233 0.00294879
R11402 DVDD.n9556 DVDD.n9555 0.00294879
R11403 DVDD.n8936 DVDD.n8935 0.00294879
R11404 DVDD.n12363 DVDD.n12362 0.00294857
R11405 DVDD.n6499 DVDD.n6498 0.00294857
R11406 DVDD.n8384 DVDD.n8383 0.00294857
R11407 DVDD.n19899 DVDD.n19898 0.00294837
R11408 DVDD.n12260 DVDD.n12259 0.00294798
R11409 DVDD.n13377 DVDD.n13376 0.00294798
R11410 DVDD.n12193 DVDD.n12192 0.00294798
R11411 DVDD.n12261 DVDD.n12260 0.00294798
R11412 DVDD.n13376 DVDD.n13375 0.00294798
R11413 DVDD.n15494 DVDD.n15493 0.00294798
R11414 DVDD.n15506 DVDD.n15505 0.00294798
R11415 DVDD.n14671 DVDD.n14670 0.00294798
R11416 DVDD.n14368 DVDD.n14367 0.00294798
R11417 DVDD.n14672 DVDD.n14671 0.00294798
R11418 DVDD.n15493 DVDD.n15492 0.00294798
R11419 DVDD.n15505 DVDD.n15504 0.00294798
R11420 DVDD.n19918 DVDD.n19917 0.00294798
R11421 DVDD.n5053 DVDD.n5052 0.00294798
R11422 DVDD.n11701 DVDD.n11700 0.00294798
R11423 DVDD.n18105 DVDD.n18104 0.00294798
R11424 DVDD.n18027 DVDD.n18026 0.00294798
R11425 DVDD.n18028 DVDD.n18027 0.00294798
R11426 DVDD.n18116 DVDD.n18115 0.00294798
R11427 DVDD.n18106 DVDD.n18105 0.00294798
R11428 DVDD.n6630 DVDD.n6629 0.00294798
R11429 DVDD.n4389 DVDD.n4388 0.00294798
R11430 DVDD.n6631 DVDD.n6630 0.00294798
R11431 DVDD.n4390 DVDD.n4389 0.00294798
R11432 DVDD.n13717 DVDD.n13716 0.00294798
R11433 DVDD.n17747 DVDD.n17746 0.00294798
R11434 DVDD.n14369 DVDD.n14368 0.00294798
R11435 DVDD.n12594 DVDD.n12593 0.00294798
R11436 DVDD.n5931 DVDD.n5930 0.00294798
R11437 DVDD.n9598 DVDD.n9597 0.00294798
R11438 DVDD.n8663 DVDD.n8662 0.00294798
R11439 DVDD.n9599 DVDD.n9598 0.00294798
R11440 DVDD.n8664 DVDD.n8663 0.00294798
R11441 DVDD.n8285 DVDD.n8284 0.0029477
R11442 DVDD.n8281 DVDD.n8280 0.0029477
R11443 DVDD.n7946 DVDD.n7945 0.0029477
R11444 DVDD.n7950 DVDD.n7949 0.0029477
R11445 DVDD.n8030 DVDD.n8029 0.0029477
R11446 DVDD.n8038 DVDD.n8037 0.0029477
R11447 DVDD.n7948 DVDD.n7947 0.0029119
R11448 DVDD.n8283 DVDD.n8282 0.00291179
R11449 DVDD.n3104 DVDD.n3103 0.00291071
R11450 DVDD.n15253 DVDD.n15252 0.00290128
R11451 DVDD.n15267 DVDD.n15266 0.00290128
R11452 DVDD.n15288 DVDD.n15131 0.00290128
R11453 DVDD.n16051 DVDD.n16050 0.00288206
R11454 DVDD.n15999 DVDD.n15998 0.00288206
R11455 DVDD.n16000 DVDD.n15999 0.00288206
R11456 DVDD.n16052 DVDD.n16051 0.00288206
R11457 DVDD.n15663 DVDD.n15662 0.00288206
R11458 DVDD.n15933 DVDD.n15932 0.00288206
R11459 DVDD.n15932 DVDD.n15931 0.00288206
R11460 DVDD.n15664 DVDD.n15663 0.00288206
R11461 DVDD.n8166 DVDD.n8165 0.00288206
R11462 DVDD.n8167 DVDD.n8166 0.00288206
R11463 DVDD.n8085 DVDD.n8084 0.00288206
R11464 DVDD.n15250 DVDD.n15249 0.0028625
R11465 DVDD.n1229 DVDD.n1228 0.00285947
R11466 DVDD.n1205 DVDD.n1204 0.00285947
R11467 DVDD.n1198 DVDD.n1197 0.00285947
R11468 DVDD.n1192 DVDD.n1191 0.00285947
R11469 DVDD.n1169 DVDD.n1168 0.00285947
R11470 DVDD.n1581 DVDD.n1580 0.00285947
R11471 DVDD.n11485 DVDD.n11484 0.00285947
R11472 DVDD.n12150 DVDD.n12149 0.00285947
R11473 DVDD.n12162 DVDD.n12161 0.00285947
R11474 DVDD.n12226 DVDD.n12225 0.00285947
R11475 DVDD.n13443 DVDD.n13442 0.00285947
R11476 DVDD.n13532 DVDD.n13531 0.00285947
R11477 DVDD.n13613 DVDD.n13612 0.00285947
R11478 DVDD.n12149 DVDD.n12148 0.00285947
R11479 DVDD.n11486 DVDD.n11485 0.00285947
R11480 DVDD.n1193 DVDD.n1192 0.00285947
R11481 DVDD.n1199 DVDD.n1198 0.00285947
R11482 DVDD.n1206 DVDD.n1205 0.00285947
R11483 DVDD.n1230 DVDD.n1229 0.00285947
R11484 DVDD.n12161 DVDD.n12160 0.00285947
R11485 DVDD.n1170 DVDD.n1169 0.00285947
R11486 DVDD.n12227 DVDD.n12226 0.00285947
R11487 DVDD.n13442 DVDD.n13441 0.00285947
R11488 DVDD.n13531 DVDD.n13530 0.00285947
R11489 DVDD.n13612 DVDD.n13611 0.00285947
R11490 DVDD.n2724 DVDD.n2723 0.00285947
R11491 DVDD.n2766 DVDD.n2765 0.00285947
R11492 DVDD.n14815 DVDD.n14814 0.00285947
R11493 DVDD.n15466 DVDD.n15465 0.00285947
R11494 DVDD.n14726 DVDD.n14725 0.00285947
R11495 DVDD.n14643 DVDD.n14642 0.00285947
R11496 DVDD.n14589 DVDD.n14588 0.00285947
R11497 DVDD.n14501 DVDD.n14500 0.00285947
R11498 DVDD.n14396 DVDD.n14395 0.00285947
R11499 DVDD.n14644 DVDD.n14643 0.00285947
R11500 DVDD.n15465 DVDD.n15464 0.00285947
R11501 DVDD.n14727 DVDD.n14726 0.00285947
R11502 DVDD.n14814 DVDD.n14813 0.00285947
R11503 DVDD.n2765 DVDD.n2764 0.00285947
R11504 DVDD.n2725 DVDD.n2724 0.00285947
R11505 DVDD.n14590 DVDD.n14589 0.00285947
R11506 DVDD.n14502 DVDD.n14501 0.00285947
R11507 DVDD.n4779 DVDD.n4778 0.00285947
R11508 DVDD.n5017 DVDD.n5016 0.00285947
R11509 DVDD.n5546 DVDD.n5545 0.00285947
R11510 DVDD.n5697 DVDD.n5696 0.00285947
R11511 DVDD.n5169 DVDD.n5168 0.00285947
R11512 DVDD.n5016 DVDD.n5015 0.00285947
R11513 DVDD.n4778 DVDD.n4777 0.00285947
R11514 DVDD.n5545 DVDD.n5544 0.00285947
R11515 DVDD.n5696 DVDD.n5695 0.00285947
R11516 DVDD.n11605 DVDD.n11604 0.00285947
R11517 DVDD.n11737 DVDD.n11736 0.00285947
R11518 DVDD.n12871 DVDD.n12870 0.00285947
R11519 DVDD.n12744 DVDD.n12743 0.00285947
R11520 DVDD.n11738 DVDD.n11737 0.00285947
R11521 DVDD.n11604 DVDD.n11603 0.00285947
R11522 DVDD.n11668 DVDD.n11667 0.00285947
R11523 DVDD.n12350 DVDD.n12349 0.00285947
R11524 DVDD.n12745 DVDD.n12744 0.00285947
R11525 DVDD.n12872 DVDD.n12871 0.00285947
R11526 DVDD.n763 DVDD.n762 0.00285947
R11527 DVDD.n800 DVDD.n799 0.00285947
R11528 DVDD.n18223 DVDD.n18222 0.00285947
R11529 DVDD.n18079 DVDD.n18078 0.00285947
R11530 DVDD.n18001 DVDD.n18000 0.00285947
R11531 DVDD.n17949 DVDD.n17948 0.00285947
R11532 DVDD.n17868 DVDD.n17867 0.00285947
R11533 DVDD.n18142 DVDD.n18141 0.00285947
R11534 DVDD.n18224 DVDD.n18223 0.00285947
R11535 DVDD.n17869 DVDD.n17868 0.00285947
R11536 DVDD.n17950 DVDD.n17949 0.00285947
R11537 DVDD.n6905 DVDD.n6904 0.00285947
R11538 DVDD.n6667 DVDD.n6666 0.00285947
R11539 DVDD.n6250 DVDD.n6249 0.00285947
R11540 DVDD.n6126 DVDD.n6125 0.00285947
R11541 DVDD.n4417 DVDD.n4416 0.00285947
R11542 DVDD.n6513 DVDD.n6512 0.00285947
R11543 DVDD.n6906 DVDD.n6905 0.00285947
R11544 DVDD.n6668 DVDD.n6667 0.00285947
R11545 DVDD.n6596 DVDD.n6595 0.00285947
R11546 DVDD.n6251 DVDD.n6250 0.00285947
R11547 DVDD.n6127 DVDD.n6126 0.00285947
R11548 DVDD.n4418 DVDD.n4417 0.00285947
R11549 DVDD.n13694 DVDD.n13693 0.00285947
R11550 DVDD.n17773 DVDD.n17772 0.00285947
R11551 DVDD.n5957 DVDD.n5956 0.00285947
R11552 DVDD.n14397 DVDD.n14396 0.00285947
R11553 DVDD.n12620 DVDD.n12619 0.00285947
R11554 DVDD.n7861 DVDD.n7860 0.00285947
R11555 DVDD.n9635 DVDD.n9634 0.00285947
R11556 DVDD.n8952 DVDD.n8951 0.00285947
R11557 DVDD.n8828 DVDD.n8827 0.00285947
R11558 DVDD.n8691 DVDD.n8690 0.00285947
R11559 DVDD.n9636 DVDD.n9635 0.00285947
R11560 DVDD.n8692 DVDD.n8691 0.00285947
R11561 DVDD.n8370 DVDD.n8369 0.00285947
R11562 DVDD.n7860 DVDD.n7859 0.00285947
R11563 DVDD.n9564 DVDD.n9563 0.00285947
R11564 DVDD.n8953 DVDD.n8952 0.00285947
R11565 DVDD.n8829 DVDD.n8828 0.00285947
R11566 DVDD.n10317 DVDD.n10228 0.00285
R11567 DVDD.n9783 DVDD.n9782 0.00284
R11568 DVDD.n9539 DVDD.n9538 0.00284
R11569 DVDD.n9242 DVDD.n9241 0.00284
R11570 DVDD.n9284 DVDD.n9283 0.00284
R11571 DVDD.n6832 DVDD.n6831 0.00284
R11572 DVDD.n6571 DVDD.n6570 0.00284
R11573 DVDD.n4000 DVDD.n3999 0.00284
R11574 DVDD.n3958 DVDD.n3957 0.00284
R11575 DVDD.n4869 DVDD.n4868 0.00284
R11576 DVDD.n5162 DVDD.n5161 0.00284
R11577 DVDD.n5305 DVDD.n5304 0.00284
R11578 DVDD.n5263 DVDD.n5262 0.00284
R11579 DVDD.n11884 DVDD.n11883 0.00284
R11580 DVDD.n12343 DVDD.n12342 0.00284
R11581 DVDD.n13153 DVDD.n13152 0.00284
R11582 DVDD.n13195 DVDD.n13194 0.00284
R11583 DVDD.n8220 DVDD.n8219 0.0028177
R11584 DVDD.n1827 DVDD.n1826 0.00281
R11585 DVDD.n19553 DVDD.n19552 0.00281
R11586 DVDD.n19539 DVDD.n19538 0.00281
R11587 DVDD.n19525 DVDD.n19524 0.00281
R11588 DVDD.n19511 DVDD.n19510 0.00281
R11589 DVDD.n18868 DVDD.n18867 0.00281
R11590 DVDD.n18855 DVDD.n18854 0.00281
R11591 DVDD.n18850 DVDD.n18849 0.00281
R11592 DVDD.n18845 DVDD.n18844 0.00281
R11593 DVDD.n18840 DVDD.n18839 0.00281
R11594 DVDD.n19605 DVDD.n19604 0.00281
R11595 DVDD.n20168 DVDD.n20167 0.00281
R11596 DVDD.n20154 DVDD.n20153 0.00281
R11597 DVDD.n20140 DVDD.n20139 0.00281
R11598 DVDD.n20126 DVDD.n20125 0.00281
R11599 DVDD.n19117 DVDD.n19116 0.00281
R11600 DVDD.n19103 DVDD.n19102 0.00281
R11601 DVDD.n19098 DVDD.n19097 0.00281
R11602 DVDD.n19093 DVDD.n19092 0.00281
R11603 DVDD.n19088 DVDD.n19087 0.00281
R11604 DVDD.n7520 DVDD.n7519 0.00281
R11605 DVDD.n851 DVDD.n850 0.00281
R11606 DVDD.n225 DVDD.n224 0.00281
R11607 DVDD.n191 DVDD.n190 0.00281
R11608 DVDD.n19394 DVDD.n19393 0.00281
R11609 DVDD.n19380 DVDD.n19379 0.00281
R11610 DVDD.n19375 DVDD.n19374 0.00281
R11611 DVDD.n19370 DVDD.n19369 0.00281
R11612 DVDD.n18265 DVDD.n18264 0.00281
R11613 DVDD.n10375 DVDD.n10374 0.00281
R11614 DVDD.n10512 DVDD.n10511 0.00281
R11615 DVDD.n10441 DVDD.n10440 0.00281
R11616 DVDD.n14971 DVDD.n14970 0.00281
R11617 DVDD.n15048 DVDD.n15047 0.00281
R11618 DVDD.n15386 DVDD.n15385 0.00281
R11619 DVDD.n16525 DVDD.n16524 0.00281
R11620 DVDD.n17122 DVDD.n17121 0.00281
R11621 DVDD.n17072 DVDD.n17071 0.00281
R11622 DVDD.n11029 DVDD.n11028 0.00281
R11623 DVDD.n11084 DVDD.n11083 0.00281
R11624 DVDD.n11195 DVDD.n11194 0.00281
R11625 DVDD.n16865 DVDD.n16864 0.00281
R11626 DVDD.n16326 DVDD.n16325 0.00281
R11627 DVDD.n16712 DVDD.n16711 0.00281
R11628 DVDD.n16734 DVDD.n16733 0.00281
R11629 DVDD.n15739 DVDD.n15738 0.00281
R11630 DVDD.n15695 DVDD.n15694 0.00281
R11631 DVDD.n16543 DVDD.n16542 0.00281
R11632 DVDD.n16565 DVDD.n16564 0.00281
R11633 DVDD.n16098 DVDD.n16097 0.00281
R11634 DVDD.n15907 DVDD.n15906 0.00281
R11635 DVDD.n3615 DVDD.n3614 0.00281
R11636 DVDD.n18604 DVDD.n18603 0.00281
R11637 DVDD.n18733 DVDD.n18732 0.00281
R11638 DVDD.n18401 DVDD.n18400 0.00281
R11639 DVDD.n18376 DVDD.n18375 0.00281
R11640 DVDD.n18371 DVDD.n18370 0.00281
R11641 DVDD.n18366 DVDD.n18365 0.00281
R11642 DVDD.n14790 DVDD.n14789 0.00281
R11643 DVDD.n4318 DVDD.n4317 0.00280842
R11644 DVDD.n4289 DVDD.n4288 0.00280842
R11645 DVDD.n4264 DVDD.n4263 0.00280842
R11646 DVDD.n3056 DVDD.n3055 0.00280731
R11647 DVDD.n3057 DVDD.n3056 0.00280731
R11648 DVDD.n15254 DVDD.n15253 0.00280523
R11649 DVDD.n1165 DVDD.n1164 0.00280315
R11650 DVDD.n1160 DVDD.n1159 0.00280315
R11651 DVDD.n1621 DVDD.n1620 0.00280315
R11652 DVDD.n1626 DVDD.n1625 0.00280315
R11653 DVDD.n867 DVDD.n866 0.00280315
R11654 DVDD.n19287 DVDD.n19286 0.00280315
R11655 DVDD.n19293 DVDD.n19292 0.00280315
R11656 DVDD.n19298 DVDD.n19297 0.00280315
R11657 DVDD.n19415 DVDD.n19309 0.00280315
R11658 DVDD.n19335 DVDD.n19334 0.00280315
R11659 DVDD.n11999 DVDD.n11998 0.00280315
R11660 DVDD.n12004 DVDD.n12003 0.00280315
R11661 DVDD.n12087 DVDD.n12086 0.00280315
R11662 DVDD.n12095 DVDD.n12094 0.00280315
R11663 DVDD.n13384 DVDD.n13383 0.00280315
R11664 DVDD.n13389 DVDD.n13388 0.00280315
R11665 DVDD.n18479 DVDD.n18478 0.00280315
R11666 DVDD.n14164 DVDD.n14163 0.00280315
R11667 DVDD.n14157 DVDD.n14156 0.00280315
R11668 DVDD.n14065 DVDD.n14064 0.00280315
R11669 DVDD.n14058 DVDD.n14057 0.00280315
R11670 DVDD.n13968 DVDD.n13967 0.00280315
R11671 DVDD.n13961 DVDD.n13960 0.00280315
R11672 DVDD.n19706 DVDD.n19705 0.00280315
R11673 DVDD.n19707 DVDD.n19706 0.00280315
R11674 DVDD.n19911 DVDD.n19910 0.00280315
R11675 DVDD.n19921 DVDD.n19920 0.00280315
R11676 DVDD.n20054 DVDD.n20053 0.00280315
R11677 DVDD.n20059 DVDD.n20058 0.00280315
R11678 DVDD.n20209 DVDD.n20208 0.00280315
R11679 DVDD.n20208 DVDD.n20207 0.00280315
R11680 DVDD.n20113 DVDD.n20112 0.00280315
R11681 DVDD.n20114 DVDD.n20113 0.00280315
R11682 DVDD.n19069 DVDD.n19068 0.00280315
R11683 DVDD.n4670 DVDD.n4669 0.00280315
R11684 DVDD.n4671 DVDD.n4670 0.00280315
R11685 DVDD.n4672 DVDD.n4671 0.00280315
R11686 DVDD.n4675 DVDD.n4674 0.00280315
R11687 DVDD.n4810 DVDD.n4809 0.00280315
R11688 DVDD.n5008 DVDD.n5007 0.00280315
R11689 DVDD.n5100 DVDD.n5099 0.00280315
R11690 DVDD.n5106 DVDD.n5105 0.00280315
R11691 DVDD.n5325 DVDD.n5324 0.00280315
R11692 DVDD.n5329 DVDD.n5328 0.00280315
R11693 DVDD.n5341 DVDD.n5340 0.00280315
R11694 DVDD.n5347 DVDD.n5346 0.00280315
R11695 DVDD.n5382 DVDD.n5381 0.00280315
R11696 DVDD.n5414 DVDD.n5413 0.00280315
R11697 DVDD.n5442 DVDD.n5441 0.00280315
R11698 DVDD.n1351 DVDD.n1350 0.00280315
R11699 DVDD.n1352 DVDD.n1351 0.00280315
R11700 DVDD.n1466 DVDD.n1465 0.00280315
R11701 DVDD.n1456 DVDD.n1455 0.00280315
R11702 DVDD.n1719 DVDD.n1718 0.00280315
R11703 DVDD.n1714 DVDD.n1713 0.00280315
R11704 DVDD.n287 DVDD.n286 0.00280315
R11705 DVDD.n286 DVDD.n285 0.00280315
R11706 DVDD.n19211 DVDD.n19210 0.00280315
R11707 DVDD.n19212 DVDD.n19211 0.00280315
R11708 DVDD.n19451 DVDD.n19450 0.00280315
R11709 DVDD.n11377 DVDD.n11376 0.00280315
R11710 DVDD.n11378 DVDD.n11377 0.00280315
R11711 DVDD.n11379 DVDD.n11378 0.00280315
R11712 DVDD.n11382 DVDD.n11381 0.00280315
R11713 DVDD.n11636 DVDD.n11635 0.00280315
R11714 DVDD.n11819 DVDD.n11818 0.00280315
R11715 DVDD.n11746 DVDD.n11745 0.00280315
R11716 DVDD.n11649 DVDD.n11648 0.00280315
R11717 DVDD.n13134 DVDD.n13133 0.00280315
R11718 DVDD.n13130 DVDD.n13129 0.00280315
R11719 DVDD.n13118 DVDD.n13117 0.00280315
R11720 DVDD.n13079 DVDD.n13078 0.00280315
R11721 DVDD.n13048 DVDD.n13047 0.00280315
R11722 DVDD.n13021 DVDD.n13020 0.00280315
R11723 DVDD.n19175 DVDD.n19174 0.00280315
R11724 DVDD.n17504 DVDD.n17503 0.00280315
R11725 DVDD.n17497 DVDD.n17496 0.00280315
R11726 DVDD.n17461 DVDD.n17460 0.00280315
R11727 DVDD.n17454 DVDD.n17453 0.00280315
R11728 DVDD.n17345 DVDD.n17344 0.00280315
R11729 DVDD.n17338 DVDD.n17337 0.00280315
R11730 DVDD.n1928 DVDD.n1927 0.00280315
R11731 DVDD.n1929 DVDD.n1928 0.00280315
R11732 DVDD.n2132 DVDD.n2131 0.00280315
R11733 DVDD.n2142 DVDD.n2141 0.00280315
R11734 DVDD.n2275 DVDD.n2274 0.00280315
R11735 DVDD.n2280 DVDD.n2279 0.00280315
R11736 DVDD.n19594 DVDD.n19593 0.00280315
R11737 DVDD.n19593 DVDD.n19592 0.00280315
R11738 DVDD.n19498 DVDD.n19497 0.00280315
R11739 DVDD.n19499 DVDD.n19498 0.00280315
R11740 DVDD.n18961 DVDD.n18960 0.00280315
R11741 DVDD.n7014 DVDD.n7013 0.00280315
R11742 DVDD.n7013 DVDD.n7012 0.00280315
R11743 DVDD.n7012 DVDD.n7011 0.00280315
R11744 DVDD.n7009 DVDD.n7008 0.00280315
R11745 DVDD.n6874 DVDD.n6873 0.00280315
R11746 DVDD.n6750 DVDD.n6749 0.00280315
R11747 DVDD.n6676 DVDD.n6675 0.00280315
R11748 DVDD.n6576 DVDD.n6575 0.00280315
R11749 DVDD.n6436 DVDD.n6435 0.00280315
R11750 DVDD.n6432 DVDD.n6431 0.00280315
R11751 DVDD.n6420 DVDD.n6419 0.00280315
R11752 DVDD.n6379 DVDD.n6378 0.00280315
R11753 DVDD.n6347 DVDD.n6346 0.00280315
R11754 DVDD.n6319 DVDD.n6318 0.00280315
R11755 DVDD.n3252 DVDD.n3251 0.00280315
R11756 DVDD.n3251 DVDD.n3250 0.00280315
R11757 DVDD.n3531 DVDD.n3530 0.00280315
R11758 DVDD.n3541 DVDD.n3540 0.00280315
R11759 DVDD.n3719 DVDD.n3718 0.00280315
R11760 DVDD.n3724 DVDD.n3723 0.00280315
R11761 DVDD.n3773 DVDD.n3772 0.00280315
R11762 DVDD.n3772 DVDD.n3771 0.00280315
R11763 DVDD.n18515 DVDD.n18514 0.00280315
R11764 DVDD.n18516 DVDD.n18515 0.00280315
R11765 DVDD.n18798 DVDD.n18797 0.00280315
R11766 DVDD.n10031 DVDD.n10030 0.00280315
R11767 DVDD.n10030 DVDD.n10029 0.00280315
R11768 DVDD.n10029 DVDD.n10028 0.00280315
R11769 DVDD.n10026 DVDD.n10025 0.00280315
R11770 DVDD.n7892 DVDD.n7891 0.00280315
R11771 DVDD.n9718 DVDD.n9717 0.00280315
R11772 DVDD.n9644 DVDD.n9643 0.00280315
R11773 DVDD.n9544 DVDD.n9543 0.00280315
R11774 DVDD.n9222 DVDD.n9221 0.00280315
R11775 DVDD.n9218 DVDD.n9217 0.00280315
R11776 DVDD.n9206 DVDD.n9205 0.00280315
R11777 DVDD.n9165 DVDD.n9164 0.00280315
R11778 DVDD.n9133 DVDD.n9132 0.00280315
R11779 DVDD.n9105 DVDD.n9104 0.00280315
R11780 DVDD.n8145 DVDD.n8144 0.00278799
R11781 DVDD.n8144 DVDD.n8143 0.00278799
R11782 DVDD.n16030 DVDD.n16029 0.00278799
R11783 DVDD.n16021 DVDD.n16020 0.00278799
R11784 DVDD.n16022 DVDD.n16021 0.00278799
R11785 DVDD.n16029 DVDD.n16028 0.00278799
R11786 DVDD.n15641 DVDD.n15640 0.00278799
R11787 DVDD.n15633 DVDD.n15632 0.00278799
R11788 DVDD.n15642 DVDD.n15641 0.00278799
R11789 DVDD.n15634 DVDD.n15633 0.00278799
R11790 DVDD.n8307 DVDD.n8306 0.00278799
R11791 DVDD.n8021 DVDD.n8020 0.00278799
R11792 DVDD.n18876 DVDD.n18875 0.00278
R11793 DVDD.n19125 DVDD.n19124 0.00278
R11794 DVDD.n208 DVDD.n207 0.00278
R11795 DVDD.n19404 DVDD.n19403 0.00278
R11796 DVDD.n18635 DVDD.n18634 0.00278
R11797 DVDD.n18411 DVDD.n18410 0.00278
R11798 DVDD.n5066 DVDD.n5065 0.00277163
R11799 DVDD.n19733 DVDD.n19732 0.00277109
R11800 DVDD.n1594 DVDD.n1593 0.00277096
R11801 DVDD.n1637 DVDD.n1636 0.00277096
R11802 DVDD.n12144 DVDD.n12143 0.00277096
R11803 DVDD.n13506 DVDD.n13505 0.00277096
R11804 DVDD.n13639 DVDD.n13638 0.00277096
R11805 DVDD.n12143 DVDD.n12142 0.00277096
R11806 DVDD.n13558 DVDD.n13557 0.00277096
R11807 DVDD.n13606 DVDD.n13605 0.00277096
R11808 DVDD.n13687 DVDD.n13686 0.00277096
R11809 DVDD.n2752 DVDD.n2751 0.00277096
R11810 DVDD.n2794 DVDD.n2793 0.00277096
R11811 DVDD.n15405 DVDD.n15404 0.00277096
R11812 DVDD.n15457 DVDD.n15456 0.00277096
R11813 DVDD.n14699 DVDD.n14698 0.00277096
R11814 DVDD.n14615 DVDD.n14614 0.00277096
R11815 DVDD.n14561 DVDD.n14560 0.00277096
R11816 DVDD.n14509 DVDD.n14508 0.00277096
R11817 DVDD.n14473 DVDD.n14472 0.00277096
R11818 DVDD.n14405 DVDD.n14404 0.00277096
R11819 DVDD.n14406 DVDD.n14405 0.00277096
R11820 DVDD.n14510 DVDD.n14509 0.00277096
R11821 DVDD.n14616 DVDD.n14615 0.00277096
R11822 DVDD.n15456 DVDD.n15455 0.00277096
R11823 DVDD.n15404 DVDD.n15403 0.00277096
R11824 DVDD.n2793 DVDD.n2792 0.00277096
R11825 DVDD.n2753 DVDD.n2752 0.00277096
R11826 DVDD.n14474 DVDD.n14473 0.00277096
R11827 DVDD.n14562 DVDD.n14561 0.00277096
R11828 DVDD.n14698 DVDD.n14697 0.00277096
R11829 DVDD.n5002 DVDD.n5001 0.00277096
R11830 DVDD.n5964 DVDD.n5963 0.00277096
R11831 DVDD.n5595 DVDD.n5594 0.00277096
R11832 DVDD.n5690 DVDD.n5689 0.00277096
R11833 DVDD.n5472 DVDD.n5471 0.00277096
R11834 DVDD.n5001 DVDD.n5000 0.00277096
R11835 DVDD.n19751 DVDD.n19750 0.00277096
R11836 DVDD.n6107 DVDD.n6102 0.00277096
R11837 DVDD.n12991 DVDD.n12990 0.00277096
R11838 DVDD.n11752 DVDD.n11751 0.00277096
R11839 DVDD.n12627 DVDD.n12626 0.00277096
R11840 DVDD.n12738 DVDD.n12734 0.00277096
R11841 DVDD.n12751 DVDD.n12750 0.00277096
R11842 DVDD.n12832 DVDD.n12831 0.00277096
R11843 DVDD.n826 DVDD.n825 0.00277096
R11844 DVDD.n18197 DVDD.n18196 0.00277096
R11845 DVDD.n17842 DVDD.n17841 0.00277096
R11846 DVDD.n17780 DVDD.n17779 0.00277096
R11847 DVDD.n17975 DVDD.n17974 0.00277096
R11848 DVDD.n18149 DVDD.n18148 0.00277096
R11849 DVDD.n789 DVDD.n788 0.00277096
R11850 DVDD.n18053 DVDD.n18052 0.00277096
R11851 DVDD.n17875 DVDD.n17874 0.00277096
R11852 DVDD.n17923 DVDD.n17922 0.00277096
R11853 DVDD.n6682 DVDD.n6681 0.00277096
R11854 DVDD.n6287 DVDD.n6286 0.00277096
R11855 DVDD.n6210 DVDD.n6209 0.00277096
R11856 DVDD.n6134 DVDD.n6133 0.00277096
R11857 DVDD.n4426 DVDD.n4425 0.00277096
R11858 DVDD.n4427 DVDD.n4426 0.00277096
R11859 DVDD.n6288 DVDD.n6287 0.00277096
R11860 DVDD.n6683 DVDD.n6682 0.00277096
R11861 DVDD.n6135 DVDD.n6134 0.00277096
R11862 DVDD.n6120 DVDD.n4551 0.00277096
R11863 DVDD.n6211 DVDD.n6210 0.00277096
R11864 DVDD.n9650 DVDD.n9649 0.00277096
R11865 DVDD.n9073 DVDD.n9072 0.00277096
R11866 DVDD.n8912 DVDD.n8911 0.00277096
R11867 DVDD.n8836 DVDD.n8835 0.00277096
R11868 DVDD.n8700 DVDD.n8699 0.00277096
R11869 DVDD.n9651 DVDD.n9650 0.00277096
R11870 DVDD.n8837 DVDD.n8836 0.00277096
R11871 DVDD.n8701 DVDD.n8700 0.00277096
R11872 DVDD.n9074 DVDD.n9073 0.00277096
R11873 DVDD.n8822 DVDD.n8818 0.00277096
R11874 DVDD.n8913 DVDD.n8912 0.00277096
R11875 DVDD.n15953 DVDD.n15952 0.00275941
R11876 DVDD.n9483 DVDD.n9482 0.00275941
R11877 DVDD.n9476 DVDD.n9475 0.00275941
R11878 DVDD.n8010 DVDD.n8009 0.00275941
R11879 DVDD.n8014 DVDD.n8013 0.00275941
R11880 DVDD.n7702 DVDD.n7701 0.00275
R11881 DVDD.n3694 DVDD.n3693 0.00275
R11882 DVDD.n18540 DVDD.n18539 0.00275
R11883 DVDD.n2946 DVDD.n2945 0.00275
R11884 DVDD.n2956 DVDD.n2955 0.00275
R11885 DVDD.n9804 DVDD.n9803 0.00275
R11886 DVDD.n9361 DVDD.n9360 0.00275
R11887 DVDD.n9358 DVDD.n9357 0.00275
R11888 DVDD.n9355 DVDD.n9354 0.00275
R11889 DVDD.n9352 DVDD.n9351 0.00275
R11890 DVDD.n9349 DVDD.n9348 0.00275
R11891 DVDD.n9346 DVDD.n9345 0.00275
R11892 DVDD.n9343 DVDD.n9342 0.00275
R11893 DVDD.n9340 DVDD.n9339 0.00275
R11894 DVDD.n9337 DVDD.n9336 0.00275
R11895 DVDD.n9334 DVDD.n9333 0.00275
R11896 DVDD.n9331 DVDD.n9330 0.00275
R11897 DVDD.n9328 DVDD.n9327 0.00275
R11898 DVDD.n9325 DVDD.n9324 0.00275
R11899 DVDD.n9322 DVDD.n9321 0.00275
R11900 DVDD.n9319 DVDD.n9318 0.00275
R11901 DVDD.n2184 DVDD.n2183 0.00275
R11902 DVDD.n2194 DVDD.n2193 0.00275
R11903 DVDD.n2250 DVDD.n2249 0.00275
R11904 DVDD.n18909 DVDD.n18908 0.00275
R11905 DVDD.n7067 DVDD.n7066 0.00275
R11906 DVDD.n6811 DVDD.n6810 0.00275
R11907 DVDD.n1900 DVDD.n1899 0.00275
R11908 DVDD.n3814 DVDD.n3813 0.00275
R11909 DVDD.n19963 DVDD.n19962 0.00275
R11910 DVDD.n19973 DVDD.n19972 0.00275
R11911 DVDD.n20029 DVDD.n20028 0.00275
R11912 DVDD.n19027 DVDD.n19026 0.00275
R11913 DVDD.n4647 DVDD.n4646 0.00275
R11914 DVDD.n4848 DVDD.n4847 0.00275
R11915 DVDD.n19678 DVDD.n19677 0.00275
R11916 DVDD.n982 DVDD.n981 0.00275
R11917 DVDD.n972 DVDD.n971 0.00275
R11918 DVDD.n937 DVDD.n936 0.00275
R11919 DVDD.n19236 DVDD.n19235 0.00275
R11920 DVDD.n18323 DVDD.n18322 0.00275
R11921 DVDD.n18998 DVDD.n18997 0.00275
R11922 DVDD.n7220 DVDD.n7219 0.00275
R11923 DVDD.n10077 DVDD.n10076 0.00275
R11924 DVDD.n7121 DVDD.n7120 0.00275
R11925 DVDD.n1813 DVDD.n1812 0.00275
R11926 DVDD.n1835 DVDD.n1834 0.00275
R11927 DVDD.n7578 DVDD.n7577 0.00275
R11928 DVDD.n19613 DVDD.n19612 0.00275
R11929 DVDD.n7534 DVDD.n7533 0.00275
R11930 DVDD.n2823 DVDD.n2822 0.00275
R11931 DVDD.n861 DVDD.n860 0.00275
R11932 DVDD.n11905 DVDD.n11904 0.00275
R11933 DVDD.n1323 DVDD.n1322 0.00275
R11934 DVDD.n14850 DVDD.n14849 0.00275
R11935 DVDD.n15079 DVDD.n15078 0.00275
R11936 DVDD.n10716 DVDD.n10691 0.00275
R11937 DVDD.n10484 DVDD.n10466 0.00275
R11938 DVDD.n10697 DVDD.n10696 0.00275
R11939 DVDD.n10601 DVDD.n10600 0.00275
R11940 DVDD.n10633 DVDD.n10632 0.00275
R11941 DVDD.n10451 DVDD.n10386 0.00275
R11942 DVDD.n13272 DVDD.n13271 0.00275
R11943 DVDD.n13269 DVDD.n13268 0.00275
R11944 DVDD.n13266 DVDD.n13265 0.00275
R11945 DVDD.n13263 DVDD.n13262 0.00275
R11946 DVDD.n13260 DVDD.n13259 0.00275
R11947 DVDD.n13257 DVDD.n13256 0.00275
R11948 DVDD.n13254 DVDD.n13253 0.00275
R11949 DVDD.n13251 DVDD.n13250 0.00275
R11950 DVDD.n13248 DVDD.n13247 0.00275
R11951 DVDD.n13245 DVDD.n13244 0.00275
R11952 DVDD.n13242 DVDD.n13241 0.00275
R11953 DVDD.n13239 DVDD.n13238 0.00275
R11954 DVDD.n13236 DVDD.n13235 0.00275
R11955 DVDD.n13233 DVDD.n13232 0.00275
R11956 DVDD.n13230 DVDD.n13229 0.00275
R11957 DVDD.n3444 DVDD.n3443 0.00275
R11958 DVDD.n3420 DVDD.n3419 0.00275
R11959 DVDD.n3416 DVDD.n3415 0.00275
R11960 DVDD.n3583 DVDD.n3582 0.00275
R11961 DVDD.n3601 DVDD.n3600 0.00275
R11962 DVDD.n7810 DVDD.n7809 0.00275
R11963 DVDD.n3280 DVDD.n3279 0.00275
R11964 DVDD.n3625 DVDD.n3624 0.00275
R11965 DVDD.n7291 DVDD.n7290 0.00275
R11966 DVDD.n4319 DVDD.n4318 0.00274945
R11967 DVDD.n4290 DVDD.n4289 0.00274945
R11968 DVDD.n4265 DVDD.n4264 0.00274945
R11969 DVDD.n3117 DVDD.n3116 0.00270694
R11970 DVDD.n3118 DVDD.n3117 0.00270694
R11971 DVDD.n16059 DVDD.n16058 0.00269392
R11972 DVDD.n16060 DVDD.n16059 0.00269392
R11973 DVDD.n15671 DVDD.n15670 0.00269392
R11974 DVDD.n15672 DVDD.n15671 0.00269392
R11975 DVDD.n9398 DVDD.n9397 0.00269392
R11976 DVDD.n8356 DVDD.n8355 0.00269392
R11977 DVDD.n9399 DVDD.n9398 0.00269392
R11978 DVDD.n8355 DVDD.n8354 0.00269392
R11979 DVDD.n8138 DVDD.n8137 0.00269392
R11980 DVDD.n8137 DVDD.n8136 0.00269392
R11981 DVDD.n7957 DVDD.n7956 0.00269392
R11982 DVDD.n1842 DVDD.n1841 0.00269
R11983 DVDD.n7571 DVDD.n7570 0.00269
R11984 DVDD.n19620 DVDD.n19619 0.00269
R11985 DVDD.n7527 DVDD.n7526 0.00269
R11986 DVDD.n18256 DVDD.n18255 0.00269
R11987 DVDD.n16259 DVDD.n16258 0.00269
R11988 DVDD.n16196 DVDD.n16195 0.00269
R11989 DVDD.n15561 DVDD.n15560 0.00269
R11990 DVDD.n15776 DVDD.n15775 0.00269
R11991 DVDD.n15839 DVDD.n15838 0.00269
R11992 DVDD.n14781 DVDD.n14780 0.00269
R11993 DVDD.n12078 DVDD.n12077 0.00268244
R11994 DVDD.n13361 DVDD.n13360 0.00268244
R11995 DVDD.n12077 DVDD.n12076 0.00268244
R11996 DVDD.n13360 DVDD.n13359 0.00268244
R11997 DVDD.n13527 DVDD.n13526 0.00268244
R11998 DVDD.n13579 DVDD.n13578 0.00268244
R11999 DVDD.n13585 DVDD.n13584 0.00268244
R12000 DVDD.n13660 DVDD.n13659 0.00268244
R12001 DVDD.n13666 DVDD.n13665 0.00268244
R12002 DVDD.n15427 DVDD.n15426 0.00268244
R12003 DVDD.n15435 DVDD.n15434 0.00268244
R12004 DVDD.n14676 DVDD.n14675 0.00268244
R12005 DVDD.n14594 DVDD.n14593 0.00268244
R12006 DVDD.n14539 DVDD.n14538 0.00268244
R12007 DVDD.n14531 DVDD.n14530 0.00268244
R12008 DVDD.n14451 DVDD.n14450 0.00268244
R12009 DVDD.n14429 DVDD.n14428 0.00268244
R12010 DVDD.n14452 DVDD.n14451 0.00268244
R12011 DVDD.n14540 DVDD.n14539 0.00268244
R12012 DVDD.n14677 DVDD.n14676 0.00268244
R12013 DVDD.n15426 DVDD.n15425 0.00268244
R12014 DVDD.n15434 DVDD.n15433 0.00268244
R12015 DVDD.n14593 DVDD.n14592 0.00268244
R12016 DVDD.n14430 DVDD.n14429 0.00268244
R12017 DVDD.n14532 DVDD.n14531 0.00268244
R12018 DVDD.n5493 DVDD.n5492 0.00268244
R12019 DVDD.n5672 DVDD.n5671 0.00268244
R12020 DVDD.n6095 DVDD.n6094 0.00268244
R12021 DVDD.n6019 DVDD.n6018 0.00268244
R12022 DVDD.n5987 DVDD.n5986 0.00268244
R12023 DVDD.n5640 DVDD.n5639 0.00268244
R12024 DVDD.n5646 DVDD.n5645 0.00268244
R12025 DVDD.n5671 DVDD.n5670 0.00268244
R12026 DVDD.n6094 DVDD.n6093 0.00268244
R12027 DVDD.n6020 DVDD.n6019 0.00268244
R12028 DVDD.n5988 DVDD.n5987 0.00268244
R12029 DVDD.n12970 DVDD.n12969 0.00268244
R12030 DVDD.n12776 DVDD.n12775 0.00268244
R12031 DVDD.n12726 DVDD.n12725 0.00268244
R12032 DVDD.n12670 DVDD.n12669 0.00268244
R12033 DVDD.n12650 DVDD.n12649 0.00268244
R12034 DVDD.n12651 DVDD.n12650 0.00268244
R12035 DVDD.n12671 DVDD.n12670 0.00268244
R12036 DVDD.n12727 DVDD.n12726 0.00268244
R12037 DVDD.n12797 DVDD.n12796 0.00268244
R12038 DVDD.n12791 DVDD.n12790 0.00268244
R12039 DVDD.n12775 DVDD.n12768 0.00268244
R12040 DVDD.n18170 DVDD.n18169 0.00268244
R12041 DVDD.n17953 DVDD.n17952 0.00268244
R12042 DVDD.n17820 DVDD.n17819 0.00268244
R12043 DVDD.n17803 DVDD.n17802 0.00268244
R12044 DVDD.n18032 DVDD.n18031 0.00268244
R12045 DVDD.n18176 DVDD.n18175 0.00268244
R12046 DVDD.n17821 DVDD.n17820 0.00268244
R12047 DVDD.n17804 DVDD.n17803 0.00268244
R12048 DVDD.n17896 DVDD.n17895 0.00268244
R12049 DVDD.n17902 DVDD.n17901 0.00268244
R12050 DVDD.n17954 DVDD.n17953 0.00268244
R12051 DVDD.n6265 DVDD.n6264 0.00268244
R12052 DVDD.n6176 DVDD.n6175 0.00268244
R12053 DVDD.n6168 DVDD.n6167 0.00268244
R12054 DVDD.n6152 DVDD.n6151 0.00268244
R12055 DVDD.n4544 DVDD.n4543 0.00268244
R12056 DVDD.n4470 DVDD.n4469 0.00268244
R12057 DVDD.n4450 DVDD.n4449 0.00268244
R12058 DVDD.n4471 DVDD.n4470 0.00268244
R12059 DVDD.n6266 DVDD.n6265 0.00268244
R12060 DVDD.n6177 DVDD.n6176 0.00268244
R12061 DVDD.n6153 DVDD.n6152 0.00268244
R12062 DVDD.n4451 DVDD.n4450 0.00268244
R12063 DVDD.n4545 DVDD.n4544 0.00268244
R12064 DVDD.n6169 DVDD.n6168 0.00268244
R12065 DVDD.n9052 DVDD.n9051 0.00268244
R12066 DVDD.n8878 DVDD.n8877 0.00268244
R12067 DVDD.n8870 DVDD.n8869 0.00268244
R12068 DVDD.n8854 DVDD.n8853 0.00268244
R12069 DVDD.n8811 DVDD.n8810 0.00268244
R12070 DVDD.n8756 DVDD.n8755 0.00268244
R12071 DVDD.n8724 DVDD.n8723 0.00268244
R12072 DVDD.n8879 DVDD.n8878 0.00268244
R12073 DVDD.n8855 DVDD.n8854 0.00268244
R12074 DVDD.n8757 DVDD.n8756 0.00268244
R12075 DVDD.n9051 DVDD.n9050 0.00268244
R12076 DVDD.n8725 DVDD.n8724 0.00268244
R12077 DVDD.n8812 DVDD.n8811 0.00268244
R12078 DVDD.n8871 DVDD.n8870 0.00268244
R12079 DVDD.n7739 DVDD.n7738 0.00266
R12080 DVDD.n7735 DVDD.n7734 0.00266
R12081 DVDD.n7764 DVDD.n7763 0.00266
R12082 DVDD.n3455 DVDD.n3454 0.00266
R12083 DVDD.n3572 DVDD.n3571 0.00266
R12084 DVDD.n2903 DVDD.n2902 0.00266
R12085 DVDD.n2900 DVDD.n2899 0.00266
R12086 DVDD.n2897 DVDD.n2896 0.00266
R12087 DVDD.n2894 DVDD.n2893 0.00266
R12088 DVDD.n2891 DVDD.n2890 0.00266
R12089 DVDD.n2888 DVDD.n2887 0.00266
R12090 DVDD.n2885 DVDD.n2884 0.00266
R12091 DVDD.n2882 DVDD.n2881 0.00266
R12092 DVDD.n2879 DVDD.n2878 0.00266
R12093 DVDD.n2876 DVDD.n2875 0.00266
R12094 DVDD.n2873 DVDD.n2872 0.00266
R12095 DVDD.n9961 DVDD.n9960 0.00266
R12096 DVDD.n9762 DVDD.n9761 0.00266
R12097 DVDD.n9774 DVDD.n9773 0.00266
R12098 DVDD.n9793 DVDD.n9792 0.00266
R12099 DVDD.n7912 DVDD.n7911 0.00266
R12100 DVDD.n9252 DVDD.n9251 0.00266
R12101 DVDD.n9275 DVDD.n9274 0.00266
R12102 DVDD.n9294 DVDD.n9293 0.00266
R12103 DVDD.n9306 DVDD.n9305 0.00266
R12104 DVDD.n2056 DVDD.n2055 0.00266
R12105 DVDD.n2210 DVDD.n2209 0.00266
R12106 DVDD.n7101 DVDD.n7100 0.00266
R12107 DVDD.n7034 DVDD.n7033 0.00266
R12108 DVDD.n6944 DVDD.n6943 0.00266
R12109 DVDD.n6853 DVDD.n6852 0.00266
R12110 DVDD.n6841 DVDD.n6840 0.00266
R12111 DVDD.n6822 DVDD.n6821 0.00266
R12112 DVDD.n6543 DVDD.n6542 0.00266
R12113 DVDD.n1863 DVDD.n1862 0.00266
R12114 DVDD.n3990 DVDD.n3989 0.00266
R12115 DVDD.n3967 DVDD.n3966 0.00266
R12116 DVDD.n3948 DVDD.n3947 0.00266
R12117 DVDD.n3936 DVDD.n3935 0.00266
R12118 DVDD.n19834 DVDD.n19833 0.00266
R12119 DVDD.n19989 DVDD.n19988 0.00266
R12120 DVDD.n3880 DVDD.n3879 0.00266
R12121 DVDD.n4614 DVDD.n4613 0.00266
R12122 DVDD.n4718 DVDD.n4717 0.00266
R12123 DVDD.n4890 DVDD.n4889 0.00266
R12124 DVDD.n4878 DVDD.n4877 0.00266
R12125 DVDD.n4859 DVDD.n4858 0.00266
R12126 DVDD.n5134 DVDD.n5133 0.00266
R12127 DVDD.n19641 DVDD.n19640 0.00266
R12128 DVDD.n5295 DVDD.n5294 0.00266
R12129 DVDD.n5272 DVDD.n5271 0.00266
R12130 DVDD.n5253 DVDD.n5252 0.00266
R12131 DVDD.n5241 DVDD.n5240 0.00266
R12132 DVDD.n1542 DVDD.n1541 0.00266
R12133 DVDD.n1677 DVDD.n1676 0.00266
R12134 DVDD.n1025 DVDD.n1024 0.00266
R12135 DVDD.n1028 DVDD.n1027 0.00266
R12136 DVDD.n1031 DVDD.n1030 0.00266
R12137 DVDD.n1034 DVDD.n1033 0.00266
R12138 DVDD.n1037 DVDD.n1036 0.00266
R12139 DVDD.n1040 DVDD.n1039 0.00266
R12140 DVDD.n1043 DVDD.n1042 0.00266
R12141 DVDD.n1046 DVDD.n1045 0.00266
R12142 DVDD.n1049 DVDD.n1048 0.00266
R12143 DVDD.n1052 DVDD.n1051 0.00266
R12144 DVDD.n1055 DVDD.n1054 0.00266
R12145 DVDD.n11544 DVDD.n11543 0.00266
R12146 DVDD.n18279 DVDD.n18278 0.00266
R12147 DVDD.n18290 DVDD.n18289 0.00266
R12148 DVDD.n18276 DVDD.n18275 0.00266
R12149 DVDD.n18883 DVDD.n18882 0.00266
R12150 DVDD.n19132 DVDD.n19131 0.00266
R12151 DVDD.n19413 DVDD.n19412 0.00266
R12152 DVDD.n11863 DVDD.n11862 0.00266
R12153 DVDD.n11875 DVDD.n11874 0.00266
R12154 DVDD.n11894 DVDD.n11893 0.00266
R12155 DVDD.n1286 DVDD.n1285 0.00266
R12156 DVDD.n11314 DVDD.n11313 0.00266
R12157 DVDD.n14951 DVDD.n14950 0.00266
R12158 DVDD.n13163 DVDD.n13162 0.00266
R12159 DVDD.n13186 DVDD.n13185 0.00266
R12160 DVDD.n13205 DVDD.n13204 0.00266
R12161 DVDD.n13217 DVDD.n13216 0.00266
R12162 DVDD.n11009 DVDD.n11008 0.00266
R12163 DVDD.n16139 DVDD.n16138 0.00266
R12164 DVDD.n3317 DVDD.n3316 0.00266
R12165 DVDD.n18420 DVDD.n18419 0.00266
R12166 DVDD.n12357 DVDD.n12356 0.00265142
R12167 DVDD.n7662 DVDD.n7624 0.00263
R12168 DVDD.n10339 DVDD.n10338 0.00263
R12169 DVDD.n10733 DVDD.n10382 0.00263
R12170 DVDD.n10503 DVDD.n10502 0.00263
R12171 DVDD.n10431 DVDD.n10430 0.00263
R12172 DVDD.n16495 DVDD.n16494 0.00263
R12173 DVDD.n17160 DVDD.n17159 0.00263
R12174 DVDD.n17114 DVDD.n17113 0.00263
R12175 DVDD.n17064 DVDD.n17063 0.00263
R12176 DVDD.n16839 DVDD.n16838 0.00263
R12177 DVDD.n16871 DVDD.n16870 0.00263
R12178 DVDD.n16717 DVDD.n16716 0.00263
R12179 DVDD.n16741 DVDD.n16740 0.00263
R12180 DVDD.n16548 DVDD.n16547 0.00263
R12181 DVDD.n16573 DVDD.n16572 0.00263
R12182 DVDD.n8316 DVDD.n8315 0.0026295
R12183 DVDD.n1225 DVDD.n1224 0.00262598
R12184 DVDD.n1565 DVDD.n1564 0.00262598
R12185 DVDD.n922 DVDD.n921 0.00262598
R12186 DVDD.n10161 DVDD.n10160 0.00262598
R12187 DVDD.n11440 DVDD.n11439 0.00262598
R12188 DVDD.n12065 DVDD.n12064 0.00262598
R12189 DVDD.n12070 DVDD.n12069 0.00262598
R12190 DVDD.n12288 DVDD.n12287 0.00262598
R12191 DVDD.n12281 DVDD.n12280 0.00262598
R12192 DVDD.n13709 DVDD.n13708 0.00262598
R12193 DVDD.n2806 DVDD.n2805 0.00262598
R12194 DVDD.n18470 DVDD.n18469 0.00262598
R12195 DVDD.n10065 DVDD.n10064 0.00262598
R12196 DVDD.n15503 DVDD.n15502 0.00262598
R12197 DVDD.n14359 DVDD.n14358 0.00262598
R12198 DVDD.n19687 DVDD.n19686 0.00262598
R12199 DVDD.n19912 DVDD.n19911 0.00262598
R12200 DVDD.n20064 DVDD.n20063 0.00262598
R12201 DVDD.n20065 DVDD.n20064 0.00262598
R12202 DVDD.n20210 DVDD.n20176 0.00262598
R12203 DVDD.n19064 DVDD.n19063 0.00262598
R12204 DVDD.n3866 DVDD.n3865 0.00262598
R12205 DVDD.n4652 DVDD.n4610 0.00262598
R12206 DVDD.n4811 DVDD.n4810 0.00262598
R12207 DVDD.n4817 DVDD.n4816 0.00262598
R12208 DVDD.n4938 DVDD.n4937 0.00262598
R12209 DVDD.n4941 DVDD.n4940 0.00262598
R12210 DVDD.n5005 DVDD.n5004 0.00262598
R12211 DVDD.n5007 DVDD.n5006 0.00262598
R12212 DVDD.n5171 DVDD.n5170 0.00262598
R12213 DVDD.n5181 DVDD.n5180 0.00262598
R12214 DVDD.n5198 DVDD.n5197 0.00262598
R12215 DVDD.n5200 DVDD.n5199 0.00262598
R12216 DVDD.n5350 DVDD.n5349 0.00262598
R12217 DVDD.n5374 DVDD.n5373 0.00262598
R12218 DVDD.n5441 DVDD.n5440 0.00262598
R12219 DVDD.n5465 DVDD.n5464 0.00262598
R12220 DVDD.n6100 DVDD.n6099 0.00262598
R12221 DVDD.n5923 DVDD.n5922 0.00262598
R12222 DVDD.n1332 DVDD.n1331 0.00262598
R12223 DVDD.n1465 DVDD.n1464 0.00262598
R12224 DVDD.n1709 DVDD.n1708 0.00262598
R12225 DVDD.n1708 DVDD.n1707 0.00262598
R12226 DVDD.n289 DVDD.n288 0.00262598
R12227 DVDD.n19446 DVDD.n19445 0.00262598
R12228 DVDD.n10113 DVDD.n10112 0.00262598
R12229 DVDD.n11359 DVDD.n11358 0.00262598
R12230 DVDD.n11637 DVDD.n11636 0.00262598
R12231 DVDD.n11643 DVDD.n11642 0.00262598
R12232 DVDD.n11815 DVDD.n11814 0.00262598
R12233 DVDD.n11812 DVDD.n11811 0.00262598
R12234 DVDD.n11749 DVDD.n11748 0.00262598
R12235 DVDD.n11747 DVDD.n11746 0.00262598
R12236 DVDD.n12352 DVDD.n12351 0.00262598
R12237 DVDD.n12361 DVDD.n12360 0.00262598
R12238 DVDD.n12378 DVDD.n12377 0.00262598
R12239 DVDD.n12380 DVDD.n12379 0.00262598
R12240 DVDD.n13110 DVDD.n13109 0.00262598
R12241 DVDD.n13086 DVDD.n13085 0.00262598
R12242 DVDD.n13022 DVDD.n13021 0.00262598
R12243 DVDD.n12998 DVDD.n12997 0.00262598
R12244 DVDD.n12732 DVDD.n12731 0.00262598
R12245 DVDD.n12586 DVDD.n12585 0.00262598
R12246 DVDD.n838 DVDD.n837 0.00262598
R12247 DVDD.n19166 DVDD.n19165 0.00262598
R12248 DVDD.n10097 DVDD.n10096 0.00262598
R12249 DVDD.n18108 DVDD.n18107 0.00262598
R12250 DVDD.n17739 DVDD.n17738 0.00262598
R12251 DVDD.n1909 DVDD.n1908 0.00262598
R12252 DVDD.n2133 DVDD.n2132 0.00262598
R12253 DVDD.n2285 DVDD.n2284 0.00262598
R12254 DVDD.n2286 DVDD.n2285 0.00262598
R12255 DVDD.n19595 DVDD.n19561 0.00262598
R12256 DVDD.n18956 DVDD.n18955 0.00262598
R12257 DVDD.n7087 DVDD.n7086 0.00262598
R12258 DVDD.n7073 DVDD.n7072 0.00262598
R12259 DVDD.n6873 DVDD.n6872 0.00262598
R12260 DVDD.n6867 DVDD.n6866 0.00262598
R12261 DVDD.n6746 DVDD.n6745 0.00262598
R12262 DVDD.n6743 DVDD.n6742 0.00262598
R12263 DVDD.n6679 DVDD.n6678 0.00262598
R12264 DVDD.n6677 DVDD.n6676 0.00262598
R12265 DVDD.n6511 DVDD.n6510 0.00262598
R12266 DVDD.n6501 DVDD.n6500 0.00262598
R12267 DVDD.n6484 DVDD.n6483 0.00262598
R12268 DVDD.n6482 DVDD.n6481 0.00262598
R12269 DVDD.n6411 DVDD.n6410 0.00262598
R12270 DVDD.n6387 DVDD.n6386 0.00262598
R12271 DVDD.n6320 DVDD.n6319 0.00262598
R12272 DVDD.n6296 DVDD.n6295 0.00262598
R12273 DVDD.n4380 DVDD.n4379 0.00262598
R12274 DVDD.n3271 DVDD.n3270 0.00262598
R12275 DVDD.n3532 DVDD.n3531 0.00262598
R12276 DVDD.n3729 DVDD.n3728 0.00262598
R12277 DVDD.n3730 DVDD.n3729 0.00262598
R12278 DVDD.n3775 DVDD.n3774 0.00262598
R12279 DVDD.n18793 DVDD.n18792 0.00262598
R12280 DVDD.n7145 DVDD.n7144 0.00262598
R12281 DVDD.n10049 DVDD.n10048 0.00262598
R12282 DVDD.n7893 DVDD.n7892 0.00262598
R12283 DVDD.n7899 DVDD.n7898 0.00262598
R12284 DVDD.n9714 DVDD.n9713 0.00262598
R12285 DVDD.n9711 DVDD.n9710 0.00262598
R12286 DVDD.n9647 DVDD.n9646 0.00262598
R12287 DVDD.n9645 DVDD.n9644 0.00262598
R12288 DVDD.n8372 DVDD.n8371 0.00262598
R12289 DVDD.n8382 DVDD.n8381 0.00262598
R12290 DVDD.n8399 DVDD.n8398 0.00262598
R12291 DVDD.n8401 DVDD.n8400 0.00262598
R12292 DVDD.n9197 DVDD.n9196 0.00262598
R12293 DVDD.n9173 DVDD.n9172 0.00262598
R12294 DVDD.n9106 DVDD.n9105 0.00262598
R12295 DVDD.n9082 DVDD.n9081 0.00262598
R12296 DVDD.n8654 DVDD.n8653 0.00262598
R12297 DVDD.n15265 DVDD.n15264 0.00261313
R12298 DVDD.n19518 DVDD.n19517 0.0026
R12299 DVDD.n20133 DVDD.n20132 0.0026
R12300 DVDD.n182 DVDD.n181 0.0026
R12301 DVDD.n173 DVDD.n172 0.0026
R12302 DVDD.n14959 DVDD.n14958 0.0026
R12303 DVDD.n15038 DVDD.n15037 0.0026
R12304 DVDD.n15323 DVDD.n15322 0.0026
R12305 DVDD.n15368 DVDD.n15366 0.0026
R12306 DVDD.n15344 DVDD.n15343 0.0026
R12307 DVDD.n11019 DVDD.n11018 0.0026
R12308 DVDD.n11075 DVDD.n11074 0.0026
R12309 DVDD.n15526 DVDD.n15525 0.0026
R12310 DVDD.n11177 DVDD.n11172 0.0026
R12311 DVDD.n11149 DVDD.n11148 0.0026
R12312 DVDD.n16320 DVDD.n16319 0.0026
R12313 DVDD.n16376 DVDD.n16375 0.0026
R12314 DVDD.n16354 DVDD.n16353 0.0026
R12315 DVDD.n15746 DVDD.n15745 0.0026
R12316 DVDD.n15710 DVDD.n15709 0.0026
R12317 DVDD.n16106 DVDD.n16105 0.0026
R12318 DVDD.n16068 DVDD.n15919 0.0026
R12319 DVDD.n18717 DVDD.n18716 0.0026
R12320 DVDD.n18701 DVDD.n18700 0.0026
R12321 DVDD.n15982 DVDD.n15981 0.00259985
R12322 DVDD.n15983 DVDD.n15982 0.00259985
R12323 DVDD.n9430 DVDD.n9429 0.00259985
R12324 DVDD.n9431 DVDD.n9430 0.00259985
R12325 DVDD.n8112 DVDD.n8111 0.00259985
R12326 DVDD.n8111 DVDD.n8110 0.00259985
R12327 DVDD.n19712 DVDD.n19711 0.00259415
R12328 DVDD.n5029 DVDD.n5028 0.00259404
R12329 DVDD.n13056 DVDD.n13055 0.00259404
R12330 DVDD.n6355 DVDD.n6354 0.00259404
R12331 DVDD.n9141 DVDD.n9140 0.00259404
R12332 DVDD.n12012 DVDD.n12011 0.00259392
R12333 DVDD.n13310 DVDD.n13309 0.00259392
R12334 DVDD.n13552 DVDD.n13551 0.00259392
R12335 DVDD.n13633 DVDD.n13632 0.00259392
R12336 DVDD.n12011 DVDD.n12010 0.00259392
R12337 DVDD.n1178 DVDD.n1177 0.00259392
R12338 DVDD.n13309 DVDD.n13308 0.00259392
R12339 DVDD.n12204 DVDD.n12203 0.00259392
R12340 DVDD.n13551 DVDD.n13550 0.00259392
R12341 DVDD.n13632 DVDD.n13631 0.00259392
R12342 DVDD.n2745 DVDD.n2744 0.00259392
R12343 DVDD.n2786 DVDD.n2785 0.00259392
R12344 DVDD.n15397 DVDD.n15396 0.00259392
R12345 DVDD.n14706 DVDD.n14705 0.00259392
R12346 DVDD.n14623 DVDD.n14622 0.00259392
R12347 DVDD.n14569 DVDD.n14568 0.00259392
R12348 DVDD.n14481 DVDD.n14480 0.00259392
R12349 DVDD.n14482 DVDD.n14481 0.00259392
R12350 DVDD.n14570 DVDD.n14569 0.00259392
R12351 DVDD.n14624 DVDD.n14623 0.00259392
R12352 DVDD.n15396 DVDD.n15395 0.00259392
R12353 DVDD.n2785 DVDD.n2784 0.00259392
R12354 DVDD.n14707 DVDD.n14706 0.00259392
R12355 DVDD.n2744 DVDD.n2743 0.00259392
R12356 DVDD.n5219 DVDD.n5218 0.00259392
R12357 DVDD.n5462 DVDD.n5461 0.00259392
R12358 DVDD.n6077 DVDD.n6076 0.00259392
R12359 DVDD.n6078 DVDD.n6077 0.00259392
R12360 DVDD.n5461 DVDD.n5460 0.00259392
R12361 DVDD.n19734 DVDD.n19733 0.00259392
R12362 DVDD.n5218 DVDD.n5217 0.00259392
R12363 DVDD.n12399 DVDD.n12398 0.00259392
R12364 DVDD.n13002 DVDD.n13001 0.00259392
R12365 DVDD.n12709 DVDD.n12708 0.00259392
R12366 DVDD.n11732 DVDD.n11731 0.00259392
R12367 DVDD.n12398 DVDD.n12397 0.00259392
R12368 DVDD.n13001 DVDD.n13000 0.00259392
R12369 DVDD.n12710 DVDD.n12709 0.00259392
R12370 DVDD.n783 DVDD.n782 0.00259392
R12371 DVDD.n820 DVDD.n819 0.00259392
R12372 DVDD.n18203 DVDD.n18202 0.00259392
R12373 DVDD.n18059 DVDD.n18058 0.00259392
R12374 DVDD.n17981 DVDD.n17980 0.00259392
R12375 DVDD.n17929 DVDD.n17928 0.00259392
R12376 DVDD.n17848 DVDD.n17847 0.00259392
R12377 DVDD.n17982 DVDD.n17981 0.00259392
R12378 DVDD.n18204 DVDD.n18203 0.00259392
R12379 DVDD.n819 DVDD.n818 0.00259392
R12380 DVDD.n782 DVDD.n781 0.00259392
R12381 DVDD.n18060 DVDD.n18059 0.00259392
R12382 DVDD.n17930 DVDD.n17929 0.00259392
R12383 DVDD.n17849 DVDD.n17848 0.00259392
R12384 DVDD.n6662 DVDD.n6661 0.00259392
R12385 DVDD.n6463 DVDD.n6462 0.00259392
R12386 DVDD.n6299 DVDD.n6298 0.00259392
R12387 DVDD.n4527 DVDD.n4526 0.00259392
R12388 DVDD.n6300 DVDD.n6299 0.00259392
R12389 DVDD.n6464 DVDD.n6463 0.00259392
R12390 DVDD.n4528 DVDD.n4527 0.00259392
R12391 DVDD.n8420 DVDD.n8419 0.00259392
R12392 DVDD.n9085 DVDD.n9084 0.00259392
R12393 DVDD.n8794 DVDD.n8793 0.00259392
R12394 DVDD.n8419 DVDD.n8418 0.00259392
R12395 DVDD.n9086 DVDD.n9085 0.00259392
R12396 DVDD.n8795 DVDD.n8794 0.00259392
R12397 DVDD.n9630 DVDD.n9629 0.00259392
R12398 DVDD.n3839 DVDD.n3838 0.00258575
R12399 DVDD.n124 DVDD.n123 0.00258575
R12400 DVDD.n3371 DVDD.n3370 0.00257472
R12401 DVDD.n15981 DVDD.n15980 0.00257113
R12402 DVDD.n8247 DVDD.n8246 0.00257113
R12403 DVDD.n9432 DVDD.n9431 0.00257113
R12404 DVDD.n8113 DVDD.n8112 0.00257113
R12405 DVDD.n7937 DVDD.n7814 0.00257113
R12406 DVDD.n8074 DVDD.n8073 0.00257113
R12407 DVDD.n8078 DVDD.n8077 0.00257113
R12408 DVDD.n3677 DVDD.n3676 0.00257
R12409 DVDD.n3706 DVDD.n3705 0.00257
R12410 DVDD.n18552 DVDD.n18551 0.00257
R12411 DVDD.n2998 DVDD.n2997 0.00257
R12412 DVDD.n2919 DVDD.n2918 0.00257
R12413 DVDD.n2934 DVDD.n2933 0.00257
R12414 DVDD.n2936 DVDD.n2935 0.00257
R12415 DVDD.n7159 DVDD.n7158 0.00257
R12416 DVDD.n9387 DVDD.n9386 0.00257
R12417 DVDD.n9384 DVDD.n9383 0.00257
R12418 DVDD.n9381 DVDD.n9380 0.00257
R12419 DVDD.n9378 DVDD.n9377 0.00257
R12420 DVDD.n9375 DVDD.n9374 0.00257
R12421 DVDD.n9372 DVDD.n9371 0.00257
R12422 DVDD.n9369 DVDD.n9368 0.00257
R12423 DVDD.n9366 DVDD.n9365 0.00257
R12424 DVDD.n2025 DVDD.n2024 0.00257
R12425 DVDD.n2157 DVDD.n2156 0.00257
R12426 DVDD.n2172 DVDD.n2171 0.00257
R12427 DVDD.n2174 DVDD.n2173 0.00257
R12428 DVDD.n2233 DVDD.n2232 0.00257
R12429 DVDD.n2262 DVDD.n2261 0.00257
R12430 DVDD.n18921 DVDD.n18920 0.00257
R12431 DVDD.n6939 DVDD.n6938 0.00257
R12432 DVDD.n1888 DVDD.n1887 0.00257
R12433 DVDD.n19803 DVDD.n19802 0.00257
R12434 DVDD.n19936 DVDD.n19935 0.00257
R12435 DVDD.n19951 DVDD.n19950 0.00257
R12436 DVDD.n19953 DVDD.n19952 0.00257
R12437 DVDD.n20012 DVDD.n20011 0.00257
R12438 DVDD.n20041 DVDD.n20040 0.00257
R12439 DVDD.n19039 DVDD.n19038 0.00257
R12440 DVDD.n4713 DVDD.n4712 0.00257
R12441 DVDD.n19666 DVDD.n19665 0.00257
R12442 DVDD.n1092 DVDD.n1091 0.00257
R12443 DVDD.n1009 DVDD.n1008 0.00257
R12444 DVDD.n994 DVDD.n993 0.00257
R12445 DVDD.n992 DVDD.n991 0.00257
R12446 DVDD.n1730 DVDD.n1729 0.00257
R12447 DVDD.n949 DVDD.n948 0.00257
R12448 DVDD.n19248 DVDD.n19247 0.00257
R12449 DVDD.n11420 DVDD.n11419 0.00257
R12450 DVDD.n19546 DVDD.n19545 0.00257
R12451 DVDD.n20161 DVDD.n20160 0.00257
R12452 DVDD.n217 DVDD.n216 0.00257
R12453 DVDD.n1311 DVDD.n1310 0.00257
R12454 DVDD.n14958 DVDD.n14957 0.00257
R12455 DVDD.n15037 DVDD.n15036 0.00257
R12456 DVDD.n15322 DVDD.n15321 0.00257
R12457 DVDD.n13298 DVDD.n13297 0.00257
R12458 DVDD.n13295 DVDD.n13294 0.00257
R12459 DVDD.n13292 DVDD.n13291 0.00257
R12460 DVDD.n13289 DVDD.n13288 0.00257
R12461 DVDD.n13286 DVDD.n13285 0.00257
R12462 DVDD.n13283 DVDD.n13282 0.00257
R12463 DVDD.n13280 DVDD.n13279 0.00257
R12464 DVDD.n13277 DVDD.n13276 0.00257
R12465 DVDD.n11018 DVDD.n11017 0.00257
R12466 DVDD.n11074 DVDD.n11073 0.00257
R12467 DVDD.n15527 DVDD.n15526 0.00257
R12468 DVDD.n16994 DVDD.n16993 0.00257
R12469 DVDD.n16319 DVDD.n16318 0.00257
R12470 DVDD.n16769 DVDD.n16768 0.00257
R12471 DVDD.n16892 DVDD.n16891 0.00257
R12472 DVDD.n15747 DVDD.n15746 0.00257
R12473 DVDD.n15711 DVDD.n15710 0.00257
R12474 DVDD.n16646 DVDD.n16645 0.00257
R12475 DVDD.n16589 DVDD.n16588 0.00257
R12476 DVDD.n16107 DVDD.n16106 0.00257
R12477 DVDD.n16069 DVDD.n16068 0.00257
R12478 DVDD.n3292 DVDD.n3291 0.00257
R12479 DVDD.n18619 DVDD.n18618 0.00257
R12480 DVDD.n2468 DVDD.n2467 0.00255714
R12481 DVDD.n1787 DVDD.n1786 0.00254
R12482 DVDD DVDD.n15338 0.00254
R12483 DVDD DVDD.n11138 0.00254
R12484 DVDD DVDD.n16348 0.00254
R12485 DVDD DVDD.n15703 0.00254
R12486 DVDD.n15908 DVDD 0.00254
R12487 DVDD.n3647 DVDD.n3646 0.00254
R12488 DVDD.n3820 DVDD.n3819 0.002525
R12489 DVDD.n19003 DVDD.n19002 0.002525
R12490 DVDD.n7224 DVDD.n7223 0.002525
R12491 DVDD.n7125 DVDD.n7124 0.002525
R12492 DVDD.n2827 DVDD.n2826 0.002525
R12493 DVDD.n14856 DVDD.n14855 0.002525
R12494 DVDD.n15083 DVDD.n15082 0.002525
R12495 DVDD.n10701 DVDD.n10700 0.002525
R12496 DVDD.n10606 DVDD.n10605 0.002525
R12497 DVDD.n7295 DVDD.n7294 0.002525
R12498 DVDD.n15195 DVDD.n15194 0.00251708
R12499 DVDD.n15262 DVDD.n15261 0.00251708
R12500 DVDD.n15281 DVDD.n15279 0.00251708
R12501 DVDD.n1856 DVDD.n1855 0.00251
R12502 DVDD.n19634 DVDD.n19633 0.00251
R12503 DVDD.n7301 DVDD.n7259 0.00251
R12504 DVDD.n10733 DVDD.n10732 0.00251
R12505 DVDD.n10502 DVDD.n10501 0.00251
R12506 DVDD.n10430 DVDD.n10429 0.00251
R12507 DVDD.n10426 DVDD.n10425 0.00251
R12508 DVDD.n17159 DVDD.n17158 0.00251
R12509 DVDD.n17113 DVDD.n17112 0.00251
R12510 DVDD.n17063 DVDD.n17062 0.00251
R12511 DVDD.n17058 DVDD.n17057 0.00251
R12512 DVDD.n16879 DVDD.n16871 0.00251
R12513 DVDD.n17002 DVDD.n17001 0.00251
R12514 DVDD.n16944 DVDD.n16943 0.00251
R12515 DVDD.n16934 DVDD.n16933 0.00251
R12516 DVDD.n16718 DVDD.n16717 0.00251
R12517 DVDD.n16744 DVDD.n16741 0.00251
R12518 DVDD.n16777 DVDD.n16776 0.00251
R12519 DVDD.n16900 DVDD.n16899 0.00251
R12520 DVDD.n16549 DVDD.n16548 0.00251
R12521 DVDD.n16576 DVDD.n16573 0.00251
R12522 DVDD.n16654 DVDD.n16653 0.00251
R12523 DVDD.n16597 DVDD.n16596 0.00251
R12524 DVDD.n20339 DVDD.n20338 0.00251
R12525 DVDD.n15955 DVDD.n15954 0.00250577
R12526 DVDD.n15954 DVDD.n15953 0.00250577
R12527 DVDD.n8180 DVDD.n8179 0.00250577
R12528 DVDD.n8181 DVDD.n8180 0.00250577
R12529 DVDD.n5093 DVDD.n5092 0.00250576
R12530 DVDD.n12171 DVDD.n12170 0.0025054
R12531 DVDD.n12235 DVDD.n12234 0.0025054
R12532 DVDD.n13701 DVDD.n13700 0.0025054
R12533 DVDD.n12170 DVDD.n12169 0.0025054
R12534 DVDD.n1238 DVDD.n1237 0.0025054
R12535 DVDD.n12236 DVDD.n12235 0.0025054
R12536 DVDD.n2717 DVDD.n2716 0.0025054
R12537 DVDD.n2757 DVDD.n2756 0.0025054
R12538 DVDD.n15474 DVDD.n15473 0.0025054
R12539 DVDD.n14734 DVDD.n14733 0.0025054
R12540 DVDD.n14651 DVDD.n14650 0.0025054
R12541 DVDD.n14388 DVDD.n14387 0.0025054
R12542 DVDD.n14652 DVDD.n14651 0.0025054
R12543 DVDD.n14735 DVDD.n14734 0.0025054
R12544 DVDD.n15473 DVDD.n15472 0.0025054
R12545 DVDD.n2716 DVDD.n2715 0.0025054
R12546 DVDD.n2758 DVDD.n2757 0.0025054
R12547 DVDD.n5497 DVDD.n5496 0.0025054
R12548 DVDD.n5501 DVDD.n5500 0.0025054
R12549 DVDD.n5626 DVDD.n5625 0.0025054
R12550 DVDD.n5950 DVDD.n5949 0.0025054
R12551 DVDD.n5496 DVDD.n5495 0.0025054
R12552 DVDD.n5625 DVDD.n5624 0.0025054
R12553 DVDD.n5393 DVDD.n5392 0.0025054
R12554 DVDD.n5500 DVDD.n5499 0.0025054
R12555 DVDD.n12966 DVDD.n12965 0.0025054
R12556 DVDD.n12963 DVDD.n12962 0.0025054
R12557 DVDD.n12811 DVDD.n12810 0.0025054
R12558 DVDD.n12613 DVDD.n12612 0.0025054
R12559 DVDD.n13096 DVDD.n13095 0.0025054
R12560 DVDD.n13068 DVDD.n13067 0.0025054
R12561 DVDD.n12967 DVDD.n12966 0.0025054
R12562 DVDD.n12962 DVDD.n12961 0.0025054
R12563 DVDD.n12812 DVDD.n12811 0.0025054
R12564 DVDD.n756 DVDD.n755 0.0025054
R12565 DVDD.n794 DVDD.n793 0.0025054
R12566 DVDD.n18135 DVDD.n18134 0.0025054
R12567 DVDD.n18085 DVDD.n18084 0.0025054
R12568 DVDD.n18007 DVDD.n18006 0.0025054
R12569 DVDD.n17766 DVDD.n17765 0.0025054
R12570 DVDD.n18008 DVDD.n18007 0.0025054
R12571 DVDD.n18086 DVDD.n18085 0.0025054
R12572 DVDD.n793 DVDD.n792 0.0025054
R12573 DVDD.n18136 DVDD.n18135 0.0025054
R12574 DVDD.n757 DVDD.n756 0.0025054
R12575 DVDD.n6261 DVDD.n6260 0.0025054
R12576 DVDD.n6257 DVDD.n6256 0.0025054
R12577 DVDD.n6190 DVDD.n6189 0.0025054
R12578 DVDD.n4409 DVDD.n4408 0.0025054
R12579 DVDD.n6258 DVDD.n6257 0.0025054
R12580 DVDD.n6397 DVDD.n6396 0.0025054
R12581 DVDD.n6384 DVDD.n6383 0.0025054
R12582 DVDD.n6368 DVDD.n6367 0.0025054
R12583 DVDD.n6262 DVDD.n6261 0.0025054
R12584 DVDD.n6191 DVDD.n6190 0.0025054
R12585 DVDD.n14389 DVDD.n14388 0.0025054
R12586 DVDD.n4410 DVDD.n4409 0.0025054
R12587 DVDD.n5951 DVDD.n5950 0.0025054
R12588 DVDD.n12614 DVDD.n12613 0.0025054
R12589 DVDD.n17767 DVDD.n17766 0.0025054
R12590 DVDD.n13700 DVDD.n13699 0.0025054
R12591 DVDD.n9047 DVDD.n9046 0.0025054
R12592 DVDD.n9043 DVDD.n9042 0.0025054
R12593 DVDD.n8892 DVDD.n8891 0.0025054
R12594 DVDD.n8683 DVDD.n8682 0.0025054
R12595 DVDD.n9048 DVDD.n9047 0.0025054
R12596 DVDD.n8893 DVDD.n8892 0.0025054
R12597 DVDD.n9044 DVDD.n9043 0.0025054
R12598 DVDD.n9183 DVDD.n9182 0.0025054
R12599 DVDD.n9170 DVDD.n9169 0.0025054
R12600 DVDD.n9154 DVDD.n9153 0.0025054
R12601 DVDD.n8684 DVDD.n8683 0.0025054
R12602 DVDD.n18980 DVDD.n18979 0.00248146
R12603 DVDD.n10547 DVDD.n10546 0.00248146
R12604 DVDD.n3671 DVDD.n3670 0.00248
R12605 DVDD.n2864 DVDD.n2863 0.00248
R12606 DVDD.n2861 DVDD.n2860 0.00248
R12607 DVDD.n2858 DVDD.n2857 0.00248
R12608 DVDD.n2855 DVDD.n2854 0.00248
R12609 DVDD.n2852 DVDD.n2851 0.00248
R12610 DVDD.n2849 DVDD.n2848 0.00248
R12611 DVDD.n2846 DVDD.n2845 0.00248
R12612 DVDD.n2843 DVDD.n2842 0.00248
R12613 DVDD.n2840 DVDD.n2839 0.00248
R12614 DVDD.n2837 DVDD.n2836 0.00248
R12615 DVDD.n3004 DVDD.n3003 0.00248
R12616 DVDD.n2913 DVDD.n2912 0.00248
R12617 DVDD.n7165 DVDD.n7164 0.00248
R12618 DVDD.n7823 DVDD.n7822 0.00248
R12619 DVDD.n9772 DVDD.n9771 0.00248
R12620 DVDD.n9795 DVDD.n9794 0.00248
R12621 DVDD.n9530 DVDD.n9529 0.00248
R12622 DVDD.n9527 DVDD.n9526 0.00248
R12623 DVDD.n9254 DVDD.n9253 0.00248
R12624 DVDD.n9273 DVDD.n9272 0.00248
R12625 DVDD.n9296 DVDD.n9295 0.00248
R12626 DVDD.n6792 DVDD.n6791 0.00248
R12627 DVDD.n6843 DVDD.n6842 0.00248
R12628 DVDD.n6820 DVDD.n6819 0.00248
R12629 DVDD.n6562 DVDD.n6561 0.00248
R12630 DVDD.n6559 DVDD.n6558 0.00248
R12631 DVDD.n3988 DVDD.n3987 0.00248
R12632 DVDD.n3969 DVDD.n3968 0.00248
R12633 DVDD.n3946 DVDD.n3945 0.00248
R12634 DVDD.n4829 DVDD.n4828 0.00248
R12635 DVDD.n4880 DVDD.n4879 0.00248
R12636 DVDD.n4857 DVDD.n4856 0.00248
R12637 DVDD.n5153 DVDD.n5152 0.00248
R12638 DVDD.n5150 DVDD.n5149 0.00248
R12639 DVDD.n5293 DVDD.n5292 0.00248
R12640 DVDD.n5274 DVDD.n5273 0.00248
R12641 DVDD.n5251 DVDD.n5250 0.00248
R12642 DVDD.n1086 DVDD.n1085 0.00248
R12643 DVDD.n1015 DVDD.n1014 0.00248
R12644 DVDD.n1736 DVDD.n1735 0.00248
R12645 DVDD.n1740 DVDD.n1739 0.00248
R12646 DVDD.n1743 DVDD.n1742 0.00248
R12647 DVDD.n1780 DVDD.n1779 0.00248
R12648 DVDD.n1777 DVDD.n1776 0.00248
R12649 DVDD.n1774 DVDD.n1773 0.00248
R12650 DVDD.n1771 DVDD.n1770 0.00248
R12651 DVDD.n1768 DVDD.n1767 0.00248
R12652 DVDD.n1765 DVDD.n1764 0.00248
R12653 DVDD.n1762 DVDD.n1761 0.00248
R12654 DVDD.n1759 DVDD.n1758 0.00248
R12655 DVDD.n1756 DVDD.n1755 0.00248
R12656 DVDD.n11426 DVDD.n11425 0.00248
R12657 DVDD.n18897 DVDD.n18896 0.00248
R12658 DVDD.n19146 DVDD.n19145 0.00248
R12659 DVDD.n11348 DVDD.n11347 0.00248
R12660 DVDD.n11873 DVDD.n11872 0.00248
R12661 DVDD.n11896 DVDD.n11895 0.00248
R12662 DVDD.n12334 DVDD.n12333 0.00248
R12663 DVDD.n12331 DVDD.n12330 0.00248
R12664 DVDD.n10358 DVDD.n10356 0.00248
R12665 DVDD.n13165 DVDD.n13164 0.00248
R12666 DVDD.n13184 DVDD.n13183 0.00248
R12667 DVDD.n13207 DVDD.n13206 0.00248
R12668 DVDD.n16511 DVDD.n16510 0.00248
R12669 DVDD.n16853 DVDD.n16852 0.00248
R12670 DVDD.n16154 DVDD.n16153 0.00248
R12671 DVDD.n16272 DVDD.n16271 0.00248
R12672 DVDD.n16210 DVDD.n16209 0.00248
R12673 DVDD.n15575 DVDD.n15574 0.00248
R12674 DVDD.n15789 DVDD.n15788 0.00248
R12675 DVDD.n15852 DVDD.n15851 0.00248
R12676 DVDD.n3921 DVDD.n3920 0.00245
R12677 DVDD.n4608 DVDD.n4607 0.00245
R12678 DVDD.n18241 DVDD.n18240 0.00245
R12679 DVDD.n14797 DVDD.n14796 0.00245
R12680 DVDD.n1566 DVDD.n1565 0.00244882
R12681 DVDD.n1625 DVDD.n1624 0.00244882
R12682 DVDD.n1660 DVDD.n1659 0.00244882
R12683 DVDD.n892 DVDD.n891 0.00244882
R12684 DVDD.n19271 DVDD.n19270 0.00244882
R12685 DVDD.n19274 DVDD.n19273 0.00244882
R12686 DVDD.n19280 DVDD.n19279 0.00244882
R12687 DVDD.n19317 DVDD.n19316 0.00244882
R12688 DVDD.n19315 DVDD.n19314 0.00244882
R12689 DVDD.n11990 DVDD.n11989 0.00244882
R12690 DVDD.n12131 DVDD.n12130 0.00244882
R12691 DVDD.n12136 DVDD.n12135 0.00244882
R12692 DVDD.n12172 DVDD.n12171 0.00244882
R12693 DVDD.n12237 DVDD.n12236 0.00244882
R12694 DVDD.n13424 DVDD.n13423 0.00244882
R12695 DVDD.n13702 DVDD.n13701 0.00244882
R12696 DVDD.n2715 DVDD.n2714 0.00244882
R12697 DVDD.n2756 DVDD.n2755 0.00244882
R12698 DVDD.n2797 DVDD.n2796 0.00244882
R12699 DVDD.n18677 DVDD.n18676 0.00244882
R12700 DVDD.n10056 DVDD.n10055 0.00244882
R12701 DVDD.n15475 DVDD.n15474 0.00244882
R12702 DVDD.n14736 DVDD.n14735 0.00244882
R12703 DVDD.n14653 DVDD.n14652 0.00244882
R12704 DVDD.n14387 DVDD.n14386 0.00244882
R12705 DVDD.n19686 DVDD.n19685 0.00244882
R12706 DVDD.n19699 DVDD.n19698 0.00244882
R12707 DVDD.n19731 DVDD.n19730 0.00244882
R12708 DVDD.n19754 DVDD.n19753 0.00244882
R12709 DVDD.n19755 DVDD.n19754 0.00244882
R12710 DVDD.n19854 DVDD.n19853 0.00244882
R12711 DVDD.n19875 DVDD.n19874 0.00244882
R12712 DVDD.n20002 DVDD.n20001 0.00244882
R12713 DVDD.n20061 DVDD.n20060 0.00244882
R12714 DVDD.n19066 DVDD.n19065 0.00244882
R12715 DVDD.n19105 DVDD.n19104 0.00244882
R12716 DVDD.n4957 DVDD.n4956 0.00244882
R12717 DVDD.n4986 DVDD.n4985 0.00244882
R12718 DVDD.n5031 DVDD.n5030 0.00244882
R12719 DVDD.n5103 DVDD.n5102 0.00244882
R12720 DVDD.n5182 DVDD.n5181 0.00244882
R12721 DVDD.n5226 DVDD.n5225 0.00244882
R12722 DVDD.n5392 DVDD.n5391 0.00244882
R12723 DVDD.n5405 DVDD.n5404 0.00244882
R12724 DVDD.n5424 DVDD.n5423 0.00244882
R12725 DVDD.n5498 DVDD.n5497 0.00244882
R12726 DVDD.n6046 DVDD.n6045 0.00244882
R12727 DVDD.n6045 DVDD.n6044 0.00244882
R12728 DVDD.n6042 DVDD.n6041 0.00244882
R12729 DVDD.n5949 DVDD.n5948 0.00244882
R12730 DVDD.n1331 DVDD.n1330 0.00244882
R12731 DVDD.n1344 DVDD.n1343 0.00244882
R12732 DVDD.n1376 DVDD.n1375 0.00244882
R12733 DVDD.n1399 DVDD.n1398 0.00244882
R12734 DVDD.n1400 DVDD.n1399 0.00244882
R12735 DVDD.n1522 DVDD.n1521 0.00244882
R12736 DVDD.n1501 DVDD.n1500 0.00244882
R12737 DVDD.n1690 DVDD.n1689 0.00244882
R12738 DVDD.n1712 DVDD.n1711 0.00244882
R12739 DVDD.n19448 DVDD.n19447 0.00244882
R12740 DVDD.n10104 DVDD.n10103 0.00244882
R12741 DVDD.n11837 DVDD.n11836 0.00244882
R12742 DVDD.n11796 DVDD.n11795 0.00244882
R12743 DVDD.n11771 DVDD.n11770 0.00244882
R12744 DVDD.n11767 DVDD.n11766 0.00244882
R12745 DVDD.n11723 DVDD.n11722 0.00244882
R12746 DVDD.n11652 DVDD.n11651 0.00244882
R12747 DVDD.n12362 DVDD.n12361 0.00244882
R12748 DVDD.n12406 DVDD.n12405 0.00244882
R12749 DVDD.n13069 DVDD.n13068 0.00244882
R12750 DVDD.n13057 DVDD.n13056 0.00244882
R12751 DVDD.n12965 DVDD.n12964 0.00244882
R12752 DVDD.n12692 DVDD.n12691 0.00244882
R12753 DVDD.n12691 DVDD.n12690 0.00244882
R12754 DVDD.n12688 DVDD.n12687 0.00244882
R12755 DVDD.n12612 DVDD.n12611 0.00244882
R12756 DVDD.n755 DVDD.n754 0.00244882
R12757 DVDD.n792 DVDD.n791 0.00244882
R12758 DVDD.n829 DVDD.n828 0.00244882
R12759 DVDD.n156 DVDD.n155 0.00244882
R12760 DVDD.n10088 DVDD.n10087 0.00244882
R12761 DVDD.n18134 DVDD.n18133 0.00244882
R12762 DVDD.n18087 DVDD.n18086 0.00244882
R12763 DVDD.n18009 DVDD.n18008 0.00244882
R12764 DVDD.n17765 DVDD.n17764 0.00244882
R12765 DVDD.n1908 DVDD.n1907 0.00244882
R12766 DVDD.n1921 DVDD.n1920 0.00244882
R12767 DVDD.n1953 DVDD.n1952 0.00244882
R12768 DVDD.n1976 DVDD.n1975 0.00244882
R12769 DVDD.n1977 DVDD.n1976 0.00244882
R12770 DVDD.n2076 DVDD.n2075 0.00244882
R12771 DVDD.n2097 DVDD.n2096 0.00244882
R12772 DVDD.n2223 DVDD.n2222 0.00244882
R12773 DVDD.n2282 DVDD.n2281 0.00244882
R12774 DVDD.n18958 DVDD.n18957 0.00244882
R12775 DVDD.n6768 DVDD.n6767 0.00244882
R12776 DVDD.n6727 DVDD.n6726 0.00244882
R12777 DVDD.n6702 DVDD.n6701 0.00244882
R12778 DVDD.n6698 DVDD.n6697 0.00244882
R12779 DVDD.n6653 DVDD.n6652 0.00244882
R12780 DVDD.n6579 DVDD.n6578 0.00244882
R12781 DVDD.n6500 DVDD.n6499 0.00244882
R12782 DVDD.n6456 DVDD.n6455 0.00244882
R12783 DVDD.n6369 DVDD.n6368 0.00244882
R12784 DVDD.n6356 DVDD.n6355 0.00244882
R12785 DVDD.n6260 DVDD.n6259 0.00244882
R12786 DVDD.n4496 DVDD.n4495 0.00244882
R12787 DVDD.n4493 DVDD.n4492 0.00244882
R12788 DVDD.n4408 DVDD.n4407 0.00244882
R12789 DVDD.n3272 DVDD.n3271 0.00244882
R12790 DVDD.n3259 DVDD.n3258 0.00244882
R12791 DVDD.n3227 DVDD.n3226 0.00244882
R12792 DVDD.n3204 DVDD.n3203 0.00244882
R12793 DVDD.n3203 DVDD.n3202 0.00244882
R12794 DVDD.n3475 DVDD.n3474 0.00244882
R12795 DVDD.n3496 DVDD.n3495 0.00244882
R12796 DVDD.n3559 DVDD.n3558 0.00244882
R12797 DVDD.n3726 DVDD.n3725 0.00244882
R12798 DVDD.n18795 DVDD.n18794 0.00244882
R12799 DVDD.n7136 DVDD.n7135 0.00244882
R12800 DVDD.n9736 DVDD.n9735 0.00244882
R12801 DVDD.n9695 DVDD.n9694 0.00244882
R12802 DVDD.n9670 DVDD.n9669 0.00244882
R12803 DVDD.n9666 DVDD.n9665 0.00244882
R12804 DVDD.n9621 DVDD.n9620 0.00244882
R12805 DVDD.n9547 DVDD.n9546 0.00244882
R12806 DVDD.n8383 DVDD.n8382 0.00244882
R12807 DVDD.n8427 DVDD.n8426 0.00244882
R12808 DVDD.n9155 DVDD.n9154 0.00244882
R12809 DVDD.n9142 DVDD.n9141 0.00244882
R12810 DVDD.n9046 DVDD.n9045 0.00244882
R12811 DVDD.n8777 DVDD.n8776 0.00244882
R12812 DVDD.n8774 DVDD.n8773 0.00244882
R12813 DVDD.n8682 DVDD.n8681 0.00244882
R12814 DVDD.n9473 DVDD.n9472 0.00244595
R12815 DVDD.n15208 DVDD.n15207 0.00242102
R12816 DVDD.n15315 DVDD.n15314 0.00242
R12817 DVDD.n15535 DVDD.n15534 0.00242
R12818 DVDD.n16313 DVDD.n16312 0.00242
R12819 DVDD.n16118 DVDD.n15755 0.00242
R12820 DVDD.n16117 DVDD.n16116 0.00242
R12821 DVDD.n5577 DVDD.n5576 0.00241726
R12822 DVDD.n12850 DVDD.n12849 0.00241726
R12823 DVDD.n6230 DVDD.n6229 0.00241726
R12824 DVDD.n8932 DVDD.n8931 0.00241726
R12825 DVDD.n13493 DVDD.n13492 0.00241688
R12826 DVDD.n13494 DVDD.n13493 0.00241688
R12827 DVDD.n15502 DVDD.n15501 0.00241688
R12828 DVDD.n15501 DVDD.n15500 0.00241688
R12829 DVDD.n19879 DVDD.n19878 0.00241688
R12830 DVDD.n5030 DVDD.n5029 0.00241688
R12831 DVDD.n5064 DVDD.n5063 0.00241688
R12832 DVDD.n5924 DVDD.n5923 0.00241688
R12833 DVDD.n5063 DVDD.n5062 0.00241688
R12834 DVDD.n19900 DVDD.n19899 0.00241688
R12835 DVDD.n19878 DVDD.n19877 0.00241688
R12836 DVDD.n11690 DVDD.n11689 0.00241688
R12837 DVDD.n12587 DVDD.n12586 0.00241688
R12838 DVDD.n13055 DVDD.n13054 0.00241688
R12839 DVDD.n11691 DVDD.n11690 0.00241688
R12840 DVDD.n18109 DVDD.n18108 0.00241688
R12841 DVDD.n17740 DVDD.n17739 0.00241688
R12842 DVDD.n18110 DVDD.n18109 0.00241688
R12843 DVDD.n4381 DVDD.n4380 0.00241688
R12844 DVDD.n6354 DVDD.n6353 0.00241688
R12845 DVDD.n5925 DVDD.n5924 0.00241688
R12846 DVDD.n12588 DVDD.n12587 0.00241688
R12847 DVDD.n17741 DVDD.n17740 0.00241688
R12848 DVDD.n4382 DVDD.n4381 0.00241688
R12849 DVDD.n9586 DVDD.n9585 0.00241688
R12850 DVDD.n9140 DVDD.n9139 0.00241688
R12851 DVDD.n9587 DVDD.n9586 0.00241688
R12852 DVDD.n13710 DVDD.n13709 0.00241688
R12853 DVDD.n14361 DVDD.n14360 0.00241688
R12854 DVDD.n6618 DVDD.n6617 0.00241688
R12855 DVDD.n6619 DVDD.n6618 0.00241688
R12856 DVDD.n13711 DVDD.n13710 0.00241688
R12857 DVDD.n14360 DVDD.n14359 0.00241688
R12858 DVDD.n8655 DVDD.n8654 0.00241688
R12859 DVDD.n8656 DVDD.n8655 0.00241688
R12860 DVDD.n17245 DVDD.n17244 0.00241489
R12861 DVDD.n17412 DVDD.n17411 0.00241489
R12862 DVDD.n17595 DVDD.n17594 0.00241489
R12863 DVDD DVDD.n2651 0.00241429
R12864 DVDD.n8244 DVDD.n8243 0.00241169
R12865 DVDD.n8243 DVDD.n8242 0.00241169
R12866 DVDD.n16476 DVDD.n16475 0.00239333
R12867 DVDD.n16475 DVDD.n16474 0.00239333
R12868 DVDD.n16474 DVDD.n16473 0.00239333
R12869 DVDD.n16473 DVDD.n16472 0.00239333
R12870 DVDD.n16472 DVDD.n16471 0.00239333
R12871 DVDD.n16471 DVDD.n16470 0.00239333
R12872 DVDD.n16470 DVDD.n16469 0.00239333
R12873 DVDD.n16469 DVDD.n16468 0.00239333
R12874 DVDD.n16468 DVDD.n16467 0.00239333
R12875 DVDD.n16467 DVDD.n16466 0.00239333
R12876 DVDD.n16464 DVDD.n16463 0.00239333
R12877 DVDD.n16463 DVDD.n16462 0.00239333
R12878 DVDD.n16462 DVDD.n16461 0.00239333
R12879 DVDD.n16461 DVDD.n16460 0.00239333
R12880 DVDD.n16460 DVDD.n16459 0.00239333
R12881 DVDD.n16459 DVDD.n16458 0.00239333
R12882 DVDD.n16458 DVDD.n16457 0.00239333
R12883 DVDD.n16457 DVDD.n16456 0.00239333
R12884 DVDD.n16456 DVDD.n16455 0.00239333
R12885 DVDD.n16455 DVDD.n16454 0.00239333
R12886 DVDD.n16454 DVDD.n16453 0.00239333
R12887 DVDD.n16453 DVDD.n16452 0.00239333
R12888 DVDD.n16452 DVDD.n16451 0.00239333
R12889 DVDD.n16451 DVDD.n16450 0.00239333
R12890 DVDD.n16450 DVDD.n16449 0.00239333
R12891 DVDD.n16449 DVDD.n16448 0.00239333
R12892 DVDD.n16448 DVDD.n16447 0.00239333
R12893 DVDD.n16447 DVDD.n16446 0.00239333
R12894 DVDD.n16446 DVDD.n16445 0.00239333
R12895 DVDD.n16445 DVDD.n16444 0.00239333
R12896 DVDD.n16444 DVDD.n16443 0.00239333
R12897 DVDD.n16443 DVDD.n16442 0.00239333
R12898 DVDD.n16442 DVDD.n16441 0.00239333
R12899 DVDD.n16439 DVDD.n16438 0.00239333
R12900 DVDD.n16438 DVDD.n16437 0.00239333
R12901 DVDD.n16437 DVDD.n16436 0.00239333
R12902 DVDD.n16436 DVDD.n16435 0.00239333
R12903 DVDD.n16435 DVDD.n16434 0.00239333
R12904 DVDD.n16434 DVDD.n16433 0.00239333
R12905 DVDD.n16433 DVDD.n16432 0.00239333
R12906 DVDD.n16432 DVDD.n16431 0.00239333
R12907 DVDD.n16431 DVDD.n16430 0.00239333
R12908 DVDD.n16430 DVDD.n16429 0.00239333
R12909 DVDD.n16429 DVDD.n16428 0.00239333
R12910 DVDD.n16428 DVDD.n16427 0.00239333
R12911 DVDD.n16427 DVDD.n16426 0.00239333
R12912 DVDD.n16426 DVDD.n16425 0.00239333
R12913 DVDD.n16425 DVDD.n16424 0.00239333
R12914 DVDD.n16424 DVDD.n16423 0.00239333
R12915 DVDD.n16423 DVDD.n16422 0.00239333
R12916 DVDD.n16422 DVDD.n16421 0.00239333
R12917 DVDD.n16421 DVDD.n16420 0.00239333
R12918 DVDD.n16420 DVDD.n16419 0.00239333
R12919 DVDD.n16419 DVDD.n16418 0.00239333
R12920 DVDD.n16418 DVDD.n16417 0.00239333
R12921 DVDD.n16417 DVDD.n16416 0.00239333
R12922 DVDD.n16414 DVDD.n16413 0.00239333
R12923 DVDD.n16413 DVDD.n16412 0.00239333
R12924 DVDD.n16412 DVDD.n16411 0.00239333
R12925 DVDD.n16411 DVDD.n16410 0.00239333
R12926 DVDD.n16410 DVDD.n16409 0.00239333
R12927 DVDD.n16409 DVDD.n16408 0.00239333
R12928 DVDD.n16408 DVDD.n16407 0.00239333
R12929 DVDD.n16407 DVDD.n16406 0.00239333
R12930 DVDD.n16406 DVDD.n16405 0.00239333
R12931 DVDD.n16405 DVDD.n16404 0.00239333
R12932 DVDD.n16404 DVDD.n16403 0.00239333
R12933 DVDD.n16403 DVDD.n16402 0.00239333
R12934 DVDD.n16402 DVDD.n16401 0.00239333
R12935 DVDD.n16401 DVDD.n16400 0.00239333
R12936 DVDD.n16400 DVDD.n16399 0.00239333
R12937 DVDD.n16399 DVDD.n16398 0.00239333
R12938 DVDD.n16398 DVDD.n16397 0.00239333
R12939 DVDD.n16397 DVDD.n16396 0.00239333
R12940 DVDD.n16396 DVDD.n16395 0.00239333
R12941 DVDD.n16395 DVDD.n16394 0.00239333
R12942 DVDD.n16394 DVDD.n16393 0.00239333
R12943 DVDD.n16393 DVDD.n16392 0.00239333
R12944 DVDD.n16392 DVDD.n16391 0.00239333
R12945 DVDD.n11126 DVDD.n10988 0.00239333
R12946 DVDD.n11127 DVDD.n11126 0.00239333
R12947 DVDD.n11128 DVDD.n11127 0.00239333
R12948 DVDD.n11129 DVDD.n11128 0.00239333
R12949 DVDD.n11130 DVDD.n11129 0.00239333
R12950 DVDD.n11131 DVDD.n11130 0.00239333
R12951 DVDD.n11132 DVDD.n11131 0.00239333
R12952 DVDD.n11133 DVDD.n11132 0.00239333
R12953 DVDD.n11134 DVDD.n11133 0.00239333
R12954 DVDD.n11135 DVDD.n11134 0.00239333
R12955 DVDD.n11143 DVDD.n11135 0.00239333
R12956 DVDD.n11143 DVDD.n11142 0.00239333
R12957 DVDD.n16820 DVDD.n16819 0.00239333
R12958 DVDD.n16819 DVDD.n16818 0.00239333
R12959 DVDD.n16818 DVDD.n16817 0.00239333
R12960 DVDD.n10807 DVDD.n10806 0.00239333
R12961 DVDD.n10808 DVDD.n10807 0.00239333
R12962 DVDD.n10809 DVDD.n10808 0.00239333
R12963 DVDD.n10810 DVDD.n10809 0.00239333
R12964 DVDD.n10811 DVDD.n10810 0.00239333
R12965 DVDD.n10812 DVDD.n10811 0.00239333
R12966 DVDD.n10836 DVDD.n10835 0.00239333
R12967 DVDD.n10835 DVDD.n10834 0.00239333
R12968 DVDD.n10834 DVDD.n10833 0.00239333
R12969 DVDD.n10833 DVDD.n10832 0.00239333
R12970 DVDD.n10832 DVDD.n10831 0.00239333
R12971 DVDD.n10831 DVDD.n10830 0.00239333
R12972 DVDD.n10830 DVDD.n10829 0.00239333
R12973 DVDD.n10829 DVDD.n10828 0.00239333
R12974 DVDD.n10828 DVDD.n10827 0.00239333
R12975 DVDD.n10827 DVDD.n10826 0.00239333
R12976 DVDD.n10826 DVDD.n10825 0.00239333
R12977 DVDD.n10825 DVDD.n10824 0.00239333
R12978 DVDD.n10824 DVDD.n10823 0.00239333
R12979 DVDD.n10823 DVDD.n10822 0.00239333
R12980 DVDD.n10822 DVDD.n10821 0.00239333
R12981 DVDD.n10821 DVDD.n10820 0.00239333
R12982 DVDD.n10820 DVDD.n10819 0.00239333
R12983 DVDD.n10819 DVDD.n10818 0.00239333
R12984 DVDD.n10818 DVDD.n10817 0.00239333
R12985 DVDD.n10817 DVDD.n10816 0.00239333
R12986 DVDD.n10816 DVDD.n10815 0.00239333
R12987 DVDD.n10815 DVDD.n10814 0.00239333
R12988 DVDD.n10814 DVDD.n10813 0.00239333
R12989 DVDD.n10911 DVDD.n10910 0.00239333
R12990 DVDD.n10910 DVDD.n10909 0.00239333
R12991 DVDD.n10909 DVDD.n10908 0.00239333
R12992 DVDD.n10908 DVDD.n10907 0.00239333
R12993 DVDD.n10907 DVDD.n10906 0.00239333
R12994 DVDD.n10906 DVDD.n10905 0.00239333
R12995 DVDD.n10905 DVDD.n10904 0.00239333
R12996 DVDD.n10904 DVDD.n10903 0.00239333
R12997 DVDD.n10903 DVDD.n10902 0.00239333
R12998 DVDD.n10902 DVDD.n10901 0.00239333
R12999 DVDD.n10901 DVDD.n10900 0.00239333
R13000 DVDD.n10900 DVDD.n10899 0.00239333
R13001 DVDD.n10899 DVDD.n10898 0.00239333
R13002 DVDD.n10898 DVDD.n10897 0.00239333
R13003 DVDD.n10897 DVDD.n10896 0.00239333
R13004 DVDD.n10896 DVDD.n10895 0.00239333
R13005 DVDD.n10895 DVDD.n10894 0.00239333
R13006 DVDD.n10894 DVDD.n10893 0.00239333
R13007 DVDD.n10893 DVDD.n10892 0.00239333
R13008 DVDD.n10892 DVDD.n10891 0.00239333
R13009 DVDD.n10891 DVDD.n10890 0.00239333
R13010 DVDD.n10890 DVDD.n10889 0.00239333
R13011 DVDD.n10889 DVDD.n10888 0.00239333
R13012 DVDD.n10936 DVDD.n10935 0.00239333
R13013 DVDD.n10935 DVDD.n10934 0.00239333
R13014 DVDD.n10934 DVDD.n10933 0.00239333
R13015 DVDD.n10933 DVDD.n10932 0.00239333
R13016 DVDD.n10932 DVDD.n10931 0.00239333
R13017 DVDD.n10931 DVDD.n10930 0.00239333
R13018 DVDD.n10930 DVDD.n10929 0.00239333
R13019 DVDD.n10929 DVDD.n10928 0.00239333
R13020 DVDD.n10928 DVDD.n10927 0.00239333
R13021 DVDD.n10927 DVDD.n10926 0.00239333
R13022 DVDD.n10926 DVDD.n10925 0.00239333
R13023 DVDD.n10925 DVDD.n10924 0.00239333
R13024 DVDD.n10924 DVDD.n10923 0.00239333
R13025 DVDD.n10923 DVDD.n10922 0.00239333
R13026 DVDD.n10922 DVDD.n10921 0.00239333
R13027 DVDD.n10921 DVDD.n10920 0.00239333
R13028 DVDD.n10920 DVDD.n10919 0.00239333
R13029 DVDD.n10919 DVDD.n10918 0.00239333
R13030 DVDD.n10918 DVDD.n10917 0.00239333
R13031 DVDD.n10917 DVDD.n10916 0.00239333
R13032 DVDD.n10916 DVDD.n10915 0.00239333
R13033 DVDD.n10915 DVDD.n10914 0.00239333
R13034 DVDD.n10914 DVDD.n10913 0.00239333
R13035 DVDD.n16388 DVDD.n16387 0.00239333
R13036 DVDD.n16387 DVDD.n16386 0.00239333
R13037 DVDD.n16386 DVDD.n16385 0.00239333
R13038 DVDD.n16385 DVDD.n16384 0.00239333
R13039 DVDD.n16384 DVDD.n16383 0.00239333
R13040 DVDD.n16383 DVDD.n16382 0.00239333
R13041 DVDD.n16381 DVDD.n10990 0.00239333
R13042 DVDD.n16344 DVDD.n10990 0.00239333
R13043 DVDD.n16345 DVDD.n16344 0.00239333
R13044 DVDD.n10771 DVDD.n10770 0.00239333
R13045 DVDD.n10772 DVDD.n10771 0.00239333
R13046 DVDD.n10773 DVDD.n10772 0.00239333
R13047 DVDD.n10774 DVDD.n10773 0.00239333
R13048 DVDD.n10775 DVDD.n10774 0.00239333
R13049 DVDD.n10776 DVDD.n10775 0.00239333
R13050 DVDD.n10777 DVDD.n10776 0.00239333
R13051 DVDD.n10778 DVDD.n10777 0.00239333
R13052 DVDD.n10779 DVDD.n10778 0.00239333
R13053 DVDD.n10780 DVDD.n10779 0.00239333
R13054 DVDD.n10804 DVDD.n10803 0.00239333
R13055 DVDD.n10803 DVDD.n10802 0.00239333
R13056 DVDD.n10802 DVDD.n10801 0.00239333
R13057 DVDD.n10801 DVDD.n10800 0.00239333
R13058 DVDD.n10800 DVDD.n10799 0.00239333
R13059 DVDD.n10799 DVDD.n10798 0.00239333
R13060 DVDD.n10798 DVDD.n10797 0.00239333
R13061 DVDD.n10797 DVDD.n10796 0.00239333
R13062 DVDD.n10796 DVDD.n10795 0.00239333
R13063 DVDD.n10795 DVDD.n10794 0.00239333
R13064 DVDD.n10794 DVDD.n10793 0.00239333
R13065 DVDD.n10793 DVDD.n10792 0.00239333
R13066 DVDD.n10792 DVDD.n10791 0.00239333
R13067 DVDD.n10791 DVDD.n10790 0.00239333
R13068 DVDD.n10790 DVDD.n10789 0.00239333
R13069 DVDD.n10789 DVDD.n10788 0.00239333
R13070 DVDD.n10788 DVDD.n10787 0.00239333
R13071 DVDD.n10787 DVDD.n10786 0.00239333
R13072 DVDD.n10786 DVDD.n10785 0.00239333
R13073 DVDD.n10785 DVDD.n10784 0.00239333
R13074 DVDD.n10784 DVDD.n10783 0.00239333
R13075 DVDD.n10783 DVDD.n10782 0.00239333
R13076 DVDD.n10782 DVDD.n10781 0.00239333
R13077 DVDD.n10886 DVDD.n10885 0.00239333
R13078 DVDD.n10885 DVDD.n10884 0.00239333
R13079 DVDD.n10884 DVDD.n10883 0.00239333
R13080 DVDD.n10883 DVDD.n10882 0.00239333
R13081 DVDD.n10882 DVDD.n10881 0.00239333
R13082 DVDD.n10881 DVDD.n10880 0.00239333
R13083 DVDD.n10880 DVDD.n10879 0.00239333
R13084 DVDD.n10879 DVDD.n10878 0.00239333
R13085 DVDD.n10878 DVDD.n10877 0.00239333
R13086 DVDD.n10877 DVDD.n10876 0.00239333
R13087 DVDD.n10876 DVDD.n10875 0.00239333
R13088 DVDD.n10875 DVDD.n10874 0.00239333
R13089 DVDD.n10874 DVDD.n10873 0.00239333
R13090 DVDD.n10873 DVDD.n10872 0.00239333
R13091 DVDD.n10872 DVDD.n10871 0.00239333
R13092 DVDD.n10871 DVDD.n10870 0.00239333
R13093 DVDD.n10870 DVDD.n10869 0.00239333
R13094 DVDD.n10869 DVDD.n10868 0.00239333
R13095 DVDD.n10868 DVDD.n10867 0.00239333
R13096 DVDD.n10867 DVDD.n10866 0.00239333
R13097 DVDD.n10866 DVDD.n10865 0.00239333
R13098 DVDD.n10865 DVDD.n10864 0.00239333
R13099 DVDD.n10864 DVDD.n10863 0.00239333
R13100 DVDD.n10985 DVDD.n10984 0.00239333
R13101 DVDD.n10984 DVDD.n10983 0.00239333
R13102 DVDD.n10983 DVDD.n10982 0.00239333
R13103 DVDD.n10982 DVDD.n10981 0.00239333
R13104 DVDD.n10981 DVDD.n10980 0.00239333
R13105 DVDD.n10980 DVDD.n10979 0.00239333
R13106 DVDD.n10979 DVDD.n10978 0.00239333
R13107 DVDD.n10978 DVDD.n10977 0.00239333
R13108 DVDD.n10977 DVDD.n10976 0.00239333
R13109 DVDD.n10976 DVDD.n10975 0.00239333
R13110 DVDD.n10975 DVDD.n10974 0.00239333
R13111 DVDD.n10974 DVDD.n10973 0.00239333
R13112 DVDD.n10973 DVDD.n10972 0.00239333
R13113 DVDD.n10972 DVDD.n10971 0.00239333
R13114 DVDD.n10971 DVDD.n10970 0.00239333
R13115 DVDD.n10970 DVDD.n10969 0.00239333
R13116 DVDD.n10969 DVDD.n10968 0.00239333
R13117 DVDD.n10968 DVDD.n10967 0.00239333
R13118 DVDD.n10967 DVDD.n10966 0.00239333
R13119 DVDD.n10966 DVDD.n10965 0.00239333
R13120 DVDD.n10965 DVDD.n10964 0.00239333
R13121 DVDD.n10964 DVDD.n10963 0.00239333
R13122 DVDD.n10963 DVDD.n10962 0.00239333
R13123 DVDD.n15616 DVDD.n15615 0.00239333
R13124 DVDD.n15617 DVDD.n15616 0.00239333
R13125 DVDD.n15618 DVDD.n15617 0.00239333
R13126 DVDD.n15619 DVDD.n15618 0.00239333
R13127 DVDD.n15620 DVDD.n15619 0.00239333
R13128 DVDD.n15621 DVDD.n15620 0.00239333
R13129 DVDD.n15622 DVDD.n15621 0.00239333
R13130 DVDD.n15623 DVDD.n15622 0.00239333
R13131 DVDD.n15706 DVDD.n15705 0.00239333
R13132 DVDD.n10735 DVDD.n10734 0.00239333
R13133 DVDD.n10736 DVDD.n10735 0.00239333
R13134 DVDD.n10737 DVDD.n10736 0.00239333
R13135 DVDD.n10738 DVDD.n10737 0.00239333
R13136 DVDD.n10739 DVDD.n10738 0.00239333
R13137 DVDD.n10740 DVDD.n10739 0.00239333
R13138 DVDD.n10741 DVDD.n10740 0.00239333
R13139 DVDD.n10742 DVDD.n10741 0.00239333
R13140 DVDD.n10743 DVDD.n10742 0.00239333
R13141 DVDD.n10744 DVDD.n10743 0.00239333
R13142 DVDD.n10768 DVDD.n10767 0.00239333
R13143 DVDD.n10767 DVDD.n10766 0.00239333
R13144 DVDD.n10766 DVDD.n10765 0.00239333
R13145 DVDD.n10765 DVDD.n10764 0.00239333
R13146 DVDD.n10764 DVDD.n10763 0.00239333
R13147 DVDD.n10763 DVDD.n10762 0.00239333
R13148 DVDD.n10762 DVDD.n10761 0.00239333
R13149 DVDD.n10761 DVDD.n10760 0.00239333
R13150 DVDD.n10760 DVDD.n10759 0.00239333
R13151 DVDD.n10759 DVDD.n10758 0.00239333
R13152 DVDD.n10758 DVDD.n10757 0.00239333
R13153 DVDD.n10757 DVDD.n10756 0.00239333
R13154 DVDD.n10756 DVDD.n10755 0.00239333
R13155 DVDD.n10755 DVDD.n10754 0.00239333
R13156 DVDD.n10754 DVDD.n10753 0.00239333
R13157 DVDD.n10753 DVDD.n10752 0.00239333
R13158 DVDD.n10752 DVDD.n10751 0.00239333
R13159 DVDD.n10751 DVDD.n10750 0.00239333
R13160 DVDD.n10750 DVDD.n10749 0.00239333
R13161 DVDD.n10749 DVDD.n10748 0.00239333
R13162 DVDD.n10748 DVDD.n10747 0.00239333
R13163 DVDD.n10747 DVDD.n10746 0.00239333
R13164 DVDD.n10746 DVDD.n10745 0.00239333
R13165 DVDD.n10861 DVDD.n10860 0.00239333
R13166 DVDD.n10860 DVDD.n10859 0.00239333
R13167 DVDD.n10859 DVDD.n10858 0.00239333
R13168 DVDD.n10858 DVDD.n10857 0.00239333
R13169 DVDD.n10857 DVDD.n10856 0.00239333
R13170 DVDD.n10856 DVDD.n10855 0.00239333
R13171 DVDD.n10855 DVDD.n10854 0.00239333
R13172 DVDD.n10854 DVDD.n10853 0.00239333
R13173 DVDD.n10853 DVDD.n10852 0.00239333
R13174 DVDD.n10852 DVDD.n10851 0.00239333
R13175 DVDD.n10851 DVDD.n10850 0.00239333
R13176 DVDD.n10850 DVDD.n10849 0.00239333
R13177 DVDD.n10849 DVDD.n10848 0.00239333
R13178 DVDD.n10848 DVDD.n10847 0.00239333
R13179 DVDD.n10847 DVDD.n10846 0.00239333
R13180 DVDD.n10846 DVDD.n10845 0.00239333
R13181 DVDD.n10845 DVDD.n10844 0.00239333
R13182 DVDD.n10844 DVDD.n10843 0.00239333
R13183 DVDD.n10843 DVDD.n10842 0.00239333
R13184 DVDD.n10842 DVDD.n10841 0.00239333
R13185 DVDD.n10841 DVDD.n10840 0.00239333
R13186 DVDD.n10840 DVDD.n10839 0.00239333
R13187 DVDD.n10839 DVDD.n10838 0.00239333
R13188 DVDD.n10960 DVDD.n10959 0.00239333
R13189 DVDD.n10959 DVDD.n10958 0.00239333
R13190 DVDD.n10958 DVDD.n10957 0.00239333
R13191 DVDD.n10957 DVDD.n10956 0.00239333
R13192 DVDD.n10956 DVDD.n10955 0.00239333
R13193 DVDD.n10955 DVDD.n10954 0.00239333
R13194 DVDD.n10954 DVDD.n10953 0.00239333
R13195 DVDD.n10953 DVDD.n10952 0.00239333
R13196 DVDD.n10952 DVDD.n10951 0.00239333
R13197 DVDD.n10951 DVDD.n10950 0.00239333
R13198 DVDD.n10950 DVDD.n10949 0.00239333
R13199 DVDD.n10949 DVDD.n10948 0.00239333
R13200 DVDD.n10948 DVDD.n10947 0.00239333
R13201 DVDD.n10947 DVDD.n10946 0.00239333
R13202 DVDD.n10946 DVDD.n10945 0.00239333
R13203 DVDD.n10945 DVDD.n10944 0.00239333
R13204 DVDD.n10944 DVDD.n10943 0.00239333
R13205 DVDD.n10943 DVDD.n10942 0.00239333
R13206 DVDD.n10942 DVDD.n10941 0.00239333
R13207 DVDD.n10941 DVDD.n10940 0.00239333
R13208 DVDD.n10940 DVDD.n10939 0.00239333
R13209 DVDD.n10939 DVDD.n10938 0.00239333
R13210 DVDD.n10938 DVDD.n10937 0.00239333
R13211 DVDD.n15896 DVDD.n15895 0.00239333
R13212 DVDD.n15897 DVDD.n15896 0.00239333
R13213 DVDD.n15898 DVDD.n15897 0.00239333
R13214 DVDD.n15899 DVDD.n15898 0.00239333
R13215 DVDD.n15900 DVDD.n15899 0.00239333
R13216 DVDD.n15901 DVDD.n15900 0.00239333
R13217 DVDD.n15902 DVDD.n15901 0.00239333
R13218 DVDD.n15903 DVDD.n15902 0.00239333
R13219 DVDD.n15916 DVDD.n15915 0.00239333
R13220 DVDD.n16 DVDD.n12 0.00239333
R13221 DVDD.n20 DVDD.n16 0.00239333
R13222 DVDD.n24 DVDD.n20 0.00239333
R13223 DVDD.n7356 DVDD.n108 0.00239333
R13224 DVDD.n7360 DVDD.n7356 0.00239333
R13225 DVDD.n7364 DVDD.n7360 0.00239333
R13226 DVDD.n7368 DVDD.n7364 0.00239333
R13227 DVDD.n7376 DVDD.n7372 0.00239333
R13228 DVDD.n7380 DVDD.n7376 0.00239333
R13229 DVDD.n7384 DVDD.n7380 0.00239333
R13230 DVDD.n7386 DVDD.n7384 0.00239333
R13231 DVDD.n7426 DVDD.n7422 0.00239333
R13232 DVDD.n7422 DVDD.n7418 0.00239333
R13233 DVDD.n7418 DVDD.n7414 0.00239333
R13234 DVDD.n7414 DVDD.n7410 0.00239333
R13235 DVDD.n7406 DVDD.n7402 0.00239333
R13236 DVDD.n7402 DVDD.n7398 0.00239333
R13237 DVDD.n7398 DVDD.n7394 0.00239333
R13238 DVDD.n7394 DVDD.n7390 0.00239333
R13239 DVDD.n7597 DVDD.n7595 0.00239333
R13240 DVDD.n7595 DVDD.n7591 0.00239333
R13241 DVDD.n7591 DVDD.n7587 0.00239333
R13242 DVDD.n98 DVDD.n94 0.00239333
R13243 DVDD.n102 DVDD.n98 0.00239333
R13244 DVDD.n106 DVDD.n102 0.00239333
R13245 DVDD.n88 DVDD.n86 0.00239333
R13246 DVDD.n86 DVDD.n82 0.00239333
R13247 DVDD.n82 DVDD.n78 0.00239333
R13248 DVDD.n78 DVDD.n74 0.00239333
R13249 DVDD.n70 DVDD.n66 0.00239333
R13250 DVDD.n66 DVDD.n62 0.00239333
R13251 DVDD.n62 DVDD.n58 0.00239333
R13252 DVDD.n58 DVDD.n54 0.00239333
R13253 DVDD.n7474 DVDD.n7470 0.00239333
R13254 DVDD.n7470 DVDD.n7466 0.00239333
R13255 DVDD.n7466 DVDD.n7462 0.00239333
R13256 DVDD.n7462 DVDD.n7458 0.00239333
R13257 DVDD.n7454 DVDD.n7450 0.00239333
R13258 DVDD.n7450 DVDD.n7446 0.00239333
R13259 DVDD.n7446 DVDD.n7442 0.00239333
R13260 DVDD.n7442 DVDD.n7438 0.00239333
R13261 DVDD.n7553 DVDD.n7551 0.00239333
R13262 DVDD.n7551 DVDD.n7547 0.00239333
R13263 DVDD.n7547 DVDD.n7543 0.00239333
R13264 DVDD.n44 DVDD.n40 0.00239333
R13265 DVDD.n48 DVDD.n44 0.00239333
R13266 DVDD.n52 DVDD.n48 0.00239333
R13267 DVDD.n7229 DVDD.n34 0.00239333
R13268 DVDD.n7233 DVDD.n7229 0.00239333
R13269 DVDD.n7237 DVDD.n7233 0.00239333
R13270 DVDD.n7241 DVDD.n7237 0.00239333
R13271 DVDD.n7249 DVDD.n7245 0.00239333
R13272 DVDD.n7253 DVDD.n7249 0.00239333
R13273 DVDD.n7257 DVDD.n7253 0.00239333
R13274 DVDD.n7258 DVDD.n7257 0.00239333
R13275 DVDD.n7483 DVDD.n7479 0.00239333
R13276 DVDD.n7487 DVDD.n7483 0.00239333
R13277 DVDD.n7491 DVDD.n7487 0.00239333
R13278 DVDD.n7495 DVDD.n7491 0.00239333
R13279 DVDD.n7503 DVDD.n7499 0.00239333
R13280 DVDD.n7507 DVDD.n7503 0.00239333
R13281 DVDD.n7511 DVDD.n7507 0.00239333
R13282 DVDD.n7512 DVDD.n7511 0.00239333
R13283 DVDD.n7199 DVDD.n7197 0.00239333
R13284 DVDD.n7197 DVDD.n7193 0.00239333
R13285 DVDD.n7193 DVDD.n7189 0.00239333
R13286 DVDD.n10328 DVDD.n10327 0.00239333
R13287 DVDD.n10327 DVDD.n10326 0.00239333
R13288 DVDD.n10326 DVDD.n10325 0.00239333
R13289 DVDD.n10325 DVDD.n10324 0.00239333
R13290 DVDD.n10324 DVDD.n10323 0.00239333
R13291 DVDD.n10323 DVDD.n10322 0.00239333
R13292 DVDD.n10322 DVDD.n10321 0.00239333
R13293 DVDD.n10321 DVDD.n10320 0.00239333
R13294 DVDD.n10320 DVDD.n10319 0.00239333
R13295 DVDD.n10319 DVDD.n10318 0.00239333
R13296 DVDD.n10316 DVDD.n10315 0.00239333
R13297 DVDD.n10315 DVDD.n10314 0.00239333
R13298 DVDD.n10314 DVDD.n10313 0.00239333
R13299 DVDD.n10313 DVDD.n10312 0.00239333
R13300 DVDD.n10312 DVDD.n10311 0.00239333
R13301 DVDD.n10311 DVDD.n10310 0.00239333
R13302 DVDD.n10310 DVDD.n10309 0.00239333
R13303 DVDD.n10309 DVDD.n10308 0.00239333
R13304 DVDD.n10308 DVDD.n10307 0.00239333
R13305 DVDD.n10307 DVDD.n10306 0.00239333
R13306 DVDD.n10306 DVDD.n10305 0.00239333
R13307 DVDD.n10305 DVDD.n10304 0.00239333
R13308 DVDD.n10304 DVDD.n10303 0.00239333
R13309 DVDD.n10303 DVDD.n10302 0.00239333
R13310 DVDD.n10302 DVDD.n10301 0.00239333
R13311 DVDD.n10301 DVDD.n10300 0.00239333
R13312 DVDD.n10300 DVDD.n10299 0.00239333
R13313 DVDD.n10299 DVDD.n10298 0.00239333
R13314 DVDD.n10298 DVDD.n10297 0.00239333
R13315 DVDD.n10297 DVDD.n10296 0.00239333
R13316 DVDD.n10296 DVDD.n10295 0.00239333
R13317 DVDD.n10295 DVDD.n10294 0.00239333
R13318 DVDD.n10294 DVDD.n10293 0.00239333
R13319 DVDD.n10269 DVDD.n10268 0.00239333
R13320 DVDD.n10268 DVDD.n10267 0.00239333
R13321 DVDD.n10267 DVDD.n10266 0.00239333
R13322 DVDD.n10266 DVDD.n10265 0.00239333
R13323 DVDD.n10265 DVDD.n10264 0.00239333
R13324 DVDD.n10264 DVDD.n10263 0.00239333
R13325 DVDD.n10263 DVDD.n10262 0.00239333
R13326 DVDD.n10262 DVDD.n10261 0.00239333
R13327 DVDD.n10261 DVDD.n10260 0.00239333
R13328 DVDD.n10260 DVDD.n10259 0.00239333
R13329 DVDD.n10259 DVDD.n10258 0.00239333
R13330 DVDD.n10258 DVDD.n10257 0.00239333
R13331 DVDD.n10257 DVDD.n10256 0.00239333
R13332 DVDD.n10256 DVDD.n10255 0.00239333
R13333 DVDD.n10255 DVDD.n10254 0.00239333
R13334 DVDD.n10254 DVDD.n10253 0.00239333
R13335 DVDD.n10253 DVDD.n10252 0.00239333
R13336 DVDD.n10252 DVDD.n10251 0.00239333
R13337 DVDD.n10251 DVDD.n10250 0.00239333
R13338 DVDD.n10250 DVDD.n10249 0.00239333
R13339 DVDD.n10249 DVDD.n10248 0.00239333
R13340 DVDD.n10248 DVDD.n10247 0.00239333
R13341 DVDD.n10247 DVDD.n10246 0.00239333
R13342 DVDD.n10230 DVDD.n10229 0.00239333
R13343 DVDD.n15160 DVDD.n15159 0.00239333
R13344 DVDD.n15161 DVDD.n15160 0.00239333
R13345 DVDD.n15162 DVDD.n15161 0.00239333
R13346 DVDD.n15163 DVDD.n15162 0.00239333
R13347 DVDD.n15164 DVDD.n15163 0.00239333
R13348 DVDD.n15165 DVDD.n15164 0.00239333
R13349 DVDD.n15166 DVDD.n15165 0.00239333
R13350 DVDD.n15167 DVDD.n15166 0.00239333
R13351 DVDD.n15168 DVDD.n15167 0.00239333
R13352 DVDD.n15169 DVDD.n15168 0.00239333
R13353 DVDD.n15170 DVDD.n15169 0.00239333
R13354 DVDD.n15171 DVDD.n15170 0.00239333
R13355 DVDD.n15172 DVDD.n15171 0.00239333
R13356 DVDD.n15173 DVDD.n15172 0.00239333
R13357 DVDD.n15174 DVDD.n15173 0.00239333
R13358 DVDD.n15175 DVDD.n15174 0.00239333
R13359 DVDD.n15176 DVDD.n15175 0.00239333
R13360 DVDD.n15177 DVDD.n15176 0.00239333
R13361 DVDD.n15178 DVDD.n15177 0.00239333
R13362 DVDD.n15179 DVDD.n15178 0.00239333
R13363 DVDD.n15180 DVDD.n15179 0.00239333
R13364 DVDD.n15326 DVDD.n14829 0.00239333
R13365 DVDD.n15327 DVDD.n15326 0.00239333
R13366 DVDD.n15328 DVDD.n15327 0.00239333
R13367 DVDD.n15329 DVDD.n15328 0.00239333
R13368 DVDD.n15330 DVDD.n15329 0.00239333
R13369 DVDD.n15331 DVDD.n15330 0.00239333
R13370 DVDD.n15332 DVDD.n15331 0.00239333
R13371 DVDD.n15333 DVDD.n15332 0.00239333
R13372 DVDD.n15334 DVDD.n15333 0.00239333
R13373 DVDD.n15335 DVDD.n15334 0.00239333
R13374 DVDD.n20234 DVDD.n20230 0.00239333
R13375 DVDD.n20238 DVDD.n20234 0.00239333
R13376 DVDD.n20242 DVDD.n20238 0.00239333
R13377 DVDD.n20340 DVDD.n20276 0.00239333
R13378 DVDD.n20276 DVDD.n20272 0.00239333
R13379 DVDD.n20272 DVDD.n20268 0.00239333
R13380 DVDD.n20268 DVDD.n20264 0.00239333
R13381 DVDD.n20260 DVDD.n20256 0.00239333
R13382 DVDD.n20256 DVDD.n20252 0.00239333
R13383 DVDD.n20252 DVDD.n20248 0.00239333
R13384 DVDD.n20248 DVDD.n20244 0.00239333
R13385 DVDD.n7342 DVDD.n7338 0.00239333
R13386 DVDD.n7338 DVDD.n7334 0.00239333
R13387 DVDD.n7334 DVDD.n7330 0.00239333
R13388 DVDD.n7330 DVDD.n7326 0.00239333
R13389 DVDD.n7322 DVDD.n7318 0.00239333
R13390 DVDD.n7318 DVDD.n7314 0.00239333
R13391 DVDD.n7314 DVDD.n7310 0.00239333
R13392 DVDD.n7310 DVDD.n7306 0.00239333
R13393 DVDD.n7680 DVDD.n7676 0.00239333
R13394 DVDD.n7684 DVDD.n7680 0.00239333
R13395 DVDD.n7688 DVDD.n7684 0.00239333
R13396 DVDD.n7704 DVDD.n7703 0.00239
R13397 DVDD.n7711 DVDD.n7710 0.00239
R13398 DVDD.n7771 DVDD.n7770 0.00239
R13399 DVDD.n3703 DVDD.n3702 0.00239
R13400 DVDD.n3696 DVDD.n3695 0.00239
R13401 DVDD.n18542 DVDD.n18541 0.00239
R13402 DVDD.n18549 DVDD.n18548 0.00239
R13403 DVDD.n3449 DVDD.n3448 0.00239
R13404 DVDD.n2958 DVDD.n2957 0.00239
R13405 DVDD.n3578 DVDD.n3577 0.00239
R13406 DVDD.n9955 DVDD.n9954 0.00239
R13407 DVDD.n9818 DVDD.n9817 0.00239
R13408 DVDD.n9516 DVDD.n9515 0.00239
R13409 DVDD.n2196 DVDD.n2195 0.00239
R13410 DVDD.n2259 DVDD.n2258 0.00239
R13411 DVDD.n2252 DVDD.n2251 0.00239
R13412 DVDD.n18911 DVDD.n18910 0.00239
R13413 DVDD.n18918 DVDD.n18917 0.00239
R13414 DVDD.n7065 DVDD.n7064 0.00239
R13415 DVDD.n7058 DVDD.n7057 0.00239
R13416 DVDD.n1898 DVDD.n1897 0.00239
R13417 DVDD.n1891 DVDD.n1890 0.00239
R13418 DVDD.n19975 DVDD.n19974 0.00239
R13419 DVDD.n20038 DVDD.n20037 0.00239
R13420 DVDD.n20031 DVDD.n20030 0.00239
R13421 DVDD.n19029 DVDD.n19028 0.00239
R13422 DVDD.n19036 DVDD.n19035 0.00239
R13423 DVDD.n4645 DVDD.n4644 0.00239
R13424 DVDD.n4638 DVDD.n4637 0.00239
R13425 DVDD.n19676 DVDD.n19675 0.00239
R13426 DVDD.n19669 DVDD.n19668 0.00239
R13427 DVDD.n1548 DVDD.n1547 0.00239
R13428 DVDD.n970 DVDD.n969 0.00239
R13429 DVDD.n1672 DVDD.n1671 0.00239
R13430 DVDD.n946 DVDD.n945 0.00239
R13431 DVDD.n939 DVDD.n938 0.00239
R13432 DVDD.n19238 DVDD.n19237 0.00239
R13433 DVDD.n19245 DVDD.n19244 0.00239
R13434 DVDD.n11539 DVDD.n11538 0.00239
R13435 DVDD.n18321 DVDD.n18320 0.00239
R13436 DVDD.n18314 DVDD.n18313 0.00239
R13437 DVDD.n10127 DVDD.n10126 0.00239
R13438 DVDD.n11919 DVDD.n11918 0.00239
R13439 DVDD.n1321 DVDD.n1320 0.00239
R13440 DVDD.n1314 DVDD.n1313 0.00239
R13441 DVDD.n1281 DVDD.n1280 0.00239
R13442 DVDD.n12321 DVDD.n12320 0.00239
R13443 DVDD.n3323 DVDD.n3322 0.00239
R13444 DVDD.n3282 DVDD.n3281 0.00239
R13445 DVDD.n3289 DVDD.n3288 0.00239
R13446 DVDD.n16061 DVDD.n16060 0.00238285
R13447 DVDD.n15673 DVDD.n15672 0.00238285
R13448 DVDD.n8184 DVDD.n8183 0.00238285
R13449 DVDD.n9400 DVDD.n9399 0.00238285
R13450 DVDD.n19504 DVDD.n19503 0.00236
R13451 DVDD.n20119 DVDD.n20118 0.00236
R13452 DVDD.n10349 DVDD.n10348 0.00236
R13453 DVDD.n16504 DVDD.n16503 0.00236
R13454 DVDD.n16846 DVDD.n16845 0.00236
R13455 DVDD.n19560 DVDD.n19559 0.00233
R13456 DVDD.n20175 DVDD.n20174 0.00233
R13457 DVDD.n234 DVDD.n233 0.00233
R13458 DVDD.n164 DVDD.n163 0.00233
R13459 DVDD.n19365 DVDD.n19364 0.00233
R13460 DVDD.n15354 DVDD.n15353 0.00233
R13461 DVDD.n11161 DVDD.n11160 0.00233
R13462 DVDD.n16365 DVDD.n16364 0.00233
R13463 DVDD.n18588 DVDD.n18587 0.00233
R13464 DVDD.n18685 DVDD.n18684 0.00233
R13465 DVDD.n18361 DVDD.n18360 0.00233
R13466 DVDD.n4983 DVDD.n4982 0.00232835
R13467 DVDD.n13427 DVDD.n13426 0.00232835
R13468 DVDD.n13428 DVDD.n13427 0.00232835
R13469 DVDD.n5579 DVDD.n5578 0.00232835
R13470 DVDD.n5578 DVDD.n5577 0.00232835
R13471 DVDD.n5328 DVDD.n5327 0.00232835
R13472 DVDD.n5443 DVDD.n5442 0.00232835
R13473 DVDD.n5418 DVDD.n5417 0.00232835
R13474 DVDD.n5353 DVDD.n5352 0.00232835
R13475 DVDD.n12848 DVDD.n12847 0.00232835
R13476 DVDD.n13131 DVDD.n13130 0.00232835
R13477 DVDD.n13020 DVDD.n13019 0.00232835
R13478 DVDD.n12849 DVDD.n12848 0.00232835
R13479 DVDD.n6228 DVDD.n6227 0.00232835
R13480 DVDD.n6433 DVDD.n6432 0.00232835
R13481 DVDD.n6318 DVDD.n6317 0.00232835
R13482 DVDD.n6229 DVDD.n6228 0.00232835
R13483 DVDD.n8930 DVDD.n8929 0.00232835
R13484 DVDD.n8931 DVDD.n8930 0.00232835
R13485 DVDD.n9219 DVDD.n9218 0.00232835
R13486 DVDD.n9104 DVDD.n9103 0.00232835
R13487 DVDD.n15209 DVDD.n15208 0.00232497
R13488 DVDD.n15128 DVDD.n15127 0.00232497
R13489 DVDD.n7970 DVDD.n7969 0.00231761
R13490 DVDD.n7969 DVDD.n7968 0.00231761
R13491 DVDD.n7760 DVDD.n7759 0.0023
R13492 DVDD.n7757 DVDD.n7756 0.0023
R13493 DVDD.n7754 DVDD.n7753 0.0023
R13494 DVDD.n7751 DVDD.n7750 0.0023
R13495 DVDD.n7748 DVDD.n7747 0.0023
R13496 DVDD.n7745 DVDD.n7694 0.0023
R13497 DVDD.n7830 DVDD.n7829 0.0023
R13498 DVDD.n9765 DVDD.n9764 0.0023
R13499 DVDD.n7934 DVDD.n7933 0.0023
R13500 DVDD.n7932 DVDD.n7931 0.0023
R13501 DVDD.n9537 DVDD.n9536 0.0023
R13502 DVDD.n9261 DVDD.n9260 0.0023
R13503 DVDD.n9266 DVDD.n9265 0.0023
R13504 DVDD.n9303 DVDD.n9302 0.0023
R13505 DVDD.n9317 DVDD.n9316 0.0023
R13506 DVDD DVDD.n13832 0.0023
R13507 DVDD.n6799 DVDD.n6798 0.0023
R13508 DVDD.n6850 DVDD.n6849 0.0023
R13509 DVDD.n6521 DVDD.n6520 0.0023
R13510 DVDD.n6523 DVDD.n6522 0.0023
R13511 DVDD.n6569 DVDD.n6568 0.0023
R13512 DVDD.n3981 DVDD.n3980 0.0023
R13513 DVDD.n3976 DVDD.n3975 0.0023
R13514 DVDD.n3939 DVDD.n3938 0.0023
R13515 DVDD.n3817 DVDD.n3816 0.0023
R13516 DVDD.n4836 DVDD.n4835 0.0023
R13517 DVDD.n4887 DVDD.n4886 0.0023
R13518 DVDD.n5112 DVDD.n5111 0.0023
R13519 DVDD.n5114 DVDD.n5113 0.0023
R13520 DVDD.n5160 DVDD.n5159 0.0023
R13521 DVDD.n5286 DVDD.n5285 0.0023
R13522 DVDD.n5281 DVDD.n5280 0.0023
R13523 DVDD.n5244 DVDD.n5243 0.0023
R13524 DVDD.n12465 DVDD.n12463 0.0023
R13525 DVDD.n12472 DVDD.n12471 0.0023
R13526 DVDD.n5707 DVDD.n5705 0.0023
R13527 DVDD.n4553 DVDD.n4552 0.0023
R13528 DVDD.n6112 DVDD.n4068 0.0023
R13529 DVDD.n4075 DVDD.n4074 0.0023
R13530 DVDD.n8490 DVDD.n8488 0.0023
R13531 DVDD.n8497 DVDD.n8496 0.0023
R13532 DVDD.n12458 DVDD.n12457 0.0023
R13533 DVDD.n5664 DVDD.n5663 0.0023
R13534 DVDD.n4570 DVDD.n4569 0.0023
R13535 DVDD.n4560 DVDD.n4559 0.0023
R13536 DVDD.n4066 DVDD.n4065 0.0023
R13537 DVDD.n8470 DVDD.n8469 0.0023
R13538 DVDD.n8482 DVDD.n8481 0.0023
R13539 DVDD.n12433 DVDD.n12432 0.0023
R13540 DVDD.n12445 DVDD.n12444 0.0023
R13541 DVDD.n5618 DVDD.n5617 0.0023
R13542 DVDD.n4585 DVDD.n4584 0.0023
R13543 DVDD.n4575 DVDD.n4574 0.0023
R13544 DVDD.n4056 DVDD.n4055 0.0023
R13545 DVDD.n8452 DVDD.n8451 0.0023
R13546 DVDD.n8464 DVDD.n8463 0.0023
R13547 DVDD.n12414 DVDD.n12413 0.0023
R13548 DVDD.n12426 DVDD.n12425 0.0023
R13549 DVDD.n5571 DVDD.n5570 0.0023
R13550 DVDD.n4600 DVDD.n4599 0.0023
R13551 DVDD.n4590 DVDD.n4589 0.0023
R13552 DVDD.n4046 DVDD.n4045 0.0023
R13553 DVDD.n8434 DVDD.n8433 0.0023
R13554 DVDD.n8446 DVDD.n8445 0.0023
R13555 DVDD.n2486 DVDD 0.0023
R13556 DVDD.n18272 DVDD.n18271 0.0023
R13557 DVDD.n18269 DVDD.n18268 0.0023
R13558 DVDD.n10156 DVDD.n10155 0.0023
R13559 DVDD.n10153 DVDD.n10152 0.0023
R13560 DVDD.n10150 DVDD.n10149 0.0023
R13561 DVDD.n10147 DVDD.n10146 0.0023
R13562 DVDD.n10083 DVDD.n10082 0.0023
R13563 DVDD.n7634 DVDD.n7633 0.0023
R13564 DVDD.n7128 DVDD.n7127 0.0023
R13565 DVDD.n7112 DVDD.n7111 0.0023
R13566 DVDD.n7658 DVDD.n7657 0.0023
R13567 DVDD.n1819 DVDD.n1818 0.0023
R13568 DVDD.n2830 DVDD.n2829 0.0023
R13569 DVDD.n2814 DVDD.n2813 0.0023
R13570 DVDD.n20300 DVDD.n20299 0.0023
R13571 DVDD.n20322 DVDD.n20321 0.0023
R13572 DVDD.n11355 DVDD.n11354 0.0023
R13573 DVDD.n11866 DVDD.n11865 0.0023
R13574 DVDD.n1244 DVDD.n1243 0.0023
R13575 DVDD.n1247 DVDD.n1246 0.0023
R13576 DVDD.n1250 DVDD.n1249 0.0023
R13577 DVDD.n1253 DVDD.n1252 0.0023
R13578 DVDD.n1256 DVDD.n1255 0.0023
R13579 DVDD.n1259 DVDD.n1258 0.0023
R13580 DVDD.n1262 DVDD.n1261 0.0023
R13581 DVDD.n1265 DVDD.n1264 0.0023
R13582 DVDD.n1268 DVDD.n1267 0.0023
R13583 DVDD.n1271 DVDD.n1270 0.0023
R13584 DVDD.n2698 DVDD 0.0023
R13585 DVDD DVDD.n2691 0.0023
R13586 DVDD.n11336 DVDD.n11335 0.0023
R13587 DVDD.n11334 DVDD.n11333 0.0023
R13588 DVDD.n12341 DVDD.n12340 0.0023
R13589 DVDD.n14981 DVDD.n14930 0.0023
R13590 DVDD.n14853 DVDD.n14852 0.0023
R13591 DVDD.n15013 DVDD.n15007 0.0023
R13592 DVDD.n13172 DVDD.n13171 0.0023
R13593 DVDD.n13177 DVDD.n13176 0.0023
R13594 DVDD.n13214 DVDD.n13213 0.0023
R13595 DVDD.n13228 DVDD.n13227 0.0023
R13596 DVDD.n3330 DVDD.n3329 0.0023
R13597 DVDD.n3442 DVDD.n3441 0.0023
R13598 DVDD.n3386 DVDD.n3385 0.0023
R13599 DVDD.n3367 DVDD.n3366 0.0023
R13600 DVDD.n3585 DVDD.n3584 0.0023
R13601 DVDD.n3664 DVDD.n3663 0.0023
R13602 DVDD.n3657 DVDD.n3656 0.0023
R13603 DVDD.n3651 DVDD.n3607 0.0023
R13604 DVDD.n3602 DVDD.n3601 0.0023
R13605 DVDD.n3595 DVDD.n3594 0.0023
R13606 DVDD.n3589 DVDD.n3588 0.0023
R13607 DVDD.n18585 DVDD.n18584 0.0023
R13608 DVDD.n18615 DVDD.n18614 0.0023
R13609 DVDD.n18631 DVDD.n18630 0.0023
R13610 DVDD.n18426 DVDD.n18425 0.0023
R13611 DVDD.n3154 DVDD.n3153 0.0023
R13612 DVDD.n3151 DVDD.n3150 0.0023
R13613 DVDD.n3148 DVDD.n3147 0.0023
R13614 DVDD.n3145 DVDD.n3144 0.0023
R13615 DVDD.n3142 DVDD.n3141 0.0023
R13616 DVDD.n3139 DVDD.n3138 0.0023
R13617 DVDD.n3136 DVDD.n3135 0.0023
R13618 DVDD.n3133 DVDD.n3132 0.0023
R13619 DVDD.n3130 DVDD.n3129 0.0023
R13620 DVDD.n3127 DVDD.n3126 0.0023
R13621 DVDD.n13061 DVDD.n13060 0.00229713
R13622 DVDD.n1569 DVDD.n1568 0.00227165
R13623 DVDD.n1622 DVDD.n1621 0.00227165
R13624 DVDD.n1661 DVDD.n1660 0.00227165
R13625 DVDD.n891 DVDD.n890 0.00227165
R13626 DVDD.n19275 DVDD.n19274 0.00227165
R13627 DVDD.n19282 DVDD.n19281 0.00227165
R13628 DVDD.n19294 DVDD.n19293 0.00227165
R13629 DVDD.n19299 DVDD.n19298 0.00227165
R13630 DVDD.n19306 DVDD.n19305 0.00227165
R13631 DVDD.n19415 DVDD.n19339 0.00227165
R13632 DVDD.n19330 DVDD.n19329 0.00227165
R13633 DVDD.n19327 DVDD.n19326 0.00227165
R13634 DVDD.n19326 DVDD.n19325 0.00227165
R13635 DVDD.n19320 DVDD.n19319 0.00227165
R13636 DVDD.n10169 DVDD.n10168 0.00227165
R13637 DVDD.n11430 DVDD.n11429 0.00227165
R13638 DVDD.n12205 DVDD.n12204 0.00227165
R13639 DVDD.n13490 DVDD.n13489 0.00227165
R13640 DVDD.n13550 DVDD.n13549 0.00227165
R13641 DVDD.n13631 DVDD.n13630 0.00227165
R13642 DVDD.n2743 DVDD.n2742 0.00227165
R13643 DVDD.n2784 DVDD.n2783 0.00227165
R13644 DVDD.n18575 DVDD.n18574 0.00227165
R13645 DVDD.n14805 DVDD.n14804 0.00227165
R13646 DVDD.n15395 DVDD.n15394 0.00227165
R13647 DVDD.n14708 DVDD.n14707 0.00227165
R13648 DVDD.n14625 DVDD.n14624 0.00227165
R13649 DVDD.n14571 DVDD.n14570 0.00227165
R13650 DVDD.n14483 DVDD.n14482 0.00227165
R13651 DVDD.n19700 DVDD.n19699 0.00227165
R13652 DVDD.n19742 DVDD.n19741 0.00227165
R13653 DVDD.n19745 DVDD.n19744 0.00227165
R13654 DVDD.n19908 DVDD.n19907 0.00227165
R13655 DVDD.n20003 DVDD.n20002 0.00227165
R13656 DVDD.n20092 DVDD.n20091 0.00227165
R13657 DVDD.n20095 DVDD.n20094 0.00227165
R13658 DVDD.n19070 DVDD.n19069 0.00227165
R13659 DVDD.n19062 DVDD.n19061 0.00227165
R13660 DVDD.n4807 DVDD.n4806 0.00227165
R13661 DVDD.n4911 DVDD.n4910 0.00227165
R13662 DVDD.n4987 DVDD.n4986 0.00227165
R13663 DVDD.n5098 DVDD.n5097 0.00227165
R13664 DVDD.n5197 DVDD.n5196 0.00227165
R13665 DVDD.n5217 DVDD.n5216 0.00227165
R13666 DVDD.n5330 DVDD.n5329 0.00227165
R13667 DVDD.n5391 DVDD.n5390 0.00227165
R13668 DVDD.n5421 DVDD.n5420 0.00227165
R13669 DVDD.n5582 DVDD.n5581 0.00227165
R13670 DVDD.n5583 DVDD.n5582 0.00227165
R13671 DVDD.n5631 DVDD.n5630 0.00227165
R13672 DVDD.n6101 DVDD.n6100 0.00227165
R13673 DVDD.n6097 DVDD.n6096 0.00227165
R13674 DVDD.n6079 DVDD.n6078 0.00227165
R13675 DVDD.n1345 DVDD.n1344 0.00227165
R13676 DVDD.n1387 DVDD.n1386 0.00227165
R13677 DVDD.n1469 DVDD.n1468 0.00227165
R13678 DVDD.n1691 DVDD.n1690 0.00227165
R13679 DVDD.n19190 DVDD.n19189 0.00227165
R13680 DVDD.n19193 DVDD.n19192 0.00227165
R13681 DVDD.n19452 DVDD.n19451 0.00227165
R13682 DVDD.n19444 DVDD.n19443 0.00227165
R13683 DVDD.n11633 DVDD.n11632 0.00227165
R13684 DVDD.n11842 DVDD.n11841 0.00227165
R13685 DVDD.n11766 DVDD.n11765 0.00227165
R13686 DVDD.n11656 DVDD.n11655 0.00227165
R13687 DVDD.n12377 DVDD.n12376 0.00227165
R13688 DVDD.n12397 DVDD.n12396 0.00227165
R13689 DVDD.n13129 DVDD.n13128 0.00227165
R13690 DVDD.n13070 DVDD.n13069 0.00227165
R13691 DVDD.n13041 DVDD.n13040 0.00227165
R13692 DVDD.n12845 DVDD.n12844 0.00227165
R13693 DVDD.n12844 DVDD.n12843 0.00227165
R13694 DVDD.n12806 DVDD.n12805 0.00227165
R13695 DVDD.n12733 DVDD.n12732 0.00227165
R13696 DVDD.n12729 DVDD.n12728 0.00227165
R13697 DVDD.n12711 DVDD.n12710 0.00227165
R13698 DVDD.n781 DVDD.n780 0.00227165
R13699 DVDD.n818 DVDD.n817 0.00227165
R13700 DVDD.n244 DVDD.n243 0.00227165
R13701 DVDD.n18233 DVDD.n18232 0.00227165
R13702 DVDD.n18205 DVDD.n18204 0.00227165
R13703 DVDD.n18061 DVDD.n18060 0.00227165
R13704 DVDD.n17983 DVDD.n17982 0.00227165
R13705 DVDD.n17931 DVDD.n17930 0.00227165
R13706 DVDD.n17850 DVDD.n17849 0.00227165
R13707 DVDD.n1922 DVDD.n1921 0.00227165
R13708 DVDD.n1964 DVDD.n1963 0.00227165
R13709 DVDD.n2129 DVDD.n2128 0.00227165
R13710 DVDD.n2224 DVDD.n2223 0.00227165
R13711 DVDD.n19477 DVDD.n19476 0.00227165
R13712 DVDD.n19480 DVDD.n19479 0.00227165
R13713 DVDD.n18962 DVDD.n18961 0.00227165
R13714 DVDD.n18954 DVDD.n18953 0.00227165
R13715 DVDD.n6877 DVDD.n6876 0.00227165
R13716 DVDD.n6773 DVDD.n6772 0.00227165
R13717 DVDD.n6697 DVDD.n6696 0.00227165
R13718 DVDD.n6584 DVDD.n6583 0.00227165
R13719 DVDD.n6485 DVDD.n6484 0.00227165
R13720 DVDD.n6465 DVDD.n6464 0.00227165
R13721 DVDD.n6431 DVDD.n6430 0.00227165
R13722 DVDD.n6370 DVDD.n6369 0.00227165
R13723 DVDD.n6340 DVDD.n6339 0.00227165
R13724 DVDD.n6225 DVDD.n6224 0.00227165
R13725 DVDD.n6224 DVDD.n6223 0.00227165
R13726 DVDD.n4550 DVDD.n4549 0.00227165
R13727 DVDD.n4547 DVDD.n4546 0.00227165
R13728 DVDD.n4529 DVDD.n4528 0.00227165
R13729 DVDD.n3258 DVDD.n3257 0.00227165
R13730 DVDD.n3216 DVDD.n3215 0.00227165
R13731 DVDD.n3528 DVDD.n3527 0.00227165
R13732 DVDD.n3558 DVDD.n3557 0.00227165
R13733 DVDD.n18494 DVDD.n18493 0.00227165
R13734 DVDD.n18497 DVDD.n18496 0.00227165
R13735 DVDD.n18799 DVDD.n18798 0.00227165
R13736 DVDD.n18791 DVDD.n18790 0.00227165
R13737 DVDD.n7889 DVDD.n7888 0.00227165
R13738 DVDD.n9741 DVDD.n9740 0.00227165
R13739 DVDD.n9665 DVDD.n9664 0.00227165
R13740 DVDD.n9552 DVDD.n9551 0.00227165
R13741 DVDD.n8398 DVDD.n8397 0.00227165
R13742 DVDD.n8418 DVDD.n8417 0.00227165
R13743 DVDD.n9217 DVDD.n9216 0.00227165
R13744 DVDD.n9156 DVDD.n9155 0.00227165
R13745 DVDD.n9126 DVDD.n9125 0.00227165
R13746 DVDD.n8927 DVDD.n8926 0.00227165
R13747 DVDD.n8926 DVDD.n8925 0.00227165
R13748 DVDD.n8817 DVDD.n8816 0.00227165
R13749 DVDD.n8814 DVDD.n8813 0.00227165
R13750 DVDD.n8796 DVDD.n8795 0.00227165
R13751 DVDD.n19341 DVDD.n19340 0.00227
R13752 DVDD.n18467 DVDD.n18463 0.00227
R13753 DVDD.n8068 DVDD.n8067 0.00225306
R13754 DVDD.n12025 DVDD.n12024 0.00223982
R13755 DVDD.n12024 DVDD.n12023 0.00223982
R13756 DVDD.n6070 DVDD.n6069 0.00223982
R13757 DVDD.n19711 DVDD.n19710 0.00223982
R13758 DVDD.n6071 DVDD.n6070 0.00223982
R13759 DVDD.n12702 DVDD.n12701 0.00223982
R13760 DVDD.n12703 DVDD.n12702 0.00223982
R13761 DVDD.n4520 DVDD.n4519 0.00223982
R13762 DVDD.n4521 DVDD.n4520 0.00223982
R13763 DVDD.n8787 DVDD.n8786 0.00223982
R13764 DVDD.n8788 DVDD.n8787 0.00223982
R13765 DVDD.n4163 DVDD.n4162 0.00223571
R13766 DVDD.n8545 DVDD.n8544 0.00223571
R13767 DVDD.n13877 DVDD.n13876 0.00223571
R13768 DVDD.n13841 DVDD.n13840 0.00223571
R13769 DVDD.n2449 DVDD.n2448 0.00223571
R13770 DVDD.n2335 DVDD.n2334 0.00223571
R13771 DVDD.n2375 DVDD.n2374 0.00223571
R13772 DVDD.n2386 DVDD.n2385 0.00223571
R13773 DVDD.n2422 DVDD.n2421 0.00223571
R13774 DVDD.n2451 DVDD.n2450 0.00223571
R13775 DVDD.n2471 DVDD.n2470 0.00223571
R13776 DVDD.n2645 DVDD.n2627 0.00223571
R13777 DVDD.n2681 DVDD.n2680 0.00223571
R13778 DVDD.n2533 DVDD.n2532 0.00223571
R13779 DVDD.n2573 DVDD.n2572 0.00223571
R13780 DVDD.n2584 DVDD.n2583 0.00223571
R13781 DVDD.n2618 DVDD.n2617 0.00223571
R13782 DVDD.n2647 DVDD.n2646 0.00223571
R13783 DVDD.n2683 DVDD.n2682 0.00223571
R13784 DVDD.n4130 DVDD.n4129 0.00223571
R13785 DVDD.n4164 DVDD.n4160 0.00223571
R13786 DVDD.n8512 DVDD.n8511 0.00223571
R13787 DVDD.n8546 DVDD.n8542 0.00223571
R13788 DVDD.n11214 DVDD.n11213 0.00223571
R13789 DVDD.n13878 DVDD.n13874 0.00223571
R13790 DVDD.n13851 DVDD.n13850 0.00223571
R13791 DVDD.n13842 DVDD.n13839 0.00223571
R13792 DVDD.n15205 DVDD.n15204 0.00222892
R13793 DVDD.n15126 DVDD.n15125 0.00222892
R13794 DVDD.n15966 DVDD.n15965 0.00222352
R13795 DVDD.n15967 DVDD.n15966 0.00222352
R13796 DVDD.n8284 DVDD.n8283 0.00222352
R13797 DVDD.n9450 DVDD.n9449 0.00222352
R13798 DVDD.n9451 DVDD.n9450 0.00222352
R13799 DVDD.n8131 DVDD.n8130 0.00222352
R13800 DVDD.n8130 DVDD.n8129 0.00222352
R13801 DVDD.n8034 DVDD.n8033 0.00222352
R13802 DVDD.n8033 DVDD.n8032 0.00222352
R13803 DVDD.n3682 DVDD.n3681 0.00221
R13804 DVDD.n3713 DVDD.n3712 0.00221
R13805 DVDD.n18559 DVDD.n18558 0.00221
R13806 DVDD.n2943 DVDD.n2942 0.00221
R13807 DVDD.n7818 DVDD.n7817 0.00221
R13808 DVDD.n7820 DVDD.n7819 0.00221
R13809 DVDD.n9811 DVDD.n9810 0.00221
R13810 DVDD.n9882 DVDD.n9881 0.00221
R13811 DVDD.n9879 DVDD.n9878 0.00221
R13812 DVDD.n9876 DVDD.n9875 0.00221
R13813 DVDD.n9873 DVDD.n9872 0.00221
R13814 DVDD.n9870 DVDD.n9869 0.00221
R13815 DVDD.n9867 DVDD.n9866 0.00221
R13816 DVDD.n9864 DVDD.n9863 0.00221
R13817 DVDD.n9861 DVDD.n9860 0.00221
R13818 DVDD.n9858 DVDD.n9857 0.00221
R13819 DVDD.n9855 DVDD.n9854 0.00221
R13820 DVDD.n9852 DVDD.n9851 0.00221
R13821 DVDD.n9849 DVDD.n9848 0.00221
R13822 DVDD.n9846 DVDD.n9845 0.00221
R13823 DVDD.n9843 DVDD.n9842 0.00221
R13824 DVDD.n9840 DVDD.n9839 0.00221
R13825 DVDD.n9837 DVDD.n9836 0.00221
R13826 DVDD.n9834 DVDD.n9833 0.00221
R13827 DVDD.n9831 DVDD.n9830 0.00221
R13828 DVDD.n9828 DVDD.n9827 0.00221
R13829 DVDD.n9825 DVDD.n9824 0.00221
R13830 DVDD.n9389 DVDD.n9388 0.00221
R13831 DVDD.n2181 DVDD.n2180 0.00221
R13832 DVDD.n2238 DVDD.n2237 0.00221
R13833 DVDD.n2269 DVDD.n2268 0.00221
R13834 DVDD.n18928 DVDD.n18927 0.00221
R13835 DVDD.n6787 DVDD.n6786 0.00221
R13836 DVDD.n6789 DVDD.n6788 0.00221
R13837 DVDD.n6804 DVDD.n6803 0.00221
R13838 DVDD.n1881 DVDD.n1880 0.00221
R13839 DVDD.n1878 DVDD.n1877 0.00221
R13840 DVDD.n19960 DVDD.n19959 0.00221
R13841 DVDD.n20017 DVDD.n20016 0.00221
R13842 DVDD.n20048 DVDD.n20047 0.00221
R13843 DVDD.n19046 DVDD.n19045 0.00221
R13844 DVDD.n4824 DVDD.n4823 0.00221
R13845 DVDD.n4826 DVDD.n4825 0.00221
R13846 DVDD.n4841 DVDD.n4840 0.00221
R13847 DVDD.n19659 DVDD.n19658 0.00221
R13848 DVDD.n19656 DVDD.n19655 0.00221
R13849 DVDD.n985 DVDD.n984 0.00221
R13850 DVDD.n1725 DVDD.n1724 0.00221
R13851 DVDD.n956 DVDD.n955 0.00221
R13852 DVDD.n19255 DVDD.n19254 0.00221
R13853 DVDD.n11343 DVDD.n11342 0.00221
R13854 DVDD.n11345 DVDD.n11344 0.00221
R13855 DVDD.n11912 DVDD.n11911 0.00221
R13856 DVDD.n11983 DVDD.n11982 0.00221
R13857 DVDD.n11980 DVDD.n11979 0.00221
R13858 DVDD.n11977 DVDD.n11976 0.00221
R13859 DVDD.n11974 DVDD.n11973 0.00221
R13860 DVDD.n11971 DVDD.n11970 0.00221
R13861 DVDD.n11968 DVDD.n11967 0.00221
R13862 DVDD.n11965 DVDD.n11964 0.00221
R13863 DVDD.n11962 DVDD.n11961 0.00221
R13864 DVDD.n11959 DVDD.n11958 0.00221
R13865 DVDD.n11956 DVDD.n11955 0.00221
R13866 DVDD.n11953 DVDD.n11952 0.00221
R13867 DVDD.n11950 DVDD.n11949 0.00221
R13868 DVDD.n11947 DVDD.n11946 0.00221
R13869 DVDD.n11944 DVDD.n11943 0.00221
R13870 DVDD.n11941 DVDD.n11940 0.00221
R13871 DVDD.n11938 DVDD.n11937 0.00221
R13872 DVDD.n11935 DVDD.n11934 0.00221
R13873 DVDD.n11932 DVDD.n11931 0.00221
R13874 DVDD.n11929 DVDD.n11928 0.00221
R13875 DVDD.n11926 DVDD.n11925 0.00221
R13876 DVDD.n1304 DVDD.n1303 0.00221
R13877 DVDD.n1301 DVDD.n1300 0.00221
R13878 DVDD.n10501 DVDD.n10499 0.00221
R13879 DVDD.n13300 DVDD.n13299 0.00221
R13880 DVDD.n17112 DVDD.n17110 0.00221
R13881 DVDD.n16719 DVDD.n16718 0.00221
R13882 DVDD.n16550 DVDD.n16549 0.00221
R13883 DVDD.n3299 DVDD.n3298 0.00221
R13884 DVDD.n3302 DVDD.n3301 0.00221
R13885 DVDD.n3063 DVDD.n3062 0.00220503
R13886 DVDD.n3064 DVDD.n3063 0.00220503
R13887 DVDD.n8097 DVDD.n8096 0.0022027
R13888 DVDD.n16031 DVDD.n16030 0.00219456
R13889 DVDD.n16020 DVDD.n16019 0.00219456
R13890 DVDD.n15643 DVDD.n15642 0.00219456
R13891 DVDD.n15632 DVDD.n15631 0.00219456
R13892 DVDD.n8146 DVDD.n8145 0.00219456
R13893 DVDD.n8342 DVDD.n8341 0.00219456
R13894 DVDD.n9475 DVDD.n9474 0.00219456
R13895 DVDD.n8037 DVDD.n8036 0.00219456
R13896 DVDD.n1849 DVDD.n1848 0.00218
R13897 DVDD.n19627 DVDD.n19626 0.00218
R13898 DVDD.n1796 DVDD.n1795 0.00218
R13899 DVDD.n17012 DVDD.n17011 0.00218
R13900 DVDD.n16954 DVDD.n16953 0.00218
R13901 DVDD.n16787 DVDD.n16786 0.00218
R13902 DVDD.n16910 DVDD.n16909 0.00218
R13903 DVDD.n16665 DVDD.n16664 0.00218
R13904 DVDD.n16608 DVDD.n16607 0.00218
R13905 DVDD.n3638 DVDD.n3637 0.00218
R13906 DVDD.n14095 DVDD.n14094 0.00217553
R13907 DVDD.n14006 DVDD.n14005 0.00217553
R13908 DVDD.n14216 DVDD.n14215 0.00217553
R13909 DVDD.n4133 DVDD.n4131 0.00217143
R13910 DVDD.n8515 DVDD.n8513 0.00217143
R13911 DVDD.n11217 DVDD.n11215 0.00217143
R13912 DVDD.n2326 DVDD.n2325 0.00217143
R13913 DVDD.n2377 DVDD.n2376 0.00217143
R13914 DVDD.n2424 DVDD.n2423 0.00217143
R13915 DVDD.n2327 DVDD.n2324 0.00217143
R13916 DVDD.n2336 DVDD.n2335 0.00217143
R13917 DVDD.n2378 DVDD.n2375 0.00217143
R13918 DVDD.n2387 DVDD.n2386 0.00217143
R13919 DVDD.n2425 DVDD.n2422 0.00217143
R13920 DVDD.n2501 DVDD.n2451 0.00217143
R13921 DVDD.n2524 DVDD.n2523 0.00217143
R13922 DVDD.n2575 DVDD.n2574 0.00217143
R13923 DVDD.n2620 DVDD.n2619 0.00217143
R13924 DVDD.n2525 DVDD.n2522 0.00217143
R13925 DVDD.n2534 DVDD.n2533 0.00217143
R13926 DVDD.n2576 DVDD.n2573 0.00217143
R13927 DVDD.n2585 DVDD.n2584 0.00217143
R13928 DVDD.n2621 DVDD.n2618 0.00217143
R13929 DVDD.n2713 DVDD.n2647 0.00217143
R13930 DVDD.n2673 DVDD.n2670 0.00217143
R13931 DVDD.n4134 DVDD.n4130 0.00217143
R13932 DVDD.n4160 DVDD.n4159 0.00217143
R13933 DVDD.n8516 DVDD.n8512 0.00217143
R13934 DVDD.n8542 DVDD.n8541 0.00217143
R13935 DVDD.n11218 DVDD.n11214 0.00217143
R13936 DVDD.n13874 DVDD.n13873 0.00217143
R13937 DVDD.n13850 DVDD.n13849 0.00217143
R13938 DVDD.n13839 DVDD.n13838 0.00217143
R13939 DVDD.n18988 DVDD.n18987 0.0021686
R13940 DVDD.n10555 DVDD.n10554 0.0021686
R13941 DVDD.n8004 DVDD.n8003 0.00215892
R13942 DVDD.n12091 DVDD.n12090 0.00215128
R13943 DVDD.n12190 DVDD.n12189 0.00215128
R13944 DVDD.n12255 DVDD.n12254 0.00215128
R13945 DVDD.n13386 DVDD.n13385 0.00215128
R13946 DVDD.n13720 DVDD.n13719 0.00215128
R13947 DVDD.n12189 DVDD.n12188 0.00215128
R13948 DVDD.n12090 DVDD.n12089 0.00215128
R13949 DVDD.n12256 DVDD.n12255 0.00215128
R13950 DVDD.n13385 DVDD.n13384 0.00215128
R13951 DVDD.n15490 DVDD.n15489 0.00215128
R13952 DVDD.n15510 DVDD.n15509 0.00215128
R13953 DVDD.n14667 DVDD.n14666 0.00215128
R13954 DVDD.n14372 DVDD.n14371 0.00215128
R13955 DVDD.n14320 DVDD.n14319 0.00215128
R13956 DVDD.n14668 DVDD.n14667 0.00215128
R13957 DVDD.n15489 DVDD.n15488 0.00215128
R13958 DVDD.n15509 DVDD.n15508 0.00215128
R13959 DVDD.n5050 DVDD.n5049 0.00215128
R13960 DVDD.n5372 DVDD.n5371 0.00215128
R13961 DVDD.n5934 DVDD.n5933 0.00215128
R13962 DVDD.n5880 DVDD.n5879 0.00215128
R13963 DVDD.n5878 DVDD.n5877 0.00215128
R13964 DVDD.n5872 DVDD.n5871 0.00215128
R13965 DVDD.n5870 DVDD.n5869 0.00215128
R13966 DVDD.n5816 DVDD.n5815 0.00215128
R13967 DVDD.n5815 DVDD.n5814 0.00215128
R13968 DVDD.n5807 DVDD.n5806 0.00215128
R13969 DVDD.n5806 DVDD.n5805 0.00215128
R13970 DVDD.n5371 DVDD.n5370 0.00215128
R13971 DVDD.n5049 DVDD.n5048 0.00215128
R13972 DVDD.n4934 DVDD.n4933 0.00215128
R13973 DVDD.n11704 DVDD.n11703 0.00215128
R13974 DVDD.n13088 DVDD.n13087 0.00215128
R13975 DVDD.n12597 DVDD.n12596 0.00215128
R13976 DVDD.n12576 DVDD.n12575 0.00215128
R13977 DVDD.n12575 DVDD.n12574 0.00215128
R13978 DVDD.n12570 DVDD.n12569 0.00215128
R13979 DVDD.n12568 DVDD.n12567 0.00215128
R13980 DVDD.n12514 DVDD.n12513 0.00215128
R13981 DVDD.n12513 DVDD.n12512 0.00215128
R13982 DVDD.n12508 DVDD.n12507 0.00215128
R13983 DVDD.n12507 DVDD.n12506 0.00215128
R13984 DVDD.n13089 DVDD.n13088 0.00215128
R13985 DVDD.n11705 DVDD.n11704 0.00215128
R13986 DVDD.n5808 DVDD.n5807 0.00215128
R13987 DVDD.n12509 DVDD.n12508 0.00215128
R13988 DVDD.n12506 DVDD.n12505 0.00215128
R13989 DVDD.n12515 DVDD.n12514 0.00215128
R13990 DVDD.n5817 DVDD.n5816 0.00215128
R13991 DVDD.n5814 DVDD.n5810 0.00215128
R13992 DVDD.n12512 DVDD.n12511 0.00215128
R13993 DVDD.n5805 DVDD.n5804 0.00215128
R13994 DVDD.n18119 DVDD.n18118 0.00215128
R13995 DVDD.n18101 DVDD.n18100 0.00215128
R13996 DVDD.n18023 DVDD.n18022 0.00215128
R13997 DVDD.n17750 DVDD.n17749 0.00215128
R13998 DVDD.n17688 DVDD.n17687 0.00215128
R13999 DVDD.n18024 DVDD.n18023 0.00215128
R14000 DVDD.n18120 DVDD.n18119 0.00215128
R14001 DVDD.n18102 DVDD.n18101 0.00215128
R14002 DVDD.n5879 DVDD.n5878 0.00215128
R14003 DVDD.n5871 DVDD.n5870 0.00215128
R14004 DVDD.n12569 DVDD.n12568 0.00215128
R14005 DVDD.n12577 DVDD.n12576 0.00215128
R14006 DVDD.n5881 DVDD.n5880 0.00215128
R14007 DVDD.n5873 DVDD.n5872 0.00215128
R14008 DVDD.n12571 DVDD.n12570 0.00215128
R14009 DVDD.n12574 DVDD.n12573 0.00215128
R14010 DVDD.n6634 DVDD.n6633 0.00215128
R14011 DVDD.n6389 DVDD.n6388 0.00215128
R14012 DVDD.n4393 DVDD.n4392 0.00215128
R14013 DVDD.n4347 DVDD.n4346 0.00215128
R14014 DVDD.n4334 DVDD.n4333 0.00215128
R14015 DVDD.n4330 DVDD.n4329 0.00215128
R14016 DVDD.n4329 DVDD.n4328 0.00215128
R14017 DVDD.n4246 DVDD.n4245 0.00215128
R14018 DVDD.n4245 DVDD.n4244 0.00215128
R14019 DVDD.n4236 DVDD.n4235 0.00215128
R14020 DVDD.n4235 DVDD.n4234 0.00215128
R14021 DVDD.n4328 DVDD.n4327 0.00215128
R14022 DVDD.n4237 DVDD.n4236 0.00215128
R14023 DVDD.n4346 DVDD.n4335 0.00215128
R14024 DVDD.n4335 DVDD.n4334 0.00215128
R14025 DVDD.n4247 DVDD.n4246 0.00215128
R14026 DVDD.n6390 DVDD.n6389 0.00215128
R14027 DVDD.n6635 DVDD.n6634 0.00215128
R14028 DVDD.n6582 DVDD.n6581 0.00215128
R14029 DVDD.n6414 DVDD.n6413 0.00215128
R14030 DVDD.n4331 DVDD.n4330 0.00215128
R14031 DVDD.n4244 DVDD.n4239 0.00215128
R14032 DVDD.n4234 DVDD.n4233 0.00215128
R14033 DVDD.n4394 DVDD.n4393 0.00215128
R14034 DVDD.n13721 DVDD.n13720 0.00215128
R14035 DVDD.n17751 DVDD.n17750 0.00215128
R14036 DVDD.n5935 DVDD.n5934 0.00215128
R14037 DVDD.n14373 DVDD.n14372 0.00215128
R14038 DVDD.n12598 DVDD.n12597 0.00215128
R14039 DVDD.n9602 DVDD.n9601 0.00215128
R14040 DVDD.n9175 DVDD.n9174 0.00215128
R14041 DVDD.n8667 DVDD.n8666 0.00215128
R14042 DVDD.n8620 DVDD.n8619 0.00215128
R14043 DVDD.n8618 DVDD.n8617 0.00215128
R14044 DVDD.n8614 DVDD.n8613 0.00215128
R14045 DVDD.n8612 DVDD.n8611 0.00215128
R14046 DVDD.n8558 DVDD.n8557 0.00215128
R14047 DVDD.n8556 DVDD.n8555 0.00215128
R14048 DVDD.n8552 DVDD.n8551 0.00215128
R14049 DVDD.n8551 DVDD.n8550 0.00215128
R14050 DVDD.n9603 DVDD.n9602 0.00215128
R14051 DVDD.n8668 DVDD.n8667 0.00215128
R14052 DVDD.n8619 DVDD.n8618 0.00215128
R14053 DVDD.n8613 DVDD.n8612 0.00215128
R14054 DVDD.n8557 DVDD.n8556 0.00215128
R14055 DVDD.n8553 DVDD.n8552 0.00215128
R14056 DVDD.n8559 DVDD.n8558 0.00215128
R14057 DVDD.n9176 DVDD.n9175 0.00215128
R14058 DVDD.n9550 DVDD.n9549 0.00215128
R14059 DVDD.n9200 DVDD.n9199 0.00215128
R14060 DVDD.n8621 DVDD.n8620 0.00215128
R14061 DVDD.n8615 DVDD.n8614 0.00215128
R14062 DVDD.n8550 DVDD.n8549 0.00215128
R14063 DVDD.n18890 DVDD.n18889 0.00215
R14064 DVDD.n19139 DVDD.n19138 0.00215
R14065 DVDD.n19350 DVDD.n19349 0.00215
R14066 DVDD.n16164 DVDD.n16163 0.00215
R14067 DVDD.n16282 DVDD.n16281 0.00215
R14068 DVDD.n16220 DVDD.n16219 0.00215
R14069 DVDD.n15585 DVDD.n15584 0.00215
R14070 DVDD.n15800 DVDD.n15799 0.00215
R14071 DVDD.n15863 DVDD.n15862 0.00215
R14072 DVDD.n18455 DVDD.n18454 0.00215
R14073 DVDD.n15202 DVDD.n15201 0.00213287
R14074 DVDD.n15945 DVDD.n15944 0.00212942
R14075 DVDD.n15944 DVDD.n15943 0.00212942
R14076 DVDD.n15685 DVDD.n15684 0.00212942
R14077 DVDD.n15684 DVDD.n15683 0.00212942
R14078 DVDD.n8221 DVDD.n8220 0.00212942
R14079 DVDD.n9414 DVDD.n9413 0.00212942
R14080 DVDD.n9415 DVDD.n9414 0.00212942
R14081 DVDD.n9897 DVDD.n9896 0.00212942
R14082 DVDD.n9898 DVDD.n9897 0.00212942
R14083 DVDD.n3430 DVDD.n3429 0.00212472
R14084 DVDD.n3423 DVDD.n3422 0.00212472
R14085 DVDD.n3410 DVDD.n3409 0.00212472
R14086 DVDD.n3396 DVDD.n3395 0.00212472
R14087 DVDD.n3390 DVDD.n3389 0.00212472
R14088 DVDD.n3377 DVDD.n3376 0.00212472
R14089 DVDD.n3370 DVDD.n3369 0.00212472
R14090 DVDD.n3363 DVDD.n3362 0.00212472
R14091 DVDD.n3384 DVDD.n3383 0.00212472
R14092 DVDD.n3403 DVDD.n3402 0.00212472
R14093 DVDD.n13138 DVDD.n13137 0.00212003
R14094 DVDD.n9755 DVDD.n9754 0.00212
R14095 DVDD.n9781 DVDD.n9780 0.00212
R14096 DVDD.n9786 DVDD.n9785 0.00212
R14097 DVDD.n7905 DVDD.n7904 0.00212
R14098 DVDD.n9490 DVDD.n9489 0.00212
R14099 DVDD.n9245 DVDD.n9244 0.00212
R14100 DVDD.n9282 DVDD.n9281 0.00212
R14101 DVDD.n9287 DVDD.n9286 0.00212
R14102 DVDD.n6860 DVDD.n6859 0.00212
R14103 DVDD.n6834 DVDD.n6833 0.00212
R14104 DVDD.n6829 DVDD.n6828 0.00212
R14105 DVDD.n6550 DVDD.n6549 0.00212
R14106 DVDD.n3997 DVDD.n3996 0.00212
R14107 DVDD.n3960 DVDD.n3959 0.00212
R14108 DVDD.n3955 DVDD.n3954 0.00212
R14109 DVDD.n4897 DVDD.n4896 0.00212
R14110 DVDD.n4871 DVDD.n4870 0.00212
R14111 DVDD.n4866 DVDD.n4865 0.00212
R14112 DVDD.n5141 DVDD.n5140 0.00212
R14113 DVDD.n5302 DVDD.n5301 0.00212
R14114 DVDD.n5265 DVDD.n5264 0.00212
R14115 DVDD.n5260 DVDD.n5259 0.00212
R14116 DVDD.n11856 DVDD.n11855 0.00212
R14117 DVDD.n11882 DVDD.n11881 0.00212
R14118 DVDD.n11887 DVDD.n11886 0.00212
R14119 DVDD.n11307 DVDD.n11305 0.00212
R14120 DVDD.n12295 DVDD.n12294 0.00212
R14121 DVDD.n13156 DVDD.n13155 0.00212
R14122 DVDD.n13193 DVDD.n13192 0.00212
R14123 DVDD.n13198 DVDD.n13197 0.00212
R14124 DVDD.n409 DVDD.n408 0.00210714
R14125 DVDD.n488 DVDD.n487 0.00210714
R14126 DVDD.n442 DVDD.n441 0.00210714
R14127 DVDD.n640 DVDD.n639 0.00210714
R14128 DVDD.n720 DVDD.n719 0.00210714
R14129 DVDD.n674 DVDD.n673 0.00210714
R14130 DVDD.n13729 DVDD.n11297 0.00210714
R14131 DVDD.n11280 DVDD.n11279 0.00210714
R14132 DVDD.n12504 DVDD.n12503 0.00210714
R14133 DVDD.n5771 DVDD.n5770 0.00210714
R14134 DVDD.n3103 DVDD.n3102 0.00210714
R14135 DVDD.n3039 DVDD.n3038 0.00210714
R14136 DVDD.n1591 DVDD.n1590 0.00209449
R14137 DVDD.n923 DVDD.n922 0.00209449
R14138 DVDD.n19302 DVDD.n19301 0.00209449
R14139 DVDD.n19305 DVDD.n19304 0.00209449
R14140 DVDD.n19337 DVDD.n19336 0.00209449
R14141 DVDD.n19334 DVDD.n19333 0.00209449
R14142 DVDD.n10166 DVDD.n10165 0.00209449
R14143 DVDD.n10173 DVDD.n10172 0.00209449
R14144 DVDD.n10178 DVDD.n10177 0.00209449
R14145 DVDD.n18266 DVDD.n10182 0.00209449
R14146 DVDD.n11429 DVDD.n11428 0.00209449
R14147 DVDD.n11431 DVDD.n11430 0.00209449
R14148 DVDD.n11438 DVDD.n11437 0.00209449
R14149 DVDD.n12094 DVDD.n12093 0.00209449
R14150 DVDD.n12280 DVDD.n12279 0.00209449
R14151 DVDD.n13323 DVDD.n13322 0.00209449
R14152 DVDD.n13526 DVDD.n13525 0.00209449
R14153 DVDD.n13578 DVDD.n13577 0.00209449
R14154 DVDD.n13586 DVDD.n13585 0.00209449
R14155 DVDD.n13659 DVDD.n13658 0.00209449
R14156 DVDD.n13667 DVDD.n13666 0.00209449
R14157 DVDD.n18577 DVDD.n18576 0.00209449
R14158 DVDD.n14803 DVDD.n14802 0.00209449
R14159 DVDD.n15425 DVDD.n15424 0.00209449
R14160 DVDD.n15436 DVDD.n15435 0.00209449
R14161 DVDD.n14678 DVDD.n14677 0.00209449
R14162 DVDD.n14595 DVDD.n14594 0.00209449
R14163 DVDD.n14541 DVDD.n14540 0.00209449
R14164 DVDD.n14530 DVDD.n14529 0.00209449
R14165 DVDD.n14453 DVDD.n14452 0.00209449
R14166 DVDD.n14428 DVDD.n14427 0.00209449
R14167 DVDD.n14319 DVDD.n14318 0.00209449
R14168 DVDD.n19867 DVDD.n19866 0.00209449
R14169 DVDD.n19897 DVDD.n19896 0.00209449
R14170 DVDD.n19904 DVDD.n19903 0.00209449
R14171 DVDD.n20191 DVDD.n20190 0.00209449
R14172 DVDD.n20190 DVDD.n20189 0.00209449
R14173 DVDD.n20187 DVDD.n20186 0.00209449
R14174 DVDD.n20185 DVDD.n20184 0.00209449
R14175 DVDD.n20090 DVDD.n20089 0.00209449
R14176 DVDD.n20096 DVDD.n20095 0.00209449
R14177 DVDD.n19012 DVDD.n19011 0.00209449
R14178 DVDD.n3886 DVDD.n3885 0.00209449
R14179 DVDD.n4653 DVDD.n4652 0.00209449
R14180 DVDD.n4815 DVDD.n4814 0.00209449
R14181 DVDD.n4907 DVDD.n4906 0.00209449
R14182 DVDD.n4942 DVDD.n4941 0.00209449
R14183 DVDD.n4958 DVDD.n4957 0.00209449
R14184 DVDD.n4963 DVDD.n4962 0.00209449
R14185 DVDD.n5027 DVDD.n5026 0.00209449
R14186 DVDD.n5172 DVDD.n5171 0.00209449
R14187 DVDD.n5342 DVDD.n5341 0.00209449
R14188 DVDD.n5352 DVDD.n5351 0.00209449
R14189 DVDD.n5383 DVDD.n5382 0.00209449
R14190 DVDD.n5429 DVDD.n5428 0.00209449
R14191 DVDD.n5492 DVDD.n5491 0.00209449
R14192 DVDD.n5499 DVDD.n5498 0.00209449
R14193 DVDD.n5563 DVDD.n5562 0.00209449
R14194 DVDD.n5639 DVDD.n5638 0.00209449
R14195 DVDD.n5647 DVDD.n5646 0.00209449
R14196 DVDD.n6021 DVDD.n6020 0.00209449
R14197 DVDD.n5986 DVDD.n5985 0.00209449
R14198 DVDD.n1509 DVDD.n1508 0.00209449
R14199 DVDD.n1480 DVDD.n1479 0.00209449
R14200 DVDD.n1473 DVDD.n1472 0.00209449
R14201 DVDD.n269 DVDD.n268 0.00209449
R14202 DVDD.n268 DVDD.n267 0.00209449
R14203 DVDD.n265 DVDD.n264 0.00209449
R14204 DVDD.n263 DVDD.n262 0.00209449
R14205 DVDD.n19188 DVDD.n19187 0.00209449
R14206 DVDD.n19194 DVDD.n19193 0.00209449
R14207 DVDD.n19221 DVDD.n19220 0.00209449
R14208 DVDD.n11356 DVDD.n10123 0.00209449
R14209 DVDD.n11360 DVDD.n11359 0.00209449
R14210 DVDD.n11641 DVDD.n11640 0.00209449
R14211 DVDD.n11846 DVDD.n11845 0.00209449
R14212 DVDD.n11811 DVDD.n11810 0.00209449
R14213 DVDD.n11795 DVDD.n11794 0.00209449
R14214 DVDD.n11790 DVDD.n11789 0.00209449
R14215 DVDD.n11787 DVDD.n11786 0.00209449
R14216 DVDD.n11786 DVDD.n11785 0.00209449
R14217 DVDD.n11727 DVDD.n11726 0.00209449
R14218 DVDD.n12353 DVDD.n12352 0.00209449
R14219 DVDD.n13117 DVDD.n13116 0.00209449
R14220 DVDD.n13108 DVDD.n13107 0.00209449
R14221 DVDD.n13078 DVDD.n13077 0.00209449
R14222 DVDD.n13034 DVDD.n13033 0.00209449
R14223 DVDD.n13003 DVDD.n13002 0.00209449
R14224 DVDD.n12971 DVDD.n12970 0.00209449
R14225 DVDD.n12964 DVDD.n12963 0.00209449
R14226 DVDD.n12854 DVDD.n12853 0.00209449
R14227 DVDD.n12798 DVDD.n12797 0.00209449
R14228 DVDD.n12790 DVDD.n12789 0.00209449
R14229 DVDD.n12672 DVDD.n12671 0.00209449
R14230 DVDD.n12649 DVDD.n12648 0.00209449
R14231 DVDD.n246 DVDD.n245 0.00209449
R14232 DVDD.n18235 DVDD.n18234 0.00209449
R14233 DVDD.n18177 DVDD.n18176 0.00209449
R14234 DVDD.n18169 DVDD.n18168 0.00209449
R14235 DVDD.n18033 DVDD.n18032 0.00209449
R14236 DVDD.n17955 DVDD.n17954 0.00209449
R14237 DVDD.n17903 DVDD.n17902 0.00209449
R14238 DVDD.n17895 DVDD.n17894 0.00209449
R14239 DVDD.n17822 DVDD.n17821 0.00209449
R14240 DVDD.n17802 DVDD.n17801 0.00209449
R14241 DVDD.n17687 DVDD.n17686 0.00209449
R14242 DVDD.n2089 DVDD.n2088 0.00209449
R14243 DVDD.n2118 DVDD.n2117 0.00209449
R14244 DVDD.n2125 DVDD.n2124 0.00209449
R14245 DVDD.n19576 DVDD.n19575 0.00209449
R14246 DVDD.n19575 DVDD.n19574 0.00209449
R14247 DVDD.n19572 DVDD.n19571 0.00209449
R14248 DVDD.n19570 DVDD.n19569 0.00209449
R14249 DVDD.n19475 DVDD.n19474 0.00209449
R14250 DVDD.n19481 DVDD.n19480 0.00209449
R14251 DVDD.n18939 DVDD.n18938 0.00209449
R14252 DVDD.n7107 DVDD.n7106 0.00209449
R14253 DVDD.n7072 DVDD.n7030 0.00209449
R14254 DVDD.n6869 DVDD.n6868 0.00209449
R14255 DVDD.n6777 DVDD.n6776 0.00209449
R14256 DVDD.n6742 DVDD.n6741 0.00209449
R14257 DVDD.n6726 DVDD.n6725 0.00209449
R14258 DVDD.n6721 DVDD.n6720 0.00209449
R14259 DVDD.n6718 DVDD.n6717 0.00209449
R14260 DVDD.n6717 DVDD.n6716 0.00209449
R14261 DVDD.n6657 DVDD.n6656 0.00209449
R14262 DVDD.n6510 DVDD.n6509 0.00209449
R14263 DVDD.n6419 DVDD.n6418 0.00209449
R14264 DVDD.n6409 DVDD.n6408 0.00209449
R14265 DVDD.n6378 DVDD.n6377 0.00209449
R14266 DVDD.n6332 DVDD.n6331 0.00209449
R14267 DVDD.n6301 DVDD.n6300 0.00209449
R14268 DVDD.n6267 DVDD.n6266 0.00209449
R14269 DVDD.n6259 DVDD.n6258 0.00209449
R14270 DVDD.n6178 DVDD.n6177 0.00209449
R14271 DVDD.n6167 DVDD.n6166 0.00209449
R14272 DVDD.n4472 DVDD.n4471 0.00209449
R14273 DVDD.n4449 DVDD.n4448 0.00209449
R14274 DVDD.n3488 DVDD.n3487 0.00209449
R14275 DVDD.n3517 DVDD.n3516 0.00209449
R14276 DVDD.n3524 DVDD.n3523 0.00209449
R14277 DVDD.n3755 DVDD.n3754 0.00209449
R14278 DVDD.n3754 DVDD.n3753 0.00209449
R14279 DVDD.n3751 DVDD.n3750 0.00209449
R14280 DVDD.n3749 DVDD.n3748 0.00209449
R14281 DVDD.n18492 DVDD.n18491 0.00209449
R14282 DVDD.n18498 DVDD.n18497 0.00209449
R14283 DVDD.n18525 DVDD.n18524 0.00209449
R14284 DVDD.n10052 DVDD.n10051 0.00209449
R14285 DVDD.n10048 DVDD.n10047 0.00209449
R14286 DVDD.n7897 DVDD.n7896 0.00209449
R14287 DVDD.n9745 DVDD.n9744 0.00209449
R14288 DVDD.n9710 DVDD.n9709 0.00209449
R14289 DVDD.n9694 DVDD.n9693 0.00209449
R14290 DVDD.n9689 DVDD.n9688 0.00209449
R14291 DVDD.n9686 DVDD.n9685 0.00209449
R14292 DVDD.n9685 DVDD.n9684 0.00209449
R14293 DVDD.n9625 DVDD.n9624 0.00209449
R14294 DVDD.n8373 DVDD.n8372 0.00209449
R14295 DVDD.n9205 DVDD.n9204 0.00209449
R14296 DVDD.n9195 DVDD.n9194 0.00209449
R14297 DVDD.n9164 DVDD.n9163 0.00209449
R14298 DVDD.n9118 DVDD.n9117 0.00209449
R14299 DVDD.n9087 DVDD.n9086 0.00209449
R14300 DVDD.n9053 DVDD.n9052 0.00209449
R14301 DVDD.n9045 DVDD.n9044 0.00209449
R14302 DVDD.n8880 DVDD.n8879 0.00209449
R14303 DVDD.n8869 DVDD.n8868 0.00209449
R14304 DVDD.n8758 DVDD.n8757 0.00209449
R14305 DVDD.n8723 DVDD.n8722 0.00209449
R14306 DVDD.n3804 DVDD.n3803 0.002075
R14307 DVDD.n18822 DVDD.n18821 0.002075
R14308 DVDD.n19154 DVDD.n19153 0.002075
R14309 DVDD.n7265 DVDD.n7264 0.002075
R14310 DVDD.n3847 DVDD.n3846 0.002075
R14311 DVDD.n3901 DVDD.n3900 0.002075
R14312 DVDD.n132 DVDD.n131 0.002075
R14313 DVDD.n3790 DVDD.n3789 0.002075
R14314 DVDD.n14840 DVDD.n14839 0.002075
R14315 DVDD.n14870 DVDD.n14869 0.002075
R14316 DVDD.n15090 DVDD.n15089 0.002075
R14317 DVDD.n10708 DVDD.n10707 0.002075
R14318 DVDD.n10616 DVDD.n10615 0.002075
R14319 DVDD.n7278 DVDD.n7277 0.002075
R14320 DVDD.n16390 DVDD.n10988 0.00207333
R14321 DVDD.n16389 DVDD.n16388 0.00207333
R14322 DVDD.n15615 DVDD.n10989 0.00207333
R14323 DVDD.n15895 DVDD.n15894 0.00207333
R14324 DVDD.n15181 DVDD.n14829 0.00207333
R14325 DVDD.n8275 DVDD.n8274 0.00206481
R14326 DVDD.n3830 DVDD.n3829 0.00206431
R14327 DVDD.n115 DVDD.n114 0.00206431
R14328 DVDD.n5624 DVDD.n5623 0.00206293
R14329 DVDD.n12813 DVDD.n12812 0.00206293
R14330 DVDD.n6192 DVDD.n6191 0.00206293
R14331 DVDD.n8894 DVDD.n8893 0.00206293
R14332 DVDD.n6148 DVDD.n6147 0.00206288
R14333 DVDD.n8850 DVDD.n8849 0.00206288
R14334 DVDD.n1588 DVDD.n1587 0.00206274
R14335 DVDD.n11481 DVDD.n11480 0.00206274
R14336 DVDD.n12219 DVDD.n12218 0.00206274
R14337 DVDD.n13451 DVDD.n13450 0.00206274
R14338 DVDD.n13536 DVDD.n13535 0.00206274
R14339 DVDD.n13617 DVDD.n13616 0.00206274
R14340 DVDD.n1184 DVDD.n1183 0.00206274
R14341 DVDD.n11482 DVDD.n11481 0.00206274
R14342 DVDD.n12220 DVDD.n12219 0.00206274
R14343 DVDD.n13452 DVDD.n13451 0.00206274
R14344 DVDD.n13535 DVDD.n13534 0.00206274
R14345 DVDD.n13616 DVDD.n13615 0.00206274
R14346 DVDD.n2729 DVDD.n2728 0.00206274
R14347 DVDD.n2770 DVDD.n2769 0.00206274
R14348 DVDD.n14819 DVDD.n14818 0.00206274
R14349 DVDD.n14722 DVDD.n14721 0.00206274
R14350 DVDD.n14639 DVDD.n14638 0.00206274
R14351 DVDD.n14585 DVDD.n14584 0.00206274
R14352 DVDD.n14497 DVDD.n14496 0.00206274
R14353 DVDD.n14723 DVDD.n14722 0.00206274
R14354 DVDD.n14818 DVDD.n14817 0.00206274
R14355 DVDD.n2728 DVDD.n2727 0.00206274
R14356 DVDD.n2769 DVDD.n2768 0.00206274
R14357 DVDD.n14640 DVDD.n14639 0.00206274
R14358 DVDD.n14498 DVDD.n14497 0.00206274
R14359 DVDD.n14586 DVDD.n14585 0.00206274
R14360 DVDD.n19710 DVDD.n19709 0.00206274
R14361 DVDD.n19877 DVDD.n19876 0.00206274
R14362 DVDD.n4783 DVDD.n4782 0.00206274
R14363 DVDD.n5203 DVDD.n5202 0.00206274
R14364 DVDD.n5426 DVDD.n5425 0.00206274
R14365 DVDD.n5550 DVDD.n5549 0.00206274
R14366 DVDD.n5425 DVDD.n5424 0.00206274
R14367 DVDD.n5202 DVDD.n5201 0.00206274
R14368 DVDD.n4782 DVDD.n4781 0.00206274
R14369 DVDD.n19709 DVDD.n19708 0.00206274
R14370 DVDD.n19876 DVDD.n19875 0.00206274
R14371 DVDD.n5549 DVDD.n5548 0.00206274
R14372 DVDD.n1355 DVDD.n1354 0.00206274
R14373 DVDD.n1499 DVDD.n1498 0.00206274
R14374 DVDD.n11609 DVDD.n11608 0.00206274
R14375 DVDD.n12383 DVDD.n12382 0.00206274
R14376 DVDD.n13037 DVDD.n13036 0.00206274
R14377 DVDD.n12868 DVDD.n12867 0.00206274
R14378 DVDD.n12382 DVDD.n12381 0.00206274
R14379 DVDD.n12364 DVDD.n12363 0.00206274
R14380 DVDD.n11608 DVDD.n11607 0.00206274
R14381 DVDD.n1354 DVDD.n1353 0.00206274
R14382 DVDD.n1500 DVDD.n1499 0.00206274
R14383 DVDD.n12867 DVDD.n12866 0.00206274
R14384 DVDD.n767 DVDD.n766 0.00206274
R14385 DVDD.n804 DVDD.n803 0.00206274
R14386 DVDD.n18219 DVDD.n18218 0.00206274
R14387 DVDD.n18075 DVDD.n18074 0.00206274
R14388 DVDD.n17997 DVDD.n17996 0.00206274
R14389 DVDD.n17945 DVDD.n17944 0.00206274
R14390 DVDD.n17864 DVDD.n17863 0.00206274
R14391 DVDD.n17998 DVDD.n17997 0.00206274
R14392 DVDD.n18076 DVDD.n18075 0.00206274
R14393 DVDD.n18220 DVDD.n18219 0.00206274
R14394 DVDD.n766 DVDD.n765 0.00206274
R14395 DVDD.n803 DVDD.n802 0.00206274
R14396 DVDD.n17865 DVDD.n17864 0.00206274
R14397 DVDD.n17946 DVDD.n17945 0.00206274
R14398 DVDD.n1932 DVDD.n1931 0.00206274
R14399 DVDD.n2099 DVDD.n2098 0.00206274
R14400 DVDD.n6901 DVDD.n6900 0.00206274
R14401 DVDD.n6498 DVDD.n6497 0.00206274
R14402 DVDD.n6479 DVDD.n6478 0.00206274
R14403 DVDD.n6335 DVDD.n6334 0.00206274
R14404 DVDD.n6246 DVDD.n6245 0.00206274
R14405 DVDD.n6480 DVDD.n6479 0.00206274
R14406 DVDD.n6902 DVDD.n6901 0.00206274
R14407 DVDD.n1931 DVDD.n1930 0.00206274
R14408 DVDD.n2098 DVDD.n2097 0.00206274
R14409 DVDD.n6336 DVDD.n6335 0.00206274
R14410 DVDD.n6247 DVDD.n6246 0.00206274
R14411 DVDD.n3248 DVDD.n3247 0.00206274
R14412 DVDD.n3498 DVDD.n3497 0.00206274
R14413 DVDD.n7865 DVDD.n7864 0.00206274
R14414 DVDD.n8404 DVDD.n8403 0.00206274
R14415 DVDD.n9121 DVDD.n9120 0.00206274
R14416 DVDD.n8948 DVDD.n8947 0.00206274
R14417 DVDD.n9122 DVDD.n9121 0.00206274
R14418 DVDD.n8403 DVDD.n8402 0.00206274
R14419 DVDD.n8385 DVDD.n8384 0.00206274
R14420 DVDD.n7864 DVDD.n7863 0.00206274
R14421 DVDD.n3249 DVDD.n3248 0.00206274
R14422 DVDD.n3497 DVDD.n3496 0.00206274
R14423 DVDD.n8949 DVDD.n8948 0.00206274
R14424 DVDD.n19357 DVDD.n19356 0.00206
R14425 DVDD.n18336 DVDD.n18335 0.00206
R14426 DVDD.n11263 DVDD.n11262 0.00204286
R14427 DVDD.n11251 DVDD.n11250 0.00204286
R14428 DVDD.n11235 DVDD.n11234 0.00204286
R14429 DVDD.n5768 DVDD.n5766 0.00204286
R14430 DVDD.n301 DVDD.n300 0.00204286
R14431 DVDD.n412 DVDD.n410 0.00204286
R14432 DVDD.n384 DVDD.n383 0.00204286
R14433 DVDD.n413 DVDD.n409 0.00204286
R14434 DVDD.n487 DVDD.n486 0.00204286
R14435 DVDD.n441 DVDD.n440 0.00204286
R14436 DVDD.n532 DVDD.n531 0.00204286
R14437 DVDD.n643 DVDD.n641 0.00204286
R14438 DVDD.n615 DVDD.n614 0.00204286
R14439 DVDD.n644 DVDD.n640 0.00204286
R14440 DVDD.n719 DVDD.n718 0.00204286
R14441 DVDD.n673 DVDD.n672 0.00204286
R14442 DVDD.n11297 DVDD.n11296 0.00204286
R14443 DVDD.n11279 DVDD.n11278 0.00204286
R14444 DVDD.n12503 DVDD.n12502 0.00204286
R14445 DVDD.n5770 DVDD.n5769 0.00204286
R14446 DVDD.n15258 DVDD.n15257 0.00203682
R14447 DVDD.n15272 DVDD.n15271 0.00203682
R14448 DVDD.n15285 DVDD.n15284 0.00203682
R14449 DVDD.n15192 DVDD 0.00203682
R14450 DVDD.n16047 DVDD.n16046 0.00203533
R14451 DVDD.n16003 DVDD.n16002 0.00203533
R14452 DVDD.n16004 DVDD.n16003 0.00203533
R14453 DVDD.n16048 DVDD.n16047 0.00203533
R14454 DVDD.n15659 DVDD.n15658 0.00203533
R14455 DVDD.n15929 DVDD.n15928 0.00203533
R14456 DVDD.n15928 DVDD.n15927 0.00203533
R14457 DVDD.n15660 DVDD.n15659 0.00203533
R14458 DVDD.n8162 DVDD.n8161 0.00203533
R14459 DVDD.n8163 DVDD.n8162 0.00203533
R14460 DVDD.n8077 DVDD.n8076 0.00203533
R14461 DVDD.n12043 DVDD.n12042 0.00203146
R14462 DVDD.n12109 DVDD.n12108 0.00203145
R14463 DVDD.n7695 DVDD.n7155 0.00203
R14464 DVDD.n7699 DVDD.n7698 0.00203
R14465 DVDD.n3691 DVDD.n3690 0.00203
R14466 DVDD.n3687 DVDD.n3686 0.00203
R14467 DVDD.n18533 DVDD.n18532 0.00203
R14468 DVDD.n18537 DVDD.n18536 0.00203
R14469 DVDD.n18781 DVDD.n18780 0.00203
R14470 DVDD.n18779 DVDD.n18778 0.00203
R14471 DVDD.n2949 DVDD.n2948 0.00203
R14472 DVDD.n2953 DVDD.n2952 0.00203
R14473 DVDD.n9807 DVDD.n9806 0.00203
R14474 DVDD.n2187 DVDD.n2186 0.00203
R14475 DVDD.n2191 DVDD.n2190 0.00203
R14476 DVDD.n2247 DVDD.n2246 0.00203
R14477 DVDD.n2243 DVDD.n2242 0.00203
R14478 DVDD.n18902 DVDD.n18901 0.00203
R14479 DVDD.n18906 DVDD.n18905 0.00203
R14480 DVDD.n18934 DVDD.n18933 0.00203
R14481 DVDD.n18932 DVDD.n18931 0.00203
R14482 DVDD.n7105 DVDD.n7104 0.00203
R14483 DVDD.n7070 DVDD.n7069 0.00203
R14484 DVDD.n6808 DVDD.n6807 0.00203
R14485 DVDD.n1903 DVDD.n1902 0.00203
R14486 DVDD.n19966 DVDD.n19965 0.00203
R14487 DVDD.n19970 DVDD.n19969 0.00203
R14488 DVDD.n20026 DVDD.n20025 0.00203
R14489 DVDD.n20022 DVDD.n20021 0.00203
R14490 DVDD.n19020 DVDD.n19019 0.00203
R14491 DVDD.n19024 DVDD.n19023 0.00203
R14492 DVDD.n19052 DVDD.n19051 0.00203
R14493 DVDD.n19050 DVDD.n19049 0.00203
R14494 DVDD.n3884 DVDD.n3883 0.00203
R14495 DVDD.n4650 DVDD.n4649 0.00203
R14496 DVDD.n4845 DVDD.n4844 0.00203
R14497 DVDD.n19681 DVDD.n19680 0.00203
R14498 DVDD.n979 DVDD.n978 0.00203
R14499 DVDD.n975 DVDD.n974 0.00203
R14500 DVDD.n934 DVDD.n933 0.00203
R14501 DVDD.n930 DVDD.n929 0.00203
R14502 DVDD.n19229 DVDD.n19228 0.00203
R14503 DVDD.n19233 DVDD.n19232 0.00203
R14504 DVDD.n19434 DVDD.n19433 0.00203
R14505 DVDD.n19432 DVDD.n19431 0.00203
R14506 DVDD.n18330 DVDD.n18329 0.00203
R14507 DVDD.n18326 DVDD.n18325 0.00203
R14508 DVDD.n11908 DVDD.n11907 0.00203
R14509 DVDD.n1326 DVDD.n1325 0.00203
R14510 DVDD.n3277 DVDD.n3276 0.00203
R14511 DVDD.n14922 DVDD.n14921 0.00201875
R14512 DVDD.n14885 DVDD.n14884 0.00201875
R14513 DVDD.n15214 DVDD.n15213 0.00201875
R14514 DVDD.n15220 DVDD.n15219 0.00201875
R14515 DVDD.n15245 DVDD.n15244 0.00201875
R14516 DVDD.n15107 DVDD.n15106 0.00201875
R14517 DVDD.n15306 DVDD.n15305 0.00201875
R14518 DVDD.n15292 DVDD.n15291 0.00201875
R14519 DVDD.n15003 DVDD.n15002 0.00201875
R14520 DVDD.n16050 DVDD.n16049 0.00200628
R14521 DVDD.n16001 DVDD.n16000 0.00200628
R14522 DVDD.n15662 DVDD.n15661 0.00200628
R14523 DVDD.n15931 DVDD.n15930 0.00200628
R14524 DVDD.n8165 DVDD.n8164 0.00200628
R14525 DVDD.n8352 DVDD.n8351 0.00200628
R14526 DVDD.n7973 DVDD.n7972 0.00200628
R14527 DVDD.n1805 DVDD.n1804 0.002
R14528 DVDD.n15357 DVDD.n15356 0.002
R14529 DVDD.n11164 DVDD.n11163 0.002
R14530 DVDD.n16368 DVDD.n16367 0.002
R14531 DVDD.n3629 DVDD.n3628 0.002
R14532 DVDD.n5459 DVDD.n5458 0.00197427
R14533 DVDD.n1586 DVDD.n1585 0.0019742
R14534 DVDD.n12135 DVDD.n12134 0.0019742
R14535 DVDD.n13510 DVDD.n13509 0.0019742
R14536 DVDD.n13562 DVDD.n13561 0.0019742
R14537 DVDD.n13603 DVDD.n13602 0.0019742
R14538 DVDD.n13643 DVDD.n13642 0.0019742
R14539 DVDD.n13684 DVDD.n13683 0.0019742
R14540 DVDD.n12134 DVDD.n12133 0.0019742
R14541 DVDD.n13509 DVDD.n13508 0.0019742
R14542 DVDD.n13602 DVDD.n13601 0.0019742
R14543 DVDD.n13561 DVDD.n13560 0.0019742
R14544 DVDD.n13683 DVDD.n13682 0.0019742
R14545 DVDD.n13642 DVDD.n13641 0.0019742
R14546 DVDD.n15409 DVDD.n15408 0.0019742
R14547 DVDD.n15453 DVDD.n15452 0.0019742
R14548 DVDD.n14694 DVDD.n14693 0.0019742
R14549 DVDD.n14611 DVDD.n14610 0.0019742
R14550 DVDD.n14557 DVDD.n14556 0.0019742
R14551 DVDD.n14513 DVDD.n14512 0.0019742
R14552 DVDD.n14469 DVDD.n14468 0.0019742
R14553 DVDD.n14409 DVDD.n14408 0.0019742
R14554 DVDD.n14410 DVDD.n14409 0.0019742
R14555 DVDD.n14514 DVDD.n14513 0.0019742
R14556 DVDD.n14695 DVDD.n14694 0.0019742
R14557 DVDD.n14612 DVDD.n14611 0.0019742
R14558 DVDD.n15452 DVDD.n15451 0.0019742
R14559 DVDD.n15408 DVDD.n15407 0.0019742
R14560 DVDD.n14558 DVDD.n14557 0.0019742
R14561 DVDD.n14470 DVDD.n14469 0.0019742
R14562 DVDD.n4916 DVDD.n4915 0.0019742
R14563 DVDD.n5315 DVDD.n5314 0.0019742
R14564 DVDD.n5476 DVDD.n5475 0.0019742
R14565 DVDD.n5599 DVDD.n5598 0.0019742
R14566 DVDD.n5687 DVDD.n5686 0.0019742
R14567 DVDD.n5967 DVDD.n5966 0.0019742
R14568 DVDD.n5686 DVDD.n5685 0.0019742
R14569 DVDD.n5968 DVDD.n5967 0.0019742
R14570 DVDD.n5314 DVDD.n5313 0.0019742
R14571 DVDD.n5475 DVDD.n5474 0.0019742
R14572 DVDD.n5195 DVDD.n5194 0.0019742
R14573 DVDD.n5598 DVDD.n5597 0.0019742
R14574 DVDD.n13143 DVDD.n13142 0.0019742
R14575 DVDD.n12987 DVDD.n12986 0.0019742
R14576 DVDD.n12828 DVDD.n12827 0.0019742
R14577 DVDD.n12754 DVDD.n12753 0.0019742
R14578 DVDD.n12630 DVDD.n12629 0.0019742
R14579 DVDD.n12988 DVDD.n12987 0.0019742
R14580 DVDD.n13144 DVDD.n13143 0.0019742
R14581 DVDD.n12631 DVDD.n12630 0.0019742
R14582 DVDD.n12755 DVDD.n12754 0.0019742
R14583 DVDD.n12829 DVDD.n12828 0.0019742
R14584 DVDD.n18193 DVDD.n18192 0.0019742
R14585 DVDD.n18152 DVDD.n18151 0.0019742
R14586 DVDD.n18049 DVDD.n18048 0.0019742
R14587 DVDD.n17971 DVDD.n17970 0.0019742
R14588 DVDD.n17919 DVDD.n17918 0.0019742
R14589 DVDD.n17878 DVDD.n17877 0.0019742
R14590 DVDD.n17838 DVDD.n17837 0.0019742
R14591 DVDD.n17783 DVDD.n17782 0.0019742
R14592 DVDD.n17784 DVDD.n17783 0.0019742
R14593 DVDD.n18050 DVDD.n18049 0.0019742
R14594 DVDD.n17972 DVDD.n17971 0.0019742
R14595 DVDD.n18153 DVDD.n18152 0.0019742
R14596 DVDD.n18194 DVDD.n18193 0.0019742
R14597 DVDD.n17879 DVDD.n17878 0.0019742
R14598 DVDD.n17920 DVDD.n17919 0.0019742
R14599 DVDD.n17839 DVDD.n17838 0.0019742
R14600 DVDD.n6446 DVDD.n6445 0.0019742
R14601 DVDD.n6283 DVDD.n6282 0.0019742
R14602 DVDD.n6206 DVDD.n6205 0.0019742
R14603 DVDD.n6138 DVDD.n6137 0.0019742
R14604 DVDD.n4430 DVDD.n4429 0.0019742
R14605 DVDD.n4431 DVDD.n4430 0.0019742
R14606 DVDD.n6284 DVDD.n6283 0.0019742
R14607 DVDD.n6447 DVDD.n6446 0.0019742
R14608 DVDD.n6337 DVDD.n6336 0.0019742
R14609 DVDD.n6139 DVDD.n6138 0.0019742
R14610 DVDD.n6207 DVDD.n6206 0.0019742
R14611 DVDD.n9232 DVDD.n9231 0.0019742
R14612 DVDD.n9069 DVDD.n9068 0.0019742
R14613 DVDD.n8908 DVDD.n8907 0.0019742
R14614 DVDD.n8840 DVDD.n8839 0.0019742
R14615 DVDD.n8704 DVDD.n8703 0.0019742
R14616 DVDD.n8841 DVDD.n8840 0.0019742
R14617 DVDD.n8705 DVDD.n8704 0.0019742
R14618 DVDD.n9233 DVDD.n9232 0.0019742
R14619 DVDD.n9070 DVDD.n9069 0.0019742
R14620 DVDD.n9123 DVDD.n9122 0.0019742
R14621 DVDD.n8909 DVDD.n8908 0.0019742
R14622 DVDD.n8212 DVDD.n8211 0.00197069
R14623 DVDD.n16415 DVDD.n16414 0.00196667
R14624 DVDD.n10987 DVDD.n10936 0.00196667
R14625 DVDD.n10986 DVDD.n10985 0.00196667
R14626 DVDD.n10961 DVDD.n10960 0.00196667
R14627 DVDD.n10245 DVDD.n10230 0.00196667
R14628 DVDD.n14917 DVDD.n14916 0.0019625
R14629 DVDD.n14923 DVDD.n14922 0.0019625
R14630 DVDD.n14886 DVDD.n14885 0.0019625
R14631 DVDD.n15215 DVDD.n15214 0.0019625
R14632 DVDD.n15221 DVDD.n15220 0.0019625
R14633 DVDD.n15238 DVDD.n15237 0.0019625
R14634 DVDD.n15310 DVDD.n15309 0.0019625
R14635 DVDD.n15296 DVDD.n15295 0.0019625
R14636 DVDD.n14999 DVDD.n14998 0.0019625
R14637 DVDD.n17198 DVDD.n17197 0.00195724
R14638 DVDD.n17197 DVDD.n17196 0.00195724
R14639 DVDD.n17365 DVDD.n17364 0.00195724
R14640 DVDD.n17364 DVDD.n17363 0.00195724
R14641 DVDD.n17525 DVDD.n17524 0.00195724
R14642 DVDD.n17526 DVDD.n17525 0.00195724
R14643 DVDD.n16033 DVDD.n16032 0.00194123
R14644 DVDD.n16017 DVDD.n16016 0.00194123
R14645 DVDD.n16034 DVDD.n16033 0.00194123
R14646 DVDD.n16018 DVDD.n16017 0.00194123
R14647 DVDD.n15645 DVDD.n15644 0.00194123
R14648 DVDD.n15629 DVDD.n15628 0.00194123
R14649 DVDD.n15646 DVDD.n15645 0.00194123
R14650 DVDD.n15630 DVDD.n15629 0.00194123
R14651 DVDD.n8148 DVDD.n8147 0.00194123
R14652 DVDD.n8149 DVDD.n8148 0.00194123
R14653 DVDD.n8315 DVDD.n8314 0.00194123
R14654 DVDD.n8013 DVDD.n8012 0.00194123
R14655 DVDD.n15259 DVDD.n15258 0.00194077
R14656 DVDD.n18744 DVDD.n18743 0.00194
R14657 DVDD.n18747 DVDD.n18746 0.00194
R14658 DVDD.n18750 DVDD.n18749 0.00194
R14659 DVDD.n18753 DVDD.n18752 0.00194
R14660 DVDD.n18756 DVDD.n18755 0.00194
R14661 DVDD.n18759 DVDD.n18758 0.00194
R14662 DVDD.n18762 DVDD.n18761 0.00194
R14663 DVDD.n18765 DVDD.n18764 0.00194
R14664 DVDD.n18768 DVDD.n18767 0.00194
R14665 DVDD.n18771 DVDD.n18770 0.00194
R14666 DVDD.n9759 DVDD.n9758 0.00194
R14667 DVDD.n9777 DVDD.n9776 0.00194
R14668 DVDD.n9790 DVDD.n9789 0.00194
R14669 DVDD.n7909 DVDD.n7908 0.00194
R14670 DVDD.n9249 DVDD.n9248 0.00194
R14671 DVDD.n9278 DVDD.n9277 0.00194
R14672 DVDD.n9291 DVDD.n9290 0.00194
R14673 DVDD.n6856 DVDD.n6855 0.00194
R14674 DVDD.n6838 DVDD.n6837 0.00194
R14675 DVDD.n6825 DVDD.n6824 0.00194
R14676 DVDD.n6546 DVDD.n6545 0.00194
R14677 DVDD.n3993 DVDD.n3992 0.00194
R14678 DVDD.n3964 DVDD.n3963 0.00194
R14679 DVDD.n3951 DVDD.n3950 0.00194
R14680 DVDD.n4893 DVDD.n4892 0.00194
R14681 DVDD.n4875 DVDD.n4874 0.00194
R14682 DVDD.n4862 DVDD.n4861 0.00194
R14683 DVDD.n5137 DVDD.n5136 0.00194
R14684 DVDD.n5298 DVDD.n5297 0.00194
R14685 DVDD.n5269 DVDD.n5268 0.00194
R14686 DVDD.n5256 DVDD.n5255 0.00194
R14687 DVDD.n1751 DVDD.n1750 0.00194
R14688 DVDD.n1748 DVDD.n1747 0.00194
R14689 DVDD.n1745 DVDD.n1744 0.00194
R14690 DVDD.n19258 DVDD.n19257 0.00194
R14691 DVDD.n19261 DVDD.n19260 0.00194
R14692 DVDD.n19264 DVDD.n19263 0.00194
R14693 DVDD.n19267 DVDD.n19266 0.00194
R14694 DVDD.n19418 DVDD.n19417 0.00194
R14695 DVDD.n19421 DVDD.n19420 0.00194
R14696 DVDD.n19424 DVDD.n19423 0.00194
R14697 DVDD.n11860 DVDD.n11859 0.00194
R14698 DVDD.n11878 DVDD.n11877 0.00194
R14699 DVDD.n11891 DVDD.n11890 0.00194
R14700 DVDD.n11311 DVDD.n11310 0.00194
R14701 DVDD.n10731 DVDD.n10730 0.00194
R14702 DVDD.n10353 DVDD.n10351 0.00194
R14703 DVDD.n10354 DVDD.n10353 0.00194
R14704 DVDD.n10732 DVDD.n10654 0.00194
R14705 DVDD.n13160 DVDD.n13159 0.00194
R14706 DVDD.n13189 DVDD.n13188 0.00194
R14707 DVDD.n13202 DVDD.n13201 0.00194
R14708 DVDD.n16507 DVDD.n16506 0.00194
R14709 DVDD.n16508 DVDD.n16507 0.00194
R14710 DVDD.n17158 DVDD.n17152 0.00194
R14711 DVDD.n16849 DVDD.n16848 0.00194
R14712 DVDD.n16850 DVDD.n16849 0.00194
R14713 DVDD.n17043 DVDD.n16879 0.00194
R14714 DVDD.n16816 DVDD.n16744 0.00194
R14715 DVDD.n16694 DVDD.n16576 0.00194
R14716 DVDD.n17157 DVDD.n17156 0.00194
R14717 DVDD.n1224 DVDD.n1223 0.00191732
R14718 DVDD.n1161 DVDD.n1160 0.00191732
R14719 DVDD.n911 DVDD.n910 0.00191732
R14720 DVDD.n869 DVDD.n868 0.00191732
R14721 DVDD.n866 DVDD.n865 0.00191732
R14722 DVDD.n19286 DVDD.n19285 0.00191732
R14723 DVDD.n11441 DVDD.n11440 0.00191732
R14724 DVDD.n11445 DVDD.n11444 0.00191732
R14725 DVDD.n12028 DVDD.n12027 0.00191732
R14726 DVDD.n12278 DVDD.n12277 0.00191732
R14727 DVDD.n13313 DVDD.n13312 0.00191732
R14728 DVDD.n13507 DVDD.n13506 0.00191732
R14729 DVDD.n13559 DVDD.n13558 0.00191732
R14730 DVDD.n13605 DVDD.n13604 0.00191732
R14731 DVDD.n13640 DVDD.n13639 0.00191732
R14732 DVDD.n13686 DVDD.n13685 0.00191732
R14733 DVDD.n2754 DVDD.n2753 0.00191732
R14734 DVDD.n2795 DVDD.n2794 0.00191732
R14735 DVDD.n18568 DVDD.n18567 0.00191732
R14736 DVDD.n18679 DVDD.n18678 0.00191732
R14737 DVDD.n14812 DVDD.n14811 0.00191732
R14738 DVDD.n15406 DVDD.n15405 0.00191732
R14739 DVDD.n15455 DVDD.n15454 0.00191732
R14740 DVDD.n14697 DVDD.n14696 0.00191732
R14741 DVDD.n14614 DVDD.n14613 0.00191732
R14742 DVDD.n14560 DVDD.n14559 0.00191732
R14743 DVDD.n14511 DVDD.n14510 0.00191732
R14744 DVDD.n14472 DVDD.n14471 0.00191732
R14745 DVDD.n14407 DVDD.n14406 0.00191732
R14746 DVDD.n19758 DVDD.n19757 0.00191732
R14747 DVDD.n19857 DVDD.n19856 0.00191732
R14748 DVDD.n19925 DVDD.n19924 0.00191732
R14749 DVDD.n20057 DVDD.n20056 0.00191732
R14750 DVDD.n20204 DVDD.n20203 0.00191732
R14751 DVDD.n20194 DVDD.n20193 0.00191732
R14752 DVDD.n20181 DVDD.n20180 0.00191732
R14753 DVDD.n19014 DVDD.n19013 0.00191732
R14754 DVDD.n19013 DVDD.n19012 0.00191732
R14755 DVDD.n19010 DVDD.n19009 0.00191732
R14756 DVDD.n3888 DVDD.n3875 0.00191732
R14757 DVDD.n4818 DVDD.n4817 0.00191732
R14758 DVDD.n4901 DVDD.n4900 0.00191732
R14759 DVDD.n4945 DVDD.n4944 0.00191732
R14760 DVDD.n4956 DVDD.n4955 0.00191732
R14761 DVDD.n4959 DVDD.n4958 0.00191732
R14762 DVDD.n4961 DVDD.n4960 0.00191732
R14763 DVDD.n4980 DVDD.n4979 0.00191732
R14764 DVDD.n5062 DVDD.n5061 0.00191732
R14765 DVDD.n5104 DVDD.n5103 0.00191732
R14766 DVDD.n5309 DVDD.n5308 0.00191732
R14767 DVDD.n5326 DVDD.n5325 0.00191732
R14768 DVDD.n5395 DVDD.n5394 0.00191732
R14769 DVDD.n5415 DVDD.n5414 0.00191732
R14770 DVDD.n5473 DVDD.n5472 0.00191732
R14771 DVDD.n5596 DVDD.n5595 0.00191732
R14772 DVDD.n5628 DVDD.n5627 0.00191732
R14773 DVDD.n5689 DVDD.n5688 0.00191732
R14774 DVDD.n6052 DVDD.n6051 0.00191732
R14775 DVDD.n5965 DVDD.n5964 0.00191732
R14776 DVDD.n1403 DVDD.n1402 0.00191732
R14777 DVDD.n1519 DVDD.n1518 0.00191732
R14778 DVDD.n1491 DVDD.n1490 0.00191732
R14779 DVDD.n1452 DVDD.n1451 0.00191732
R14780 DVDD.n1716 DVDD.n1715 0.00191732
R14781 DVDD.n282 DVDD.n281 0.00191732
R14782 DVDD.n272 DVDD.n271 0.00191732
R14783 DVDD.n259 DVDD.n258 0.00191732
R14784 DVDD.n19223 DVDD.n19222 0.00191732
R14785 DVDD.n19222 DVDD.n19221 0.00191732
R14786 DVDD.n19219 DVDD.n19218 0.00191732
R14787 DVDD.n18332 DVDD.n10122 0.00191732
R14788 DVDD.n11644 DVDD.n11643 0.00191732
R14789 DVDD.n11852 DVDD.n11851 0.00191732
R14790 DVDD.n11808 DVDD.n11807 0.00191732
R14791 DVDD.n11797 DVDD.n11796 0.00191732
R14792 DVDD.n11794 DVDD.n11793 0.00191732
R14793 DVDD.n11792 DVDD.n11791 0.00191732
R14794 DVDD.n11773 DVDD.n11772 0.00191732
R14795 DVDD.n11692 DVDD.n11691 0.00191732
R14796 DVDD.n11688 DVDD.n11687 0.00191732
R14797 DVDD.n11651 DVDD.n11650 0.00191732
R14798 DVDD.n13149 DVDD.n13148 0.00191732
R14799 DVDD.n13133 DVDD.n13132 0.00191732
R14800 DVDD.n13066 DVDD.n13065 0.00191732
R14801 DVDD.n13047 DVDD.n13046 0.00191732
R14802 DVDD.n12990 DVDD.n12989 0.00191732
R14803 DVDD.n12831 DVDD.n12830 0.00191732
R14804 DVDD.n12809 DVDD.n12808 0.00191732
R14805 DVDD.n12752 DVDD.n12751 0.00191732
R14806 DVDD.n12698 DVDD.n12697 0.00191732
R14807 DVDD.n12628 DVDD.n12627 0.00191732
R14808 DVDD.n790 DVDD.n789 0.00191732
R14809 DVDD.n827 DVDD.n826 0.00191732
R14810 DVDD.n237 DVDD.n236 0.00191732
R14811 DVDD.n158 DVDD.n157 0.00191732
R14812 DVDD.n18226 DVDD.n18225 0.00191732
R14813 DVDD.n18196 DVDD.n18195 0.00191732
R14814 DVDD.n18150 DVDD.n18149 0.00191732
R14815 DVDD.n18052 DVDD.n18051 0.00191732
R14816 DVDD.n17974 DVDD.n17973 0.00191732
R14817 DVDD.n17922 DVDD.n17921 0.00191732
R14818 DVDD.n17876 DVDD.n17875 0.00191732
R14819 DVDD.n17841 DVDD.n17840 0.00191732
R14820 DVDD.n17781 DVDD.n17780 0.00191732
R14821 DVDD.n1980 DVDD.n1979 0.00191732
R14822 DVDD.n2079 DVDD.n2078 0.00191732
R14823 DVDD.n2107 DVDD.n2106 0.00191732
R14824 DVDD.n2146 DVDD.n2145 0.00191732
R14825 DVDD.n2278 DVDD.n2277 0.00191732
R14826 DVDD.n19589 DVDD.n19588 0.00191732
R14827 DVDD.n19579 DVDD.n19578 0.00191732
R14828 DVDD.n19566 DVDD.n19565 0.00191732
R14829 DVDD.n18941 DVDD.n18940 0.00191732
R14830 DVDD.n18940 DVDD.n18939 0.00191732
R14831 DVDD.n18937 DVDD.n18936 0.00191732
R14832 DVDD.n7109 DVDD.n7096 0.00191732
R14833 DVDD.n6866 DVDD.n6865 0.00191732
R14834 DVDD.n6783 DVDD.n6782 0.00191732
R14835 DVDD.n6739 DVDD.n6738 0.00191732
R14836 DVDD.n6728 DVDD.n6727 0.00191732
R14837 DVDD.n6725 DVDD.n6724 0.00191732
R14838 DVDD.n6723 DVDD.n6722 0.00191732
R14839 DVDD.n6704 DVDD.n6703 0.00191732
R14840 DVDD.n6620 DVDD.n6619 0.00191732
R14841 DVDD.n6616 DVDD.n6615 0.00191732
R14842 DVDD.n6578 DVDD.n6577 0.00191732
R14843 DVDD.n6452 DVDD.n6451 0.00191732
R14844 DVDD.n6435 DVDD.n6434 0.00191732
R14845 DVDD.n6366 DVDD.n6365 0.00191732
R14846 DVDD.n6346 DVDD.n6345 0.00191732
R14847 DVDD.n6286 DVDD.n6285 0.00191732
R14848 DVDD.n6209 DVDD.n6208 0.00191732
R14849 DVDD.n6188 DVDD.n6187 0.00191732
R14850 DVDD.n6136 DVDD.n6135 0.00191732
R14851 DVDD.n4509 DVDD.n4508 0.00191732
R14852 DVDD.n4428 DVDD.n4427 0.00191732
R14853 DVDD.n3200 DVDD.n3199 0.00191732
R14854 DVDD.n3478 DVDD.n3477 0.00191732
R14855 DVDD.n3506 DVDD.n3505 0.00191732
R14856 DVDD.n3545 DVDD.n3544 0.00191732
R14857 DVDD.n3722 DVDD.n3721 0.00191732
R14858 DVDD.n3768 DVDD.n3767 0.00191732
R14859 DVDD.n3758 DVDD.n3757 0.00191732
R14860 DVDD.n3745 DVDD.n3744 0.00191732
R14861 DVDD.n18527 DVDD.n18526 0.00191732
R14862 DVDD.n18526 DVDD.n18525 0.00191732
R14863 DVDD.n18523 DVDD.n18522 0.00191732
R14864 DVDD.n10054 DVDD.n7154 0.00191732
R14865 DVDD.n7900 DVDD.n7899 0.00191732
R14866 DVDD.n9751 DVDD.n9750 0.00191732
R14867 DVDD.n9707 DVDD.n9706 0.00191732
R14868 DVDD.n9696 DVDD.n9695 0.00191732
R14869 DVDD.n9693 DVDD.n9692 0.00191732
R14870 DVDD.n9691 DVDD.n9690 0.00191732
R14871 DVDD.n9672 DVDD.n9671 0.00191732
R14872 DVDD.n9588 DVDD.n9587 0.00191732
R14873 DVDD.n9584 DVDD.n9583 0.00191732
R14874 DVDD.n9546 DVDD.n9545 0.00191732
R14875 DVDD.n9238 DVDD.n9237 0.00191732
R14876 DVDD.n9221 DVDD.n9220 0.00191732
R14877 DVDD.n9152 DVDD.n9151 0.00191732
R14878 DVDD.n9132 DVDD.n9131 0.00191732
R14879 DVDD.n9072 DVDD.n9071 0.00191732
R14880 DVDD.n8911 DVDD.n8910 0.00191732
R14881 DVDD.n8890 DVDD.n8889 0.00191732
R14882 DVDD.n8838 DVDD.n8837 0.00191732
R14883 DVDD.n8783 DVDD.n8782 0.00191732
R14884 DVDD.n8702 DVDD.n8701 0.00191732
R14885 DVDD.n7077 DVDD.n7076 0.00191
R14886 DVDD.n4602 DVDD.n3889 0.00191
R14887 DVDD.n10185 DVDD.n10184 0.00191
R14888 DVDD.n10429 DVDD.n10428 0.00191
R14889 DVDD.n17062 DVDD.n17060 0.00191
R14890 DVDD.n14743 DVDD.n14742 0.00191
R14891 DVDD.n10402 DVDD.n10401 0.00190625
R14892 DVDD.n10589 DVDD.n10588 0.00190625
R14893 DVDD.n10635 DVDD.n10634 0.00190625
R14894 DVDD.n3119 DVDD.n3118 0.00190625
R14895 DVDD.n3101 DVDD.n3100 0.00190625
R14896 DVDD.n3100 DVDD.n3099 0.00190625
R14897 DVDD.n3094 DVDD.n3093 0.00190625
R14898 DVDD.n3080 DVDD.n3079 0.00190625
R14899 DVDD.n3074 DVDD.n3073 0.00190625
R14900 DVDD.n3067 DVDD.n3066 0.00190625
R14901 DVDD.n3058 DVDD.n3057 0.00190625
R14902 DVDD.n3042 DVDD.n3041 0.00190625
R14903 DVDD.n3040 DVDD.n3039 0.00190625
R14904 DVDD.n3065 DVDD.n3064 0.00190384
R14905 DVDD.n3066 DVDD.n3065 0.00190384
R14906 DVDD.n15148 DVDD.n15147 0.0019
R14907 DVDD.n3328 DVDD.n3327 0.00188889
R14908 DVDD.n12069 DVDD.n12068 0.00188565
R14909 DVDD.n13352 DVDD.n13351 0.00188565
R14910 DVDD.n13524 DVDD.n13523 0.00188565
R14911 DVDD.n13576 DVDD.n13575 0.00188565
R14912 DVDD.n13589 DVDD.n13588 0.00188565
R14913 DVDD.n13657 DVDD.n13656 0.00188565
R14914 DVDD.n13670 DVDD.n13669 0.00188565
R14915 DVDD.n12068 DVDD.n12067 0.00188565
R14916 DVDD.n13351 DVDD.n13350 0.00188565
R14917 DVDD.n13523 DVDD.n13522 0.00188565
R14918 DVDD.n13575 DVDD.n13574 0.00188565
R14919 DVDD.n13588 DVDD.n13587 0.00188565
R14920 DVDD.n13656 DVDD.n13655 0.00188565
R14921 DVDD.n13669 DVDD.n13668 0.00188565
R14922 DVDD.n15423 DVDD.n15422 0.00188565
R14923 DVDD.n15439 DVDD.n15438 0.00188565
R14924 DVDD.n14680 DVDD.n14679 0.00188565
R14925 DVDD.n14597 DVDD.n14596 0.00188565
R14926 DVDD.n14543 DVDD.n14542 0.00188565
R14927 DVDD.n14527 DVDD.n14526 0.00188565
R14928 DVDD.n14455 DVDD.n14454 0.00188565
R14929 DVDD.n14424 DVDD.n14423 0.00188565
R14930 DVDD.n14456 DVDD.n14455 0.00188565
R14931 DVDD.n14544 DVDD.n14543 0.00188565
R14932 DVDD.n14598 DVDD.n14597 0.00188565
R14933 DVDD.n14681 DVDD.n14680 0.00188565
R14934 DVDD.n15422 DVDD.n15421 0.00188565
R14935 DVDD.n15438 DVDD.n15437 0.00188565
R14936 DVDD.n14425 DVDD.n14424 0.00188565
R14937 DVDD.n14528 DVDD.n14527 0.00188565
R14938 DVDD.n19728 DVDD.n19727 0.00188565
R14939 DVDD.n4936 DVDD.n4935 0.00188565
R14940 DVDD.n4965 DVDD.n4964 0.00188565
R14941 DVDD.n5346 DVDD.n5345 0.00188565
R14942 DVDD.n5490 DVDD.n5489 0.00188565
R14943 DVDD.n5630 DVDD.n5629 0.00188565
R14944 DVDD.n5650 DVDD.n5649 0.00188565
R14945 DVDD.n6023 DVDD.n6022 0.00188565
R14946 DVDD.n5982 DVDD.n5981 0.00188565
R14947 DVDD.n5629 DVDD.n5628 0.00188565
R14948 DVDD.n6024 DVDD.n6023 0.00188565
R14949 DVDD.n5345 DVDD.n5344 0.00188565
R14950 DVDD.n4964 DVDD.n4963 0.00188565
R14951 DVDD.n4935 DVDD.n4934 0.00188565
R14952 DVDD.n5983 DVDD.n5982 0.00188565
R14953 DVDD.n5649 DVDD.n5648 0.00188565
R14954 DVDD.n5489 DVDD.n5488 0.00188565
R14955 DVDD.n11817 DVDD.n11816 0.00188565
R14956 DVDD.n11788 DVDD.n11787 0.00188565
R14957 DVDD.n12973 DVDD.n12972 0.00188565
R14958 DVDD.n12807 DVDD.n12806 0.00188565
R14959 DVDD.n12787 DVDD.n12786 0.00188565
R14960 DVDD.n12674 DVDD.n12673 0.00188565
R14961 DVDD.n12645 DVDD.n12644 0.00188565
R14962 DVDD.n13114 DVDD.n13113 0.00188565
R14963 DVDD.n12974 DVDD.n12973 0.00188565
R14964 DVDD.n11818 DVDD.n11817 0.00188565
R14965 DVDD.n11789 DVDD.n11788 0.00188565
R14966 DVDD.n1373 DVDD.n1372 0.00188565
R14967 DVDD.n12374 DVDD.n12373 0.00188565
R14968 DVDD.n1390 DVDD.n1389 0.00188565
R14969 DVDD.n12646 DVDD.n12645 0.00188565
R14970 DVDD.n12675 DVDD.n12674 0.00188565
R14971 DVDD.n12808 DVDD.n12807 0.00188565
R14972 DVDD.n12788 DVDD.n12787 0.00188565
R14973 DVDD.n18179 DVDD.n18178 0.00188565
R14974 DVDD.n18166 DVDD.n18165 0.00188565
R14975 DVDD.n18035 DVDD.n18034 0.00188565
R14976 DVDD.n17957 DVDD.n17956 0.00188565
R14977 DVDD.n17905 DVDD.n17904 0.00188565
R14978 DVDD.n17892 DVDD.n17891 0.00188565
R14979 DVDD.n17824 DVDD.n17823 0.00188565
R14980 DVDD.n17798 DVDD.n17797 0.00188565
R14981 DVDD.n18036 DVDD.n18035 0.00188565
R14982 DVDD.n18180 DVDD.n18179 0.00188565
R14983 DVDD.n18167 DVDD.n18166 0.00188565
R14984 DVDD.n17825 DVDD.n17824 0.00188565
R14985 DVDD.n17799 DVDD.n17798 0.00188565
R14986 DVDD.n17906 DVDD.n17905 0.00188565
R14987 DVDD.n17893 DVDD.n17892 0.00188565
R14988 DVDD.n17958 DVDD.n17957 0.00188565
R14989 DVDD.n6748 DVDD.n6747 0.00188565
R14990 DVDD.n6719 DVDD.n6718 0.00188565
R14991 DVDD.n6415 DVDD.n6414 0.00188565
R14992 DVDD.n6269 DVDD.n6268 0.00188565
R14993 DVDD.n6164 DVDD.n6163 0.00188565
R14994 DVDD.n4474 DVDD.n4473 0.00188565
R14995 DVDD.n4445 DVDD.n4444 0.00188565
R14996 DVDD.n4475 DVDD.n4474 0.00188565
R14997 DVDD.n6416 DVDD.n6415 0.00188565
R14998 DVDD.n6488 DVDD.n6487 0.00188565
R14999 DVDD.n6720 DVDD.n6719 0.00188565
R15000 DVDD.n6749 DVDD.n6748 0.00188565
R15001 DVDD.n1950 DVDD.n1949 0.00188565
R15002 DVDD.n1967 DVDD.n1966 0.00188565
R15003 DVDD.n6270 DVDD.n6269 0.00188565
R15004 DVDD.n6187 DVDD.n6186 0.00188565
R15005 DVDD.n4446 DVDD.n4445 0.00188565
R15006 DVDD.n6165 DVDD.n6164 0.00188565
R15007 DVDD.n9716 DVDD.n9715 0.00188565
R15008 DVDD.n9687 DVDD.n9686 0.00188565
R15009 DVDD.n9201 DVDD.n9200 0.00188565
R15010 DVDD.n9055 DVDD.n9054 0.00188565
R15011 DVDD.n8866 DVDD.n8865 0.00188565
R15012 DVDD.n8760 DVDD.n8759 0.00188565
R15013 DVDD.n8719 DVDD.n8718 0.00188565
R15014 DVDD.n9717 DVDD.n9716 0.00188565
R15015 DVDD.n9202 DVDD.n9201 0.00188565
R15016 DVDD.n9056 DVDD.n9055 0.00188565
R15017 DVDD.n8889 DVDD.n8888 0.00188565
R15018 DVDD.n8761 DVDD.n8760 0.00188565
R15019 DVDD.n8395 DVDD.n8394 0.00188565
R15020 DVDD.n9688 DVDD.n9687 0.00188565
R15021 DVDD.n3230 DVDD.n3229 0.00188565
R15022 DVDD.n3213 DVDD.n3212 0.00188565
R15023 DVDD.n8720 DVDD.n8719 0.00188565
R15024 DVDD.n8867 DVDD.n8866 0.00188565
R15025 DVDD.n2469 DVDD.n2468 0.00186769
R15026 DVDD.n2470 DVDD.n2469 0.00186769
R15027 DVDD.n16440 DVDD.n16439 0.00186
R15028 DVDD.n10912 DVDD.n10911 0.00186
R15029 DVDD.n10887 DVDD.n10886 0.00186
R15030 DVDD.n10862 DVDD.n10861 0.00186
R15031 DVDD.n10292 DVDD.n10269 0.00186
R15032 DVDD.n3709 DVDD.n3708 0.00185
R15033 DVDD.n18555 DVDD.n18554 0.00185
R15034 DVDD.n18774 DVDD.n18773 0.00185
R15035 DVDD.n2931 DVDD.n2930 0.00185
R15036 DVDD.n2939 DVDD.n2938 0.00185
R15037 DVDD.n9884 DVDD.n9883 0.00185
R15038 DVDD.n8364 DVDD.n8363 0.00185
R15039 DVDD.n9240 DVDD.n8365 0.00185
R15040 DVDD.n2169 DVDD.n2168 0.00185
R15041 DVDD.n2177 DVDD.n2176 0.00185
R15042 DVDD.n2265 DVDD.n2264 0.00185
R15043 DVDD.n18924 DVDD.n18923 0.00185
R15044 DVDD.n1885 DVDD.n1884 0.00185
R15045 DVDD.n1874 DVDD.n1873 0.00185
R15046 DVDD.n3926 DVDD.n3925 0.00185
R15047 DVDD.n4001 DVDD.n3927 0.00185
R15048 DVDD.n18821 DVDD.n18820 0.00185
R15049 DVDD.n19948 DVDD.n19947 0.00185
R15050 DVDD.n19956 DVDD.n19955 0.00185
R15051 DVDD.n20044 DVDD.n20043 0.00185
R15052 DVDD.n19042 DVDD.n19041 0.00185
R15053 DVDD.n19663 DVDD.n19662 0.00185
R15054 DVDD.n19652 DVDD.n19651 0.00185
R15055 DVDD.n5231 DVDD.n5230 0.00185
R15056 DVDD.n5306 DVDD.n5232 0.00185
R15057 DVDD.n997 DVDD.n996 0.00185
R15058 DVDD.n989 DVDD.n988 0.00185
R15059 DVDD.n2474 DVDD.n2473 0.00185
R15060 DVDD.n952 DVDD.n951 0.00185
R15061 DVDD.n19251 DVDD.n19250 0.00185
R15062 DVDD.n19427 DVDD.n19426 0.00185
R15063 DVDD.n19153 DVDD.n19152 0.00185
R15064 DVDD.n3848 DVDD.n3847 0.00185
R15065 DVDD.n7614 DVDD.n7613 0.00185
R15066 DVDD.n3902 DVDD.n3901 0.00185
R15067 DVDD.n7641 DVDD.n7640 0.00185
R15068 DVDD.n133 DVDD.n132 0.00185
R15069 DVDD.n19598 DVDD.n19597 0.00185
R15070 DVDD.n19466 DVDD.n19465 0.00185
R15071 DVDD.n20213 DVDD.n20212 0.00185
R15072 DVDD.n20081 DVDD.n20080 0.00185
R15073 DVDD.n3791 DVDD.n3790 0.00185
R15074 DVDD.n20282 DVDD.n20281 0.00185
R15075 DVDD.n20329 DVDD.n20328 0.00185
R15076 DVDD.n145 DVDD.n144 0.00185
R15077 DVDD.n11985 DVDD.n11984 0.00185
R15078 DVDD.n1308 DVDD.n1307 0.00185
R15079 DVDD.n1297 DVDD.n1296 0.00185
R15080 DVDD.n15314 DVDD.n14903 0.00185
R15081 DVDD.n15311 DVDD.n15119 0.00185
R15082 DVDD.n14869 DVDD.n14868 0.00185
R15083 DVDD.n10479 DVDD.n10478 0.00185
R15084 DVDD.n10670 DVDD.n10669 0.00185
R15085 DVDD.n10682 DVDD.n10681 0.00185
R15086 DVDD.n10615 DVDD.n10614 0.00185
R15087 DVDD.n10401 DVDD.n10400 0.00185
R15088 DVDD.n10568 DVDD.n10567 0.00185
R15089 DVDD.n10590 DVDD.n10589 0.00185
R15090 DVDD.n11302 DVDD.n11301 0.00185
R15091 DVDD.n13151 DVDD.n11303 0.00185
R15092 DVDD.n16998 DVDD.n16996 0.00185
R15093 DVDD.n16940 DVDD.n16938 0.00185
R15094 DVDD.n16151 DVDD.n16150 0.00185
R15095 DVDD.n16269 DVDD.n16268 0.00185
R15096 DVDD.n16773 DVDD.n16771 0.00185
R15097 DVDD.n16896 DVDD.n16894 0.00185
R15098 DVDD.n16207 DVDD.n16206 0.00185
R15099 DVDD.n15572 DVDD.n15571 0.00185
R15100 DVDD.n16650 DVDD.n16648 0.00185
R15101 DVDD.n16593 DVDD.n16591 0.00185
R15102 DVDD.n15786 DVDD.n15785 0.00185
R15103 DVDD.n15849 DVDD.n15848 0.00185
R15104 DVDD.n3597 DVDD.n3596 0.00185
R15105 DVDD.n18647 DVDD.n18646 0.00185
R15106 DVDD.n18694 DVDD.n18693 0.00185
R15107 DVDD.n18436 DVDD.n18435 0.00185
R15108 DVDD.n18351 DVDD.n18350 0.00185
R15109 DVDD.n14764 DVDD.n14763 0.00185
R15110 DVDD.n3295 DVDD.n3294 0.00185
R15111 DVDD.n3306 DVDD.n3305 0.00185
R15112 DVDD.n18661 DVDD.n18660 0.00185
R15113 DVDD.n16063 DVDD.n16062 0.00184712
R15114 DVDD.n16064 DVDD.n16063 0.00184712
R15115 DVDD.n15675 DVDD.n15674 0.00184712
R15116 DVDD.n15676 DVDD.n15675 0.00184712
R15117 DVDD.n9402 DVDD.n9401 0.00184712
R15118 DVDD.n8346 DVDD.n8345 0.00184712
R15119 DVDD.n8347 DVDD.n8346 0.00184712
R15120 DVDD.n9403 DVDD.n9402 0.00184712
R15121 DVDD.n9479 DVDD.n9478 0.00184712
R15122 DVDD.n9480 DVDD.n9479 0.00184712
R15123 DVDD.n7949 DVDD.n7948 0.00184712
R15124 DVDD DVDD.n15623 0.00184667
R15125 DVDD.n14107 DVDD.n14106 0.00183761
R15126 DVDD.n14108 DVDD.n14107 0.00183761
R15127 DVDD.n14017 DVDD.n14016 0.00183761
R15128 DVDD.n14018 DVDD.n14017 0.00183761
R15129 DVDD.n14230 DVDD.n14229 0.00183761
R15130 DVDD.n14229 DVDD.n14228 0.00183761
R15131 DVDD DVDD.n15135 0.00182337
R15132 DVDD.n15992 DVDD.n15991 0.00181799
R15133 DVDD.n15942 DVDD.n15941 0.00181799
R15134 DVDD.n15682 DVDD.n15681 0.00181799
R15135 DVDD.n8194 DVDD.n8193 0.00181799
R15136 DVDD.n9420 DVDD.n9419 0.00181799
R15137 DVDD.n8359 DVDD.n8358 0.00181799
R15138 DVDD.n8310 DVDD.n8309 0.00181799
R15139 DVDD.n8306 DVDD.n8305 0.00181799
R15140 DVDD.n8101 DVDD.n8100 0.00181799
R15141 DVDD.n9900 DVDD.n9899 0.00181799
R15142 DVDD.n7944 DVDD.n7943 0.00181799
R15143 DVDD.n7952 DVDD.n7951 0.00181799
R15144 DVDD.n7960 DVDD.n7959 0.00181799
R15145 DVDD.n7967 DVDD.n7966 0.00181799
R15146 DVDD.n7976 DVDD.n7975 0.00181799
R15147 DVDD.n7985 DVDD.n7984 0.00181799
R15148 DVDD.n7994 DVDD.n7993 0.00181799
R15149 DVDD.n8000 DVDD.n7999 0.00181799
R15150 DVDD.n8008 DVDD.n8007 0.00181799
R15151 DVDD.n8016 DVDD.n8015 0.00181799
R15152 DVDD.n8024 DVDD.n8023 0.00181799
R15153 DVDD.n8031 DVDD.n8030 0.00181799
R15154 DVDD.n8040 DVDD.n8039 0.00181799
R15155 DVDD.n8049 DVDD.n8048 0.00181799
R15156 DVDD.n8058 DVDD.n8057 0.00181799
R15157 DVDD.n8064 DVDD.n8063 0.00181799
R15158 DVDD.n8072 DVDD.n8071 0.00181799
R15159 DVDD.n8080 DVDD.n8079 0.00181799
R15160 DVDD.n8088 DVDD.n8087 0.00181799
R15161 DVDD DVDD.n16381 0.00180667
R15162 DVDD.n12003 DVDD.n12002 0.0017971
R15163 DVDD.n12284 DVDD.n12283 0.0017971
R15164 DVDD.n12207 DVDD.n12206 0.0017971
R15165 DVDD.n13319 DVDD.n13318 0.0017971
R15166 DVDD.n13548 DVDD.n13547 0.0017971
R15167 DVDD.n13629 DVDD.n13628 0.0017971
R15168 DVDD.n1186 DVDD.n1185 0.0017971
R15169 DVDD.n12285 DVDD.n12284 0.0017971
R15170 DVDD.n12002 DVDD.n12001 0.0017971
R15171 DVDD.n13318 DVDD.n13317 0.0017971
R15172 DVDD.n12208 DVDD.n12207 0.0017971
R15173 DVDD.n13547 DVDD.n13546 0.0017971
R15174 DVDD.n13628 DVDD.n13627 0.0017971
R15175 DVDD.n2741 DVDD.n2740 0.0017971
R15176 DVDD.n2782 DVDD.n2781 0.0017971
R15177 DVDD.n15393 DVDD.n15392 0.0017971
R15178 DVDD.n14710 DVDD.n14709 0.0017971
R15179 DVDD.n14627 DVDD.n14626 0.0017971
R15180 DVDD.n14573 DVDD.n14572 0.0017971
R15181 DVDD.n14485 DVDD.n14484 0.0017971
R15182 DVDD.n14486 DVDD.n14485 0.0017971
R15183 DVDD.n14574 DVDD.n14573 0.0017971
R15184 DVDD.n14628 DVDD.n14627 0.0017971
R15185 DVDD.n2740 DVDD.n2739 0.0017971
R15186 DVDD.n15392 DVDD.n15391 0.0017971
R15187 DVDD.n2781 DVDD.n2780 0.0017971
R15188 DVDD.n14711 DVDD.n14710 0.0017971
R15189 DVDD.n19736 DVDD.n19735 0.0017971
R15190 DVDD.n19902 DVDD.n19901 0.0017971
R15191 DVDD.n4801 DVDD.n4800 0.0017971
R15192 DVDD.n4966 DVDD.n4965 0.0017971
R15193 DVDD.n5215 DVDD.n5214 0.0017971
R15194 DVDD.n5454 DVDD.n5453 0.0017971
R15195 DVDD.n6081 DVDD.n6080 0.0017971
R15196 DVDD.n6082 DVDD.n6081 0.0017971
R15197 DVDD.n5453 DVDD.n5452 0.0017971
R15198 DVDD.n5214 DVDD.n5213 0.0017971
R15199 DVDD.n19901 DVDD.n19900 0.0017971
R15200 DVDD.n19735 DVDD.n19734 0.0017971
R15201 DVDD.n4800 DVDD.n4799 0.0017971
R15202 DVDD.n5094 DVDD.n5093 0.0017971
R15203 DVDD.n5460 DVDD.n5459 0.0017971
R15204 DVDD.n1381 DVDD.n1380 0.0017971
R15205 DVDD.n1475 DVDD.n1474 0.0017971
R15206 DVDD.n11627 DVDD.n11626 0.0017971
R15207 DVDD.n12395 DVDD.n12394 0.0017971
R15208 DVDD.n13009 DVDD.n13008 0.0017971
R15209 DVDD.n12713 DVDD.n12712 0.0017971
R15210 DVDD.n13010 DVDD.n13009 0.0017971
R15211 DVDD.n1380 DVDD.n1379 0.0017971
R15212 DVDD.n1476 DVDD.n1475 0.0017971
R15213 DVDD.n11626 DVDD.n11625 0.0017971
R15214 DVDD.n12394 DVDD.n12393 0.0017971
R15215 DVDD.n12714 DVDD.n12713 0.0017971
R15216 DVDD.n779 DVDD.n778 0.0017971
R15217 DVDD.n816 DVDD.n815 0.0017971
R15218 DVDD.n18207 DVDD.n18206 0.0017971
R15219 DVDD.n18063 DVDD.n18062 0.0017971
R15220 DVDD.n17985 DVDD.n17984 0.0017971
R15221 DVDD.n17933 DVDD.n17932 0.0017971
R15222 DVDD.n17852 DVDD.n17851 0.0017971
R15223 DVDD.n17986 DVDD.n17985 0.0017971
R15224 DVDD.n18064 DVDD.n18063 0.0017971
R15225 DVDD.n18208 DVDD.n18207 0.0017971
R15226 DVDD.n815 DVDD.n814 0.0017971
R15227 DVDD.n778 DVDD.n777 0.0017971
R15228 DVDD.n17934 DVDD.n17933 0.0017971
R15229 DVDD.n17853 DVDD.n17852 0.0017971
R15230 DVDD.n1958 DVDD.n1957 0.0017971
R15231 DVDD.n2123 DVDD.n2122 0.0017971
R15232 DVDD.n6883 DVDD.n6882 0.0017971
R15233 DVDD.n6467 DVDD.n6466 0.0017971
R15234 DVDD.n6307 DVDD.n6306 0.0017971
R15235 DVDD.n4531 DVDD.n4530 0.0017971
R15236 DVDD.n6468 DVDD.n6467 0.0017971
R15237 DVDD.n6884 DVDD.n6883 0.0017971
R15238 DVDD.n1957 DVDD.n1956 0.0017971
R15239 DVDD.n2122 DVDD.n2121 0.0017971
R15240 DVDD.n6308 DVDD.n6307 0.0017971
R15241 DVDD.n4532 DVDD.n4531 0.0017971
R15242 DVDD.n3222 DVDD.n3221 0.0017971
R15243 DVDD.n3522 DVDD.n3521 0.0017971
R15244 DVDD.n7883 DVDD.n7882 0.0017971
R15245 DVDD.n8416 DVDD.n8415 0.0017971
R15246 DVDD.n9093 DVDD.n9092 0.0017971
R15247 DVDD.n8798 DVDD.n8797 0.0017971
R15248 DVDD.n3223 DVDD.n3222 0.0017971
R15249 DVDD.n3521 DVDD.n3520 0.0017971
R15250 DVDD.n7882 DVDD.n7881 0.0017971
R15251 DVDD.n8415 DVDD.n8414 0.0017971
R15252 DVDD.n9094 DVDD.n9093 0.0017971
R15253 DVDD.n8799 DVDD.n8798 0.0017971
R15254 DVDD.n19599 DVDD.n19598 0.00179
R15255 DVDD.n19467 DVDD.n19466 0.00179
R15256 DVDD.n20214 DVDD.n20213 0.00179
R15257 DVDD.n20082 DVDD.n20081 0.00179
R15258 DVDD.n253 DVDD.n252 0.00179
R15259 DVDD.n146 DVDD.n145 0.00179
R15260 DVDD.n16999 DVDD.n16998 0.00179
R15261 DVDD.n16941 DVDD.n16940 0.00179
R15262 DVDD.n16774 DVDD.n16773 0.00179
R15263 DVDD.n16897 DVDD.n16896 0.00179
R15264 DVDD.n16651 DVDD.n16650 0.00179
R15265 DVDD.n16594 DVDD.n16593 0.00179
R15266 DVDD.n18564 DVDD.n18563 0.00179
R15267 DVDD.n18662 DVDD.n18661 0.00179
R15268 DVDD.n2478 DVDD.n2477 0.00178571
R15269 DVDD.n8324 DVDD.n8323 0.00178242
R15270 DVDD.n7826 DVDD.n7825 0.00176
R15271 DVDD.n9769 DVDD.n9768 0.00176
R15272 DVDD.n9798 DVDD.n9797 0.00176
R15273 DVDD.n9533 DVDD.n9532 0.00176
R15274 DVDD.n9523 DVDD.n9522 0.00176
R15275 DVDD.n9488 DVDD.n9487 0.00176
R15276 DVDD.n9257 DVDD.n9256 0.00176
R15277 DVDD.n9270 DVDD.n9269 0.00176
R15278 DVDD.n9299 DVDD.n9298 0.00176
R15279 DVDD.n9309 DVDD.n9308 0.00176
R15280 DVDD.n9311 DVDD.n9310 0.00176
R15281 DVDD.n6795 DVDD.n6794 0.00176
R15282 DVDD.n6846 DVDD.n6845 0.00176
R15283 DVDD.n6817 DVDD.n6816 0.00176
R15284 DVDD.n6565 DVDD.n6564 0.00176
R15285 DVDD.n6555 DVDD.n6554 0.00176
R15286 DVDD.n3985 DVDD.n3984 0.00176
R15287 DVDD.n3972 DVDD.n3971 0.00176
R15288 DVDD.n3943 DVDD.n3942 0.00176
R15289 DVDD.n3933 DVDD.n3932 0.00176
R15290 DVDD.n3931 DVDD.n3930 0.00176
R15291 DVDD.n4832 DVDD.n4831 0.00176
R15292 DVDD.n4883 DVDD.n4882 0.00176
R15293 DVDD.n4854 DVDD.n4853 0.00176
R15294 DVDD.n5156 DVDD.n5155 0.00176
R15295 DVDD.n5146 DVDD.n5145 0.00176
R15296 DVDD.n5290 DVDD.n5289 0.00176
R15297 DVDD.n5277 DVDD.n5276 0.00176
R15298 DVDD.n5248 DVDD.n5247 0.00176
R15299 DVDD.n5238 DVDD.n5237 0.00176
R15300 DVDD.n5236 DVDD.n5235 0.00176
R15301 DVDD.n11351 DVDD.n11350 0.00176
R15302 DVDD.n11870 DVDD.n11869 0.00176
R15303 DVDD.n11899 DVDD.n11898 0.00176
R15304 DVDD.n12337 DVDD.n12336 0.00176
R15305 DVDD.n12327 DVDD.n12326 0.00176
R15306 DVDD.n12293 DVDD.n12292 0.00176
R15307 DVDD.n13168 DVDD.n13167 0.00176
R15308 DVDD.n13181 DVDD.n13180 0.00176
R15309 DVDD.n13210 DVDD.n13209 0.00176
R15310 DVDD.n13220 DVDD.n13219 0.00176
R15311 DVDD.n13222 DVDD.n13221 0.00176
R15312 DVDD.n16465 DVDD.n16464 0.00175333
R15313 DVDD.n10837 DVDD.n10836 0.00175333
R15314 DVDD.n10805 DVDD.n10804 0.00175333
R15315 DVDD.n10769 DVDD.n10768 0.00175333
R15316 DVDD.n10317 DVDD.n10316 0.00175333
R15317 DVDD.n15978 DVDD.n15977 0.00175301
R15318 DVDD.n15979 DVDD.n15978 0.00175301
R15319 DVDD.n9435 DVDD.n9434 0.00175301
R15320 DVDD.n9436 DVDD.n9435 0.00175301
R15321 DVDD.n8119 DVDD.n8118 0.00175301
R15322 DVDD.n8118 DVDD.n8117 0.00175301
R15323 DVDD.n15260 DVDD.n15259 0.00174867
R15324 DVDD.n1239 DVDD.n1238 0.00174016
R15325 DVDD.n1222 DVDD.n1221 0.00174016
R15326 DVDD.n1221 DVDD.n1220 0.00174016
R15327 DVDD.n1215 DVDD.n1214 0.00174016
R15328 DVDD.n1200 DVDD.n1199 0.00174016
R15329 DVDD.n1194 DVDD.n1193 0.00174016
R15330 DVDD.n1187 DVDD.n1186 0.00174016
R15331 DVDD.n1179 DVDD.n1178 0.00174016
R15332 DVDD.n1164 DVDD.n1163 0.00174016
R15333 DVDD.n1162 DVDD.n1161 0.00174016
R15334 DVDD.n1659 DVDD.n1658 0.00174016
R15335 DVDD.n1652 DVDD.n1651 0.00174016
R15336 DVDD.n1649 DVDD.n1648 0.00174016
R15337 DVDD.n1782 DVDD.n864 0.00174016
R15338 DVDD.n921 DVDD.n920 0.00174016
R15339 DVDD.n914 DVDD.n913 0.00174016
R15340 DVDD.n908 DVDD.n907 0.00174016
R15341 DVDD.n903 DVDD.n902 0.00174016
R15342 DVDD.n897 DVDD.n896 0.00174016
R15343 DVDD.n890 DVDD.n889 0.00174016
R15344 DVDD.n888 DVDD.n887 0.00174016
R15345 DVDD.n883 DVDD.n882 0.00174016
R15346 DVDD.n876 DVDD.n875 0.00174016
R15347 DVDD.n868 DVDD.n867 0.00174016
R15348 DVDD.n19285 DVDD.n19284 0.00174016
R15349 DVDD.n19288 DVDD.n19287 0.00174016
R15350 DVDD.n10159 DVDD.n10158 0.00174016
R15351 DVDD.n11484 DVDD.n11483 0.00174016
R15352 DVDD.n11997 DVDD.n11996 0.00174016
R15353 DVDD.n12006 DVDD.n12005 0.00174016
R15354 DVDD.n12015 DVDD.n12014 0.00174016
R15355 DVDD.n12022 DVDD.n12021 0.00174016
R15356 DVDD.n12031 DVDD.n12030 0.00174016
R15357 DVDD.n12040 DVDD.n12039 0.00174016
R15358 DVDD.n12048 DVDD.n12047 0.00174016
R15359 DVDD.n12054 DVDD.n12053 0.00174016
R15360 DVDD.n12063 DVDD.n12062 0.00174016
R15361 DVDD.n12072 DVDD.n12071 0.00174016
R15362 DVDD.n12081 DVDD.n12080 0.00174016
R15363 DVDD.n12088 DVDD.n12087 0.00174016
R15364 DVDD.n12097 DVDD.n12096 0.00174016
R15365 DVDD.n12106 DVDD.n12105 0.00174016
R15366 DVDD.n12114 DVDD.n12113 0.00174016
R15367 DVDD.n12120 DVDD.n12119 0.00174016
R15368 DVDD.n12129 DVDD.n12128 0.00174016
R15369 DVDD.n12138 DVDD.n12137 0.00174016
R15370 DVDD.n12147 DVDD.n12146 0.00174016
R15371 DVDD.n12156 DVDD.n12155 0.00174016
R15372 DVDD.n12160 DVDD.n12159 0.00174016
R15373 DVDD.n12225 DVDD.n12224 0.00174016
R15374 DVDD.n13306 DVDD.n13305 0.00174016
R15375 DVDD.n13357 DVDD.n13356 0.00174016
R15376 DVDD.n13362 DVDD.n13361 0.00174016
R15377 DVDD.n13480 DVDD.n13479 0.00174016
R15378 DVDD.n13533 DVDD.n13532 0.00174016
R15379 DVDD.n13614 DVDD.n13613 0.00174016
R15380 DVDD.n13693 DVDD.n13692 0.00174016
R15381 DVDD.n2726 DVDD.n2725 0.00174016
R15382 DVDD.n2767 DVDD.n2766 0.00174016
R15383 DVDD.n2804 DVDD.n2803 0.00174016
R15384 DVDD.n18670 DVDD.n18669 0.00174016
R15385 DVDD.n10063 DVDD.n10062 0.00174016
R15386 DVDD.n14816 DVDD.n14815 0.00174016
R15387 DVDD.n15464 DVDD.n15463 0.00174016
R15388 DVDD.n14725 DVDD.n14724 0.00174016
R15389 DVDD.n14642 DVDD.n14641 0.00174016
R15390 DVDD.n14588 DVDD.n14587 0.00174016
R15391 DVDD.n14500 DVDD.n14499 0.00174016
R15392 DVDD.n14398 DVDD.n14397 0.00174016
R15393 DVDD.n19703 DVDD.n19702 0.00174016
R15394 DVDD.n19738 DVDD.n19737 0.00174016
R15395 DVDD.n19748 DVDD.n19747 0.00174016
R15396 DVDD.n19749 DVDD.n19748 0.00174016
R15397 DVDD.n19871 DVDD.n19870 0.00174016
R15398 DVDD.n19881 DVDD.n19880 0.00174016
R15399 DVDD.n19922 DVDD.n19921 0.00174016
R15400 DVDD.n20001 DVDD.n20000 0.00174016
R15401 DVDD.n20004 DVDD.n20003 0.00174016
R15402 DVDD.n20056 DVDD.n20055 0.00174016
R15403 DVDD.n20058 DVDD.n20057 0.00174016
R15404 DVDD.n20198 DVDD.n20197 0.00174016
R15405 DVDD.n20086 DVDD.n20085 0.00174016
R15406 DVDD.n20099 DVDD.n20098 0.00174016
R15407 DVDD.n19061 DVDD.n19060 0.00174016
R15408 DVDD.n3864 DVDD.n3863 0.00174016
R15409 DVDD.n4780 DVDD.n4779 0.00174016
R15410 DVDD.n4792 DVDD.n4791 0.00174016
R15411 DVDD.n4820 DVDD.n4819 0.00174016
R15412 DVDD.n4943 DVDD.n4942 0.00174016
R15413 DVDD.n5015 DVDD.n5014 0.00174016
R15414 DVDD.n5018 DVDD.n5017 0.00174016
R15415 DVDD.n5033 DVDD.n5032 0.00174016
R15416 DVDD.n5035 DVDD.n5034 0.00174016
R15417 DVDD.n5168 DVDD.n5167 0.00174016
R15418 DVDD.n5196 DVDD.n5195 0.00174016
R15419 DVDD.n5380 DVDD.n5379 0.00174016
R15420 DVDD.n5419 DVDD.n5418 0.00174016
R15421 DVDD.n5547 DVDD.n5546 0.00174016
R15422 DVDD.n5698 DVDD.n5697 0.00174016
R15423 DVDD.n5958 DVDD.n5957 0.00174016
R15424 DVDD.n1348 DVDD.n1347 0.00174016
R15425 DVDD.n1383 DVDD.n1382 0.00174016
R15426 DVDD.n1393 DVDD.n1392 0.00174016
R15427 DVDD.n1394 DVDD.n1393 0.00174016
R15428 DVDD.n1505 DVDD.n1504 0.00174016
R15429 DVDD.n1496 DVDD.n1495 0.00174016
R15430 DVDD.n1455 DVDD.n1454 0.00174016
R15431 DVDD.n1689 DVDD.n1688 0.00174016
R15432 DVDD.n1692 DVDD.n1691 0.00174016
R15433 DVDD.n1717 DVDD.n1716 0.00174016
R15434 DVDD.n1715 DVDD.n1714 0.00174016
R15435 DVDD.n276 DVDD.n275 0.00174016
R15436 DVDD.n19184 DVDD.n19183 0.00174016
R15437 DVDD.n19197 DVDD.n19196 0.00174016
R15438 DVDD.n19443 DVDD.n19442 0.00174016
R15439 DVDD.n10111 DVDD.n10110 0.00174016
R15440 DVDD.n11606 DVDD.n11605 0.00174016
R15441 DVDD.n11618 DVDD.n11617 0.00174016
R15442 DVDD.n11810 DVDD.n11809 0.00174016
R15443 DVDD.n11739 DVDD.n11738 0.00174016
R15444 DVDD.n11736 DVDD.n11735 0.00174016
R15445 DVDD.n11721 DVDD.n11720 0.00174016
R15446 DVDD.n11719 DVDD.n11718 0.00174016
R15447 DVDD.n12349 DVDD.n12348 0.00174016
R15448 DVDD.n12376 DVDD.n12375 0.00174016
R15449 DVDD.n13101 DVDD.n13100 0.00174016
R15450 DVDD.n13081 DVDD.n13080 0.00174016
R15451 DVDD.n13043 DVDD.n13042 0.00174016
R15452 DVDD.n12870 DVDD.n12869 0.00174016
R15453 DVDD.n12743 DVDD.n12742 0.00174016
R15454 DVDD.n12621 DVDD.n12620 0.00174016
R15455 DVDD.n764 DVDD.n763 0.00174016
R15456 DVDD.n801 DVDD.n800 0.00174016
R15457 DVDD.n836 DVDD.n835 0.00174016
R15458 DVDD.n149 DVDD.n148 0.00174016
R15459 DVDD.n10095 DVDD.n10094 0.00174016
R15460 DVDD.n18222 DVDD.n18221 0.00174016
R15461 DVDD.n18143 DVDD.n18142 0.00174016
R15462 DVDD.n18078 DVDD.n18077 0.00174016
R15463 DVDD.n18000 DVDD.n17999 0.00174016
R15464 DVDD.n17948 DVDD.n17947 0.00174016
R15465 DVDD.n17867 DVDD.n17866 0.00174016
R15466 DVDD.n17774 DVDD.n17773 0.00174016
R15467 DVDD.n1925 DVDD.n1924 0.00174016
R15468 DVDD.n1960 DVDD.n1959 0.00174016
R15469 DVDD.n1970 DVDD.n1969 0.00174016
R15470 DVDD.n1971 DVDD.n1970 0.00174016
R15471 DVDD.n2093 DVDD.n2092 0.00174016
R15472 DVDD.n2102 DVDD.n2101 0.00174016
R15473 DVDD.n2143 DVDD.n2142 0.00174016
R15474 DVDD.n2222 DVDD.n2221 0.00174016
R15475 DVDD.n2225 DVDD.n2224 0.00174016
R15476 DVDD.n2277 DVDD.n2276 0.00174016
R15477 DVDD.n2279 DVDD.n2278 0.00174016
R15478 DVDD.n19583 DVDD.n19582 0.00174016
R15479 DVDD.n19471 DVDD.n19470 0.00174016
R15480 DVDD.n19484 DVDD.n19483 0.00174016
R15481 DVDD.n18953 DVDD.n18952 0.00174016
R15482 DVDD.n7085 DVDD.n7084 0.00174016
R15483 DVDD.n6904 DVDD.n6903 0.00174016
R15484 DVDD.n6892 DVDD.n6891 0.00174016
R15485 DVDD.n6741 DVDD.n6740 0.00174016
R15486 DVDD.n6669 DVDD.n6668 0.00174016
R15487 DVDD.n6666 DVDD.n6665 0.00174016
R15488 DVDD.n6651 DVDD.n6650 0.00174016
R15489 DVDD.n6649 DVDD.n6648 0.00174016
R15490 DVDD.n6514 DVDD.n6513 0.00174016
R15491 DVDD.n6486 DVDD.n6485 0.00174016
R15492 DVDD.n6402 DVDD.n6401 0.00174016
R15493 DVDD.n6381 DVDD.n6380 0.00174016
R15494 DVDD.n6342 DVDD.n6341 0.00174016
R15495 DVDD.n6249 DVDD.n6248 0.00174016
R15496 DVDD.n6125 DVDD.n6124 0.00174016
R15497 DVDD.n4419 DVDD.n4418 0.00174016
R15498 DVDD.n3255 DVDD.n3254 0.00174016
R15499 DVDD.n3220 DVDD.n3219 0.00174016
R15500 DVDD.n3210 DVDD.n3209 0.00174016
R15501 DVDD.n3209 DVDD.n3208 0.00174016
R15502 DVDD.n3492 DVDD.n3491 0.00174016
R15503 DVDD.n3501 DVDD.n3500 0.00174016
R15504 DVDD.n3542 DVDD.n3541 0.00174016
R15505 DVDD.n3560 DVDD.n3559 0.00174016
R15506 DVDD.n3557 DVDD.n3556 0.00174016
R15507 DVDD.n3721 DVDD.n3720 0.00174016
R15508 DVDD.n3723 DVDD.n3722 0.00174016
R15509 DVDD.n3762 DVDD.n3761 0.00174016
R15510 DVDD.n18488 DVDD.n18487 0.00174016
R15511 DVDD.n18501 DVDD.n18500 0.00174016
R15512 DVDD.n18790 DVDD.n18789 0.00174016
R15513 DVDD.n7143 DVDD.n7142 0.00174016
R15514 DVDD.n7862 DVDD.n7861 0.00174016
R15515 DVDD.n7874 DVDD.n7873 0.00174016
R15516 DVDD.n9709 DVDD.n9708 0.00174016
R15517 DVDD.n9637 DVDD.n9636 0.00174016
R15518 DVDD.n9634 DVDD.n9633 0.00174016
R15519 DVDD.n9619 DVDD.n9618 0.00174016
R15520 DVDD.n9617 DVDD.n9616 0.00174016
R15521 DVDD.n8369 DVDD.n8368 0.00174016
R15522 DVDD.n8397 DVDD.n8396 0.00174016
R15523 DVDD.n9188 DVDD.n9187 0.00174016
R15524 DVDD.n9167 DVDD.n9166 0.00174016
R15525 DVDD.n9128 DVDD.n9127 0.00174016
R15526 DVDD.n8951 DVDD.n8950 0.00174016
R15527 DVDD.n8827 DVDD.n8826 0.00174016
R15528 DVDD.n8693 DVDD.n8692 0.00174016
R15529 DVDD.n7076 DVDD.n7075 0.00173
R15530 DVDD.n4603 DVDD.n4602 0.00173
R15531 DVDD.n382 DVDD.n381 0.00172143
R15532 DVDD.n388 DVDD.n387 0.00172143
R15533 DVDD.n392 DVDD.n391 0.00172143
R15534 DVDD.n2480 DVDD.n2479 0.00172143
R15535 DVDD.n613 DVDD.n612 0.00172143
R15536 DVDD.n619 DVDD.n618 0.00172143
R15537 DVDD.n623 DVDD.n622 0.00172143
R15538 DVDD.n2676 DVDD.n2675 0.00172143
R15539 DVDD.n2685 DVDD.n2684 0.00172143
R15540 DVDD.n9904 DVDD.n9903 0.00171622
R15541 DVDD.n5670 DVDD.n5669 0.0017086
R15542 DVDD.n12777 DVDD.n12776 0.0017086
R15543 DVDD.n6154 DVDD.n6153 0.0017086
R15544 DVDD.n8856 DVDD.n8855 0.0017086
R15545 DVDD.n12178 DVDD.n12177 0.00170855
R15546 DVDD.n12240 DVDD.n12239 0.00170855
R15547 DVDD.n13705 DVDD.n13704 0.00170855
R15548 DVDD.n12177 DVDD.n12176 0.00170855
R15549 DVDD.n12241 DVDD.n12240 0.00170855
R15550 DVDD.n15478 DVDD.n15477 0.00170855
R15551 DVDD.n14738 DVDD.n14737 0.00170855
R15552 DVDD.n14655 DVDD.n14654 0.00170855
R15553 DVDD.n14384 DVDD.n14383 0.00170855
R15554 DVDD.n14656 DVDD.n14655 0.00170855
R15555 DVDD.n14739 DVDD.n14738 0.00170855
R15556 DVDD.n15477 DVDD.n15476 0.00170855
R15557 DVDD.n5038 DVDD.n5037 0.00170855
R15558 DVDD.n5176 DVDD.n5175 0.00170855
R15559 DVDD.n5400 DVDD.n5399 0.00170855
R15560 DVDD.n5676 DVDD.n5675 0.00170855
R15561 DVDD.n5946 DVDD.n5945 0.00170855
R15562 DVDD.n5675 DVDD.n5674 0.00170855
R15563 DVDD.n5399 DVDD.n5398 0.00170855
R15564 DVDD.n5175 DVDD.n5174 0.00170855
R15565 DVDD.n5037 DVDD.n5036 0.00170855
R15566 DVDD.n5023 DVDD.n5022 0.00170855
R15567 DVDD.n19894 DVDD.n19893 0.00170855
R15568 DVDD.n19886 DVDD.n19885 0.00170855
R15569 DVDD.n11716 DVDD.n11715 0.00170855
R15570 DVDD.n12765 DVDD.n12764 0.00170855
R15571 DVDD.n12609 DVDD.n12608 0.00170855
R15572 DVDD.n13062 DVDD.n13061 0.00170855
R15573 DVDD.n12356 DVDD.n12355 0.00170855
R15574 DVDD.n11717 DVDD.n11716 0.00170855
R15575 DVDD.n1483 DVDD.n1482 0.00170855
R15576 DVDD.n12766 DVDD.n12765 0.00170855
R15577 DVDD.n18131 DVDD.n18130 0.00170855
R15578 DVDD.n18089 DVDD.n18088 0.00170855
R15579 DVDD.n18011 DVDD.n18010 0.00170855
R15580 DVDD.n17762 DVDD.n17761 0.00170855
R15581 DVDD.n18012 DVDD.n18011 0.00170855
R15582 DVDD.n18090 DVDD.n18089 0.00170855
R15583 DVDD.n18132 DVDD.n18131 0.00170855
R15584 DVDD.n6646 DVDD.n6645 0.00170855
R15585 DVDD.n6506 DVDD.n6505 0.00170855
R15586 DVDD.n6361 DVDD.n6360 0.00170855
R15587 DVDD.n4405 DVDD.n4404 0.00170855
R15588 DVDD.n6362 DVDD.n6361 0.00170855
R15589 DVDD.n6647 DVDD.n6646 0.00170855
R15590 DVDD.n2115 DVDD.n2114 0.00170855
R15591 DVDD.n6507 DVDD.n6506 0.00170855
R15592 DVDD.n6149 DVDD.n6148 0.00170855
R15593 DVDD.n14385 DVDD.n14384 0.00170855
R15594 DVDD.n4406 DVDD.n4405 0.00170855
R15595 DVDD.n5947 DVDD.n5946 0.00170855
R15596 DVDD.n12610 DVDD.n12609 0.00170855
R15597 DVDD.n17763 DVDD.n17762 0.00170855
R15598 DVDD.n13704 DVDD.n13703 0.00170855
R15599 DVDD.n9614 DVDD.n9613 0.00170855
R15600 DVDD.n8377 DVDD.n8376 0.00170855
R15601 DVDD.n9147 DVDD.n9146 0.00170855
R15602 DVDD.n8679 DVDD.n8678 0.00170855
R15603 DVDD.n8376 DVDD.n8375 0.00170855
R15604 DVDD.n9148 DVDD.n9147 0.00170855
R15605 DVDD.n8851 DVDD.n8850 0.00170855
R15606 DVDD.n9615 DVDD.n9614 0.00170855
R15607 DVDD.n3514 DVDD.n3513 0.00170855
R15608 DVDD.n8680 DVDD.n8679 0.00170855
R15609 DVDD.n3112 DVDD.n3111 0.00170536
R15610 DVDD.n3102 DVDD.n3101 0.00170536
R15611 DVDD.n3089 DVDD.n3088 0.00170536
R15612 DVDD.n3081 DVDD.n3080 0.00170536
R15613 DVDD.n3075 DVDD.n3074 0.00170536
R15614 DVDD.n3069 DVDD.n3068 0.00170536
R15615 DVDD.n3068 DVDD.n3067 0.00170536
R15616 DVDD.n3051 DVDD.n3050 0.00170536
R15617 DVDD.n3050 DVDD.n3049 0.00170536
R15618 DVDD.n3041 DVDD.n3040 0.00170536
R15619 DVDD.n10317 DVDD.n10205 0.0017
R15620 DVDD.n10281 DVDD.n10280 0.0017
R15621 DVDD.n10485 DVDD.n10484 0.0017
R15622 DVDD.n10452 DVDD.n10451 0.0017
R15623 DVDD.n17087 DVDD.n17079 0.0017
R15624 DVDD.n16967 DVDD.n16966 0.0017
R15625 DVDD.n16623 DVDD.n16620 0.0017
R15626 DVDD.n16622 DVDD.n16621 0.0017
R15627 DVDD.n16971 DVDD.n16970 0.0017
R15628 DVDD.n17086 DVDD.n17085 0.0017
R15629 DVDD.n3365 DVDD.n3364 0.0016749
R15630 DVDD.n7707 DVDD.n7706 0.00167
R15631 DVDD.n7708 DVDD.n7707 0.00167
R15632 DVDD.n3700 DVDD.n3699 0.00167
R15633 DVDD.n3699 DVDD.n3698 0.00167
R15634 DVDD.n18545 DVDD.n18544 0.00167
R15635 DVDD.n18546 DVDD.n18545 0.00167
R15636 DVDD.n2961 DVDD.n2960 0.00167
R15637 DVDD.n2962 DVDD.n2961 0.00167
R15638 DVDD.n2199 DVDD.n2198 0.00167
R15639 DVDD.n2200 DVDD.n2199 0.00167
R15640 DVDD.n2256 DVDD.n2255 0.00167
R15641 DVDD.n2255 DVDD.n2254 0.00167
R15642 DVDD.n18914 DVDD.n18913 0.00167
R15643 DVDD.n18915 DVDD.n18914 0.00167
R15644 DVDD.n7062 DVDD.n7061 0.00167
R15645 DVDD.n7061 DVDD.n7060 0.00167
R15646 DVDD.n1895 DVDD.n1894 0.00167
R15647 DVDD.n1894 DVDD.n1893 0.00167
R15648 DVDD.n19978 DVDD.n19977 0.00167
R15649 DVDD.n19979 DVDD.n19978 0.00167
R15650 DVDD.n20035 DVDD.n20034 0.00167
R15651 DVDD.n20034 DVDD.n20033 0.00167
R15652 DVDD.n19032 DVDD.n19031 0.00167
R15653 DVDD.n19033 DVDD.n19032 0.00167
R15654 DVDD.n4642 DVDD.n4641 0.00167
R15655 DVDD.n4641 DVDD.n4640 0.00167
R15656 DVDD.n19673 DVDD.n19672 0.00167
R15657 DVDD.n19672 DVDD.n19671 0.00167
R15658 DVDD.n967 DVDD.n966 0.00167
R15659 DVDD.n966 DVDD.n965 0.00167
R15660 DVDD.n943 DVDD.n942 0.00167
R15661 DVDD.n942 DVDD.n941 0.00167
R15662 DVDD.n19241 DVDD.n19240 0.00167
R15663 DVDD.n19242 DVDD.n19241 0.00167
R15664 DVDD.n18318 DVDD.n18317 0.00167
R15665 DVDD.n18317 DVDD.n18316 0.00167
R15666 DVDD.n1318 DVDD.n1317 0.00167
R15667 DVDD.n1317 DVDD.n1316 0.00167
R15668 DVDD.n3285 DVDD.n3284 0.00167
R15669 DVDD.n3286 DVDD.n3285 0.00167
R15670 DVDD.n8189 DVDD.n8188 0.0016589
R15671 DVDD.n8190 DVDD.n8189 0.0016589
R15672 DVDD.n8140 DVDD.n8139 0.0016589
R15673 DVDD.n9477 DVDD.n9476 0.0016589
R15674 DVDD.n9478 DVDD.n9477 0.0016589
R15675 DVDD.n8139 DVDD.n8138 0.0016589
R15676 DVDD.n4155 DVDD.n4154 0.00165714
R15677 DVDD.n8537 DVDD.n8536 0.00165714
R15678 DVDD.n13869 DVDD.n13868 0.00165714
R15679 DVDD.n13834 DVDD.n13833 0.00165714
R15680 DVDD.n2497 DVDD.n2454 0.00165714
R15681 DVDD.n432 DVDD.n431 0.00165714
R15682 DVDD.n2343 DVDD.n2342 0.00165714
R15683 DVDD.n2394 DVDD.n2393 0.00165714
R15684 DVDD.n2498 DVDD.n2452 0.00165714
R15685 DVDD.n2709 DVDD.n2650 0.00165714
R15686 DVDD.n2697 DVDD.n2696 0.00165714
R15687 DVDD.n664 DVDD.n663 0.00165714
R15688 DVDD.n2541 DVDD.n2540 0.00165714
R15689 DVDD.n2592 DVDD.n2591 0.00165714
R15690 DVDD.n2710 DVDD.n2648 0.00165714
R15691 DVDD.n2667 DVDD.n2666 0.00165714
R15692 DVDD.n2670 DVDD.n2669 0.00165714
R15693 DVDD.n2695 DVDD.n2694 0.00165714
R15694 DVDD.n4156 DVDD.n4149 0.00165714
R15695 DVDD.n8538 DVDD.n8532 0.00165714
R15696 DVDD.n13870 DVDD.n13864 0.00165714
R15697 DVDD.n13835 DVDD.n11220 0.00165714
R15698 DVDD DVDD.n15250 0.00165261
R15699 DVDD.n15257 DVDD.n15256 0.00165261
R15700 DVDD.n15273 DVDD.n15272 0.00165261
R15701 DVDD.n15290 DVDD 0.00165261
R15702 DVDD.n15285 DVDD.n15283 0.00165261
R15703 DVDD.n3837 DVDD.n3836 0.00164716
R15704 DVDD.n122 DVDD.n121 0.00164716
R15705 DVDD.n10186 DVDD.n10185 0.00164
R15706 DVDD.n14744 DVDD.n14743 0.00164
R15707 DVDD.n15964 DVDD.n15963 0.00162971
R15708 DVDD.n8257 DVDD.n8256 0.00162971
R15709 DVDD.n8177 DVDD.n8176 0.00162971
R15710 DVDD.n9454 DVDD.n9453 0.00162971
R15711 DVDD.n8133 DVDD.n8132 0.00162971
R15712 DVDD.n8029 DVDD.n8028 0.00162971
R15713 DVDD DVDD.n15335 0.00162
R15714 DVDD.n12197 DVDD.n12196 0.00161999
R15715 DVDD.n12283 DVDD.n12282 0.00161999
R15716 DVDD.n13484 DVDD.n13483 0.00161999
R15717 DVDD.n12282 DVDD.n12281 0.00161999
R15718 DVDD.n12198 DVDD.n12197 0.00161999
R15719 DVDD.n13485 DVDD.n13484 0.00161999
R15720 DVDD.n6092 DVDD.n6091 0.00161999
R15721 DVDD.n6093 DVDD.n6092 0.00161999
R15722 DVDD.n5359 DVDD.n5358 0.00161999
R15723 DVDD.n4977 DVDD.n4976 0.00161999
R15724 DVDD.n5448 DVDD.n5447 0.00161999
R15725 DVDD.n5681 DVDD.n5680 0.00161999
R15726 DVDD.n5635 DVDD.n5634 0.00161999
R15727 DVDD.n5587 DVDD.n5586 0.00161999
R15728 DVDD.n1397 DVDD.n1396 0.00161999
R15729 DVDD.n12724 DVDD.n12723 0.00161999
R15730 DVDD.n11646 DVDD.n11645 0.00161999
R15731 DVDD.n11776 DVDD.n11775 0.00161999
R15732 DVDD.n13015 DVDD.n13014 0.00161999
R15733 DVDD.n12725 DVDD.n12724 0.00161999
R15734 DVDD.n12760 DVDD.n12759 0.00161999
R15735 DVDD.n12802 DVDD.n12801 0.00161999
R15736 DVDD.n12840 DVDD.n12839 0.00161999
R15737 DVDD.n1974 DVDD.n1973 0.00161999
R15738 DVDD.n6864 DVDD.n6863 0.00161999
R15739 DVDD.n6707 DVDD.n6706 0.00161999
R15740 DVDD.n4542 DVDD.n4541 0.00161999
R15741 DVDD.n6313 DVDD.n6312 0.00161999
R15742 DVDD.n4543 DVDD.n4542 0.00161999
R15743 DVDD.n6144 DVDD.n6143 0.00161999
R15744 DVDD.n6182 DVDD.n6181 0.00161999
R15745 DVDD.n6220 DVDD.n6219 0.00161999
R15746 DVDD.n8809 DVDD.n8808 0.00161999
R15747 DVDD.n8810 DVDD.n8809 0.00161999
R15748 DVDD.n7902 DVDD.n7901 0.00161999
R15749 DVDD.n9675 DVDD.n9674 0.00161999
R15750 DVDD.n3206 DVDD.n3205 0.00161999
R15751 DVDD.n9099 DVDD.n9098 0.00161999
R15752 DVDD.n8846 DVDD.n8845 0.00161999
R15753 DVDD.n8884 DVDD.n8883 0.00161999
R15754 DVDD.n8922 DVDD.n8921 0.00161999
R15755 DVDD DVDD.n15903 0.00160667
R15756 DVDD.n3046 DVDD.n3045 0.0016026
R15757 DVDD.n3045 DVDD.n3044 0.0016026
R15758 DVDD.n2344 DVDD.n2343 0.00159286
R15759 DVDD.n2455 DVDD.n2452 0.00159286
R15760 DVDD.n2542 DVDD.n2541 0.00159286
R15761 DVDD.n2653 DVDD.n2648 0.00159286
R15762 DVDD.n2694 DVDD.n2693 0.00159286
R15763 DVDD.n4149 DVDD.n4148 0.00159286
R15764 DVDD.n8532 DVDD.n8531 0.00159286
R15765 DVDD.n13864 DVDD.n13863 0.00159286
R15766 DVDD.n11222 DVDD.n11220 0.00159286
R15767 DVDD.n7827 DVDD.n7826 0.00158
R15768 DVDD.n9768 DVDD.n9767 0.00158
R15769 DVDD.n9799 DVDD.n9798 0.00158
R15770 DVDD.n9534 DVDD.n9533 0.00158
R15771 DVDD.n9524 DVDD.n9523 0.00158
R15772 DVDD.n9522 DVDD.n9521 0.00158
R15773 DVDD.n9487 DVDD.n9486 0.00158
R15774 DVDD.n9258 DVDD.n9257 0.00158
R15775 DVDD.n9269 DVDD.n9268 0.00158
R15776 DVDD.n9300 DVDD.n9299 0.00158
R15777 DVDD.n9310 DVDD.n9309 0.00158
R15778 DVDD.n6796 DVDD.n6795 0.00158
R15779 DVDD.n6847 DVDD.n6846 0.00158
R15780 DVDD.n6816 DVDD.n6815 0.00158
R15781 DVDD.n6566 DVDD.n6565 0.00158
R15782 DVDD.n6556 DVDD.n6555 0.00158
R15783 DVDD.n6554 DVDD.n6553 0.00158
R15784 DVDD.n3984 DVDD.n3983 0.00158
R15785 DVDD.n3973 DVDD.n3972 0.00158
R15786 DVDD.n3942 DVDD.n3941 0.00158
R15787 DVDD.n3932 DVDD.n3931 0.00158
R15788 DVDD.n4833 DVDD.n4832 0.00158
R15789 DVDD.n4884 DVDD.n4883 0.00158
R15790 DVDD.n4853 DVDD.n4852 0.00158
R15791 DVDD.n5157 DVDD.n5156 0.00158
R15792 DVDD.n5147 DVDD.n5146 0.00158
R15793 DVDD.n5145 DVDD.n5144 0.00158
R15794 DVDD.n5289 DVDD.n5288 0.00158
R15795 DVDD.n5278 DVDD.n5277 0.00158
R15796 DVDD.n5247 DVDD.n5246 0.00158
R15797 DVDD.n5237 DVDD.n5236 0.00158
R15798 DVDD.n252 DVDD.n251 0.00158
R15799 DVDD.n11352 DVDD.n11351 0.00158
R15800 DVDD.n11869 DVDD.n11868 0.00158
R15801 DVDD.n11900 DVDD.n11899 0.00158
R15802 DVDD.n12338 DVDD.n12337 0.00158
R15803 DVDD.n12328 DVDD.n12327 0.00158
R15804 DVDD.n12326 DVDD.n12325 0.00158
R15805 DVDD.n12292 DVDD.n12291 0.00158
R15806 DVDD.n13169 DVDD.n13168 0.00158
R15807 DVDD.n13180 DVDD.n13179 0.00158
R15808 DVDD.n13211 DVDD.n13210 0.00158
R15809 DVDD.n13221 DVDD.n13220 0.00158
R15810 DVDD.n18565 DVDD.n18564 0.00158
R15811 DVDD.n15241 DVDD.n15240 0.00156875
R15812 DVDD.n15247 DVDD.n15246 0.00156875
R15813 DVDD.n10566 DVDD.n10565 0.00156875
R15814 DVDD.n10572 DVDD.n10571 0.00156875
R15815 DVDD.n10576 DVDD.n10575 0.00156875
R15816 DVDD.n8253 DVDD.n8252 0.00156478
R15817 DVDD.n8252 DVDD.n8251 0.00156478
R15818 DVDD.n9889 DVDD.n9888 0.00156478
R15819 DVDD.n7941 DVDD.n7940 0.00156478
R15820 DVDD.n7972 DVDD.n7971 0.00156478
R15821 DVDD.n7981 DVDD.n7980 0.00156478
R15822 DVDD.n7997 DVDD.n7996 0.00156478
R15823 DVDD.n8027 DVDD.n8026 0.00156478
R15824 DVDD.n8036 DVDD.n8035 0.00156478
R15825 DVDD.n8045 DVDD.n8044 0.00156478
R15826 DVDD.n8061 DVDD.n8060 0.00156478
R15827 DVDD.n8093 DVDD.n8092 0.00156478
R15828 DVDD.n9890 DVDD.n9889 0.00156478
R15829 DVDD.n7940 DVDD.n7939 0.00156478
R15830 DVDD.n7947 DVDD.n7946 0.00156478
R15831 DVDD.n7955 DVDD.n7954 0.00156478
R15832 DVDD.n7971 DVDD.n7970 0.00156478
R15833 DVDD.n7980 DVDD.n7979 0.00156478
R15834 DVDD.n7996 DVDD.n7995 0.00156478
R15835 DVDD.n8003 DVDD.n8002 0.00156478
R15836 DVDD.n8011 DVDD.n8010 0.00156478
R15837 DVDD.n8019 DVDD.n8018 0.00156478
R15838 DVDD.n8026 DVDD.n8025 0.00156478
R15839 DVDD.n8035 DVDD.n8034 0.00156478
R15840 DVDD.n8044 DVDD.n8043 0.00156478
R15841 DVDD.n8060 DVDD.n8059 0.00156478
R15842 DVDD.n8067 DVDD.n8066 0.00156478
R15843 DVDD.n8075 DVDD.n8074 0.00156478
R15844 DVDD.n8083 DVDD.n8082 0.00156478
R15845 DVDD.n8092 DVDD.n8091 0.00156478
R15846 DVDD.n1233 DVDD.n1232 0.00156299
R15847 DVDD.n1223 DVDD.n1222 0.00156299
R15848 DVDD.n1210 DVDD.n1209 0.00156299
R15849 DVDD.n1201 DVDD.n1200 0.00156299
R15850 DVDD.n1195 DVDD.n1194 0.00156299
R15851 DVDD.n1189 DVDD.n1188 0.00156299
R15852 DVDD.n1188 DVDD.n1187 0.00156299
R15853 DVDD.n1173 DVDD.n1172 0.00156299
R15854 DVDD.n1172 DVDD.n1171 0.00156299
R15855 DVDD.n1163 DVDD.n1162 0.00156299
R15856 DVDD.n1600 DVDD.n1599 0.00156299
R15857 DVDD.n1657 DVDD.n1656 0.00156299
R15858 DVDD.n880 DVDD.n879 0.00156299
R15859 DVDD.n19336 DVDD.n19335 0.00156299
R15860 DVDD.n10174 DVDD.n10173 0.00156299
R15861 DVDD.n10179 DVDD.n10178 0.00156299
R15862 DVDD.n18266 DVDD.n10183 0.00156299
R15863 DVDD.n11432 DVDD.n11431 0.00156299
R15864 DVDD.n11439 DVDD.n11438 0.00156299
R15865 DVDD.n11447 DVDD.n11446 0.00156299
R15866 DVDD.n12086 DVDD.n12085 0.00156299
R15867 DVDD.n12192 DVDD.n12191 0.00156299
R15868 DVDD.n12259 DVDD.n12258 0.00156299
R15869 DVDD.n13414 DVDD.n13413 0.00156299
R15870 DVDD.n13497 DVDD.n13496 0.00156299
R15871 DVDD.n13718 DVDD.n13717 0.00156299
R15872 DVDD.n18477 DVDD.n18476 0.00156299
R15873 DVDD.n15492 DVDD.n15491 0.00156299
R15874 DVDD.n15507 DVDD.n15506 0.00156299
R15875 DVDD.n14670 DVDD.n14669 0.00156299
R15876 DVDD.n14370 DVDD.n14369 0.00156299
R15877 DVDD.n19702 DVDD.n19701 0.00156299
R15878 DVDD.n19862 DVDD.n19861 0.00156299
R15879 DVDD.n19865 DVDD.n19864 0.00156299
R15880 DVDD.n19923 DVDD.n19922 0.00156299
R15881 DVDD.n19926 DVDD.n19925 0.00156299
R15882 DVDD.n20055 DVDD.n20054 0.00156299
R15883 DVDD.n20103 DVDD.n20102 0.00156299
R15884 DVDD.n20109 DVDD.n20108 0.00156299
R15885 DVDD.n19081 DVDD.n19080 0.00156299
R15886 DVDD.n19063 DVDD.n19062 0.00156299
R15887 DVDD.n4666 DVDD.n4665 0.00156299
R15888 DVDD.n4681 DVDD.n4680 0.00156299
R15889 DVDD.n4816 DVDD.n4815 0.00156299
R15890 DVDD.n4905 DVDD.n4904 0.00156299
R15891 DVDD.n4931 DVDD.n4930 0.00156299
R15892 DVDD.n4990 DVDD.n4989 0.00156299
R15893 DVDD.n5052 DVDD.n5051 0.00156299
R15894 DVDD.n5060 DVDD.n5059 0.00156299
R15895 DVDD.n5088 DVDD.n5087 0.00156299
R15896 DVDD.n5167 DVDD.n5166 0.00156299
R15897 DVDD.n5356 DVDD.n5355 0.00156299
R15898 DVDD.n5366 DVDD.n5365 0.00156299
R15899 DVDD.n5369 DVDD.n5368 0.00156299
R15900 DVDD.n5420 DVDD.n5419 0.00156299
R15901 DVDD.n5445 DVDD.n5444 0.00156299
R15902 DVDD.n5584 DVDD.n5583 0.00156299
R15903 DVDD.n6069 DVDD.n6054 0.00156299
R15904 DVDD.n6054 DVDD.n6053 0.00156299
R15905 DVDD.n6051 DVDD.n6050 0.00156299
R15906 DVDD.n5932 DVDD.n5931 0.00156299
R15907 DVDD.n1347 DVDD.n1346 0.00156299
R15908 DVDD.n1364 DVDD.n1363 0.00156299
R15909 DVDD.n1514 DVDD.n1513 0.00156299
R15910 DVDD.n1511 DVDD.n1510 0.00156299
R15911 DVDD.n1454 DVDD.n1453 0.00156299
R15912 DVDD.n1451 DVDD.n1450 0.00156299
R15913 DVDD.n1718 DVDD.n1717 0.00156299
R15914 DVDD.n19201 DVDD.n19200 0.00156299
R15915 DVDD.n19207 DVDD.n19206 0.00156299
R15916 DVDD.n19463 DVDD.n19462 0.00156299
R15917 DVDD.n19445 DVDD.n19444 0.00156299
R15918 DVDD.n11373 DVDD.n11372 0.00156299
R15919 DVDD.n11388 DVDD.n11387 0.00156299
R15920 DVDD.n11642 DVDD.n11641 0.00156299
R15921 DVDD.n11848 DVDD.n11847 0.00156299
R15922 DVDD.n11822 DVDD.n11821 0.00156299
R15923 DVDD.n11763 DVDD.n11762 0.00156299
R15924 DVDD.n11702 DVDD.n11701 0.00156299
R15925 DVDD.n11694 DVDD.n11693 0.00156299
R15926 DVDD.n11666 DVDD.n11665 0.00156299
R15927 DVDD.n12348 DVDD.n12347 0.00156299
R15928 DVDD.n13104 DVDD.n13103 0.00156299
R15929 DVDD.n13094 DVDD.n13093 0.00156299
R15930 DVDD.n13091 DVDD.n13090 0.00156299
R15931 DVDD.n13042 DVDD.n13041 0.00156299
R15932 DVDD.n13018 DVDD.n13017 0.00156299
R15933 DVDD.n12843 DVDD.n12842 0.00156299
R15934 DVDD.n12701 DVDD.n12700 0.00156299
R15935 DVDD.n12700 DVDD.n12699 0.00156299
R15936 DVDD.n12697 DVDD.n12696 0.00156299
R15937 DVDD.n12595 DVDD.n12594 0.00156299
R15938 DVDD.n19173 DVDD.n19172 0.00156299
R15939 DVDD.n18117 DVDD.n18116 0.00156299
R15940 DVDD.n18104 DVDD.n18103 0.00156299
R15941 DVDD.n18026 DVDD.n18025 0.00156299
R15942 DVDD.n17748 DVDD.n17747 0.00156299
R15943 DVDD.n1924 DVDD.n1923 0.00156299
R15944 DVDD.n1941 DVDD.n1940 0.00156299
R15945 DVDD.n2084 DVDD.n2083 0.00156299
R15946 DVDD.n2087 DVDD.n2086 0.00156299
R15947 DVDD.n2144 DVDD.n2143 0.00156299
R15948 DVDD.n2147 DVDD.n2146 0.00156299
R15949 DVDD.n2276 DVDD.n2275 0.00156299
R15950 DVDD.n19488 DVDD.n19487 0.00156299
R15951 DVDD.n19494 DVDD.n19493 0.00156299
R15952 DVDD.n18973 DVDD.n18972 0.00156299
R15953 DVDD.n18955 DVDD.n18954 0.00156299
R15954 DVDD.n7018 DVDD.n7017 0.00156299
R15955 DVDD.n7003 DVDD.n7002 0.00156299
R15956 DVDD.n6868 DVDD.n6867 0.00156299
R15957 DVDD.n6779 DVDD.n6778 0.00156299
R15958 DVDD.n6753 DVDD.n6752 0.00156299
R15959 DVDD.n6694 DVDD.n6693 0.00156299
R15960 DVDD.n6632 DVDD.n6631 0.00156299
R15961 DVDD.n6622 DVDD.n6621 0.00156299
R15962 DVDD.n6594 DVDD.n6593 0.00156299
R15963 DVDD.n6515 DVDD.n6514 0.00156299
R15964 DVDD.n6405 DVDD.n6404 0.00156299
R15965 DVDD.n6395 DVDD.n6394 0.00156299
R15966 DVDD.n6392 DVDD.n6391 0.00156299
R15967 DVDD.n6341 DVDD.n6340 0.00156299
R15968 DVDD.n6316 DVDD.n6315 0.00156299
R15969 DVDD.n6223 DVDD.n6222 0.00156299
R15970 DVDD.n4519 DVDD.n4511 0.00156299
R15971 DVDD.n4511 DVDD.n4510 0.00156299
R15972 DVDD.n4508 DVDD.n4507 0.00156299
R15973 DVDD.n4391 DVDD.n4390 0.00156299
R15974 DVDD.n3256 DVDD.n3255 0.00156299
R15975 DVDD.n3239 DVDD.n3238 0.00156299
R15976 DVDD.n3483 DVDD.n3482 0.00156299
R15977 DVDD.n3486 DVDD.n3485 0.00156299
R15978 DVDD.n3543 DVDD.n3542 0.00156299
R15979 DVDD.n3546 DVDD.n3545 0.00156299
R15980 DVDD.n3720 DVDD.n3719 0.00156299
R15981 DVDD.n18505 DVDD.n18504 0.00156299
R15982 DVDD.n18511 DVDD.n18510 0.00156299
R15983 DVDD.n18810 DVDD.n18809 0.00156299
R15984 DVDD.n18792 DVDD.n18791 0.00156299
R15985 DVDD.n10035 DVDD.n10034 0.00156299
R15986 DVDD.n10020 DVDD.n10019 0.00156299
R15987 DVDD.n7898 DVDD.n7897 0.00156299
R15988 DVDD.n9747 DVDD.n9746 0.00156299
R15989 DVDD.n9721 DVDD.n9720 0.00156299
R15990 DVDD.n9662 DVDD.n9661 0.00156299
R15991 DVDD.n9600 DVDD.n9599 0.00156299
R15992 DVDD.n9590 DVDD.n9589 0.00156299
R15993 DVDD.n9562 DVDD.n9561 0.00156299
R15994 DVDD.n8368 DVDD.n8367 0.00156299
R15995 DVDD.n9191 DVDD.n9190 0.00156299
R15996 DVDD.n9181 DVDD.n9180 0.00156299
R15997 DVDD.n9178 DVDD.n9177 0.00156299
R15998 DVDD.n9127 DVDD.n9126 0.00156299
R15999 DVDD.n9102 DVDD.n9101 0.00156299
R16000 DVDD.n8925 DVDD.n8924 0.00156299
R16001 DVDD.n8786 DVDD.n8785 0.00156299
R16002 DVDD.n8785 DVDD.n8784 0.00156299
R16003 DVDD.n8782 DVDD.n8781 0.00156299
R16004 DVDD.n8665 DVDD.n8664 0.00156299
R16005 DVDD.n15203 DVDD.n15202 0.00155656
R16006 DVDD.n18978 DVDD.n18977 0.00154287
R16007 DVDD.n10545 DVDD.n10544 0.00154287
R16008 DVDD.n1167 DVDD.n1166 0.00153143
R16009 DVDD.n11474 DVDD.n11473 0.00153143
R16010 DVDD.n11994 DVDD.n11993 0.00153143
R16011 DVDD.n12001 DVDD.n12000 0.00153143
R16012 DVDD.n12010 DVDD.n12009 0.00153143
R16013 DVDD.n12027 DVDD.n12026 0.00153143
R16014 DVDD.n12036 DVDD.n12035 0.00153143
R16015 DVDD.n12051 DVDD.n12050 0.00153143
R16016 DVDD.n12058 DVDD.n12057 0.00153143
R16017 DVDD.n12067 DVDD.n12066 0.00153143
R16018 DVDD.n12076 DVDD.n12075 0.00153143
R16019 DVDD.n12084 DVDD.n12083 0.00153143
R16020 DVDD.n12093 DVDD.n12092 0.00153143
R16021 DVDD.n12102 DVDD.n12101 0.00153143
R16022 DVDD.n12117 DVDD.n12116 0.00153143
R16023 DVDD.n12124 DVDD.n12123 0.00153143
R16024 DVDD.n12133 DVDD.n12132 0.00153143
R16025 DVDD.n12142 DVDD.n12141 0.00153143
R16026 DVDD.n12152 DVDD.n12151 0.00153143
R16027 DVDD.n13418 DVDD.n13417 0.00153143
R16028 DVDD.n11473 DVDD.n11339 0.00153143
R16029 DVDD.n12000 DVDD.n11999 0.00153143
R16030 DVDD.n12009 DVDD.n12008 0.00153143
R16031 DVDD.n12026 DVDD.n12025 0.00153143
R16032 DVDD.n12035 DVDD.n12034 0.00153143
R16033 DVDD.n12050 DVDD.n12049 0.00153143
R16034 DVDD.n12057 DVDD.n12056 0.00153143
R16035 DVDD.n12066 DVDD.n12065 0.00153143
R16036 DVDD.n12075 DVDD.n12074 0.00153143
R16037 DVDD.n12083 DVDD.n12082 0.00153143
R16038 DVDD.n12092 DVDD.n12091 0.00153143
R16039 DVDD.n12101 DVDD.n12100 0.00153143
R16040 DVDD.n12116 DVDD.n12115 0.00153143
R16041 DVDD.n12123 DVDD.n12122 0.00153143
R16042 DVDD.n12132 DVDD.n12131 0.00153143
R16043 DVDD.n12141 DVDD.n12140 0.00153143
R16044 DVDD.n12151 DVDD.n12150 0.00153143
R16045 DVDD.n11993 DVDD.n11992 0.00153143
R16046 DVDD.n1168 DVDD.n1167 0.00153143
R16047 DVDD.n13419 DVDD.n13418 0.00153143
R16048 DVDD.n5589 DVDD.n5588 0.00153143
R16049 DVDD.n6098 DVDD.n6097 0.00153143
R16050 DVDD.n6048 DVDD.n6047 0.00153143
R16051 DVDD.n6043 DVDD.n6042 0.00153143
R16052 DVDD.n19719 DVDD.n19718 0.00153143
R16053 DVDD.n6099 DVDD.n6098 0.00153143
R16054 DVDD.n5623 DVDD.n5612 0.00153143
R16055 DVDD.n5588 DVDD.n5587 0.00153143
R16056 DVDD.n5576 DVDD.n5565 0.00153143
R16057 DVDD.n5669 DVDD.n5658 0.00153143
R16058 DVDD.n6044 DVDD.n6043 0.00153143
R16059 DVDD.n6049 DVDD.n6048 0.00153143
R16060 DVDD.n12838 DVDD.n12837 0.00153143
R16061 DVDD.n12730 DVDD.n12729 0.00153143
R16062 DVDD.n12694 DVDD.n12693 0.00153143
R16063 DVDD.n12689 DVDD.n12688 0.00153143
R16064 DVDD.n13045 DVDD.n13044 0.00153143
R16065 DVDD.n12778 DVDD.n12777 0.00153143
R16066 DVDD.n12814 DVDD.n12813 0.00153143
R16067 DVDD.n12839 DVDD.n12838 0.00153143
R16068 DVDD.n12851 DVDD.n12850 0.00153143
R16069 DVDD.n12731 DVDD.n12730 0.00153143
R16070 DVDD.n12695 DVDD.n12694 0.00153143
R16071 DVDD.n12690 DVDD.n12689 0.00153143
R16072 DVDD.n6218 DVDD.n6217 0.00153143
R16073 DVDD.n4548 DVDD.n4547 0.00153143
R16074 DVDD.n4506 DVDD.n4505 0.00153143
R16075 DVDD.n4494 DVDD.n4493 0.00153143
R16076 DVDD.n6344 DVDD.n6343 0.00153143
R16077 DVDD.n6193 DVDD.n6192 0.00153143
R16078 DVDD.n6219 DVDD.n6218 0.00153143
R16079 DVDD.n6231 DVDD.n6230 0.00153143
R16080 DVDD.n6155 DVDD.n6154 0.00153143
R16081 DVDD.n4505 DVDD.n4497 0.00153143
R16082 DVDD.n8920 DVDD.n8919 0.00153143
R16083 DVDD.n8815 DVDD.n8814 0.00153143
R16084 DVDD.n8779 DVDD.n8778 0.00153143
R16085 DVDD.n8775 DVDD.n8774 0.00153143
R16086 DVDD.n8780 DVDD.n8779 0.00153143
R16087 DVDD.n9130 DVDD.n9129 0.00153143
R16088 DVDD.n8895 DVDD.n8894 0.00153143
R16089 DVDD.n8921 DVDD.n8920 0.00153143
R16090 DVDD.n8933 DVDD.n8932 0.00153143
R16091 DVDD.n8857 DVDD.n8856 0.00153143
R16092 DVDD.n376 DVDD.n375 0.00152857
R16093 DVDD.n401 DVDD.n400 0.00152857
R16094 DVDD.n451 DVDD.n450 0.00152857
R16095 DVDD.n2319 DVDD.n2318 0.00152857
R16096 DVDD.n2324 DVDD.n2323 0.00152857
R16097 DVDD.n607 DVDD.n606 0.00152857
R16098 DVDD.n632 DVDD.n631 0.00152857
R16099 DVDD.n683 DVDD.n682 0.00152857
R16100 DVDD.n2519 DVDD.n2518 0.00152857
R16101 DVDD.n2522 DVDD.n2521 0.00152857
R16102 DVDD.n13734 DVDD.n13733 0.00152857
R16103 DVDD.n11285 DVDD.n11284 0.00152857
R16104 DVDD.n12489 DVDD.n12488 0.00152857
R16105 DVDD.n5740 DVDD.n5739 0.00152857
R16106 DVDD.n14927 DVDD.n14926 0.0015125
R16107 DVDD.n14890 DVDD.n14889 0.0015125
R16108 DVDD.n15225 DVDD.n15224 0.0015125
R16109 DVDD.n15234 DVDD.n15233 0.0015125
R16110 DVDD.n15237 DVDD.n15236 0.0015125
R16111 DVDD.n15110 DVDD.n15109 0.0015125
R16112 DVDD.n15303 DVDD.n15302 0.0015125
R16113 DVDD.n15006 DVDD.n15005 0.0015125
R16114 DVDD.n10395 DVDD.n10394 0.0015125
R16115 DVDD.n3111 DVDD.n3110 0.00150446
R16116 DVDD.n3095 DVDD.n3094 0.00150446
R16117 DVDD.n3092 DVDD.n3091 0.00150446
R16118 DVDD.n3107 DVDD.n3106 0.00150218
R16119 DVDD.n3106 DVDD.n3105 0.00150218
R16120 DVDD.n20341 DVDD.n24 0.0015
R16121 DVDD.n7475 DVDD.n7426 0.0015
R16122 DVDD.n20341 DVDD.n106 0.0015
R16123 DVDD.n7475 DVDD.n7474 0.0015
R16124 DVDD.n20341 DVDD.n52 0.0015
R16125 DVDD.n7479 DVDD.n7475 0.0015
R16126 DVDD.n7674 DVDD.n7512 0.0015
R16127 DVDD.n10218 DVDD.n10213 0.0015
R16128 DVDD.n10292 DVDD.n10276 0.0015
R16129 DVDD.n20341 DVDD.n20242 0.0015
R16130 DVDD.n7475 DVDD.n7342 0.0015
R16131 DVDD.n3710 DVDD.n3709 0.00149
R16132 DVDD.n18556 DVDD.n18555 0.00149
R16133 DVDD.n18773 DVDD.n18772 0.00149
R16134 DVDD.n2930 DVDD.n2929 0.00149
R16135 DVDD.n2940 DVDD.n2939 0.00149
R16136 DVDD.n9885 DVDD.n9884 0.00149
R16137 DVDD.n8365 DVDD.n8364 0.00149
R16138 DVDD.n2168 DVDD.n2167 0.00149
R16139 DVDD.n2178 DVDD.n2177 0.00149
R16140 DVDD.n2266 DVDD.n2265 0.00149
R16141 DVDD.n18925 DVDD.n18924 0.00149
R16142 DVDD.n1884 DVDD.n1883 0.00149
R16143 DVDD.n1875 DVDD.n1874 0.00149
R16144 DVDD.n3927 DVDD.n3926 0.00149
R16145 DVDD.n19947 DVDD.n19946 0.00149
R16146 DVDD.n19957 DVDD.n19956 0.00149
R16147 DVDD.n20045 DVDD.n20044 0.00149
R16148 DVDD.n19043 DVDD.n19042 0.00149
R16149 DVDD.n19662 DVDD.n19661 0.00149
R16150 DVDD.n19653 DVDD.n19652 0.00149
R16151 DVDD.n5232 DVDD.n5231 0.00149
R16152 DVDD.n998 DVDD.n997 0.00149
R16153 DVDD.n988 DVDD.n987 0.00149
R16154 DVDD.n953 DVDD.n952 0.00149
R16155 DVDD.n19252 DVDD.n19251 0.00149
R16156 DVDD.n19426 DVDD.n19425 0.00149
R16157 DVDD.n11986 DVDD.n11985 0.00149
R16158 DVDD.n1307 DVDD.n1306 0.00149
R16159 DVDD.n1298 DVDD.n1297 0.00149
R16160 DVDD.n11303 DVDD.n11302 0.00149
R16161 DVDD.n3296 DVDD.n3295 0.00149
R16162 DVDD.n3305 DVDD.n3304 0.00149
R16163 DVDD.n12931 DVDD.n12928 0.00147826
R16164 DVDD.n12950 DVDD.n12947 0.00147826
R16165 DVDD.n5515 DVDD.n5512 0.00147826
R16166 DVDD.n5541 DVDD.n5538 0.00147826
R16167 DVDD.n4013 DVDD.n4010 0.00147826
R16168 DVDD.n4036 DVDD.n4033 0.00147826
R16169 DVDD.n8969 DVDD.n8966 0.00147826
R16170 DVDD.n9038 DVDD.n9035 0.00147826
R16171 DVDD.n12904 DVDD.n12903 0.00147826
R16172 DVDD.n12891 DVDD.n12888 0.00147826
R16173 DVDD.n5723 DVDD.n5716 0.00147826
R16174 DVDD.n6061 DVDD.n6058 0.00147826
R16175 DVDD.n4094 DVDD.n4087 0.00147826
R16176 DVDD.n4504 DVDD.n4501 0.00147826
R16177 DVDD.n8996 DVDD.n8993 0.00147826
R16178 DVDD.n9011 DVDD.n9010 0.00147826
R16179 DVDD.n7812 DVDD.n7811 0.00147297
R16180 DVDD.n7979 DVDD.n7978 0.00147066
R16181 DVDD.n8051 DVDD.n8050 0.00147066
R16182 DVDD.n7978 DVDD.n7977 0.00147066
R16183 DVDD.n8052 DVDD.n8051 0.00147066
R16184 DVDD.n11266 DVDD.n11265 0.00146429
R16185 DVDD.n11254 DVDD.n11253 0.00146429
R16186 DVDD.n11238 DVDD.n11237 0.00146429
R16187 DVDD.n5743 DVDD.n5741 0.00146429
R16188 DVDD.n304 DVDD.n303 0.00146429
R16189 DVDD.n404 DVDD.n402 0.00146429
R16190 DVDD.n494 DVDD.n491 0.00146429
R16191 DVDD.n448 DVDD.n445 0.00146429
R16192 DVDD.n377 DVDD.n376 0.00146429
R16193 DVDD.n405 DVDD.n401 0.00146429
R16194 DVDD.n496 DVDD.n495 0.00146429
R16195 DVDD.n450 DVDD.n449 0.00146429
R16196 DVDD.n535 DVDD.n534 0.00146429
R16197 DVDD.n635 DVDD.n633 0.00146429
R16198 DVDD.n726 DVDD.n723 0.00146429
R16199 DVDD.n680 DVDD.n677 0.00146429
R16200 DVDD.n608 DVDD.n607 0.00146429
R16201 DVDD.n636 DVDD.n632 0.00146429
R16202 DVDD.n728 DVDD.n727 0.00146429
R16203 DVDD.n682 DVDD.n681 0.00146429
R16204 DVDD.n13733 DVDD.n13732 0.00146429
R16205 DVDD.n11284 DVDD.n11283 0.00146429
R16206 DVDD.n12490 DVDD.n12489 0.00146429
R16207 DVDD.n5744 DVDD.n5740 0.00146429
R16208 DVDD.n15204 DVDD.n15203 0.00146051
R16209 DVDD.n15125 DVDD.n15124 0.00146051
R16210 DVDD.n15013 DVDD.n15012 0.00146
R16211 DVDD.n14981 DVDD.n14980 0.00146
R16212 DVDD.n11040 DVDD.n11039 0.00146
R16213 DVDD.n16233 DVDD.n16175 0.00146
R16214 DVDD.n16232 DVDD.n16231 0.00146
R16215 DVDD.n15814 DVDD.n15813 0.00146
R16216 DVDD.n15812 DVDD.n15811 0.00146
R16217 DVDD.n14928 DVDD.n14927 0.00145625
R16218 DVDD.n15226 DVDD.n15225 0.00145625
R16219 DVDD.n10666 DVDD.n10665 0.00145625
R16220 DVDD.n3418 DVDD.n3417 0.00144995
R16221 DVDD.n1228 DVDD.n1227 0.00144287
R16222 DVDD.n12034 DVDD.n12033 0.00144287
R16223 DVDD.n12033 DVDD.n12032 0.00144287
R16224 DVDD.n12108 DVDD.n12107 0.00144287
R16225 DVDD.n1227 DVDD.n1226 0.00144287
R16226 DVDD.n4795 DVDD.n4794 0.00144287
R16227 DVDD.n5365 DVDD.n5364 0.00144287
R16228 DVDD.n5183 DVDD.n5182 0.00144287
R16229 DVDD.n4926 DVDD.n4925 0.00144287
R16230 DVDD.n11621 DVDD.n11620 0.00144287
R16231 DVDD.n1458 DVDD.n1457 0.00144287
R16232 DVDD.n2140 DVDD.n2139 0.00144287
R16233 DVDD.n6505 DVDD.n6504 0.00144287
R16234 DVDD.n6441 DVDD.n6440 0.00144287
R16235 DVDD.n6889 DVDD.n6888 0.00144287
R16236 DVDD.n9227 DVDD.n9226 0.00144287
R16237 DVDD.n8378 DVDD.n8377 0.00144287
R16238 DVDD.n7877 DVDD.n7876 0.00144287
R16239 DVDD.n3539 DVDD.n3538 0.00144287
R16240 DVDD.n8230 DVDD.n8229 0.00144142
R16241 DVDD.n8226 DVDD.n8225 0.00144142
R16242 DVDD.n9417 DVDD.n9416 0.00144142
R16243 DVDD.n8116 DVDD.n8115 0.00144142
R16244 DVDD.n7962 DVDD.n7961 0.00144142
R16245 DVDD.n7965 DVDD.n7964 0.00144142
R16246 DVDD.n7983 DVDD.n7982 0.00144142
R16247 DVDD.n8056 DVDD.n8055 0.00144142
R16248 DVDD.n11069 DVDD.n11068 0.00140496
R16249 DVDD.n15532 DVDD.n15531 0.00140496
R16250 DVDD.n16114 DVDD.n16113 0.00140496
R16251 DVDD.n16076 DVDD.n16075 0.00140496
R16252 DVDD.n16115 DVDD.n16114 0.00140496
R16253 DVDD.n15533 DVDD.n15532 0.00140496
R16254 DVDD.n16077 DVDD.n16076 0.00140496
R16255 DVDD.n11068 DVDD.n11067 0.00140496
R16256 DVDD.n3115 DVDD.n3114 0.00140175
R16257 DVDD.n3116 DVDD.n3115 0.00140175
R16258 DVDD.n18743 DVDD.n18742 0.0014
R16259 DVDD.n18746 DVDD.n18745 0.0014
R16260 DVDD.n18749 DVDD.n18748 0.0014
R16261 DVDD.n18752 DVDD.n18751 0.0014
R16262 DVDD.n18755 DVDD.n18754 0.0014
R16263 DVDD.n18758 DVDD.n18757 0.0014
R16264 DVDD.n18761 DVDD.n18760 0.0014
R16265 DVDD.n18764 DVDD.n18763 0.0014
R16266 DVDD.n18767 DVDD.n18766 0.0014
R16267 DVDD.n18770 DVDD.n18769 0.0014
R16268 DVDD.n9758 DVDD.n9757 0.0014
R16269 DVDD.n9778 DVDD.n9777 0.0014
R16270 DVDD.n9789 DVDD.n9788 0.0014
R16271 DVDD.n7908 DVDD.n7907 0.0014
R16272 DVDD.n9248 DVDD.n9247 0.0014
R16273 DVDD.n9279 DVDD.n9278 0.0014
R16274 DVDD.n9290 DVDD.n9289 0.0014
R16275 DVDD.n6857 DVDD.n6856 0.0014
R16276 DVDD.n6837 DVDD.n6836 0.0014
R16277 DVDD.n6826 DVDD.n6825 0.0014
R16278 DVDD.n6547 DVDD.n6546 0.0014
R16279 DVDD.n3994 DVDD.n3993 0.0014
R16280 DVDD.n3963 DVDD.n3962 0.0014
R16281 DVDD.n3952 DVDD.n3951 0.0014
R16282 DVDD.n18830 DVDD.n18829 0.0014
R16283 DVDD.n4894 DVDD.n4893 0.0014
R16284 DVDD.n4874 DVDD.n4873 0.0014
R16285 DVDD.n4863 DVDD.n4862 0.0014
R16286 DVDD.n5138 DVDD.n5137 0.0014
R16287 DVDD.n5299 DVDD.n5298 0.0014
R16288 DVDD.n5268 DVDD.n5267 0.0014
R16289 DVDD.n5257 DVDD.n5256 0.0014
R16290 DVDD.n2476 DVDD.n2475 0.0014
R16291 DVDD.n1752 DVDD.n1751 0.0014
R16292 DVDD.n1749 DVDD.n1748 0.0014
R16293 DVDD.n1746 DVDD.n1745 0.0014
R16294 DVDD.n19257 DVDD.n19256 0.0014
R16295 DVDD.n19260 DVDD.n19259 0.0014
R16296 DVDD.n19263 DVDD.n19262 0.0014
R16297 DVDD.n19266 DVDD.n19265 0.0014
R16298 DVDD.n19417 DVDD.n19416 0.0014
R16299 DVDD.n19420 DVDD.n19419 0.0014
R16300 DVDD.n19423 DVDD.n19422 0.0014
R16301 DVDD.n3857 DVDD.n3856 0.0014
R16302 DVDD.n7621 DVDD.n7620 0.0014
R16303 DVDD.n3913 DVDD.n3912 0.0014
R16304 DVDD.n7648 DVDD.n7647 0.0014
R16305 DVDD.n142 DVDD.n141 0.0014
R16306 DVDD.n3802 DVDD.n3801 0.0014
R16307 DVDD.n20289 DVDD.n20288 0.0014
R16308 DVDD.n20336 DVDD.n20335 0.0014
R16309 DVDD.n11859 DVDD.n11858 0.0014
R16310 DVDD.n11879 DVDD.n11878 0.0014
R16311 DVDD.n11890 DVDD.n11889 0.0014
R16312 DVDD.n11310 DVDD.n11309 0.0014
R16313 DVDD.n14913 DVDD.n14912 0.0014
R16314 DVDD.n14916 DVDD.n14915 0.0014
R16315 DVDD.n14878 DVDD.n14877 0.0014
R16316 DVDD.n10407 DVDD.n10406 0.0014
R16317 DVDD.n10560 DVDD.n10559 0.0014
R16318 DVDD.n10584 DVDD.n10583 0.0014
R16319 DVDD.n13159 DVDD.n13158 0.0014
R16320 DVDD.n13190 DVDD.n13189 0.0014
R16321 DVDD.n13201 DVDD.n13200 0.0014
R16322 DVDD.n3429 DVDD.n3428 0.0014
R16323 DVDD.n3422 DVDD.n3421 0.0014
R16324 DVDD.n3415 DVDD.n3414 0.0014
R16325 DVDD.n3409 DVDD.n3408 0.0014
R16326 DVDD.n3402 DVDD.n3401 0.0014
R16327 DVDD.n3395 DVDD.n3394 0.0014
R16328 DVDD.n3389 DVDD.n3388 0.0014
R16329 DVDD.n3383 DVDD.n3382 0.0014
R16330 DVDD.n3382 DVDD.n3381 0.0014
R16331 DVDD.n3376 DVDD.n3375 0.0014
R16332 DVDD.n3369 DVDD.n3368 0.0014
R16333 DVDD.n3362 DVDD.n3361 0.0014
R16334 DVDD.n3659 DVDD.n3658 0.0014
R16335 DVDD.n18595 DVDD.n18594 0.0014
R16336 DVDD.n18600 DVDD.n18599 0.0014
R16337 DVDD.n18599 DVDD.n18598 0.0014
R16338 DVDD.n18562 DVDD.n18561 0.0014
R16339 DVDD.n18721 DVDD.n18720 0.0014
R16340 DVDD.n18704 DVDD.n18703 0.0014
R16341 DVDD.n18709 DVDD.n18706 0.0014
R16342 DVDD.n18387 DVDD.n18386 0.0014
R16343 DVDD.n18341 DVDD.n18340 0.0014
R16344 DVDD.n18356 DVDD.n18355 0.0014
R16345 DVDD.n18353 DVDD.n18352 0.0014
R16346 DVDD.n20341 DVDD.n108 0.00139333
R16347 DVDD.n7475 DVDD.n7386 0.00139333
R16348 DVDD.n7674 DVDD.n7597 0.00139333
R16349 DVDD.n20341 DVDD.n88 0.00139333
R16350 DVDD.n7674 DVDD.n7553 0.00139333
R16351 DVDD.n20341 DVDD.n34 0.00139333
R16352 DVDD.n7674 DVDD.n7199 0.00139333
R16353 DVDD.n20341 DVDD.n20340 0.00139333
R16354 DVDD.n7676 DVDD.n7674 0.00139333
R16355 DVDD.n16324 DVDD.n16323 0.00138997
R16356 DVDD.n16323 DVDD.n16322 0.00138997
R16357 DVDD.n15045 DVDD.n15044 0.00138997
R16358 DVDD.n11026 DVDD.n11025 0.00138997
R16359 DVDD.n11081 DVDD.n11080 0.00138997
R16360 DVDD.n11027 DVDD.n11026 0.00138997
R16361 DVDD.n15046 DVDD.n15045 0.00138997
R16362 DVDD.n11082 DVDD.n11081 0.00138997
R16363 DVDD.n1232 DVDD.n1231 0.00138583
R16364 DVDD.n1216 DVDD.n1215 0.00138583
R16365 DVDD.n1213 DVDD.n1212 0.00138583
R16366 DVDD.n1150 DVDD.n1149 0.00138583
R16367 DVDD.n1553 DVDD.n1552 0.00138583
R16368 DVDD.n1567 DVDD.n1566 0.00138583
R16369 DVDD.n1574 DVDD.n1573 0.00138583
R16370 DVDD.n1577 DVDD.n1576 0.00138583
R16371 DVDD.n1582 DVDD.n1581 0.00138583
R16372 DVDD.n1589 DVDD.n1588 0.00138583
R16373 DVDD.n1597 DVDD.n1596 0.00138583
R16374 DVDD.n1604 DVDD.n1603 0.00138583
R16375 DVDD.n1610 DVDD.n1609 0.00138583
R16376 DVDD.n1616 DVDD.n1615 0.00138583
R16377 DVDD.n1623 DVDD.n1622 0.00138583
R16378 DVDD.n1630 DVDD.n1629 0.00138583
R16379 DVDD.n1638 DVDD.n1637 0.00138583
R16380 DVDD.n1667 DVDD.n1666 0.00138583
R16381 DVDD.n919 DVDD.n918 0.00138583
R16382 DVDD.n11469 DVDD.n11468 0.00138583
R16383 DVDD.n11488 DVDD.n11487 0.00138583
R16384 DVDD.n12017 DVDD.n12016 0.00138583
R16385 DVDD.n12020 DVDD.n12019 0.00138583
R16386 DVDD.n12038 DVDD.n12037 0.00138583
R16387 DVDD.n12112 DVDD.n12111 0.00138583
R16388 DVDD.n12175 DVDD.n12174 0.00138583
R16389 DVDD.n12222 DVDD.n12221 0.00138583
R16390 DVDD.n13441 DVDD.n13440 0.00138583
R16391 DVDD.n13446 DVDD.n13445 0.00138583
R16392 DVDD.n13883 DVDD.n13882 0.00138583
R16393 DVDD.n19685 DVDD.n19684 0.00138583
R16394 DVDD.n19688 DVDD.n19687 0.00138583
R16395 DVDD.n19701 DVDD.n19700 0.00138583
R16396 DVDD.n19714 DVDD.n19713 0.00138583
R16397 DVDD.n19915 DVDD.n19914 0.00138583
R16398 DVDD.n19916 DVDD.n19915 0.00138583
R16399 DVDD.n20077 DVDD.n20076 0.00138583
R16400 DVDD.n19007 DVDD.n19006 0.00138583
R16401 DVDD.n19071 DVDD.n19070 0.00138583
R16402 DVDD.n19068 DVDD.n19067 0.00138583
R16403 DVDD.n19060 DVDD.n19059 0.00138583
R16404 DVDD.n4656 DVDD.n4655 0.00138583
R16405 DVDD.n4677 DVDD.n4676 0.00138583
R16406 DVDD.n4937 DVDD.n4936 0.00138583
R16407 DVDD.n4992 DVDD.n4991 0.00138583
R16408 DVDD.n5000 DVDD.n4999 0.00138583
R16409 DVDD.n5105 DVDD.n5104 0.00138583
R16410 DVDD.n5173 DVDD.n5172 0.00138583
R16411 DVDD.n5177 DVDD.n5176 0.00138583
R16412 DVDD.n5320 DVDD.n5319 0.00138583
R16413 DVDD.n5324 DVDD.n5323 0.00138583
R16414 DVDD.n5344 DVDD.n5343 0.00138583
R16415 DVDD.n5410 DVDD.n5409 0.00138583
R16416 DVDD.n5413 DVDD.n5412 0.00138583
R16417 DVDD.n5427 DVDD.n5426 0.00138583
R16418 DVDD.n1330 DVDD.n1329 0.00138583
R16419 DVDD.n1333 DVDD.n1332 0.00138583
R16420 DVDD.n1346 DVDD.n1345 0.00138583
R16421 DVDD.n1359 DVDD.n1358 0.00138583
R16422 DVDD.n1462 DVDD.n1461 0.00138583
R16423 DVDD.n1461 DVDD.n1460 0.00138583
R16424 DVDD.n291 DVDD.n290 0.00138583
R16425 DVDD.n19216 DVDD.n19215 0.00138583
R16426 DVDD.n19453 DVDD.n19452 0.00138583
R16427 DVDD.n19450 DVDD.n19449 0.00138583
R16428 DVDD.n19442 DVDD.n19441 0.00138583
R16429 DVDD.n11363 DVDD.n11362 0.00138583
R16430 DVDD.n11384 DVDD.n11383 0.00138583
R16431 DVDD.n11827 DVDD.n11826 0.00138583
R16432 DVDD.n11820 DVDD.n11819 0.00138583
R16433 DVDD.n11816 DVDD.n11815 0.00138583
R16434 DVDD.n11761 DVDD.n11760 0.00138583
R16435 DVDD.n11753 DVDD.n11752 0.00138583
R16436 DVDD.n11650 DVDD.n11649 0.00138583
R16437 DVDD.n12354 DVDD.n12353 0.00138583
R16438 DVDD.n13135 DVDD.n13134 0.00138583
R16439 DVDD.n13115 DVDD.n13114 0.00138583
R16440 DVDD.n13052 DVDD.n13051 0.00138583
R16441 DVDD.n13049 DVDD.n13048 0.00138583
R16442 DVDD.n13036 DVDD.n13035 0.00138583
R16443 DVDD.n17261 DVDD.n17260 0.00138583
R16444 DVDD.n1907 DVDD.n1906 0.00138583
R16445 DVDD.n1910 DVDD.n1909 0.00138583
R16446 DVDD.n1923 DVDD.n1922 0.00138583
R16447 DVDD.n1936 DVDD.n1935 0.00138583
R16448 DVDD.n2136 DVDD.n2135 0.00138583
R16449 DVDD.n2137 DVDD.n2136 0.00138583
R16450 DVDD.n2298 DVDD.n2297 0.00138583
R16451 DVDD.n18899 DVDD.n18898 0.00138583
R16452 DVDD.n18963 DVDD.n18962 0.00138583
R16453 DVDD.n18960 DVDD.n18959 0.00138583
R16454 DVDD.n18952 DVDD.n18951 0.00138583
R16455 DVDD.n7028 DVDD.n7027 0.00138583
R16456 DVDD.n7007 DVDD.n7006 0.00138583
R16457 DVDD.n6758 DVDD.n6757 0.00138583
R16458 DVDD.n6751 DVDD.n6750 0.00138583
R16459 DVDD.n6747 DVDD.n6746 0.00138583
R16460 DVDD.n6692 DVDD.n6691 0.00138583
R16461 DVDD.n6684 DVDD.n6683 0.00138583
R16462 DVDD.n6577 DVDD.n6576 0.00138583
R16463 DVDD.n6509 DVDD.n6508 0.00138583
R16464 DVDD.n6437 DVDD.n6436 0.00138583
R16465 DVDD.n6417 DVDD.n6416 0.00138583
R16466 DVDD.n6351 DVDD.n6350 0.00138583
R16467 DVDD.n6348 DVDD.n6347 0.00138583
R16468 DVDD.n6334 DVDD.n6333 0.00138583
R16469 DVDD.n3273 DVDD.n3272 0.00138583
R16470 DVDD.n3270 DVDD.n3269 0.00138583
R16471 DVDD.n3257 DVDD.n3256 0.00138583
R16472 DVDD.n3244 DVDD.n3243 0.00138583
R16473 DVDD.n3535 DVDD.n3534 0.00138583
R16474 DVDD.n3536 DVDD.n3535 0.00138583
R16475 DVDD.n3777 DVDD.n3776 0.00138583
R16476 DVDD.n18520 DVDD.n18519 0.00138583
R16477 DVDD.n18800 DVDD.n18799 0.00138583
R16478 DVDD.n18797 DVDD.n18796 0.00138583
R16479 DVDD.n18789 DVDD.n18788 0.00138583
R16480 DVDD.n10045 DVDD.n10044 0.00138583
R16481 DVDD.n10024 DVDD.n10023 0.00138583
R16482 DVDD.n9726 DVDD.n9725 0.00138583
R16483 DVDD.n9719 DVDD.n9718 0.00138583
R16484 DVDD.n9715 DVDD.n9714 0.00138583
R16485 DVDD.n9660 DVDD.n9659 0.00138583
R16486 DVDD.n9652 DVDD.n9651 0.00138583
R16487 DVDD.n9545 DVDD.n9544 0.00138583
R16488 DVDD.n8374 DVDD.n8373 0.00138583
R16489 DVDD.n9223 DVDD.n9222 0.00138583
R16490 DVDD.n9203 DVDD.n9202 0.00138583
R16491 DVDD.n9137 DVDD.n9136 0.00138583
R16492 DVDD.n9134 DVDD.n9133 0.00138583
R16493 DVDD.n9120 DVDD.n9119 0.00138583
R16494 DVDD.n501 DVDD.n500 0.00138568
R16495 DVDD.n500 DVDD.n499 0.00138568
R16496 DVDD.n15970 DVDD.n15969 0.00137654
R16497 DVDD.n15971 DVDD.n15970 0.00137654
R16498 DVDD.n8276 DVDD.n8275 0.00137654
R16499 DVDD.n9445 DVDD.n9444 0.00137654
R16500 DVDD.n9446 DVDD.n9445 0.00137654
R16501 DVDD.n8127 DVDD.n8126 0.00137654
R16502 DVDD.n8126 DVDD.n8125 0.00137654
R16503 DVDD.n7987 DVDD.n7986 0.00137654
R16504 DVDD.n8043 DVDD.n8042 0.00137654
R16505 DVDD.n7988 DVDD.n7987 0.00137654
R16506 DVDD.n8042 DVDD.n8041 0.00137654
R16507 DVDD.n10509 DVDD.n10508 0.00137497
R16508 DVDD.n17166 DVDD.n17165 0.00137497
R16509 DVDD.n17119 DVDD.n17118 0.00137497
R16510 DVDD.n17069 DVDD.n17068 0.00137497
R16511 DVDD.n17070 DVDD.n17069 0.00137497
R16512 DVDD.n17120 DVDD.n17119 0.00137497
R16513 DVDD.n10510 DVDD.n10509 0.00137497
R16514 DVDD.n17167 DVDD.n17166 0.00137497
R16515 DVDD.n15210 DVDD.n15209 0.00136446
R16516 DVDD.n15129 DVDD.n15128 0.00136446
R16517 DVDD.n6196 DVDD.n6195 0.00135432
R16518 DVDD.n8898 DVDD.n8897 0.00135432
R16519 DVDD.n1236 DVDD.n1235 0.0013543
R16520 DVDD.n12100 DVDD.n12099 0.0013543
R16521 DVDD.n12186 DVDD.n12185 0.0013543
R16522 DVDD.n12250 DVDD.n12249 0.0013543
R16523 DVDD.n13395 DVDD.n13394 0.0013543
R16524 DVDD.n13724 DVDD.n13723 0.0013543
R16525 DVDD.n12185 DVDD.n12184 0.0013543
R16526 DVDD.n12099 DVDD.n12098 0.0013543
R16527 DVDD.n12042 DVDD.n12041 0.0013543
R16528 DVDD.n12251 DVDD.n12250 0.0013543
R16529 DVDD.n13394 DVDD.n13393 0.0013543
R16530 DVDD.n15486 DVDD.n15485 0.0013543
R16531 DVDD.n15514 DVDD.n15513 0.0013543
R16532 DVDD.n14663 DVDD.n14662 0.0013543
R16533 DVDD.n14376 DVDD.n14375 0.0013543
R16534 DVDD.n14664 DVDD.n14663 0.0013543
R16535 DVDD.n15485 DVDD.n15484 0.0013543
R16536 DVDD.n15513 DVDD.n15512 0.0013543
R16537 DVDD.n5046 DVDD.n5045 0.0013543
R16538 DVDD.n5065 DVDD.n5064 0.0013543
R16539 DVDD.n5102 DVDD.n5101 0.0013543
R16540 DVDD.n5379 DVDD.n5378 0.0013543
R16541 DVDD.n5562 DVDD.n5561 0.0013543
R16542 DVDD.n5637 DVDD.n5636 0.0013543
R16543 DVDD.n5938 DVDD.n5937 0.0013543
R16544 DVDD.n5561 DVDD.n5560 0.0013543
R16545 DVDD.n5378 DVDD.n5377 0.0013543
R16546 DVDD.n5045 DVDD.n5044 0.0013543
R16547 DVDD.n5101 DVDD.n5100 0.0013543
R16548 DVDD.n5636 DVDD.n5635 0.0013543
R16549 DVDD.n11708 DVDD.n11707 0.0013543
R16550 DVDD.n11653 DVDD.n11652 0.0013543
R16551 DVDD.n13082 DVDD.n13081 0.0013543
R16552 DVDD.n12855 DVDD.n12854 0.0013543
R16553 DVDD.n12800 DVDD.n12799 0.0013543
R16554 DVDD.n12601 DVDD.n12600 0.0013543
R16555 DVDD.n11709 DVDD.n11708 0.0013543
R16556 DVDD.n11661 DVDD.n11660 0.0013543
R16557 DVDD.n13106 DVDD.n13105 0.0013543
R16558 DVDD.n12856 DVDD.n12855 0.0013543
R16559 DVDD.n12801 DVDD.n12800 0.0013543
R16560 DVDD.n18123 DVDD.n18122 0.0013543
R16561 DVDD.n18097 DVDD.n18096 0.0013543
R16562 DVDD.n18019 DVDD.n18018 0.0013543
R16563 DVDD.n17754 DVDD.n17753 0.0013543
R16564 DVDD.n18020 DVDD.n18019 0.0013543
R16565 DVDD.n18124 DVDD.n18123 0.0013543
R16566 DVDD.n18098 DVDD.n18097 0.0013543
R16567 DVDD.n6638 DVDD.n6637 0.0013543
R16568 DVDD.n6580 DVDD.n6579 0.0013543
R16569 DVDD.n6382 DVDD.n6381 0.0013543
R16570 DVDD.n6180 DVDD.n6179 0.0013543
R16571 DVDD.n4397 DVDD.n4396 0.0013543
R16572 DVDD.n6407 DVDD.n6406 0.0013543
R16573 DVDD.n6383 DVDD.n6382 0.0013543
R16574 DVDD.n6639 DVDD.n6638 0.0013543
R16575 DVDD.n6589 DVDD.n6588 0.0013543
R16576 DVDD.n6581 DVDD.n6580 0.0013543
R16577 DVDD.n6235 DVDD.n6234 0.0013543
R16578 DVDD.n6181 DVDD.n6180 0.0013543
R16579 DVDD.n4398 DVDD.n4397 0.0013543
R16580 DVDD.n13725 DVDD.n13724 0.0013543
R16581 DVDD.n17755 DVDD.n17754 0.0013543
R16582 DVDD.n5939 DVDD.n5938 0.0013543
R16583 DVDD.n14377 DVDD.n14376 0.0013543
R16584 DVDD.n12602 DVDD.n12601 0.0013543
R16585 DVDD.n9606 DVDD.n9605 0.0013543
R16586 DVDD.n9548 DVDD.n9547 0.0013543
R16587 DVDD.n9168 DVDD.n9167 0.0013543
R16588 DVDD.n8882 DVDD.n8881 0.0013543
R16589 DVDD.n8671 DVDD.n8670 0.0013543
R16590 DVDD.n9607 DVDD.n9606 0.0013543
R16591 DVDD.n8937 DVDD.n8936 0.0013543
R16592 DVDD.n8672 DVDD.n8671 0.0013543
R16593 DVDD.n9193 DVDD.n9192 0.0013543
R16594 DVDD.n9169 DVDD.n9168 0.0013543
R16595 DVDD.n9557 DVDD.n9556 0.0013543
R16596 DVDD.n9549 DVDD.n9548 0.0013543
R16597 DVDD.n8883 DVDD.n8882 0.0013543
R16598 DVDD.n498 DVDD.n497 0.00135354
R16599 DVDD.n2323 DVDD.n2322 0.00135354
R16600 DVDD.n2399 DVDD.n2398 0.00135354
R16601 DVDD.n499 DVDD.n498 0.00135354
R16602 DVDD.n2322 DVDD.n2321 0.00135354
R16603 DVDD.n2398 DVDD.n2397 0.00135354
R16604 DVDD.n10482 DVDD.n10481 0.00134375
R16605 DVDD.n10667 DVDD.n10666 0.00134375
R16606 DVDD.n10679 DVDD.n10678 0.00134375
R16607 DVDD.n10720 DVDD.n10719 0.00134375
R16608 DVDD.n10406 DVDD.n10405 0.00134375
R16609 DVDD.n10561 DVDD.n10560 0.00134375
R16610 DVDD.n10585 DVDD.n10584 0.00134375
R16611 DVDD.n10639 DVDD.n10638 0.00134375
R16612 DVDD.n11139 DVDD 0.00134
R16613 DVDD DVDD.n11144 0.00134
R16614 DVDD.n11265 DVDD.n11264 0.00133571
R16615 DVDD.n11253 DVDD.n11252 0.00133571
R16616 DVDD.n11237 DVDD.n11236 0.00133571
R16617 DVDD.n5743 DVDD.n5742 0.00133571
R16618 DVDD.n303 DVDD.n302 0.00133571
R16619 DVDD.n404 DVDD.n403 0.00133571
R16620 DVDD.n494 DVDD.n493 0.00133571
R16621 DVDD.n448 DVDD.n447 0.00133571
R16622 DVDD.n378 DVDD.n377 0.00133571
R16623 DVDD.n406 DVDD.n405 0.00133571
R16624 DVDD.n495 DVDD.n490 0.00133571
R16625 DVDD.n449 DVDD.n444 0.00133571
R16626 DVDD.n534 DVDD.n533 0.00133571
R16627 DVDD.n635 DVDD.n634 0.00133571
R16628 DVDD.n726 DVDD.n725 0.00133571
R16629 DVDD.n680 DVDD.n679 0.00133571
R16630 DVDD.n609 DVDD.n608 0.00133571
R16631 DVDD.n637 DVDD.n636 0.00133571
R16632 DVDD.n727 DVDD.n722 0.00133571
R16633 DVDD.n681 DVDD.n676 0.00133571
R16634 DVDD.n13732 DVDD.n13731 0.00133571
R16635 DVDD.n11283 DVDD.n11282 0.00133571
R16636 DVDD.n12491 DVDD.n12490 0.00133571
R16637 DVDD.n5745 DVDD.n5744 0.00133571
R16638 DVDD.n11142 DVDD 0.00132667
R16639 DVDD.n2396 DVDD.n2395 0.00132141
R16640 DVDD.n2397 DVDD.n2396 0.00132141
R16641 DVDD.n7696 DVDD.n7695 0.00131
R16642 DVDD.n7698 DVDD.n7697 0.00131
R16643 DVDD.n3690 DVDD.n3689 0.00131
R16644 DVDD.n3688 DVDD.n3687 0.00131
R16645 DVDD.n18534 DVDD.n18533 0.00131
R16646 DVDD.n18536 DVDD.n18535 0.00131
R16647 DVDD.n18780 DVDD.n18779 0.00131
R16648 DVDD.n2950 DVDD.n2949 0.00131
R16649 DVDD.n2952 DVDD.n2951 0.00131
R16650 DVDD.n9808 DVDD.n9807 0.00131
R16651 DVDD.n2188 DVDD.n2187 0.00131
R16652 DVDD.n2190 DVDD.n2189 0.00131
R16653 DVDD.n2246 DVDD.n2245 0.00131
R16654 DVDD.n2244 DVDD.n2243 0.00131
R16655 DVDD.n18903 DVDD.n18902 0.00131
R16656 DVDD.n18905 DVDD.n18904 0.00131
R16657 DVDD.n18933 DVDD.n18932 0.00131
R16658 DVDD.n7104 DVDD.n7103 0.00131
R16659 DVDD.n7071 DVDD.n7070 0.00131
R16660 DVDD.n6807 DVDD.n6806 0.00131
R16661 DVDD.n1904 DVDD.n1903 0.00131
R16662 DVDD.n19967 DVDD.n19966 0.00131
R16663 DVDD.n19969 DVDD.n19968 0.00131
R16664 DVDD.n20025 DVDD.n20024 0.00131
R16665 DVDD.n20023 DVDD.n20022 0.00131
R16666 DVDD.n19021 DVDD.n19020 0.00131
R16667 DVDD.n19023 DVDD.n19022 0.00131
R16668 DVDD.n19051 DVDD.n19050 0.00131
R16669 DVDD.n3883 DVDD.n3882 0.00131
R16670 DVDD.n4651 DVDD.n4650 0.00131
R16671 DVDD.n4844 DVDD.n4843 0.00131
R16672 DVDD.n19682 DVDD.n19681 0.00131
R16673 DVDD.n978 DVDD.n977 0.00131
R16674 DVDD.n976 DVDD.n975 0.00131
R16675 DVDD.n933 DVDD.n932 0.00131
R16676 DVDD.n931 DVDD.n930 0.00131
R16677 DVDD.n19230 DVDD.n19229 0.00131
R16678 DVDD.n19232 DVDD.n19231 0.00131
R16679 DVDD.n19433 DVDD.n19432 0.00131
R16680 DVDD.n18329 DVDD.n18328 0.00131
R16681 DVDD.n18327 DVDD.n18326 0.00131
R16682 DVDD.n7375 DVDD.n7374 0.00131
R16683 DVDD.n65 DVDD.n64 0.00131
R16684 DVDD.n7248 DVDD.n7247 0.00131
R16685 DVDD.n11909 DVDD.n11908 0.00131
R16686 DVDD.n1327 DVDD.n1326 0.00131
R16687 DVDD.n14965 DVDD.n14964 0.00131
R16688 DVDD.n15042 DVDD.n15041 0.00131
R16689 DVDD.n15325 DVDD.n14832 0.00131
R16690 DVDD.n15351 DVDD.n15350 0.00131
R16691 DVDD.n14967 DVDD.n14966 0.00131
R16692 DVDD.n15032 DVDD.n15031 0.00131
R16693 DVDD.n15044 DVDD.n15043 0.00131
R16694 DVDD.n15317 DVDD.n15316 0.00131
R16695 DVDD.n15324 DVDD.n14826 0.00131
R16696 DVDD.n15352 DVDD.n15348 0.00131
R16697 DVDD.n11025 DVDD.n11024 0.00131
R16698 DVDD.n11080 DVDD.n11079 0.00131
R16699 DVDD.n15524 DVDD.n15519 0.00131
R16700 DVDD.n11159 DVDD.n11155 0.00131
R16701 DVDD.n16159 DVDD.n16158 0.00131
R16702 DVDD.n16277 DVDD.n16276 0.00131
R16703 DVDD.n16316 DVDD.n16315 0.00131
R16704 DVDD.n16322 DVDD.n16321 0.00131
R16705 DVDD.n16363 DVDD.n16359 0.00131
R16706 DVDD.n16215 DVDD.n16214 0.00131
R16707 DVDD.n15580 DVDD.n15579 0.00131
R16708 DVDD.n15754 DVDD.n15753 0.00131
R16709 DVDD.n15744 DVDD.n15741 0.00131
R16710 DVDD.n15718 DVDD.n15717 0.00131
R16711 DVDD.n15708 DVDD.n15613 0.00131
R16712 DVDD.n15794 DVDD.n15793 0.00131
R16713 DVDD.n15857 DVDD.n15856 0.00131
R16714 DVDD.n16104 DVDD.n16101 0.00131
R16715 DVDD.n15918 DVDD.n15892 0.00131
R16716 DVDD.n15792 DVDD.n15791 0.00131
R16717 DVDD.n15855 DVDD.n15854 0.00131
R16718 DVDD.n16103 DVDD.n16102 0.00131
R16719 DVDD.n15917 DVDD.n15893 0.00131
R16720 DVDD.n16213 DVDD.n16212 0.00131
R16721 DVDD.n15578 DVDD.n15577 0.00131
R16722 DVDD.n15743 DVDD.n15742 0.00131
R16723 DVDD.n15707 DVDD.n15614 0.00131
R16724 DVDD.n16157 DVDD.n16156 0.00131
R16725 DVDD.n16275 DVDD.n16274 0.00131
R16726 DVDD.n11115 DVDD.n11114 0.00131
R16727 DVDD.n16362 DVDD.n16361 0.00131
R16728 DVDD.n11023 DVDD.n11022 0.00131
R16729 DVDD.n15523 DVDD.n15522 0.00131
R16730 DVDD.n11158 DVDD.n11157 0.00131
R16731 DVDD.n3276 DVDD.n3275 0.00131
R16732 DVDD.n20255 DVDD.n20254 0.00131
R16733 DVDD.n3120 DVDD.n3119 0.00130357
R16734 DVDD.n3088 DVDD.n3087 0.00130357
R16735 DVDD.n3084 DVDD.n3083 0.00130357
R16736 DVDD.n3054 DVDD.n3053 0.00130132
R16737 DVDD.n3087 DVDD.n3086 0.00130132
R16738 DVDD.n3055 DVDD.n3054 0.00130132
R16739 DVDD.n10195 DVDD.n10194 0.0013
R16740 DVDD.n10245 DVDD.n10237 0.0013
R16741 DVDD.n15916 DVDD 0.00128667
R16742 DVDD.n15949 DVDD.n15948 0.00128241
R16743 DVDD.n15948 DVDD.n15947 0.00128241
R16744 DVDD.n15689 DVDD.n15688 0.00128241
R16745 DVDD.n15688 DVDD.n15687 0.00128241
R16746 DVDD.n8213 DVDD.n8212 0.00128241
R16747 DVDD.n9410 DVDD.n9409 0.00128241
R16748 DVDD.n9411 DVDD.n9410 0.00128241
R16749 DVDD.n9893 DVDD.n9892 0.00128241
R16750 DVDD.n9894 DVDD.n9893 0.00128241
R16751 DVDD.n18851 DVDD.n18850 0.00128
R16752 DVDD.n19099 DVDD.n19098 0.00128
R16753 DVDD.n7363 DVDD.n7361 0.00128
R16754 DVDD.n7413 DVDD.n7412 0.00128
R16755 DVDD.n7586 DVDD.n7584 0.00128
R16756 DVDD.n77 DVDD.n75 0.00128
R16757 DVDD.n7461 DVDD.n7460 0.00128
R16758 DVDD.n7542 DVDD.n7540 0.00128
R16759 DVDD.n7236 DVDD.n7234 0.00128
R16760 DVDD.n7490 DVDD.n7489 0.00128
R16761 DVDD.n7188 DVDD.n7186 0.00128
R16762 DVDD.n19376 DVDD.n19375 0.00128
R16763 DVDD.n14961 DVDD.n14960 0.00128
R16764 DVDD.n15034 DVDD.n15033 0.00128
R16765 DVDD.n15319 DVDD.n15318 0.00128
R16766 DVDD.n15360 DVDD.n15358 0.00128
R16767 DVDD.n14956 DVDD.n14955 0.00128
R16768 DVDD.n14968 DVDD.n14967 0.00128
R16769 DVDD.n15035 DVDD.n15032 0.00128
R16770 DVDD.n15320 DVDD.n15317 0.00128
R16771 DVDD.n15387 DVDD.n14826 0.00128
R16772 DVDD.n15362 DVDD.n15361 0.00128
R16773 DVDD.n11016 DVDD.n11013 0.00128
R16774 DVDD.n11072 DVDD.n11069 0.00128
R16775 DVDD.n15531 DVDD.n15530 0.00128
R16776 DVDD.n15519 DVDD.n15518 0.00128
R16777 DVDD.n11166 DVDD.n11165 0.00128
R16778 DVDD.n16149 DVDD.n16145 0.00128
R16779 DVDD.n16267 DVDD.n16263 0.00128
R16780 DVDD.n16317 DVDD.n16316 0.00128
R16781 DVDD.n16370 DVDD.n16369 0.00128
R16782 DVDD.n16205 DVDD.n16201 0.00128
R16783 DVDD.n15570 DVDD.n15566 0.00128
R16784 DVDD.n15753 DVDD.n15752 0.00128
R16785 DVDD.n15741 DVDD.n15740 0.00128
R16786 DVDD.n15717 DVDD.n15716 0.00128
R16787 DVDD.n15693 DVDD.n15613 0.00128
R16788 DVDD.n15784 DVDD.n15780 0.00128
R16789 DVDD.n15847 DVDD.n15843 0.00128
R16790 DVDD.n16113 DVDD.n16112 0.00128
R16791 DVDD.n16101 DVDD.n16100 0.00128
R16792 DVDD.n16075 DVDD.n16074 0.00128
R16793 DVDD.n15905 DVDD.n15892 0.00128
R16794 DVDD.n15783 DVDD.n15781 0.00128
R16795 DVDD.n15846 DVDD.n15844 0.00128
R16796 DVDD.n16111 DVDD.n16108 0.00128
R16797 DVDD.n16073 DVDD.n16070 0.00128
R16798 DVDD.n16204 DVDD.n16202 0.00128
R16799 DVDD.n15569 DVDD.n15567 0.00128
R16800 DVDD.n15751 DVDD.n15748 0.00128
R16801 DVDD.n15715 DVDD.n15712 0.00128
R16802 DVDD.n16148 DVDD.n16146 0.00128
R16803 DVDD.n16266 DVDD.n16264 0.00128
R16804 DVDD.n11119 DVDD.n11118 0.00128
R16805 DVDD.n16379 DVDD.n16378 0.00128
R16806 DVDD.n11015 DVDD.n11014 0.00128
R16807 DVDD.n11071 DVDD.n11070 0.00128
R16808 DVDD.n15529 DVDD.n15528 0.00128
R16809 DVDD.n11175 DVDD.n11174 0.00128
R16810 DVDD.n18372 DVDD.n18371 0.00128
R16811 DVDD.n20267 DVDD.n20265 0.00128
R16812 DVDD.n7329 DVDD.n7328 0.00128
R16813 DVDD.n7687 DVDD.n7685 0.00128
R16814 DVDD.n375 DVDD.n374 0.00127143
R16815 DVDD.n400 DVDD.n399 0.00127143
R16816 DVDD.n452 DVDD.n451 0.00127143
R16817 DVDD.n606 DVDD.n605 0.00127143
R16818 DVDD.n631 DVDD.n630 0.00127143
R16819 DVDD.n731 DVDD.n730 0.00127143
R16820 DVDD.n684 DVDD.n683 0.00127143
R16821 DVDD.n13735 DVDD.n13734 0.00127143
R16822 DVDD.n11286 DVDD.n11285 0.00127143
R16823 DVDD.n12488 DVDD.n12487 0.00127143
R16824 DVDD.n5739 DVDD.n5738 0.00127143
R16825 DVDD.n11172 DVDD.n11171 0.00126998
R16826 DVDD.n11168 DVDD.n11167 0.00126998
R16827 DVDD.n11167 DVDD.n11166 0.00126998
R16828 DVDD.n11171 DVDD.n11170 0.00126998
R16829 DVDD.n15207 DVDD.n15206 0.00126841
R16830 DVDD.n1207 DVDD.n1206 0.00126573
R16831 DVDD.n1596 DVDD.n1595 0.00126573
R16832 DVDD.n11477 DVDD.n11476 0.00126573
R16833 DVDD.n12215 DVDD.n12214 0.00126573
R16834 DVDD.n13460 DVDD.n13459 0.00126573
R16835 DVDD.n13540 DVDD.n13539 0.00126573
R16836 DVDD.n13621 DVDD.n13620 0.00126573
R16837 DVDD.n11478 DVDD.n11477 0.00126573
R16838 DVDD.n1635 DVDD.n1634 0.00126573
R16839 DVDD.n1208 DVDD.n1207 0.00126573
R16840 DVDD.n1176 DVDD.n1175 0.00126573
R16841 DVDD.n12216 DVDD.n12215 0.00126573
R16842 DVDD.n13461 DVDD.n13460 0.00126573
R16843 DVDD.n13539 DVDD.n13538 0.00126573
R16844 DVDD.n13620 DVDD.n13619 0.00126573
R16845 DVDD.n2733 DVDD.n2732 0.00126573
R16846 DVDD.n2774 DVDD.n2773 0.00126573
R16847 DVDD.n14823 DVDD.n14822 0.00126573
R16848 DVDD.n14718 DVDD.n14717 0.00126573
R16849 DVDD.n14635 DVDD.n14634 0.00126573
R16850 DVDD.n14581 DVDD.n14580 0.00126573
R16851 DVDD.n14493 DVDD.n14492 0.00126573
R16852 DVDD.n14719 DVDD.n14718 0.00126573
R16853 DVDD.n14822 DVDD.n14821 0.00126573
R16854 DVDD.n2732 DVDD.n2731 0.00126573
R16855 DVDD.n2773 DVDD.n2772 0.00126573
R16856 DVDD.n14636 DVDD.n14635 0.00126573
R16857 DVDD.n14582 DVDD.n14581 0.00126573
R16858 DVDD.n14494 DVDD.n14493 0.00126573
R16859 DVDD.n19718 DVDD.n19717 0.00126573
R16860 DVDD.n19885 DVDD.n19884 0.00126573
R16861 DVDD.n4787 DVDD.n4786 0.00126573
R16862 DVDD.n4922 DVDD.n4921 0.00126573
R16863 DVDD.n5207 DVDD.n5206 0.00126573
R16864 DVDD.n5436 DVDD.n5435 0.00126573
R16865 DVDD.n5554 DVDD.n5553 0.00126573
R16866 DVDD.n6089 DVDD.n6088 0.00126573
R16867 DVDD.n5206 DVDD.n5205 0.00126573
R16868 DVDD.n4799 DVDD.n4798 0.00126573
R16869 DVDD.n4786 DVDD.n4785 0.00126573
R16870 DVDD.n19717 DVDD.n19716 0.00126573
R16871 DVDD.n19884 DVDD.n19883 0.00126573
R16872 DVDD.n5435 DVDD.n5434 0.00126573
R16873 DVDD.n5553 DVDD.n5552 0.00126573
R16874 DVDD.n6090 DVDD.n6089 0.00126573
R16875 DVDD.n1363 DVDD.n1362 0.00126573
R16876 DVDD.n1492 DVDD.n1491 0.00126573
R16877 DVDD.n11613 DVDD.n11612 0.00126573
R16878 DVDD.n12387 DVDD.n12386 0.00126573
R16879 DVDD.n13027 DVDD.n13026 0.00126573
R16880 DVDD.n12863 DVDD.n12862 0.00126573
R16881 DVDD.n12721 DVDD.n12720 0.00126573
R16882 DVDD.n12386 DVDD.n12385 0.00126573
R16883 DVDD.n11831 DVDD.n11830 0.00126573
R16884 DVDD.n11801 DVDD.n11800 0.00126573
R16885 DVDD.n11612 DVDD.n11611 0.00126573
R16886 DVDD.n1362 DVDD.n1361 0.00126573
R16887 DVDD.n1493 DVDD.n1492 0.00126573
R16888 DVDD.n13028 DVDD.n13027 0.00126573
R16889 DVDD.n12864 DVDD.n12863 0.00126573
R16890 DVDD.n12722 DVDD.n12721 0.00126573
R16891 DVDD.n771 DVDD.n770 0.00126573
R16892 DVDD.n808 DVDD.n807 0.00126573
R16893 DVDD.n18215 DVDD.n18214 0.00126573
R16894 DVDD.n18071 DVDD.n18070 0.00126573
R16895 DVDD.n17993 DVDD.n17992 0.00126573
R16896 DVDD.n17941 DVDD.n17940 0.00126573
R16897 DVDD.n17860 DVDD.n17859 0.00126573
R16898 DVDD.n18072 DVDD.n18071 0.00126573
R16899 DVDD.n18216 DVDD.n18215 0.00126573
R16900 DVDD.n770 DVDD.n769 0.00126573
R16901 DVDD.n807 DVDD.n806 0.00126573
R16902 DVDD.n17994 DVDD.n17993 0.00126573
R16903 DVDD.n17942 DVDD.n17941 0.00126573
R16904 DVDD.n17861 DVDD.n17860 0.00126573
R16905 DVDD.n1940 DVDD.n1939 0.00126573
R16906 DVDD.n2106 DVDD.n2105 0.00126573
R16907 DVDD.n6897 DVDD.n6896 0.00126573
R16908 DVDD.n6732 DVDD.n6731 0.00126573
R16909 DVDD.n6681 DVDD.n6680 0.00126573
R16910 DVDD.n6475 DVDD.n6474 0.00126573
R16911 DVDD.n6325 DVDD.n6324 0.00126573
R16912 DVDD.n6242 DVDD.n6241 0.00126573
R16913 DVDD.n4539 DVDD.n4538 0.00126573
R16914 DVDD.n6476 DVDD.n6475 0.00126573
R16915 DVDD.n6762 DVDD.n6761 0.00126573
R16916 DVDD.n6898 DVDD.n6897 0.00126573
R16917 DVDD.n1939 DVDD.n1938 0.00126573
R16918 DVDD.n2105 DVDD.n2104 0.00126573
R16919 DVDD.n6326 DVDD.n6325 0.00126573
R16920 DVDD.n6243 DVDD.n6242 0.00126573
R16921 DVDD.n4540 DVDD.n4539 0.00126573
R16922 DVDD.n3240 DVDD.n3239 0.00126573
R16923 DVDD.n3505 DVDD.n3504 0.00126573
R16924 DVDD.n7869 DVDD.n7868 0.00126573
R16925 DVDD.n8408 DVDD.n8407 0.00126573
R16926 DVDD.n9111 DVDD.n9110 0.00126573
R16927 DVDD.n8944 DVDD.n8943 0.00126573
R16928 DVDD.n8806 DVDD.n8805 0.00126573
R16929 DVDD.n8407 DVDD.n8406 0.00126573
R16930 DVDD.n9730 DVDD.n9729 0.00126573
R16931 DVDD.n9700 DVDD.n9699 0.00126573
R16932 DVDD.n9649 DVDD.n9648 0.00126573
R16933 DVDD.n7868 DVDD.n7867 0.00126573
R16934 DVDD.n3241 DVDD.n3240 0.00126573
R16935 DVDD.n3504 DVDD.n3503 0.00126573
R16936 DVDD.n9112 DVDD.n9111 0.00126573
R16937 DVDD.n8945 DVDD.n8944 0.00126573
R16938 DVDD.n8807 DVDD.n8806 0.00126573
R16939 DVDD.n11032 DVDD.n11031 0.00125499
R16940 DVDD.n11189 DVDD.n11188 0.00125499
R16941 DVDD.n11136 DVDD.n11124 0.00125499
R16942 DVDD.n16332 DVDD.n16331 0.00125499
R16943 DVDD.n16347 DVDD.n16346 0.00125499
R16944 DVDD.n11188 DVDD.n11187 0.00125499
R16945 DVDD.n16331 DVDD.n16330 0.00125499
R16946 DVDD.n11033 DVDD.n11032 0.00125499
R16947 DVDD.n16346 DVDD.n16342 0.00125499
R16948 DVDD.n11137 DVDD.n11136 0.00125499
R16949 DVDD.n8293 DVDD.n8292 0.00125314
R16950 DVDD.n8289 DVDD.n8288 0.00125314
R16951 DVDD.n7954 DVDD.n7953 0.00125314
R16952 DVDD.n7958 DVDD.n7957 0.00125314
R16953 DVDD.n7992 DVDD.n7991 0.00125314
R16954 DVDD.n8047 DVDD.n8046 0.00125314
R16955 DVDD.n1833 DVDD.n1832 0.00125
R16956 DVDD.n18895 DVDD.n18894 0.00125
R16957 DVDD.n18874 DVDD.n18873 0.00125
R16958 DVDD.n18854 DVDD.n18853 0.00125
R16959 DVDD.n18838 DVDD.n18837 0.00125
R16960 DVDD.n19611 DVDD.n19610 0.00125
R16961 DVDD.n19144 DVDD.n19143 0.00125
R16962 DVDD.n19123 DVDD.n19122 0.00125
R16963 DVDD.n19102 DVDD.n19101 0.00125
R16964 DVDD.n19086 DVDD.n19085 0.00125
R16965 DVDD.n11 DVDD.n9 0.00125
R16966 DVDD.n7425 DVDD.n7424 0.00125
R16967 DVDD.n7401 DVDD.n7399 0.00125
R16968 DVDD.n93 DVDD.n91 0.00125
R16969 DVDD.n7473 DVDD.n7472 0.00125
R16970 DVDD.n7449 DVDD.n7447 0.00125
R16971 DVDD.n39 DVDD.n37 0.00125
R16972 DVDD.n7478 DVDD.n7477 0.00125
R16973 DVDD.n7502 DVDD.n7500 0.00125
R16974 DVDD.n19343 DVDD.n19342 0.00125
R16975 DVDD.n19379 DVDD.n19378 0.00125
R16976 DVDD.n10377 DVDD.n10376 0.00125
R16977 DVDD.n10438 DVDD.n10437 0.00125
R16978 DVDD.n16868 DVDD.n16867 0.00125
R16979 DVDD.n16714 DVDD.n16713 0.00125
R16980 DVDD.n16736 DVDD.n16735 0.00125
R16981 DVDD.n16545 DVDD.n16544 0.00125
R16982 DVDD.n16568 DVDD.n16567 0.00125
R16983 DVDD.n18462 DVDD.n18461 0.00125
R16984 DVDD.n18375 DVDD.n18374 0.00125
R16985 DVDD.n20229 DVDD.n20227 0.00125
R16986 DVDD.n7341 DVDD.n7340 0.00125
R16987 DVDD.n7317 DVDD.n7315 0.00125
R16988 DVDD.n10447 DVDD.n10446 0.00123999
R16989 DVDD.n17075 DVDD.n17074 0.00123999
R16990 DVDD.n17076 DVDD.n17075 0.00123999
R16991 DVDD.n10448 DVDD.n10447 0.00123999
R16992 DVDD.n10481 DVDD.n10480 0.00123125
R16993 DVDD.n10668 DVDD.n10667 0.00123125
R16994 DVDD.n10680 DVDD.n10679 0.00123125
R16995 DVDD.n10719 DVDD.n10718 0.00123125
R16996 DVDD.n10405 DVDD.n10404 0.00123125
R16997 DVDD.n10562 DVDD.n10561 0.00123125
R16998 DVDD.n10586 DVDD.n10585 0.00123125
R16999 DVDD.n10638 DVDD.n10637 0.00123125
R17000 DVDD.n18986 DVDD.n18985 0.00123001
R17001 DVDD.n10553 DVDD.n10552 0.00123001
R17002 DVDD.n8298 DVDD.n8297 0.00122973
R17003 DVDD.n9756 DVDD.n9755 0.00122
R17004 DVDD.n9780 DVDD.n9779 0.00122
R17005 DVDD.n9787 DVDD.n9786 0.00122
R17006 DVDD.n7906 DVDD.n7905 0.00122
R17007 DVDD.n9491 DVDD.n9490 0.00122
R17008 DVDD.n9246 DVDD.n9245 0.00122
R17009 DVDD.n9281 DVDD.n9280 0.00122
R17010 DVDD.n9288 DVDD.n9287 0.00122
R17011 DVDD.n6859 DVDD.n6858 0.00122
R17012 DVDD.n6835 DVDD.n6834 0.00122
R17013 DVDD.n6828 DVDD.n6827 0.00122
R17014 DVDD.n6549 DVDD.n6548 0.00122
R17015 DVDD.n3996 DVDD.n3995 0.00122
R17016 DVDD.n3961 DVDD.n3960 0.00122
R17017 DVDD.n3954 DVDD.n3953 0.00122
R17018 DVDD.n4896 DVDD.n4895 0.00122
R17019 DVDD.n4872 DVDD.n4871 0.00122
R17020 DVDD.n4865 DVDD.n4864 0.00122
R17021 DVDD.n5140 DVDD.n5139 0.00122
R17022 DVDD.n5301 DVDD.n5300 0.00122
R17023 DVDD.n5266 DVDD.n5265 0.00122
R17024 DVDD.n5259 DVDD.n5258 0.00122
R17025 DVDD.n1854 DVDD.n1853 0.00122
R17026 DVDD.n20215 DVDD.n19599 0.00122
R17027 DVDD.n19632 DVDD.n19631 0.00122
R17028 DVDD.n20215 DVDD.n20214 0.00122
R17029 DVDD.n23 DVDD.n21 0.00122
R17030 DVDD.n7389 DVDD.n7387 0.00122
R17031 DVDD.n105 DVDD.n103 0.00122
R17032 DVDD.n7437 DVDD.n7435 0.00122
R17033 DVDD.n51 DVDD.n49 0.00122
R17034 DVDD.n7623 DVDD.n7622 0.00122
R17035 DVDD.n1803 DVDD.n1802 0.00122
R17036 DVDD.n11857 DVDD.n11856 0.00122
R17037 DVDD.n11881 DVDD.n11880 0.00122
R17038 DVDD.n11888 DVDD.n11887 0.00122
R17039 DVDD.n11308 DVDD.n11307 0.00122
R17040 DVDD.n12296 DVDD.n12295 0.00122
R17041 DVDD.n10346 DVDD.n10344 0.00122
R17042 DVDD.n10380 DVDD.n10378 0.00122
R17043 DVDD.n10506 DVDD.n10504 0.00122
R17044 DVDD.n10435 DVDD.n10432 0.00122
R17045 DVDD.n15312 DVDD.n15311 0.00122
R17046 DVDD.n10347 DVDD.n10343 0.00122
R17047 DVDD.n10381 DVDD.n10377 0.00122
R17048 DVDD.n10508 DVDD.n10507 0.00122
R17049 DVDD.n10437 DVDD.n10436 0.00122
R17050 DVDD.n15314 DVDD.n15313 0.00122
R17051 DVDD.n13157 DVDD.n13156 0.00122
R17052 DVDD.n13192 DVDD.n13191 0.00122
R17053 DVDD.n13199 DVDD.n13198 0.00122
R17054 DVDD.n16502 DVDD.n16501 0.00122
R17055 DVDD.n17165 DVDD.n17164 0.00122
R17056 DVDD.n17118 DVDD.n17117 0.00122
R17057 DVDD.n17068 DVDD.n17067 0.00122
R17058 DVDD.n15535 DVDD.n11123 0.00122
R17059 DVDD.n16844 DVDD.n16843 0.00122
R17060 DVDD.n16869 DVDD.n16868 0.00122
R17061 DVDD.n17007 DVDD.n17006 0.00122
R17062 DVDD.n17000 DVDD.n16999 0.00122
R17063 DVDD.n16949 DVDD.n16948 0.00122
R17064 DVDD.n16942 DVDD.n16941 0.00122
R17065 DVDD.n16152 DVDD.n16151 0.00122
R17066 DVDD.n16270 DVDD.n16269 0.00122
R17067 DVDD.n16312 DVDD.n16311 0.00122
R17068 DVDD.n16715 DVDD.n16714 0.00122
R17069 DVDD.n16739 DVDD.n16736 0.00122
R17070 DVDD.n16782 DVDD.n16781 0.00122
R17071 DVDD.n16775 DVDD.n16774 0.00122
R17072 DVDD.n16905 DVDD.n16904 0.00122
R17073 DVDD.n16898 DVDD.n16897 0.00122
R17074 DVDD.n16208 DVDD.n16207 0.00122
R17075 DVDD.n15573 DVDD.n15572 0.00122
R17076 DVDD.n16118 DVDD.n15612 0.00122
R17077 DVDD.n16546 DVDD.n16545 0.00122
R17078 DVDD.n16571 DVDD.n16568 0.00122
R17079 DVDD.n16659 DVDD.n16658 0.00122
R17080 DVDD.n16652 DVDD.n16651 0.00122
R17081 DVDD.n16602 DVDD.n16601 0.00122
R17082 DVDD.n16595 DVDD.n16594 0.00122
R17083 DVDD.n15787 DVDD.n15786 0.00122
R17084 DVDD.n15850 DVDD.n15849 0.00122
R17085 DVDD.n16117 DVDD.n15891 0.00122
R17086 DVDD.n16533 DVDD.n16532 0.00122
R17087 DVDD.n16570 DVDD.n16569 0.00122
R17088 DVDD.n16657 DVDD.n16655 0.00122
R17089 DVDD.n16600 DVDD.n16598 0.00122
R17090 DVDD.n16702 DVDD.n16701 0.00122
R17091 DVDD.n16738 DVDD.n16737 0.00122
R17092 DVDD.n16780 DVDD.n16778 0.00122
R17093 DVDD.n16903 DVDD.n16901 0.00122
R17094 DVDD.n16828 DVDD.n16827 0.00122
R17095 DVDD.n16876 DVDD.n16875 0.00122
R17096 DVDD.n17005 DVDD.n17003 0.00122
R17097 DVDD.n16947 DVDD.n16945 0.00122
R17098 DVDD.n16484 DVDD.n16483 0.00122
R17099 DVDD.n17163 DVDD.n17161 0.00122
R17100 DVDD.n11122 DVDD.n11121 0.00122
R17101 DVDD.n3631 DVDD.n3630 0.00122
R17102 DVDD.n20241 DVDD.n20239 0.00122
R17103 DVDD.n7305 DVDD.n7303 0.00122
R17104 DVDD.n1240 DVDD.n1239 0.00120866
R17105 DVDD.n1209 DVDD.n1208 0.00120866
R17106 DVDD.n1204 DVDD.n1203 0.00120866
R17107 DVDD.n1148 DVDD.n1147 0.00120866
R17108 DVDD.n1555 DVDD.n1554 0.00120866
R17109 DVDD.n1614 DVDD.n1613 0.00120866
R17110 DVDD.n1633 DVDD.n1632 0.00120866
R17111 DVDD.n1665 DVDD.n1664 0.00120866
R17112 DVDD.n1658 DVDD.n1657 0.00120866
R17113 DVDD.n1651 DVDD.n1650 0.00120866
R17114 DVDD.n1782 DVDD.n925 0.00120866
R17115 DVDD.n920 DVDD.n919 0.00120866
R17116 DVDD.n913 DVDD.n912 0.00120866
R17117 DVDD.n907 DVDD.n906 0.00120866
R17118 DVDD.n902 DVDD.n901 0.00120866
R17119 DVDD.n889 DVDD.n888 0.00120866
R17120 DVDD.n882 DVDD.n881 0.00120866
R17121 DVDD.n19304 DVDD.n19303 0.00120866
R17122 DVDD.n11471 DVDD.n11470 0.00120866
R17123 DVDD.n12008 DVDD.n12007 0.00120866
R17124 DVDD.n12013 DVDD.n12012 0.00120866
R17125 DVDD.n12046 DVDD.n12045 0.00120866
R17126 DVDD.n12104 DVDD.n12103 0.00120866
R17127 DVDD.n13375 DVDD.n13374 0.00120866
R17128 DVDD.n13380 DVDD.n13379 0.00120866
R17129 DVDD.n18482 DVDD.n18481 0.00120866
R17130 DVDD.n14318 DVDD.n14317 0.00120866
R17131 DVDD.n19689 DVDD.n19688 0.00120866
R17132 DVDD.n19694 DVDD.n19693 0.00120866
R17133 DVDD.n19697 DVDD.n19696 0.00120866
R17134 DVDD.n19756 DVDD.n19755 0.00120866
R17135 DVDD.n19759 DVDD.n19758 0.00120866
R17136 DVDD.n19870 DVDD.n19869 0.00120866
R17137 DVDD.n19909 DVDD.n19908 0.00120866
R17138 DVDD.n20063 DVDD.n20062 0.00120866
R17139 DVDD.n20066 DVDD.n20065 0.00120866
R17140 DVDD.n20072 DVDD.n20071 0.00120866
R17141 DVDD.n20079 DVDD.n20075 0.00120866
R17142 DVDD.n20202 DVDD.n20201 0.00120866
R17143 DVDD.n20101 DVDD.n20100 0.00120866
R17144 DVDD.n19076 DVDD.n19075 0.00120866
R17145 DVDD.n4658 DVDD.n4657 0.00120866
R17146 DVDD.n4660 DVDD.n4659 0.00120866
R17147 DVDD.n4665 DVDD.n4664 0.00120866
R17148 DVDD.n4668 DVDD.n4667 0.00120866
R17149 DVDD.n4804 DVDD.n4803 0.00120866
R17150 DVDD.n4944 DVDD.n4943 0.00120866
R17151 DVDD.n4994 DVDD.n4993 0.00120866
R17152 DVDD.n5096 DVDD.n5095 0.00120866
R17153 DVDD.n5179 DVDD.n5178 0.00120866
R17154 DVDD.n5192 DVDD.n5191 0.00120866
R17155 DVDD.n5337 DVDD.n5336 0.00120866
R17156 DVDD.n5343 DVDD.n5342 0.00120866
R17157 DVDD.n5351 DVDD.n5350 0.00120866
R17158 DVDD.n5381 DVDD.n5380 0.00120866
R17159 DVDD.n5433 DVDD.n5432 0.00120866
R17160 DVDD.n5632 DVDD.n5631 0.00120866
R17161 DVDD.n5633 DVDD.n5632 0.00120866
R17162 DVDD.n1334 DVDD.n1333 0.00120866
R17163 DVDD.n1339 DVDD.n1338 0.00120866
R17164 DVDD.n1342 DVDD.n1341 0.00120866
R17165 DVDD.n1401 DVDD.n1400 0.00120866
R17166 DVDD.n1404 DVDD.n1403 0.00120866
R17167 DVDD.n1506 DVDD.n1505 0.00120866
R17168 DVDD.n1468 DVDD.n1467 0.00120866
R17169 DVDD.n1710 DVDD.n1709 0.00120866
R17170 DVDD.n1707 DVDD.n1706 0.00120866
R17171 DVDD.n1701 DVDD.n1700 0.00120866
R17172 DVDD.n1697 DVDD.n293 0.00120866
R17173 DVDD.n280 DVDD.n279 0.00120866
R17174 DVDD.n19199 DVDD.n19198 0.00120866
R17175 DVDD.n19458 DVDD.n19457 0.00120866
R17176 DVDD.n11365 DVDD.n11364 0.00120866
R17177 DVDD.n11367 DVDD.n11366 0.00120866
R17178 DVDD.n11372 DVDD.n11371 0.00120866
R17179 DVDD.n11375 DVDD.n11374 0.00120866
R17180 DVDD.n11630 DVDD.n11629 0.00120866
R17181 DVDD.n11809 DVDD.n11808 0.00120866
R17182 DVDD.n11759 DVDD.n11758 0.00120866
R17183 DVDD.n11689 DVDD.n11688 0.00120866
R17184 DVDD.n11658 DVDD.n11657 0.00120866
R17185 DVDD.n12359 DVDD.n12358 0.00120866
R17186 DVDD.n12372 DVDD.n12371 0.00120866
R17187 DVDD.n13126 DVDD.n13125 0.00120866
R17188 DVDD.n13122 DVDD.n13121 0.00120866
R17189 DVDD.n13116 DVDD.n13115 0.00120866
R17190 DVDD.n13109 DVDD.n13108 0.00120866
R17191 DVDD.n13080 DVDD.n13079 0.00120866
R17192 DVDD.n13030 DVDD.n13029 0.00120866
R17193 DVDD.n12805 DVDD.n12804 0.00120866
R17194 DVDD.n12804 DVDD.n12803 0.00120866
R17195 DVDD.n19178 DVDD.n19177 0.00120866
R17196 DVDD.n17686 DVDD.n17685 0.00120866
R17197 DVDD.n1911 DVDD.n1910 0.00120866
R17198 DVDD.n1916 DVDD.n1915 0.00120866
R17199 DVDD.n1919 DVDD.n1918 0.00120866
R17200 DVDD.n1978 DVDD.n1977 0.00120866
R17201 DVDD.n1981 DVDD.n1980 0.00120866
R17202 DVDD.n2092 DVDD.n2091 0.00120866
R17203 DVDD.n2130 DVDD.n2129 0.00120866
R17204 DVDD.n2284 DVDD.n2283 0.00120866
R17205 DVDD.n2287 DVDD.n2286 0.00120866
R17206 DVDD.n2293 DVDD.n2292 0.00120866
R17207 DVDD.n2300 DVDD.n2296 0.00120866
R17208 DVDD.n19587 DVDD.n19586 0.00120866
R17209 DVDD.n19486 DVDD.n19485 0.00120866
R17210 DVDD.n18968 DVDD.n18967 0.00120866
R17211 DVDD.n7026 DVDD.n7025 0.00120866
R17212 DVDD.n7024 DVDD.n7023 0.00120866
R17213 DVDD.n7019 DVDD.n7018 0.00120866
R17214 DVDD.n7016 DVDD.n7015 0.00120866
R17215 DVDD.n6880 DVDD.n6879 0.00120866
R17216 DVDD.n6740 DVDD.n6739 0.00120866
R17217 DVDD.n6690 DVDD.n6689 0.00120866
R17218 DVDD.n6617 DVDD.n6616 0.00120866
R17219 DVDD.n6586 DVDD.n6585 0.00120866
R17220 DVDD.n6503 DVDD.n6502 0.00120866
R17221 DVDD.n6490 DVDD.n6489 0.00120866
R17222 DVDD.n6428 DVDD.n6427 0.00120866
R17223 DVDD.n6424 DVDD.n6423 0.00120866
R17224 DVDD.n6418 DVDD.n6417 0.00120866
R17225 DVDD.n6410 DVDD.n6409 0.00120866
R17226 DVDD.n6380 DVDD.n6379 0.00120866
R17227 DVDD.n6328 DVDD.n6327 0.00120866
R17228 DVDD.n6185 DVDD.n6184 0.00120866
R17229 DVDD.n6184 DVDD.n6183 0.00120866
R17230 DVDD.n3269 DVDD.n3268 0.00120866
R17231 DVDD.n3264 DVDD.n3263 0.00120866
R17232 DVDD.n3261 DVDD.n3260 0.00120866
R17233 DVDD.n3202 DVDD.n3201 0.00120866
R17234 DVDD.n3199 DVDD.n3198 0.00120866
R17235 DVDD.n3491 DVDD.n3490 0.00120866
R17236 DVDD.n3529 DVDD.n3528 0.00120866
R17237 DVDD.n3728 DVDD.n3727 0.00120866
R17238 DVDD.n3731 DVDD.n3730 0.00120866
R17239 DVDD.n3737 DVDD.n3736 0.00120866
R17240 DVDD.n3779 DVDD.n3740 0.00120866
R17241 DVDD.n3766 DVDD.n3765 0.00120866
R17242 DVDD.n18503 DVDD.n18502 0.00120866
R17243 DVDD.n18805 DVDD.n18804 0.00120866
R17244 DVDD.n10043 DVDD.n10042 0.00120866
R17245 DVDD.n10041 DVDD.n10040 0.00120866
R17246 DVDD.n10036 DVDD.n10035 0.00120866
R17247 DVDD.n10033 DVDD.n10032 0.00120866
R17248 DVDD.n7886 DVDD.n7885 0.00120866
R17249 DVDD.n9708 DVDD.n9707 0.00120866
R17250 DVDD.n9658 DVDD.n9657 0.00120866
R17251 DVDD.n9585 DVDD.n9584 0.00120866
R17252 DVDD.n9554 DVDD.n9553 0.00120866
R17253 DVDD.n8380 DVDD.n8379 0.00120866
R17254 DVDD.n8393 DVDD.n8392 0.00120866
R17255 DVDD.n9214 DVDD.n9213 0.00120866
R17256 DVDD.n9210 DVDD.n9209 0.00120866
R17257 DVDD.n9204 DVDD.n9203 0.00120866
R17258 DVDD.n9196 DVDD.n9195 0.00120866
R17259 DVDD.n9166 DVDD.n9165 0.00120866
R17260 DVDD.n9114 DVDD.n9113 0.00120866
R17261 DVDD.n8887 DVDD.n8886 0.00120866
R17262 DVDD.n8886 DVDD.n8885 0.00120866
R17263 DVDD.n2345 DVDD.n2344 0.00120714
R17264 DVDD.n2456 DVDD.n2455 0.00120714
R17265 DVDD.n730 DVDD.n729 0.00120714
R17266 DVDD.n2521 DVDD.n2520 0.00120714
R17267 DVDD.n2543 DVDD.n2542 0.00120714
R17268 DVDD.n2595 DVDD.n2594 0.00120714
R17269 DVDD.n2654 DVDD.n2653 0.00120714
R17270 DVDD.n2693 DVDD.n2692 0.00120714
R17271 DVDD.n4148 DVDD.n4147 0.00120714
R17272 DVDD.n8531 DVDD.n8530 0.00120714
R17273 DVDD.n13863 DVDD.n13862 0.00120714
R17274 DVDD.n11223 DVDD.n11222 0.00120714
R17275 DVDD.n17179 DVDD.n17176 0.0011923
R17276 DVDD.n17702 DVDD.n17699 0.0011923
R17277 DVDD.n17699 DVDD.n17698 0.0011923
R17278 DVDD.n17176 DVDD.n17175 0.0011923
R17279 DVDD.n18870 DVDD.n18869 0.00119
R17280 DVDD.n19119 DVDD.n19118 0.00119
R17281 DVDD.n16043 DVDD.n16042 0.00118828
R17282 DVDD.n16007 DVDD.n16006 0.00118828
R17283 DVDD.n16008 DVDD.n16007 0.00118828
R17284 DVDD.n16044 DVDD.n16043 0.00118828
R17285 DVDD.n15655 DVDD.n15654 0.00118828
R17286 DVDD.n15925 DVDD.n15924 0.00118828
R17287 DVDD.n15924 DVDD.n15923 0.00118828
R17288 DVDD.n15656 DVDD.n15655 0.00118828
R17289 DVDD.n8290 DVDD.n8289 0.00118828
R17290 DVDD.n8282 DVDD.n8281 0.00118828
R17291 DVDD.n8274 DVDD.n8273 0.00118828
R17292 DVDD.n8267 DVDD.n8266 0.00118828
R17293 DVDD.n8261 DVDD.n8260 0.00118828
R17294 DVDD.n8254 DVDD.n8253 0.00118828
R17295 DVDD.n8245 DVDD.n8244 0.00118828
R17296 DVDD.n8236 DVDD.n8235 0.00118828
R17297 DVDD.n8227 DVDD.n8226 0.00118828
R17298 DVDD.n8219 DVDD.n8218 0.00118828
R17299 DVDD.n8211 DVDD.n8210 0.00118828
R17300 DVDD.n8204 DVDD.n8203 0.00118828
R17301 DVDD.n8198 DVDD.n8197 0.00118828
R17302 DVDD.n8191 DVDD.n8190 0.00118828
R17303 DVDD.n8183 DVDD.n8182 0.00118828
R17304 DVDD.n8172 DVDD.n8171 0.00118828
R17305 DVDD.n8158 DVDD.n8157 0.00118828
R17306 DVDD.n8159 DVDD.n8158 0.00118828
R17307 DVDD.n8192 DVDD.n8191 0.00118828
R17308 DVDD.n8205 DVDD.n8204 0.00118828
R17309 DVDD.n8268 DVDD.n8267 0.00118828
R17310 DVDD.n8262 DVDD.n8261 0.00118828
R17311 DVDD.n8255 DVDD.n8254 0.00118828
R17312 DVDD.n8246 DVDD.n8245 0.00118828
R17313 DVDD.n8237 DVDD.n8236 0.00118828
R17314 DVDD.n8199 DVDD.n8198 0.00118828
R17315 DVDD.n8182 DVDD.n8181 0.00118828
R17316 DVDD.n8173 DVDD.n8172 0.00118828
R17317 DVDD.n8353 DVDD.n8352 0.00118828
R17318 DVDD.n8344 DVDD.n8343 0.00118828
R17319 DVDD.n8338 DVDD.n8337 0.00118828
R17320 DVDD.n8331 DVDD.n8330 0.00118828
R17321 DVDD.n8301 DVDD.n8300 0.00118828
R17322 DVDD.n8345 DVDD.n8344 0.00118828
R17323 DVDD.n8332 DVDD.n8331 0.00118828
R17324 DVDD.n8325 DVDD.n8324 0.00118828
R17325 DVDD.n8317 DVDD.n8316 0.00118828
R17326 DVDD.n8309 DVDD.n8308 0.00118828
R17327 DVDD.n8302 DVDD.n8301 0.00118828
R17328 DVDD.n8337 DVDD.n8336 0.00118828
R17329 DVDD.n8354 DVDD.n8353 0.00118828
R17330 DVDD.n7990 DVDD.n7989 0.00118828
R17331 DVDD.n8069 DVDD.n8068 0.00118828
R17332 DVDD.n7989 DVDD.n7988 0.00118828
R17333 DVDD.n10331 DVDD.n10330 0.00117999
R17334 DVDD.n10332 DVDD.n10331 0.00117999
R17335 DVDD.n16490 DVDD.n16489 0.00117999
R17336 DVDD.n16491 DVDD.n16490 0.00117999
R17337 DVDD.n16834 DVDD.n16833 0.00117999
R17338 DVDD.n16860 DVDD.n16859 0.00117999
R17339 DVDD.n16835 DVDD.n16834 0.00117999
R17340 DVDD.n16861 DVDD.n16860 0.00117999
R17341 DVDD.n1579 DVDD.n1578 0.00117716
R17342 DVDD.n12126 DVDD.n12125 0.00117716
R17343 DVDD.n13312 DVDD.n13311 0.00117716
R17344 DVDD.n13321 DVDD.n13320 0.00117716
R17345 DVDD.n13327 DVDD.n13326 0.00117716
R17346 DVDD.n13334 DVDD.n13333 0.00117716
R17347 DVDD.n13341 DVDD.n13340 0.00117716
R17348 DVDD.n13350 DVDD.n13349 0.00117716
R17349 DVDD.n13359 DVDD.n13358 0.00117716
R17350 DVDD.n13367 DVDD.n13366 0.00117716
R17351 DVDD.n13379 DVDD.n13378 0.00117716
R17352 DVDD.n13388 DVDD.n13387 0.00117716
R17353 DVDD.n13397 DVDD.n13396 0.00117716
R17354 DVDD.n13404 DVDD.n13403 0.00117716
R17355 DVDD.n13410 DVDD.n13409 0.00117716
R17356 DVDD.n13417 DVDD.n13416 0.00117716
R17357 DVDD.n13426 DVDD.n13425 0.00117716
R17358 DVDD.n13435 DVDD.n13434 0.00117716
R17359 DVDD.n13445 DVDD.n13444 0.00117716
R17360 DVDD.n13454 DVDD.n13453 0.00117716
R17361 DVDD.n13463 DVDD.n13462 0.00117716
R17362 DVDD.n13470 DVDD.n13469 0.00117716
R17363 DVDD.n13476 DVDD.n13475 0.00117716
R17364 DVDD.n13483 DVDD.n13482 0.00117716
R17365 DVDD.n13492 DVDD.n13491 0.00117716
R17366 DVDD.n13502 DVDD.n13501 0.00117716
R17367 DVDD.n13514 DVDD.n13513 0.00117716
R17368 DVDD.n13566 DVDD.n13565 0.00117716
R17369 DVDD.n13599 DVDD.n13598 0.00117716
R17370 DVDD.n13647 DVDD.n13646 0.00117716
R17371 DVDD.n13680 DVDD.n13679 0.00117716
R17372 DVDD.n12044 DVDD.n12043 0.00117716
R17373 DVDD.n12125 DVDD.n12124 0.00117716
R17374 DVDD.n13311 DVDD.n13310 0.00117716
R17375 DVDD.n13320 DVDD.n13319 0.00117716
R17376 DVDD.n13333 DVDD.n13332 0.00117716
R17377 DVDD.n13340 DVDD.n13339 0.00117716
R17378 DVDD.n13349 DVDD.n13348 0.00117716
R17379 DVDD.n13358 DVDD.n13357 0.00117716
R17380 DVDD.n13366 DVDD.n13365 0.00117716
R17381 DVDD.n13328 DVDD.n13327 0.00117716
R17382 DVDD.n13513 DVDD.n13512 0.00117716
R17383 DVDD.n13482 DVDD.n13481 0.00117716
R17384 DVDD.n13469 DVDD.n13468 0.00117716
R17385 DVDD.n13453 DVDD.n13452 0.00117716
R17386 DVDD.n13378 DVDD.n13377 0.00117716
R17387 DVDD.n13387 DVDD.n13386 0.00117716
R17388 DVDD.n13396 DVDD.n13395 0.00117716
R17389 DVDD.n13403 DVDD.n13402 0.00117716
R17390 DVDD.n13409 DVDD.n13408 0.00117716
R17391 DVDD.n13416 DVDD.n13415 0.00117716
R17392 DVDD.n13425 DVDD.n13424 0.00117716
R17393 DVDD.n13434 DVDD.n13433 0.00117716
R17394 DVDD.n13444 DVDD.n13443 0.00117716
R17395 DVDD.n13462 DVDD.n13461 0.00117716
R17396 DVDD.n13475 DVDD.n13474 0.00117716
R17397 DVDD.n13491 DVDD.n13490 0.00117716
R17398 DVDD.n13501 DVDD.n13500 0.00117716
R17399 DVDD.n13598 DVDD.n13597 0.00117716
R17400 DVDD.n13565 DVDD.n13564 0.00117716
R17401 DVDD.n13679 DVDD.n13678 0.00117716
R17402 DVDD.n13646 DVDD.n13645 0.00117716
R17403 DVDD.n15413 DVDD.n15412 0.00117716
R17404 DVDD.n15449 DVDD.n15448 0.00117716
R17405 DVDD.n14690 DVDD.n14689 0.00117716
R17406 DVDD.n14607 DVDD.n14606 0.00117716
R17407 DVDD.n14553 DVDD.n14552 0.00117716
R17408 DVDD.n14517 DVDD.n14516 0.00117716
R17409 DVDD.n14465 DVDD.n14464 0.00117716
R17410 DVDD.n14413 DVDD.n14412 0.00117716
R17411 DVDD.n14414 DVDD.n14413 0.00117716
R17412 DVDD.n14518 DVDD.n14517 0.00117716
R17413 DVDD.n14608 DVDD.n14607 0.00117716
R17414 DVDD.n14691 DVDD.n14690 0.00117716
R17415 DVDD.n15448 DVDD.n15447 0.00117716
R17416 DVDD.n15412 DVDD.n15411 0.00117716
R17417 DVDD.n14554 DVDD.n14553 0.00117716
R17418 DVDD.n14466 DVDD.n14465 0.00117716
R17419 DVDD.n19723 DVDD.n19722 0.00117716
R17420 DVDD.n4915 DVDD.n4914 0.00117716
R17421 DVDD.n4985 DVDD.n4984 0.00117716
R17422 DVDD.n5322 DVDD.n5321 0.00117716
R17423 DVDD.n5480 DVDD.n5479 0.00117716
R17424 DVDD.n5603 DVDD.n5602 0.00117716
R17425 DVDD.n5609 DVDD.n5608 0.00117716
R17426 DVDD.n5683 DVDD.n5682 0.00117716
R17427 DVDD.n6033 DVDD.n6032 0.00117716
R17428 DVDD.n5971 DVDD.n5970 0.00117716
R17429 DVDD.n5865 DVDD.n5864 0.00117716
R17430 DVDD.n5848 DVDD.n5847 0.00117716
R17431 DVDD.n5831 DVDD.n5830 0.00117716
R17432 DVDD.n5608 DVDD.n5607 0.00117716
R17433 DVDD.n5972 DVDD.n5971 0.00117716
R17434 DVDD.n5479 DVDD.n5478 0.00117716
R17435 DVDD.n5321 DVDD.n5320 0.00117716
R17436 DVDD.n4914 DVDD.n4913 0.00117716
R17437 DVDD.n4984 DVDD.n4983 0.00117716
R17438 DVDD.n5682 DVDD.n5681 0.00117716
R17439 DVDD.n5602 DVDD.n5601 0.00117716
R17440 DVDD.n6034 DVDD.n6033 0.00117716
R17441 DVDD.n11838 DVDD.n11837 0.00117716
R17442 DVDD.n11768 DVDD.n11767 0.00117716
R17443 DVDD.n13137 DVDD.n13136 0.00117716
R17444 DVDD.n12983 DVDD.n12982 0.00117716
R17445 DVDD.n12824 DVDD.n12823 0.00117716
R17446 DVDD.n12818 DVDD.n12817 0.00117716
R17447 DVDD.n12758 DVDD.n12757 0.00117716
R17448 DVDD.n12684 DVDD.n12683 0.00117716
R17449 DVDD.n12634 DVDD.n12633 0.00117716
R17450 DVDD.n12564 DVDD.n12563 0.00117716
R17451 DVDD.n12546 DVDD.n12545 0.00117716
R17452 DVDD.n12529 DVDD.n12528 0.00117716
R17453 DVDD.n12984 DVDD.n12983 0.00117716
R17454 DVDD.n11769 DVDD.n11768 0.00117716
R17455 DVDD.n11839 DVDD.n11838 0.00117716
R17456 DVDD.n1368 DVDD.n1367 0.00117716
R17457 DVDD.n12635 DVDD.n12634 0.00117716
R17458 DVDD.n12759 DVDD.n12758 0.00117716
R17459 DVDD.n12819 DVDD.n12818 0.00117716
R17460 DVDD.n12825 DVDD.n12824 0.00117716
R17461 DVDD.n12685 DVDD.n12684 0.00117716
R17462 DVDD.n18189 DVDD.n18188 0.00117716
R17463 DVDD.n18156 DVDD.n18155 0.00117716
R17464 DVDD.n18045 DVDD.n18044 0.00117716
R17465 DVDD.n17967 DVDD.n17966 0.00117716
R17466 DVDD.n17915 DVDD.n17914 0.00117716
R17467 DVDD.n17882 DVDD.n17881 0.00117716
R17468 DVDD.n17834 DVDD.n17833 0.00117716
R17469 DVDD.n17787 DVDD.n17786 0.00117716
R17470 DVDD.n17788 DVDD.n17787 0.00117716
R17471 DVDD.n17968 DVDD.n17967 0.00117716
R17472 DVDD.n18157 DVDD.n18156 0.00117716
R17473 DVDD.n18190 DVDD.n18189 0.00117716
R17474 DVDD.n18046 DVDD.n18045 0.00117716
R17475 DVDD.n17883 DVDD.n17882 0.00117716
R17476 DVDD.n17916 DVDD.n17915 0.00117716
R17477 DVDD.n17835 DVDD.n17834 0.00117716
R17478 DVDD.n5849 DVDD.n5848 0.00117716
R17479 DVDD.n12547 DVDD.n12546 0.00117716
R17480 DVDD.n5832 DVDD.n5831 0.00117716
R17481 DVDD.n12530 DVDD.n12529 0.00117716
R17482 DVDD.n5866 DVDD.n5865 0.00117716
R17483 DVDD.n12563 DVDD.n12562 0.00117716
R17484 DVDD.n6769 DVDD.n6768 0.00117716
R17485 DVDD.n6699 DVDD.n6698 0.00117716
R17486 DVDD.n6439 DVDD.n6438 0.00117716
R17487 DVDD.n6279 DVDD.n6278 0.00117716
R17488 DVDD.n6202 DVDD.n6201 0.00117716
R17489 DVDD.n6142 DVDD.n6141 0.00117716
R17490 DVDD.n4484 DVDD.n4483 0.00117716
R17491 DVDD.n4434 DVDD.n4433 0.00117716
R17492 DVDD.n4323 DVDD.n4322 0.00117716
R17493 DVDD.n4294 DVDD.n4293 0.00117716
R17494 DVDD.n4269 DVDD.n4268 0.00117716
R17495 DVDD.n4270 DVDD.n4269 0.00117716
R17496 DVDD.n4295 DVDD.n4294 0.00117716
R17497 DVDD.n4324 DVDD.n4323 0.00117716
R17498 DVDD.n4435 DVDD.n4434 0.00117716
R17499 DVDD.n6280 DVDD.n6279 0.00117716
R17500 DVDD.n6440 DVDD.n6439 0.00117716
R17501 DVDD.n6770 DVDD.n6769 0.00117716
R17502 DVDD.n6700 DVDD.n6699 0.00117716
R17503 DVDD.n1945 DVDD.n1944 0.00117716
R17504 DVDD.n6197 DVDD.n6196 0.00117716
R17505 DVDD.n6143 DVDD.n6142 0.00117716
R17506 DVDD.n6203 DVDD.n6202 0.00117716
R17507 DVDD.n4485 DVDD.n4484 0.00117716
R17508 DVDD.n9737 DVDD.n9736 0.00117716
R17509 DVDD.n9667 DVDD.n9666 0.00117716
R17510 DVDD.n9225 DVDD.n9224 0.00117716
R17511 DVDD.n9065 DVDD.n9064 0.00117716
R17512 DVDD.n8904 DVDD.n8903 0.00117716
R17513 DVDD.n8844 DVDD.n8843 0.00117716
R17514 DVDD.n8770 DVDD.n8769 0.00117716
R17515 DVDD.n8708 DVDD.n8707 0.00117716
R17516 DVDD.n8607 DVDD.n8606 0.00117716
R17517 DVDD.n8590 DVDD.n8589 0.00117716
R17518 DVDD.n8573 DVDD.n8572 0.00117716
R17519 DVDD.n9668 DVDD.n9667 0.00117716
R17520 DVDD.n8899 DVDD.n8898 0.00117716
R17521 DVDD.n8709 DVDD.n8708 0.00117716
R17522 DVDD.n8608 DVDD.n8607 0.00117716
R17523 DVDD.n8591 DVDD.n8590 0.00117716
R17524 DVDD.n8574 DVDD.n8573 0.00117716
R17525 DVDD.n9066 DVDD.n9065 0.00117716
R17526 DVDD.n9226 DVDD.n9225 0.00117716
R17527 DVDD.n9738 DVDD.n9737 0.00117716
R17528 DVDD.n3235 DVDD.n3234 0.00117716
R17529 DVDD.n8845 DVDD.n8844 0.00117716
R17530 DVDD.n8905 DVDD.n8904 0.00117716
R17531 DVDD.n8771 DVDD.n8770 0.00117716
R17532 DVDD.n18833 DVDD.n18832 0.001175
R17533 DVDD.n18817 DVDD.n18816 0.001175
R17534 DVDD.n19163 DVDD.n19162 0.001175
R17535 DVDD.n19151 DVDD.n19150 0.001175
R17536 DVDD.n7272 DVDD.n7271 0.001175
R17537 DVDD.n3844 DVDD.n3843 0.001175
R17538 DVDD.n7612 DVDD.n7611 0.001175
R17539 DVDD.n3896 DVDD.n3895 0.001175
R17540 DVDD.n3910 DVDD.n3909 0.001175
R17541 DVDD.n7639 DVDD.n7638 0.001175
R17542 DVDD.n129 DVDD.n128 0.001175
R17543 DVDD.n3785 DVDD.n3784 0.001175
R17544 DVDD.n3799 DVDD.n3798 0.001175
R17545 DVDD.n20280 DVDD.n20279 0.001175
R17546 DVDD.n20327 DVDD.n20326 0.001175
R17547 DVDD.n14881 DVDD.n14880 0.001175
R17548 DVDD.n14865 DVDD.n14864 0.001175
R17549 DVDD.n15097 DVDD.n15096 0.001175
R17550 DVDD.n10715 DVDD.n10714 0.001175
R17551 DVDD.n10625 DVDD.n10624 0.001175
R17552 DVDD.n10613 DVDD.n10612 0.001175
R17553 DVDD.n10408 DVDD.n10407 0.001175
R17554 DVDD.n10583 DVDD.n10582 0.001175
R17555 DVDD.n10642 DVDD.n10641 0.001175
R17556 DVDD.n7285 DVDD.n7284 0.001175
R17557 DVDD.n15194 DVDD.n15193 0.00117236
R17558 DVDD.n15263 DVDD.n15262 0.00117236
R17559 DVDD.n15281 DVDD.n15280 0.00117236
R17560 DVDD.n14979 DVDD.n14978 0.00116499
R17561 DVDD.n15378 DVDD.n15377 0.00116499
R17562 DVDD.n15338 DVDD.n15337 0.00116499
R17563 DVDD.n15731 DVDD.n15730 0.00116499
R17564 DVDD.n15703 DVDD.n15702 0.00116499
R17565 DVDD.n15809 DVDD.n15808 0.00116499
R17566 DVDD.n15872 DVDD.n15871 0.00116499
R17567 DVDD.n16090 DVDD.n16089 0.00116499
R17568 DVDD.n16091 DVDD.n16090 0.00116499
R17569 DVDD.n15732 DVDD.n15731 0.00116499
R17570 DVDD.n15379 DVDD.n15378 0.00116499
R17571 DVDD.n15808 DVDD.n15807 0.00116499
R17572 DVDD.n14978 DVDD.n14977 0.00116499
R17573 DVDD.n15702 DVDD.n15701 0.00116499
R17574 DVDD.n15337 DVDD.n15336 0.00116499
R17575 DVDD.n15871 DVDD.n15870 0.00116499
R17576 DVDD.n19465 DVDD.n19464 0.00116
R17577 DVDD.n18894 DVDD.n18893 0.00116
R17578 DVDD.n18891 DVDD.n18890 0.00116
R17579 DVDD.n18846 DVDD.n18845 0.00116
R17580 DVDD.n19143 DVDD.n19142 0.00116
R17581 DVDD.n19140 DVDD.n19139 0.00116
R17582 DVDD.n19094 DVDD.n19093 0.00116
R17583 DVDD.n15 DVDD.n14 0.00116
R17584 DVDD.n7397 DVDD.n7396 0.00116
R17585 DVDD.n97 DVDD.n96 0.00116
R17586 DVDD.n7445 DVDD.n7444 0.00116
R17587 DVDD.n43 DVDD.n42 0.00116
R17588 DVDD.n7506 DVDD.n7505 0.00116
R17589 DVDD.n19371 DVDD.n19370 0.00116
R17590 DVDD.n16160 DVDD.n16159 0.00116
R17591 DVDD.n16163 DVDD.n16162 0.00116
R17592 DVDD.n16278 DVDD.n16277 0.00116
R17593 DVDD.n16281 DVDD.n16280 0.00116
R17594 DVDD.n16216 DVDD.n16215 0.00116
R17595 DVDD.n16219 DVDD.n16218 0.00116
R17596 DVDD.n15581 DVDD.n15580 0.00116
R17597 DVDD.n15584 DVDD.n15583 0.00116
R17598 DVDD.n15795 DVDD.n15794 0.00116
R17599 DVDD.n15799 DVDD.n15798 0.00116
R17600 DVDD.n15858 DVDD.n15857 0.00116
R17601 DVDD.n15862 DVDD.n15861 0.00116
R17602 DVDD.n18367 DVDD.n18366 0.00116
R17603 DVDD.n20233 DVDD.n20232 0.00116
R17604 DVDD.n7313 DVDD.n7312 0.00116
R17605 DVDD.n4155 DVDD.n4150 0.00114286
R17606 DVDD.n8537 DVDD.n8533 0.00114286
R17607 DVDD.n13869 DVDD.n13865 0.00114286
R17608 DVDD.n13834 DVDD.n11221 0.00114286
R17609 DVDD.n2341 DVDD.n2340 0.00114286
R17610 DVDD.n2392 DVDD.n2391 0.00114286
R17611 DVDD.n2497 DVDD.n2453 0.00114286
R17612 DVDD.n433 DVDD.n432 0.00114286
R17613 DVDD.n2342 DVDD.n2338 0.00114286
R17614 DVDD.n2393 DVDD.n2389 0.00114286
R17615 DVDD.n2499 DVDD.n2498 0.00114286
R17616 DVDD.n2539 DVDD.n2538 0.00114286
R17617 DVDD.n2590 DVDD.n2589 0.00114286
R17618 DVDD.n2709 DVDD.n2649 0.00114286
R17619 DVDD.n2696 DVDD.n2652 0.00114286
R17620 DVDD.n665 DVDD.n664 0.00114286
R17621 DVDD.n2540 DVDD.n2536 0.00114286
R17622 DVDD.n2591 DVDD.n2587 0.00114286
R17623 DVDD.n2594 DVDD.n2593 0.00114286
R17624 DVDD.n2711 DVDD.n2710 0.00114286
R17625 DVDD.n2695 DVDD.n2688 0.00114286
R17626 DVDD.n4157 DVDD.n4156 0.00114286
R17627 DVDD.n8539 DVDD.n8538 0.00114286
R17628 DVDD.n13871 DVDD.n13870 0.00114286
R17629 DVDD.n13836 DVDD.n13835 0.00114286
R17630 DVDD.n16466 DVDD.n16465 0.00114
R17631 DVDD.n10837 DVDD.n10812 0.00114
R17632 DVDD.n10805 DVDD.n10780 0.00114
R17633 DVDD.n10769 DVDD.n10744 0.00114
R17634 DVDD.n10318 DVDD.n10317 0.00114
R17635 DVDD.n3681 DVDD.n3680 0.00113
R17636 DVDD.n3712 DVDD.n3711 0.00113
R17637 DVDD.n18558 DVDD.n18557 0.00113
R17638 DVDD.n2942 DVDD.n2941 0.00113
R17639 DVDD.n7819 DVDD.n7818 0.00113
R17640 DVDD.n9810 DVDD.n9809 0.00113
R17641 DVDD.n9812 DVDD.n9811 0.00113
R17642 DVDD.n9881 DVDD.n9880 0.00113
R17643 DVDD.n9878 DVDD.n9877 0.00113
R17644 DVDD.n9875 DVDD.n9874 0.00113
R17645 DVDD.n9872 DVDD.n9871 0.00113
R17646 DVDD.n9869 DVDD.n9868 0.00113
R17647 DVDD.n9866 DVDD.n9865 0.00113
R17648 DVDD.n9863 DVDD.n9862 0.00113
R17649 DVDD.n9860 DVDD.n9859 0.00113
R17650 DVDD.n9857 DVDD.n9856 0.00113
R17651 DVDD.n9854 DVDD.n9853 0.00113
R17652 DVDD.n9851 DVDD.n9850 0.00113
R17653 DVDD.n9848 DVDD.n9847 0.00113
R17654 DVDD.n9845 DVDD.n9844 0.00113
R17655 DVDD.n9842 DVDD.n9841 0.00113
R17656 DVDD.n9839 DVDD.n9838 0.00113
R17657 DVDD.n9836 DVDD.n9835 0.00113
R17658 DVDD.n9833 DVDD.n9832 0.00113
R17659 DVDD.n9830 DVDD.n9829 0.00113
R17660 DVDD.n9827 DVDD.n9826 0.00113
R17661 DVDD.n9824 DVDD.n9823 0.00113
R17662 DVDD.n9390 DVDD.n9389 0.00113
R17663 DVDD.n2180 DVDD.n2179 0.00113
R17664 DVDD.n2237 DVDD.n2236 0.00113
R17665 DVDD.n2268 DVDD.n2267 0.00113
R17666 DVDD.n18927 DVDD.n18926 0.00113
R17667 DVDD.n6788 DVDD.n6787 0.00113
R17668 DVDD.n6805 DVDD.n6804 0.00113
R17669 DVDD.n6803 DVDD.n6802 0.00113
R17670 DVDD.n1882 DVDD.n1881 0.00113
R17671 DVDD.n1877 DVDD.n1876 0.00113
R17672 DVDD.n19959 DVDD.n19958 0.00113
R17673 DVDD.n20016 DVDD.n20015 0.00113
R17674 DVDD.n20047 DVDD.n20046 0.00113
R17675 DVDD.n19045 DVDD.n19044 0.00113
R17676 DVDD.n4825 DVDD.n4824 0.00113
R17677 DVDD.n4842 DVDD.n4841 0.00113
R17678 DVDD.n4840 DVDD.n4839 0.00113
R17679 DVDD.n19660 DVDD.n19659 0.00113
R17680 DVDD.n19655 DVDD.n19654 0.00113
R17681 DVDD.n986 DVDD.n985 0.00113
R17682 DVDD.n1726 DVDD.n1725 0.00113
R17683 DVDD.n955 DVDD.n954 0.00113
R17684 DVDD.n19254 DVDD.n19253 0.00113
R17685 DVDD.n1829 DVDD.n1828 0.00113
R17686 DVDD.n1850 DVDD.n1849 0.00113
R17687 DVDD.n1853 DVDD.n1852 0.00113
R17688 DVDD.n19533 DVDD.n19532 0.00113
R17689 DVDD.n18849 DVDD.n18848 0.00113
R17690 DVDD.n18836 DVDD.n18835 0.00113
R17691 DVDD.n19607 DVDD.n19606 0.00113
R17692 DVDD.n19628 DVDD.n19627 0.00113
R17693 DVDD.n19631 DVDD.n19630 0.00113
R17694 DVDD.n20148 DVDD.n20147 0.00113
R17695 DVDD.n19097 DVDD.n19096 0.00113
R17696 DVDD.n19084 DVDD.n19083 0.00113
R17697 DVDD.n7367 DVDD.n7366 0.00113
R17698 DVDD.n7417 DVDD.n7415 0.00113
R17699 DVDD.n73 DVDD.n72 0.00113
R17700 DVDD.n7465 DVDD.n7463 0.00113
R17701 DVDD.n7240 DVDD.n7239 0.00113
R17702 DVDD.n7486 DVDD.n7484 0.00113
R17703 DVDD.n200 DVDD.n199 0.00113
R17704 DVDD.n19374 DVDD.n19373 0.00113
R17705 DVDD.n19359 DVDD.n19358 0.00113
R17706 DVDD.n11344 DVDD.n11343 0.00113
R17707 DVDD.n11911 DVDD.n11910 0.00113
R17708 DVDD.n11913 DVDD.n11912 0.00113
R17709 DVDD.n11982 DVDD.n11981 0.00113
R17710 DVDD.n11979 DVDD.n11978 0.00113
R17711 DVDD.n11976 DVDD.n11975 0.00113
R17712 DVDD.n11973 DVDD.n11972 0.00113
R17713 DVDD.n11970 DVDD.n11969 0.00113
R17714 DVDD.n11967 DVDD.n11966 0.00113
R17715 DVDD.n11964 DVDD.n11963 0.00113
R17716 DVDD.n11961 DVDD.n11960 0.00113
R17717 DVDD.n11958 DVDD.n11957 0.00113
R17718 DVDD.n11955 DVDD.n11954 0.00113
R17719 DVDD.n11952 DVDD.n11951 0.00113
R17720 DVDD.n11949 DVDD.n11948 0.00113
R17721 DVDD.n11946 DVDD.n11945 0.00113
R17722 DVDD.n11943 DVDD.n11942 0.00113
R17723 DVDD.n11940 DVDD.n11939 0.00113
R17724 DVDD.n11937 DVDD.n11936 0.00113
R17725 DVDD.n11934 DVDD.n11933 0.00113
R17726 DVDD.n11931 DVDD.n11930 0.00113
R17727 DVDD.n11928 DVDD.n11927 0.00113
R17728 DVDD.n11925 DVDD.n11924 0.00113
R17729 DVDD.n1305 DVDD.n1304 0.00113
R17730 DVDD.n1300 DVDD.n1299 0.00113
R17731 DVDD.n13301 DVDD.n13300 0.00113
R17732 DVDD.n17011 DVDD.n17010 0.00113
R17733 DVDD.n17008 DVDD.n17007 0.00113
R17734 DVDD.n16953 DVDD.n16952 0.00113
R17735 DVDD.n16950 DVDD.n16949 0.00113
R17736 DVDD.n16786 DVDD.n16785 0.00113
R17737 DVDD.n16783 DVDD.n16782 0.00113
R17738 DVDD.n16909 DVDD.n16908 0.00113
R17739 DVDD.n16906 DVDD.n16905 0.00113
R17740 DVDD.n16664 DVDD.n16663 0.00113
R17741 DVDD.n16660 DVDD.n16659 0.00113
R17742 DVDD.n16607 DVDD.n16606 0.00113
R17743 DVDD.n16603 DVDD.n16602 0.00113
R17744 DVDD.n3298 DVDD.n3297 0.00113
R17745 DVDD.n3303 DVDD.n3302 0.00113
R17746 DVDD.n18653 DVDD.n18652 0.00113
R17747 DVDD.n18370 DVDD.n18369 0.00113
R17748 DVDD.n18338 DVDD.n18337 0.00113
R17749 DVDD.n20263 DVDD.n20262 0.00113
R17750 DVDD.n7333 DVDD.n7331 0.00113
R17751 DVDD.n3828 DVDD.n3827 0.00112572
R17752 DVDD.n113 DVDD.n112 0.00112572
R17753 DVDD.n14915 DVDD.n14914 0.00111875
R17754 DVDD.n14929 DVDD.n14928 0.00111875
R17755 DVDD.n14893 DVDD.n14892 0.00111875
R17756 DVDD.n15227 DVDD.n15226 0.00111875
R17757 DVDD.n10641 DVDD.n10640 0.00111875
R17758 DVDD.n11154 DVDD.n11153 0.001105
R17759 DVDD.n11151 DVDD.n11150 0.001105
R17760 DVDD.n11155 DVDD.n11154 0.001105
R17761 DVDD.n11150 DVDD.n11149 0.001105
R17762 DVDD.n3060 DVDD.n3059 0.00110268
R17763 DVDD.n3059 DVDD.n3058 0.00110268
R17764 DVDD.n19531 DVDD.n19530 0.0011
R17765 DVDD.n19527 DVDD.n19526 0.0011
R17766 DVDD.n19508 DVDD.n19507 0.0011
R17767 DVDD.n18333 DVDD.n7077 0.0011
R17768 DVDD.n7580 DVDD.n7579 0.0011
R17769 DVDD.n20146 DVDD.n20145 0.0011
R17770 DVDD.n20142 DVDD.n20141 0.0011
R17771 DVDD.n20123 DVDD.n20122 0.0011
R17772 DVDD.n18333 DVDD.n3889 0.0011
R17773 DVDD.n7536 DVDD.n7535 0.0011
R17774 DVDD.n7355 DVDD.n7354 0.0011
R17775 DVDD.n7371 DVDD.n7369 0.0011
R17776 DVDD.n7594 DVDD.n7593 0.0011
R17777 DVDD.n85 DVDD.n84 0.0011
R17778 DVDD.n69 DVDD.n67 0.0011
R17779 DVDD.n7550 DVDD.n7549 0.0011
R17780 DVDD.n7228 DVDD.n7227 0.0011
R17781 DVDD.n7244 DVDD.n7242 0.0011
R17782 DVDD.n7196 DVDD.n7195 0.0011
R17783 DVDD.n198 DVDD.n197 0.0011
R17784 DVDD.n15181 DVDD.n15158 0.0011
R17785 DVDD.n18655 DVDD.n18654 0.0011
R17786 DVDD.n20275 DVDD.n20274 0.0011
R17787 DVDD.n20259 DVDD.n20257 0.0011
R17788 DVDD.n7679 DVDD.n7678 0.0011
R17789 DVDD.n11207 DVDD.n11206 0.00109615
R17790 DVDD.n11207 DVDD.n11201 0.00109615
R17791 DVDD.n14334 DVDD.n14333 0.00109615
R17792 DVDD.n14337 DVDD.n14334 0.00109615
R17793 DVDD.n16037 DVDD.n16036 0.00109414
R17794 DVDD.n16013 DVDD.n16012 0.00109414
R17795 DVDD.n16038 DVDD.n16037 0.00109414
R17796 DVDD.n16014 DVDD.n16013 0.00109414
R17797 DVDD.n15649 DVDD.n15648 0.00109414
R17798 DVDD.n15625 DVDD.n15624 0.00109414
R17799 DVDD.n15650 DVDD.n15649 0.00109414
R17800 DVDD.n15626 DVDD.n15625 0.00109414
R17801 DVDD.n8152 DVDD.n8151 0.00109414
R17802 DVDD.n8153 DVDD.n8152 0.00109414
R17803 DVDD.n8323 DVDD.n8322 0.00109414
R17804 DVDD.n8005 DVDD.n8004 0.00109414
R17805 DVDD.n8054 DVDD.n8053 0.00109414
R17806 DVDD.n8053 DVDD.n8052 0.00109414
R17807 DVDD.n16497 DVDD.n16496 0.00109
R17808 DVDD.n16501 DVDD.n16500 0.00109
R17809 DVDD.n16496 DVDD.n16495 0.00109
R17810 DVDD.n16500 DVDD.n16499 0.00109
R17811 DVDD.n14523 DVDD.n14522 0.00108858
R17812 DVDD.n14524 DVDD.n14523 0.00108858
R17813 DVDD.n6109 DVDD.n5699 0.00108858
R17814 DVDD.n6109 DVDD.n6108 0.00108858
R17815 DVDD.n12783 DVDD.n12782 0.00108858
R17816 DVDD.n12784 DVDD.n12783 0.00108858
R17817 DVDD.n6160 DVDD.n6159 0.00108858
R17818 DVDD.n6161 DVDD.n6160 0.00108858
R17819 DVDD.n8862 DVDD.n8861 0.00108858
R17820 DVDD.n8863 DVDD.n8862 0.00108858
R17821 DVDD.n12060 DVDD.n12059 0.00108858
R17822 DVDD.n13343 DVDD.n13342 0.00108858
R17823 DVDD.n13520 DVDD.n13519 0.00108858
R17824 DVDD.n13572 DVDD.n13571 0.00108858
R17825 DVDD.n13593 DVDD.n13592 0.00108858
R17826 DVDD.n13653 DVDD.n13652 0.00108858
R17827 DVDD.n13674 DVDD.n13673 0.00108858
R17828 DVDD.n12059 DVDD.n12058 0.00108858
R17829 DVDD.n12110 DVDD.n12109 0.00108858
R17830 DVDD.n13342 DVDD.n13341 0.00108858
R17831 DVDD.n13519 DVDD.n13518 0.00108858
R17832 DVDD.n13571 DVDD.n13570 0.00108858
R17833 DVDD.n13592 DVDD.n13591 0.00108858
R17834 DVDD.n13652 DVDD.n13651 0.00108858
R17835 DVDD.n13673 DVDD.n13672 0.00108858
R17836 DVDD.n15419 DVDD.n15418 0.00108858
R17837 DVDD.n15443 DVDD.n15442 0.00108858
R17838 DVDD.n14684 DVDD.n14683 0.00108858
R17839 DVDD.n14601 DVDD.n14600 0.00108858
R17840 DVDD.n14547 DVDD.n14546 0.00108858
R17841 DVDD.n14459 DVDD.n14458 0.00108858
R17842 DVDD.n14419 DVDD.n14418 0.00108858
R17843 DVDD.n14460 DVDD.n14459 0.00108858
R17844 DVDD.n14548 DVDD.n14547 0.00108858
R17845 DVDD.n14602 DVDD.n14601 0.00108858
R17846 DVDD.n14685 DVDD.n14684 0.00108858
R17847 DVDD.n15418 DVDD.n15417 0.00108858
R17848 DVDD.n15442 DVDD.n15441 0.00108858
R17849 DVDD.n14420 DVDD.n14419 0.00108858
R17850 DVDD.n4928 DVDD.n4927 0.00108858
R17851 DVDD.n4972 DVDD.n4971 0.00108858
R17852 DVDD.n4973 DVDD.n4972 0.00108858
R17853 DVDD.n5336 DVDD.n5335 0.00108858
R17854 DVDD.n5486 DVDD.n5485 0.00108858
R17855 DVDD.n5654 DVDD.n5653 0.00108858
R17856 DVDD.n6027 DVDD.n6026 0.00108858
R17857 DVDD.n5977 DVDD.n5976 0.00108858
R17858 DVDD.n5855 DVDD.n5854 0.00108858
R17859 DVDD.n5838 DVDD.n5837 0.00108858
R17860 DVDD.n5821 DVDD.n5820 0.00108858
R17861 DVDD.n6028 DVDD.n6027 0.00108858
R17862 DVDD.n5335 DVDD.n5334 0.00108858
R17863 DVDD.n5485 DVDD.n5484 0.00108858
R17864 DVDD.n5452 DVDD.n5451 0.00108858
R17865 DVDD.n5406 DVDD.n5405 0.00108858
R17866 DVDD.n4971 DVDD.n4970 0.00108858
R17867 DVDD.n4927 DVDD.n4926 0.00108858
R17868 DVDD.n5087 DVDD.n5086 0.00108858
R17869 DVDD.n5316 DVDD.n5315 0.00108858
R17870 DVDD.n5978 DVDD.n5977 0.00108858
R17871 DVDD.n5653 DVDD.n5652 0.00108858
R17872 DVDD.n11825 DVDD.n11824 0.00108858
R17873 DVDD.n11781 DVDD.n11780 0.00108858
R17874 DVDD.n13123 DVDD.n13122 0.00108858
R17875 DVDD.n12977 DVDD.n12976 0.00108858
R17876 DVDD.n12740 DVDD.n12739 0.00108858
R17877 DVDD.n12678 DVDD.n12677 0.00108858
R17878 DVDD.n12640 DVDD.n12639 0.00108858
R17879 DVDD.n12553 DVDD.n12552 0.00108858
R17880 DVDD.n12536 DVDD.n12535 0.00108858
R17881 DVDD.n12519 DVDD.n12518 0.00108858
R17882 DVDD.n13124 DVDD.n13123 0.00108858
R17883 DVDD.n12978 DVDD.n12977 0.00108858
R17884 DVDD.n11826 DVDD.n11825 0.00108858
R17885 DVDD.n11782 DVDD.n11781 0.00108858
R17886 DVDD.n11725 DVDD.n11724 0.00108858
R17887 DVDD.n12641 DVDD.n12640 0.00108858
R17888 DVDD.n12679 DVDD.n12678 0.00108858
R17889 DVDD.n12741 DVDD.n12740 0.00108858
R17890 DVDD.n18183 DVDD.n18182 0.00108858
R17891 DVDD.n18162 DVDD.n18161 0.00108858
R17892 DVDD.n18039 DVDD.n18038 0.00108858
R17893 DVDD.n17961 DVDD.n17960 0.00108858
R17894 DVDD.n17909 DVDD.n17908 0.00108858
R17895 DVDD.n17888 DVDD.n17887 0.00108858
R17896 DVDD.n17828 DVDD.n17827 0.00108858
R17897 DVDD.n17793 DVDD.n17792 0.00108858
R17898 DVDD.n18040 DVDD.n18039 0.00108858
R17899 DVDD.n18184 DVDD.n18183 0.00108858
R17900 DVDD.n18163 DVDD.n18162 0.00108858
R17901 DVDD.n17962 DVDD.n17961 0.00108858
R17902 DVDD.n17829 DVDD.n17828 0.00108858
R17903 DVDD.n17794 DVDD.n17793 0.00108858
R17904 DVDD.n17910 DVDD.n17909 0.00108858
R17905 DVDD.n17889 DVDD.n17888 0.00108858
R17906 DVDD.n5839 DVDD.n5838 0.00108858
R17907 DVDD.n12537 DVDD.n12536 0.00108858
R17908 DVDD.n5822 DVDD.n5821 0.00108858
R17909 DVDD.n12520 DVDD.n12519 0.00108858
R17910 DVDD.n5856 DVDD.n5855 0.00108858
R17911 DVDD.n12554 DVDD.n12553 0.00108858
R17912 DVDD.n6756 DVDD.n6755 0.00108858
R17913 DVDD.n6712 DVDD.n6711 0.00108858
R17914 DVDD.n6425 DVDD.n6424 0.00108858
R17915 DVDD.n6273 DVDD.n6272 0.00108858
R17916 DVDD.n6122 DVDD.n6121 0.00108858
R17917 DVDD.n4478 DVDD.n4477 0.00108858
R17918 DVDD.n4440 DVDD.n4439 0.00108858
R17919 DVDD.n4301 DVDD.n4300 0.00108858
R17920 DVDD.n4276 DVDD.n4275 0.00108858
R17921 DVDD.n4251 DVDD.n4250 0.00108858
R17922 DVDD.n4479 DVDD.n4478 0.00108858
R17923 DVDD.n4302 DVDD.n4301 0.00108858
R17924 DVDD.n4277 DVDD.n4276 0.00108858
R17925 DVDD.n4252 DVDD.n4251 0.00108858
R17926 DVDD.n6274 DVDD.n6273 0.00108858
R17927 DVDD.n6426 DVDD.n6425 0.00108858
R17928 DVDD.n6360 DVDD.n6359 0.00108858
R17929 DVDD.n6655 DVDD.n6654 0.00108858
R17930 DVDD.n6713 DVDD.n6712 0.00108858
R17931 DVDD.n6757 DVDD.n6756 0.00108858
R17932 DVDD.n4441 DVDD.n4440 0.00108858
R17933 DVDD.n6123 DVDD.n6122 0.00108858
R17934 DVDD.n9724 DVDD.n9723 0.00108858
R17935 DVDD.n9680 DVDD.n9679 0.00108858
R17936 DVDD.n9211 DVDD.n9210 0.00108858
R17937 DVDD.n9059 DVDD.n9058 0.00108858
R17938 DVDD.n8824 DVDD.n8823 0.00108858
R17939 DVDD.n8764 DVDD.n8763 0.00108858
R17940 DVDD.n8714 DVDD.n8713 0.00108858
R17941 DVDD.n8597 DVDD.n8596 0.00108858
R17942 DVDD.n8580 DVDD.n8579 0.00108858
R17943 DVDD.n8563 DVDD.n8562 0.00108858
R17944 DVDD.n9725 DVDD.n9724 0.00108858
R17945 DVDD.n9212 DVDD.n9211 0.00108858
R17946 DVDD.n9060 DVDD.n9059 0.00108858
R17947 DVDD.n8765 DVDD.n8764 0.00108858
R17948 DVDD.n8598 DVDD.n8597 0.00108858
R17949 DVDD.n8581 DVDD.n8580 0.00108858
R17950 DVDD.n8564 DVDD.n8563 0.00108858
R17951 DVDD.n9146 DVDD.n9145 0.00108858
R17952 DVDD.n9623 DVDD.n9622 0.00108858
R17953 DVDD.n9681 DVDD.n9680 0.00108858
R17954 DVDD.n8715 DVDD.n8714 0.00108858
R17955 DVDD.n8825 DVDD.n8824 0.00108858
R17956 DVDD.n16382 DVDD 0.00108667
R17957 DVDD.n387 DVDD.n386 0.00107857
R17958 DVDD.n391 DVDD.n390 0.00107857
R17959 DVDD.n618 DVDD.n617 0.00107857
R17960 DVDD.n622 DVDD.n621 0.00107857
R17961 DVDD.n2669 DVDD.n2668 0.00107857
R17962 DVDD.n2677 DVDD.n2676 0.00107857
R17963 DVDD.n15264 DVDD.n15263 0.00107631
R17964 DVDD.n19558 DVDD.n19557 0.00107
R17965 DVDD.n19556 DVDD.n19555 0.00107
R17966 DVDD.n19545 DVDD.n19544 0.00107
R17967 DVDD.n3917 DVDD.n3916 0.00107
R17968 DVDD.n20173 DVDD.n20172 0.00107
R17969 DVDD.n20171 DVDD.n20170 0.00107
R17970 DVDD.n20160 DVDD.n20159 0.00107
R17971 DVDD.n7383 DVDD.n7381 0.00107
R17972 DVDD.n57 DVDD.n55 0.00107
R17973 DVDD.n7256 DVDD.n7254 0.00107
R17974 DVDD.n859 DVDD.n858 0.00107
R17975 DVDD.n229 DVDD.n228 0.00107
R17976 DVDD.n18245 DVDD.n18244 0.00107
R17977 DVDD.n7181 DVDD.n7180 0.00107
R17978 DVDD.n10342 DVDD.n10341 0.00107
R17979 DVDD.n10351 DVDD.n10350 0.00107
R17980 DVDD.n10356 DVDD.n10355 0.00107
R17981 DVDD.n15356 DVDD.n15355 0.00107
R17982 DVDD.n15347 DVDD.n15346 0.00107
R17983 DVDD.n16499 DVDD.n16498 0.00107
R17984 DVDD.n16506 DVDD.n16505 0.00107
R17985 DVDD.n16510 DVDD.n16509 0.00107
R17986 DVDD.n11163 DVDD.n11162 0.00107
R17987 DVDD.n11153 DVDD.n11152 0.00107
R17988 DVDD.n16842 DVDD.n16841 0.00107
R17989 DVDD.n16848 DVDD.n16847 0.00107
R17990 DVDD.n16852 DVDD.n16851 0.00107
R17991 DVDD.n16367 DVDD.n16366 0.00107
R17992 DVDD.n16358 DVDD.n16357 0.00107
R17993 DVDD.n3623 DVDD.n3622 0.00107
R17994 DVDD.n18593 DVDD.n18592 0.00107
R17995 DVDD.n14793 DVDD.n14792 0.00107
R17996 DVDD.n7173 DVDD.n7172 0.00107
R17997 DVDD.n20247 DVDD.n20245 0.00107
R17998 DVDD.n15957 DVDD.n15956 0.00106485
R17999 DVDD.n8349 DVDD.n8348 0.00106485
R18000 DVDD.n8340 DVDD.n8339 0.00106485
R18001 DVDD.n8334 DVDD.n8333 0.00106485
R18002 DVDD.n8328 DVDD.n8327 0.00106485
R18003 DVDD.n8320 DVDD.n8319 0.00106485
R18004 DVDD.n8312 DVDD.n8311 0.00106485
R18005 DVDD.n8304 DVDD.n8303 0.00106485
R18006 DVDD.n8141 DVDD.n8140 0.00106485
R18007 DVDD.n8018 DVDD.n8017 0.00106485
R18008 DVDD.n8022 DVDD.n8021 0.00106485
R18009 DVDD.n14926 DVDD.n14925 0.0010625
R18010 DVDD.n14889 DVDD.n14888 0.0010625
R18011 DVDD.n14892 DVDD.n14891 0.0010625
R18012 DVDD.n15224 DVDD.n15223 0.0010625
R18013 DVDD.n15109 DVDD.n15108 0.0010625
R18014 DVDD.n15304 DVDD.n15303 0.0010625
R18015 DVDD.n15005 DVDD.n15004 0.0010625
R18016 DVDD.n10717 DVDD.n10716 0.0010625
R18017 DVDD.n10396 DVDD.n10395 0.0010625
R18018 DVDD.n10634 DVDD.n10633 0.0010625
R18019 DVDD.n7665 DVDD 0.00105496
R18020 DVDD.n15706 DVDD 0.00104667
R18021 DVDD.n10439 DVDD.n10438 0.001045
R18022 DVDD.n16866 DVDD.n16865 0.001045
R18023 DVDD.n16566 DVDD.n16565 0.001045
R18024 DVDD.n16662 DVDD.n16661 0.001045
R18025 DVDD.n16606 DVDD.n16605 0.001045
R18026 DVDD.n16605 DVDD.n16604 0.001045
R18027 DVDD.n10440 DVDD.n10439 0.001045
R18028 DVDD.n16663 DVDD.n16662 0.001045
R18029 DVDD.n16567 DVDD.n16566 0.001045
R18030 DVDD.n16867 DVDD.n16866 0.001045
R18031 DVDD.n7761 DVDD.n7760 0.00104
R18032 DVDD.n7758 DVDD.n7757 0.00104
R18033 DVDD.n7755 DVDD.n7754 0.00104
R18034 DVDD.n7752 DVDD.n7751 0.00104
R18035 DVDD.n7749 DVDD.n7748 0.00104
R18036 DVDD.n7746 DVDD.n7745 0.00104
R18037 DVDD.n7829 DVDD.n7828 0.00104
R18038 DVDD.n9766 DVDD.n9765 0.00104
R18039 DVDD.n7933 DVDD.n7932 0.00104
R18040 DVDD.n9536 DVDD.n9535 0.00104
R18041 DVDD.n9260 DVDD.n9259 0.00104
R18042 DVDD.n9267 DVDD.n9266 0.00104
R18043 DVDD.n9302 DVDD.n9301 0.00104
R18044 DVDD.n9316 DVDD.n9315 0.00104
R18045 DVDD.n6798 DVDD.n6797 0.00104
R18046 DVDD.n6849 DVDD.n6848 0.00104
R18047 DVDD.n6522 DVDD.n6521 0.00104
R18048 DVDD.n6568 DVDD.n6567 0.00104
R18049 DVDD.n3982 DVDD.n3981 0.00104
R18050 DVDD.n3975 DVDD.n3974 0.00104
R18051 DVDD.n3940 DVDD.n3939 0.00104
R18052 DVDD.n4835 DVDD.n4834 0.00104
R18053 DVDD.n4886 DVDD.n4885 0.00104
R18054 DVDD.n5113 DVDD.n5112 0.00104
R18055 DVDD.n5159 DVDD.n5158 0.00104
R18056 DVDD.n5287 DVDD.n5286 0.00104
R18057 DVDD.n5280 DVDD.n5279 0.00104
R18058 DVDD.n5245 DVDD.n5244 0.00104
R18059 DVDD.n18273 DVDD.n18272 0.00104
R18060 DVDD.n18270 DVDD.n18269 0.00104
R18061 DVDD.n18267 DVDD.n10156 0.00104
R18062 DVDD.n10154 DVDD.n10153 0.00104
R18063 DVDD.n10151 DVDD.n10150 0.00104
R18064 DVDD.n10148 DVDD.n10147 0.00104
R18065 DVDD.n19548 DVDD.n19547 0.00104
R18066 DVDD.n19541 DVDD.n19540 0.00104
R18067 DVDD.n19537 DVDD.n19536 0.00104
R18068 DVDD.n19519 DVDD.n19518 0.00104
R18069 DVDD.n19512 DVDD.n19511 0.00104
R18070 DVDD.n7569 DVDD.n7568 0.00104
R18071 DVDD.n20163 DVDD.n20162 0.00104
R18072 DVDD.n20156 DVDD.n20155 0.00104
R18073 DVDD.n20152 DVDD.n20151 0.00104
R18074 DVDD.n20134 DVDD.n20133 0.00104
R18075 DVDD.n20127 DVDD.n20126 0.00104
R18076 DVDD.n7525 DVDD.n7524 0.00104
R18077 DVDD.n7379 DVDD.n7378 0.00104
R18078 DVDD.n61 DVDD.n60 0.00104
R18079 DVDD.n7252 DVDD.n7251 0.00104
R18080 DVDD.n1798 DVDD.n1797 0.00104
R18081 DVDD.n1802 DVDD.n1801 0.00104
R18082 DVDD.n232 DVDD.n231 0.00104
R18083 DVDD.n205 DVDD.n204 0.00104
R18084 DVDD.n174 DVDD.n173 0.00104
R18085 DVDD.n11354 DVDD.n11353 0.00104
R18086 DVDD.n11867 DVDD.n11866 0.00104
R18087 DVDD.n1245 DVDD.n1244 0.00104
R18088 DVDD.n1248 DVDD.n1247 0.00104
R18089 DVDD.n1251 DVDD.n1250 0.00104
R18090 DVDD.n1254 DVDD.n1253 0.00104
R18091 DVDD.n1257 DVDD.n1256 0.00104
R18092 DVDD.n1260 DVDD.n1259 0.00104
R18093 DVDD.n1263 DVDD.n1262 0.00104
R18094 DVDD.n1266 DVDD.n1265 0.00104
R18095 DVDD.n1269 DVDD.n1268 0.00104
R18096 DVDD.n1272 DVDD.n1271 0.00104
R18097 DVDD.n11335 DVDD.n11334 0.00104
R18098 DVDD.n12340 DVDD.n12339 0.00104
R18099 DVDD.n14974 DVDD.n14973 0.00104
R18100 DVDD.n15051 DVDD.n15050 0.00104
R18101 DVDD.n15383 DVDD.n15382 0.00104
R18102 DVDD.n15341 DVDD.n15340 0.00104
R18103 DVDD.n10427 DVDD.n10426 0.00104
R18104 DVDD.n14976 DVDD.n14975 0.00104
R18105 DVDD.n15053 DVDD.n15052 0.00104
R18106 DVDD.n15384 DVDD.n15380 0.00104
R18107 DVDD.n15366 DVDD.n15365 0.00104
R18108 DVDD.n15363 DVDD.n15362 0.00104
R18109 DVDD.n15342 DVDD.n14827 0.00104
R18110 DVDD.n13171 DVDD.n13170 0.00104
R18111 DVDD.n13178 DVDD.n13177 0.00104
R18112 DVDD.n13213 DVDD.n13212 0.00104
R18113 DVDD.n13227 DVDD.n13226 0.00104
R18114 DVDD.n17059 DVDD.n17058 0.00104
R18115 DVDD.n11031 DVDD.n11030 0.00104
R18116 DVDD.n11086 DVDD.n11085 0.00104
R18117 DVDD.n11193 DVDD.n11189 0.00104
R18118 DVDD.n11147 DVDD.n11124 0.00104
R18119 DVDD.n16166 DVDD.n16165 0.00104
R18120 DVDD.n16284 DVDD.n16283 0.00104
R18121 DVDD.n16330 DVDD.n16329 0.00104
R18122 DVDD.n16375 DVDD.n16374 0.00104
R18123 DVDD.n16371 DVDD.n16370 0.00104
R18124 DVDD.n16352 DVDD.n16342 0.00104
R18125 DVDD.n16225 DVDD.n16224 0.00104
R18126 DVDD.n15590 DVDD.n15589 0.00104
R18127 DVDD.n15737 DVDD.n15733 0.00104
R18128 DVDD.n15700 DVDD.n15699 0.00104
R18129 DVDD.n15805 DVDD.n15804 0.00104
R18130 DVDD.n15868 DVDD.n15867 0.00104
R18131 DVDD.n16096 DVDD.n16092 0.00104
R18132 DVDD.n15911 DVDD.n15910 0.00104
R18133 DVDD.n15803 DVDD.n15802 0.00104
R18134 DVDD.n15866 DVDD.n15865 0.00104
R18135 DVDD.n16095 DVDD.n16094 0.00104
R18136 DVDD.n15913 DVDD.n15912 0.00104
R18137 DVDD.n16223 DVDD.n16222 0.00104
R18138 DVDD.n15588 DVDD.n15587 0.00104
R18139 DVDD.n15736 DVDD.n15735 0.00104
R18140 DVDD.n15698 DVDD.n15697 0.00104
R18141 DVDD.n16173 DVDD.n16172 0.00104
R18142 DVDD.n16293 DVDD.n16292 0.00104
R18143 DVDD.n16328 DVDD.n16327 0.00104
R18144 DVDD.n16351 DVDD.n16350 0.00104
R18145 DVDD.n11037 DVDD.n11036 0.00104
R18146 DVDD.n11094 DVDD.n11093 0.00104
R18147 DVDD.n11192 DVDD.n11191 0.00104
R18148 DVDD.n11146 DVDD.n11145 0.00104
R18149 DVDD.n3153 DVDD.n3152 0.00104
R18150 DVDD.n3150 DVDD.n3149 0.00104
R18151 DVDD.n3147 DVDD.n3146 0.00104
R18152 DVDD.n3144 DVDD.n3143 0.00104
R18153 DVDD.n3141 DVDD.n3140 0.00104
R18154 DVDD.n3138 DVDD.n3137 0.00104
R18155 DVDD.n3135 DVDD.n3134 0.00104
R18156 DVDD.n3132 DVDD.n3131 0.00104
R18157 DVDD.n3129 DVDD.n3128 0.00104
R18158 DVDD.n3126 DVDD.n3125 0.00104
R18159 DVDD.n3636 DVDD.n3635 0.00104
R18160 DVDD.n3632 DVDD.n3631 0.00104
R18161 DVDD.n18590 DVDD.n18589 0.00104
R18162 DVDD.n18638 DVDD.n18637 0.00104
R18163 DVDD.n18702 DVDD.n18701 0.00104
R18164 DVDD.n20251 DVDD.n20250 0.00104
R18165 DVDD.n16441 DVDD.n16440 0.00103333
R18166 DVDD.n10293 DVDD.n10292 0.00103333
R18167 DVDD.n2321 DVDD.n2320 0.00103214
R18168 DVDD.n2320 DVDD.n2319 0.00103214
R18169 DVDD.n1181 DVDD.n1180 0.0010315
R18170 DVDD.n1180 DVDD.n1179 0.0010315
R18171 DVDD.n915 DVDD.n914 0.0010315
R18172 DVDD.n874 DVDD.n873 0.0010315
R18173 DVDD.n19289 DVDD.n19288 0.0010315
R18174 DVDD.n19328 DVDD.n19327 0.0010315
R18175 DVDD.n10165 DVDD.n10164 0.0010315
R18176 DVDD.n11433 DVDD.n11432 0.0010315
R18177 DVDD.n12074 DVDD.n12073 0.0010315
R18178 DVDD.n12079 DVDD.n12078 0.0010315
R18179 DVDD.n12199 DVDD.n12198 0.0010315
R18180 DVDD.n13316 DVDD.n13315 0.0010315
R18181 DVDD.n13325 DVDD.n13324 0.0010315
R18182 DVDD.n13331 DVDD.n13330 0.0010315
R18183 DVDD.n13337 DVDD.n13336 0.0010315
R18184 DVDD.n13346 DVDD.n13345 0.0010315
R18185 DVDD.n13355 DVDD.n13354 0.0010315
R18186 DVDD.n13364 DVDD.n13363 0.0010315
R18187 DVDD.n13370 DVDD.n13369 0.0010315
R18188 DVDD.n13713 DVDD.n13712 0.0010315
R18189 DVDD.n2809 DVDD.n2808 0.0010315
R18190 DVDD.n18473 DVDD.n18472 0.0010315
R18191 DVDD.n10068 DVDD.n10067 0.0010315
R18192 DVDD.n15499 DVDD.n15498 0.0010315
R18193 DVDD.n14363 DVDD.n14362 0.0010315
R18194 DVDD.n19726 DVDD.n19725 0.0010315
R18195 DVDD.n19773 DVDD.n19772 0.0010315
R18196 DVDD.n19843 DVDD.n19842 0.0010315
R18197 DVDD.n19853 DVDD.n19852 0.0010315
R18198 DVDD.n19856 DVDD.n19855 0.0010315
R18199 DVDD.n19863 DVDD.n19862 0.0010315
R18200 DVDD.n19869 DVDD.n19868 0.0010315
R18201 DVDD.n19903 DVDD.n19902 0.0010315
R18202 DVDD.n19998 DVDD.n19997 0.0010315
R18203 DVDD.n20068 DVDD.n20067 0.0010315
R18204 DVDD.n20071 DVDD.n20070 0.0010315
R18205 DVDD.n20107 DVDD.n20106 0.0010315
R18206 DVDD.n19073 DVDD.n19072 0.0010315
R18207 DVDD.n19011 DVDD.n19010 0.0010315
R18208 DVDD.n3869 DVDD.n3868 0.0010315
R18209 DVDD.n3871 DVDD.n3870 0.0010315
R18210 DVDD.n4709 DVDD.n4708 0.0010315
R18211 DVDD.n4950 DVDD.n4949 0.0010315
R18212 DVDD.n4999 DVDD.n4998 0.0010315
R18213 DVDD.n5003 DVDD.n5002 0.0010315
R18214 DVDD.n5057 DVDD.n5056 0.0010315
R18215 DVDD.n5163 DVDD.n5108 0.0010315
R18216 DVDD.n5387 DVDD.n5386 0.0010315
R18217 DVDD.n5927 DVDD.n5926 0.0010315
R18218 DVDD.n1371 DVDD.n1370 0.0010315
R18219 DVDD.n1418 DVDD.n1417 0.0010315
R18220 DVDD.n1533 DVDD.n1532 0.0010315
R18221 DVDD.n1523 DVDD.n1522 0.0010315
R18222 DVDD.n1520 DVDD.n1519 0.0010315
R18223 DVDD.n1513 DVDD.n1512 0.0010315
R18224 DVDD.n1507 DVDD.n1506 0.0010315
R18225 DVDD.n1478 DVDD.n1477 0.0010315
R18226 DVDD.n1474 DVDD.n1473 0.0010315
R18227 DVDD.n1686 DVDD.n1685 0.0010315
R18228 DVDD.n1705 DVDD.n1704 0.0010315
R18229 DVDD.n1702 DVDD.n1701 0.0010315
R18230 DVDD.n19205 DVDD.n19204 0.0010315
R18231 DVDD.n19455 DVDD.n19454 0.0010315
R18232 DVDD.n19220 DVDD.n19219 0.0010315
R18233 DVDD.n10116 DVDD.n10115 0.0010315
R18234 DVDD.n10118 DVDD.n10117 0.0010315
R18235 DVDD.n11416 DVDD.n11415 0.0010315
R18236 DVDD.n11625 DVDD.n11624 0.0010315
R18237 DVDD.n11803 DVDD.n11802 0.0010315
R18238 DVDD.n11754 DVDD.n11753 0.0010315
R18239 DVDD.n11697 DVDD.n11696 0.0010315
R18240 DVDD.n12344 DVDD.n11304 0.0010315
R18241 DVDD.n13074 DVDD.n13073 0.0010315
R18242 DVDD.n12590 DVDD.n12589 0.0010315
R18243 DVDD.n841 DVDD.n840 0.0010315
R18244 DVDD.n19169 DVDD.n19168 0.0010315
R18245 DVDD.n10100 DVDD.n10099 0.0010315
R18246 DVDD.n18112 DVDD.n18111 0.0010315
R18247 DVDD.n17743 DVDD.n17742 0.0010315
R18248 DVDD.n1948 DVDD.n1947 0.0010315
R18249 DVDD.n1995 DVDD.n1994 0.0010315
R18250 DVDD.n2065 DVDD.n2064 0.0010315
R18251 DVDD.n2075 DVDD.n2074 0.0010315
R18252 DVDD.n2078 DVDD.n2077 0.0010315
R18253 DVDD.n2085 DVDD.n2084 0.0010315
R18254 DVDD.n2091 DVDD.n2090 0.0010315
R18255 DVDD.n2120 DVDD.n2119 0.0010315
R18256 DVDD.n2124 DVDD.n2123 0.0010315
R18257 DVDD.n2219 DVDD.n2218 0.0010315
R18258 DVDD.n2289 DVDD.n2288 0.0010315
R18259 DVDD.n2292 DVDD.n2291 0.0010315
R18260 DVDD.n19492 DVDD.n19491 0.0010315
R18261 DVDD.n18965 DVDD.n18964 0.0010315
R18262 DVDD.n18938 DVDD.n18937 0.0010315
R18263 DVDD.n7090 DVDD.n7089 0.0010315
R18264 DVDD.n7092 DVDD.n7091 0.0010315
R18265 DVDD.n6975 DVDD.n6974 0.0010315
R18266 DVDD.n6885 DVDD.n6884 0.0010315
R18267 DVDD.n6734 DVDD.n6733 0.0010315
R18268 DVDD.n6685 DVDD.n6684 0.0010315
R18269 DVDD.n6625 DVDD.n6624 0.0010315
R18270 DVDD.n6573 DVDD.n6572 0.0010315
R18271 DVDD.n6374 DVDD.n6373 0.0010315
R18272 DVDD.n4384 DVDD.n4383 0.0010315
R18273 DVDD.n3232 DVDD.n3231 0.0010315
R18274 DVDD.n3185 DVDD.n3184 0.0010315
R18275 DVDD.n3464 DVDD.n3463 0.0010315
R18276 DVDD.n3474 DVDD.n3473 0.0010315
R18277 DVDD.n3477 DVDD.n3476 0.0010315
R18278 DVDD.n3484 DVDD.n3483 0.0010315
R18279 DVDD.n3490 DVDD.n3489 0.0010315
R18280 DVDD.n3519 DVDD.n3518 0.0010315
R18281 DVDD.n3523 DVDD.n3522 0.0010315
R18282 DVDD.n3563 DVDD.n3562 0.0010315
R18283 DVDD.n3733 DVDD.n3732 0.0010315
R18284 DVDD.n3736 DVDD.n3735 0.0010315
R18285 DVDD.n18509 DVDD.n18508 0.0010315
R18286 DVDD.n18802 DVDD.n18801 0.0010315
R18287 DVDD.n18524 DVDD.n18523 0.0010315
R18288 DVDD.n7148 DVDD.n7147 0.0010315
R18289 DVDD.n7150 DVDD.n7149 0.0010315
R18290 DVDD.n9992 DVDD.n9991 0.0010315
R18291 DVDD.n7881 DVDD.n7880 0.0010315
R18292 DVDD.n9702 DVDD.n9701 0.0010315
R18293 DVDD.n9653 DVDD.n9652 0.0010315
R18294 DVDD.n9593 DVDD.n9592 0.0010315
R18295 DVDD.n9541 DVDD.n9540 0.0010315
R18296 DVDD.n9160 DVDD.n9159 0.0010315
R18297 DVDD.n8658 DVDD.n8657 0.0010315
R18298 DVDD.n14970 DVDD.n14969 0.00103
R18299 DVDD.n16357 DVDD.n16356 0.00103
R18300 DVDD.n15798 DVDD.n15797 0.00103
R18301 DVDD.n15861 DVDD.n15860 0.00103
R18302 DVDD.n16099 DVDD.n16098 0.00103
R18303 DVDD.n16100 DVDD.n16099 0.00103
R18304 DVDD.n15797 DVDD.n15796 0.00103
R18305 DVDD.n14969 DVDD.n14968 0.00103
R18306 DVDD.n16356 DVDD.n16355 0.00103
R18307 DVDD.n15860 DVDD.n15859 0.00103
R18308 DVDD.n15030 DVDD.n15029 0.001015
R18309 DVDD.n16315 DVDD.n16314 0.001015
R18310 DVDD.n16373 DVDD.n16372 0.001015
R18311 DVDD.n16199 DVDD.n16198 0.001015
R18312 DVDD.n15564 DVDD.n15563 0.001015
R18313 DVDD.n16314 DVDD.n16313 0.001015
R18314 DVDD.n16198 DVDD.n16197 0.001015
R18315 DVDD.n16374 DVDD.n16373 0.001015
R18316 DVDD.n15031 DVDD.n15030 0.001015
R18317 DVDD.n15563 DVDD.n15562 0.001015
R18318 DVDD.n2479 DVDD.n2478 0.00101429
R18319 DVDD.n19552 DVDD.n19551 0.00101
R18320 DVDD.n19516 DVDD.n19515 0.00101
R18321 DVDD.n19506 DVDD.n19505 0.00101
R18322 DVDD.n18862 DVDD.n18861 0.00101
R18323 DVDD.n18856 DVDD.n18855 0.00101
R18324 DVDD.n7565 DVDD.n7564 0.00101
R18325 DVDD.n20167 DVDD.n20166 0.00101
R18326 DVDD.n20131 DVDD.n20130 0.00101
R18327 DVDD.n20121 DVDD.n20120 0.00101
R18328 DVDD.n19111 DVDD.n19110 0.00101
R18329 DVDD.n19106 DVDD.n19103 0.00101
R18330 DVDD.n7521 DVDD.n7520 0.00101
R18331 DVDD.n7359 DVDD.n7357 0.00101
R18332 DVDD.n7409 DVDD.n7408 0.00101
R18333 DVDD.n7590 DVDD.n7588 0.00101
R18334 DVDD.n81 DVDD.n79 0.00101
R18335 DVDD.n7457 DVDD.n7456 0.00101
R18336 DVDD.n7546 DVDD.n7544 0.00101
R18337 DVDD.n7232 DVDD.n7230 0.00101
R18338 DVDD.n7494 DVDD.n7493 0.00101
R18339 DVDD.n7192 DVDD.n7190 0.00101
R18340 DVDD.n1806 DVDD.n1805 0.00101
R18341 DVDD.n254 DVDD.n253 0.00101
R18342 DVDD.n224 DVDD.n223 0.00101
R18343 DVDD.n183 DVDD.n182 0.00101
R18344 DVDD.n166 DVDD.n165 0.00101
R18345 DVDD.n19386 DVDD.n19385 0.00101
R18346 DVDD.n19381 DVDD.n19380 0.00101
R18347 DVDD.n18264 DVDD.n18263 0.00101
R18348 DVDD.n14977 DVDD.n14976 0.00101
R18349 DVDD.n15380 DVDD.n15379 0.00101
R18350 DVDD.n15336 DVDD.n14827 0.00101
R18351 DVDD.n15733 DVDD.n15732 0.00101
R18352 DVDD.n15701 DVDD.n15700 0.00101
R18353 DVDD.n16092 DVDD.n16091 0.00101
R18354 DVDD.n15910 DVDD.n15909 0.00101
R18355 DVDD.n3628 DVDD.n2812 0.00101
R18356 DVDD.n18563 DVDD.n2301 0.00101
R18357 DVDD.n18605 DVDD.n18604 0.00101
R18358 DVDD.n18725 DVDD.n18717 0.00101
R18359 DVDD.n18687 DVDD.n18686 0.00101
R18360 DVDD.n18382 DVDD.n18381 0.00101
R18361 DVDD.n18377 DVDD.n18376 0.00101
R18362 DVDD.n14789 DVDD.n14788 0.00101
R18363 DVDD.n20271 DVDD.n20269 0.00101
R18364 DVDD.n7325 DVDD.n7324 0.00101
R18365 DVDD.n7683 DVDD.n7681 0.00101
R18366 DVDD.n15236 DVDD.n15235 0.00100625
R18367 DVDD.n15242 DVDD.n15241 0.00100625
R18368 DVDD.n10571 DVDD.n10570 0.00100625
R18369 DVDD.n10575 DVDD.n10574 0.00100625
R18370 DVDD.n10654 DVDD.n10653 0.00100625
R18371 DVDD.n19596 DVDD.n19560 0.00098
R18372 DVDD.n19523 DVDD.n19522 0.00098
R18373 DVDD.n18888 DVDD.n18887 0.00098
R18374 DVDD.n18882 DVDD.n18881 0.00098
R18375 DVDD.n18860 DVDD.n18859 0.00098
R18376 DVDD.n18843 DVDD.n18842 0.00098
R18377 DVDD.n7075 DVDD.n7074 0.00098
R18378 DVDD.n20211 DVDD.n20175 0.00098
R18379 DVDD.n20138 DVDD.n20137 0.00098
R18380 DVDD.n19137 DVDD.n19136 0.00098
R18381 DVDD.n19131 DVDD.n19130 0.00098
R18382 DVDD.n19109 DVDD.n19108 0.00098
R18383 DVDD.n19091 DVDD.n19090 0.00098
R18384 DVDD.n4609 DVDD.n4603 0.00098
R18385 DVDD.n7421 DVDD.n7420 0.00098
R18386 DVDD.n7405 DVDD.n7403 0.00098
R18387 DVDD.n7469 DVDD.n7468 0.00098
R18388 DVDD.n7453 DVDD.n7451 0.00098
R18389 DVDD.n7482 DVDD.n7481 0.00098
R18390 DVDD.n7498 DVDD.n7496 0.00098
R18391 DVDD.n854 DVDD.n853 0.00098
R18392 DVDD.n19352 DVDD.n19351 0.00098
R18393 DVDD.n19412 DVDD.n19411 0.00098
R18394 DVDD.n19384 DVDD.n19383 0.00098
R18395 DVDD.n19368 DVDD.n19367 0.00098
R18396 DVDD.n19364 DVDD.n19363 0.00098
R18397 DVDD.n19361 DVDD.n19360 0.00098
R18398 DVDD.n18238 DVDD.n10187 0.00098
R18399 DVDD.n10333 DVDD.n10332 0.00098
R18400 DVDD.n10369 DVDD.n10368 0.00098
R18401 DVDD.n14952 DVDD.n14951 0.00098
R18402 DVDD.n14955 DVDD.n14954 0.00098
R18403 DVDD.n16492 DVDD.n16491 0.00098
R18404 DVDD.n16519 DVDD.n16518 0.00098
R18405 DVDD.n11010 DVDD.n11009 0.00098
R18406 DVDD.n11013 DVDD.n11012 0.00098
R18407 DVDD.n16836 DVDD.n16835 0.00098
R18408 DVDD.n16862 DVDD.n16861 0.00098
R18409 DVDD.n16995 DVDD.n16994 0.00098
R18410 DVDD.n16936 DVDD.n16935 0.00098
R18411 DVDD.n16709 DVDD.n16708 0.00098
R18412 DVDD.n16728 DVDD.n16727 0.00098
R18413 DVDD.n16770 DVDD.n16769 0.00098
R18414 DVDD.n16893 DVDD.n16892 0.00098
R18415 DVDD.n16540 DVDD.n16539 0.00098
R18416 DVDD.n16559 DVDD.n16558 0.00098
R18417 DVDD.n16647 DVDD.n16646 0.00098
R18418 DVDD.n16590 DVDD.n16589 0.00098
R18419 DVDD.n3618 DVDD.n3617 0.00098
R18420 DVDD.n18453 DVDD.n18452 0.00098
R18421 DVDD.n18419 DVDD.n18418 0.00098
R18422 DVDD.n18380 DVDD.n18379 0.00098
R18423 DVDD.n18364 DVDD.n18363 0.00098
R18424 DVDD.n18360 DVDD.n18359 0.00098
R18425 DVDD.n18357 DVDD.n18339 0.00098
R18426 DVDD.n14799 DVDD.n14745 0.00098
R18427 DVDD.n7337 DVDD.n7336 0.00098
R18428 DVDD.n7321 DVDD.n7319 0.00098
R18429 DVDD.n7705 DVDD.n7704 0.00095
R18430 DVDD.n7710 DVDD.n7709 0.00095
R18431 DVDD.n7770 DVDD.n7769 0.00095
R18432 DVDD.n3702 DVDD.n3701 0.00095
R18433 DVDD.n3697 DVDD.n3696 0.00095
R18434 DVDD.n18543 DVDD.n18542 0.00095
R18435 DVDD.n18548 DVDD.n18547 0.00095
R18436 DVDD.n3450 DVDD.n3449 0.00095
R18437 DVDD.n2959 DVDD.n2958 0.00095
R18438 DVDD.n3577 DVDD.n3576 0.00095
R18439 DVDD.n9956 DVDD.n9955 0.00095
R18440 DVDD.n9817 DVDD.n9816 0.00095
R18441 DVDD.n9517 DVDD.n9516 0.00095
R18442 DVDD.n2197 DVDD.n2196 0.00095
R18443 DVDD.n2258 DVDD.n2257 0.00095
R18444 DVDD.n2253 DVDD.n2252 0.00095
R18445 DVDD.n18912 DVDD.n18911 0.00095
R18446 DVDD.n18917 DVDD.n18916 0.00095
R18447 DVDD.n7064 DVDD.n7063 0.00095
R18448 DVDD.n7059 DVDD.n7058 0.00095
R18449 DVDD.n1897 DVDD.n1896 0.00095
R18450 DVDD.n1892 DVDD.n1891 0.00095
R18451 DVDD.n3808 DVDD.n3807 0.00095
R18452 DVDD.n18816 DVDD.n18815 0.00095
R18453 DVDD.n19976 DVDD.n19975 0.00095
R18454 DVDD.n20037 DVDD.n20036 0.00095
R18455 DVDD.n20032 DVDD.n20031 0.00095
R18456 DVDD.n19030 DVDD.n19029 0.00095
R18457 DVDD.n19035 DVDD.n19034 0.00095
R18458 DVDD.n4644 DVDD.n4643 0.00095
R18459 DVDD.n4639 DVDD.n4638 0.00095
R18460 DVDD.n19675 DVDD.n19674 0.00095
R18461 DVDD.n19670 DVDD.n19669 0.00095
R18462 DVDD.n1547 DVDD.n1546 0.00095
R18463 DVDD.n969 DVDD.n968 0.00095
R18464 DVDD.n1673 DVDD.n1672 0.00095
R18465 DVDD.n2395 DVDD.n2394 0.00095
R18466 DVDD.n2400 DVDD.n2399 0.00095
R18467 DVDD.n2475 DVDD.n2472 0.00095
R18468 DVDD.n2477 DVDD.n2476 0.00095
R18469 DVDD.n945 DVDD.n944 0.00095
R18470 DVDD.n940 DVDD.n939 0.00095
R18471 DVDD.n19239 DVDD.n19238 0.00095
R18472 DVDD.n19244 DVDD.n19243 0.00095
R18473 DVDD.n11540 DVDD.n11539 0.00095
R18474 DVDD.n18320 DVDD.n18319 0.00095
R18475 DVDD.n18315 DVDD.n18314 0.00095
R18476 DVDD.n10126 DVDD.n10125 0.00095
R18477 DVDD.n18993 DVDD.n18992 0.00095
R18478 DVDD.n19150 DVDD.n19149 0.00095
R18479 DVDD.n7263 DVDD.n7262 0.00095
R18480 DVDD.n3845 DVDD.n3844 0.00095
R18481 DVDD.n10074 DVDD.n10073 0.00095
R18482 DVDD.n7627 DVDD.n7626 0.00095
R18483 DVDD.n3897 DVDD.n3896 0.00095
R18484 DVDD.n7117 DVDD.n7116 0.00095
R18485 DVDD.n7651 DVDD.n7650 0.00095
R18486 DVDD.n130 DVDD.n129 0.00095
R18487 DVDD.n1810 DVDD.n1809 0.00095
R18488 DVDD.n1841 DVDD.n1840 0.00095
R18489 DVDD.n1847 DVDD.n1846 0.00095
R18490 DVDD.n18842 DVDD.n18841 0.00095
R18491 DVDD.n3919 DVDD.n3918 0.00095
R18492 DVDD.n7572 DVDD.n7571 0.00095
R18493 DVDD.n19619 DVDD.n19618 0.00095
R18494 DVDD.n19625 DVDD.n19624 0.00095
R18495 DVDD.n19090 DVDD.n19089 0.00095
R18496 DVDD.n4606 DVDD.n4605 0.00095
R18497 DVDD.n7528 DVDD.n7527 0.00095
R18498 DVDD.n3786 DVDD.n3785 0.00095
R18499 DVDD.n2819 DVDD.n2818 0.00095
R18500 DVDD.n20293 DVDD.n20292 0.00095
R18501 DVDD.n19 DVDD.n17 0.00095
R18502 DVDD.n7393 DVDD.n7391 0.00095
R18503 DVDD.n101 DVDD.n99 0.00095
R18504 DVDD.n7441 DVDD.n7439 0.00095
R18505 DVDD.n20315 DVDD.n20314 0.00095
R18506 DVDD.n47 DVDD.n45 0.00095
R18507 DVDD.n7510 DVDD.n7508 0.00095
R18508 DVDD.n1786 DVDD.n1785 0.00095
R18509 DVDD.n1794 DVDD.n1793 0.00095
R18510 DVDD.n188 DVDD.n187 0.00095
R18511 DVDD.n179 DVDD.n178 0.00095
R18512 DVDD.n19401 DVDD.n19400 0.00095
R18513 DVDD.n19396 DVDD.n19395 0.00095
R18514 DVDD.n19367 DVDD.n19366 0.00095
R18515 DVDD.n18243 DVDD.n18242 0.00095
R18516 DVDD.n11918 DVDD.n11917 0.00095
R18517 DVDD.n1320 DVDD.n1319 0.00095
R18518 DVDD.n1315 DVDD.n1314 0.00095
R18519 DVDD.n1282 DVDD.n1281 0.00095
R18520 DVDD.n2593 DVDD.n2592 0.00095
R18521 DVDD.n2596 DVDD.n2595 0.00095
R18522 DVDD.n2684 DVDD.n2683 0.00095
R18523 DVDD.n2687 DVDD.n2686 0.00095
R18524 DVDD.n12322 DVDD.n12321 0.00095
R18525 DVDD.n14844 DVDD.n14843 0.00095
R18526 DVDD.n14864 DVDD.n14863 0.00095
R18527 DVDD.n15088 DVDD.n15087 0.00095
R18528 DVDD.n10336 DVDD.n10334 0.00095
R18529 DVDD.n10372 DVDD.n10370 0.00095
R18530 DVDD.n10515 DVDD.n10513 0.00095
R18531 DVDD.n10444 DVDD.n10442 0.00095
R18532 DVDD.n10706 DVDD.n10705 0.00095
R18533 DVDD.n10596 DVDD.n10595 0.00095
R18534 DVDD.n10612 DVDD.n10611 0.00095
R18535 DVDD.n10337 DVDD.n10333 0.00095
R18536 DVDD.n10373 DVDD.n10369 0.00095
R18537 DVDD.n10517 DVDD.n10516 0.00095
R18538 DVDD.n10446 DVDD.n10445 0.00095
R18539 DVDD.n16493 DVDD.n16492 0.00095
R18540 DVDD.n16523 DVDD.n16519 0.00095
R18541 DVDD.n17124 DVDD.n17123 0.00095
R18542 DVDD.n17074 DVDD.n17073 0.00095
R18543 DVDD.n16837 DVDD.n16836 0.00095
R18544 DVDD.n16863 DVDD.n16862 0.00095
R18545 DVDD.n17014 DVDD.n17013 0.00095
R18546 DVDD.n16956 DVDD.n16955 0.00095
R18547 DVDD.n16141 DVDD.n16140 0.00095
R18548 DVDD.n16145 DVDD.n16144 0.00095
R18549 DVDD.n16260 DVDD.n16259 0.00095
R18550 DVDD.n16263 DVDD.n16262 0.00095
R18551 DVDD.n16710 DVDD.n16709 0.00095
R18552 DVDD.n16732 DVDD.n16728 0.00095
R18553 DVDD.n16792 DVDD.n16791 0.00095
R18554 DVDD.n16915 DVDD.n16914 0.00095
R18555 DVDD.n16197 DVDD.n16196 0.00095
R18556 DVDD.n16201 DVDD.n16200 0.00095
R18557 DVDD.n15562 DVDD.n15561 0.00095
R18558 DVDD.n15566 DVDD.n15565 0.00095
R18559 DVDD.n16541 DVDD.n16540 0.00095
R18560 DVDD.n16563 DVDD.n16559 0.00095
R18561 DVDD.n16670 DVDD.n16669 0.00095
R18562 DVDD.n16613 DVDD.n16612 0.00095
R18563 DVDD.n15777 DVDD.n15776 0.00095
R18564 DVDD.n15780 DVDD.n15779 0.00095
R18565 DVDD.n15840 DVDD.n15839 0.00095
R18566 DVDD.n15843 DVDD.n15842 0.00095
R18567 DVDD.n16536 DVDD.n16535 0.00095
R18568 DVDD.n16562 DVDD.n16560 0.00095
R18569 DVDD.n16668 DVDD.n16666 0.00095
R18570 DVDD.n16611 DVDD.n16609 0.00095
R18571 DVDD.n16705 DVDD.n16704 0.00095
R18572 DVDD.n16731 DVDD.n16729 0.00095
R18573 DVDD.n16790 DVDD.n16788 0.00095
R18574 DVDD.n16913 DVDD.n16911 0.00095
R18575 DVDD.n16831 DVDD.n16830 0.00095
R18576 DVDD.n16873 DVDD.n16872 0.00095
R18577 DVDD.n17023 DVDD.n17022 0.00095
R18578 DVDD.n16963 DVDD.n16962 0.00095
R18579 DVDD.n16487 DVDD.n16486 0.00095
R18580 DVDD.n16522 DVDD.n16520 0.00095
R18581 DVDD.n17132 DVDD.n17131 0.00095
R18582 DVDD.n17083 DVDD.n17082 0.00095
R18583 DVDD.n3361 DVDD.n3360 0.00095
R18584 DVDD.n18627 DVDD.n18626 0.00095
R18585 DVDD.n18640 DVDD.n18639 0.00095
R18586 DVDD.n18648 DVDD.n18647 0.00095
R18587 DVDD.n18441 DVDD.n18440 0.00095
R18588 DVDD.n18385 DVDD.n18384 0.00095
R18589 DVDD.n18394 DVDD.n18388 0.00095
R18590 DVDD.n14760 DVDD.n14759 0.00095
R18591 DVDD.n7167 DVDD.n7166 0.00095
R18592 DVDD.n7691 DVDD.n7169 0.00095
R18593 DVDD.n3322 DVDD.n3321 0.00095
R18594 DVDD.n3283 DVDD.n3282 0.00095
R18595 DVDD.n3288 DVDD.n3287 0.00095
R18596 DVDD.n3648 DVDD.n3647 0.00095
R18597 DVDD.n3640 DVDD.n3639 0.00095
R18598 DVDD.n18730 DVDD.n18729 0.00095
R18599 DVDD.n18714 DVDD.n18713 0.00095
R18600 DVDD.n18408 DVDD.n18407 0.00095
R18601 DVDD.n18403 DVDD.n18402 0.00095
R18602 DVDD.n18363 DVDD.n18362 0.00095
R18603 DVDD.n14795 DVDD.n14794 0.00095
R18604 DVDD.n7276 DVDD.n7275 0.00095
R18605 DVDD.n20237 DVDD.n20235 0.00095
R18606 DVDD.n7309 DVDD.n7307 0.00095
R18607 DVDD.n16416 DVDD.n16415 0.000926667
R18608 DVDD.n10246 DVDD.n10245 0.000926667
R18609 DVDD.n19503 DVDD.n19502 0.00092
R18610 DVDD.n19502 DVDD.n19467 0.00092
R18611 DVDD.n7576 DVDD.n7575 0.00092
R18612 DVDD.n20118 DVDD.n20117 0.00092
R18613 DVDD.n20117 DVDD.n20082 0.00092
R18614 DVDD.n7532 DVDD.n7531 0.00092
R18615 DVDD.n162 DVDD.n161 0.00092
R18616 DVDD.n18683 DVDD.n18682 0.00092
R18617 DVDD.n3110 DVDD.n3109 0.000901786
R18618 DVDD.n14891 DVDD.n14890 0.00089375
R18619 DVDD.n14894 DVDD.n14893 0.00089375
R18620 DVDD.n15246 DVDD.n15245 0.00089375
R18621 DVDD.n15249 DVDD.n15248 0.00089375
R18622 DVDD.n1836 DVDD.n1835 0.00089
R18623 DVDD.n1848 DVDD.n1847 0.00089
R18624 DVDD.n18885 DVDD.n18884 0.00089
R18625 DVDD.n18841 DVDD.n18840 0.00089
R18626 DVDD.n7577 DVDD.n7576 0.00089
R18627 DVDD.n19614 DVDD.n19613 0.00089
R18628 DVDD.n19626 DVDD.n19625 0.00089
R18629 DVDD.n19134 DVDD.n19133 0.00089
R18630 DVDD.n19089 DVDD.n19088 0.00089
R18631 DVDD.n7533 DVDD.n7532 0.00089
R18632 DVDD.n19 DVDD.n18 0.00089
R18633 DVDD.n7393 DVDD.n7392 0.00089
R18634 DVDD.n101 DVDD.n100 0.00089
R18635 DVDD.n7441 DVDD.n7440 0.00089
R18636 DVDD.n47 DVDD.n46 0.00089
R18637 DVDD.n7510 DVDD.n7509 0.00089
R18638 DVDD.n862 DVDD.n861 0.00089
R18639 DVDD.n1795 DVDD.n1794 0.00089
R18640 DVDD.n194 DVDD.n193 0.00089
R18641 DVDD.n169 DVDD.n168 0.00089
R18642 DVDD.n161 DVDD.n147 0.00089
R18643 DVDD.n19345 DVDD.n19344 0.00089
R18644 DVDD.n19349 DVDD.n19348 0.00089
R18645 DVDD.n19414 DVDD.n19354 0.00089
R18646 DVDD.n19366 DVDD.n19365 0.00089
R18647 DVDD.n18248 DVDD.n18247 0.00089
R18648 DVDD.n10336 DVDD.n10335 0.00089
R18649 DVDD.n10372 DVDD.n10371 0.00089
R18650 DVDD.n10515 DVDD.n10514 0.00089
R18651 DVDD.n10444 DVDD.n10443 0.00089
R18652 DVDD.n10338 DVDD.n10337 0.00089
R18653 DVDD.n10374 DVDD.n10373 0.00089
R18654 DVDD.n10516 DVDD.n10512 0.00089
R18655 DVDD.n10445 DVDD.n10441 0.00089
R18656 DVDD.n16494 DVDD.n16493 0.00089
R18657 DVDD.n16524 DVDD.n16523 0.00089
R18658 DVDD.n17123 DVDD.n17122 0.00089
R18659 DVDD.n17073 DVDD.n17072 0.00089
R18660 DVDD.n16838 DVDD.n16837 0.00089
R18661 DVDD.n16864 DVDD.n16863 0.00089
R18662 DVDD.n17013 DVDD.n17012 0.00089
R18663 DVDD.n16955 DVDD.n16954 0.00089
R18664 DVDD.n16711 DVDD.n16710 0.00089
R18665 DVDD.n16733 DVDD.n16732 0.00089
R18666 DVDD.n16791 DVDD.n16787 0.00089
R18667 DVDD.n16914 DVDD.n16910 0.00089
R18668 DVDD.n16542 DVDD.n16541 0.00089
R18669 DVDD.n16564 DVDD.n16563 0.00089
R18670 DVDD.n16669 DVDD.n16665 0.00089
R18671 DVDD.n16612 DVDD.n16608 0.00089
R18672 DVDD.n16535 DVDD.n16534 0.00089
R18673 DVDD.n16562 DVDD.n16561 0.00089
R18674 DVDD.n16668 DVDD.n16667 0.00089
R18675 DVDD.n16611 DVDD.n16610 0.00089
R18676 DVDD.n16704 DVDD.n16703 0.00089
R18677 DVDD.n16731 DVDD.n16730 0.00089
R18678 DVDD.n16790 DVDD.n16789 0.00089
R18679 DVDD.n16913 DVDD.n16912 0.00089
R18680 DVDD.n16830 DVDD.n16829 0.00089
R18681 DVDD.n16874 DVDD.n16873 0.00089
R18682 DVDD.n17022 DVDD.n17021 0.00089
R18683 DVDD.n16962 DVDD.n16961 0.00089
R18684 DVDD.n16486 DVDD.n16485 0.00089
R18685 DVDD.n16522 DVDD.n16521 0.00089
R18686 DVDD.n17131 DVDD.n17130 0.00089
R18687 DVDD.n17082 DVDD.n17081 0.00089
R18688 DVDD.n3626 DVDD.n3625 0.00089
R18689 DVDD.n3639 DVDD.n3638 0.00089
R18690 DVDD.n18735 DVDD.n18658 0.00089
R18691 DVDD.n18697 DVDD.n18696 0.00089
R18692 DVDD.n18682 DVDD.n18668 0.00089
R18693 DVDD.n18460 DVDD.n18459 0.00089
R18694 DVDD.n18456 DVDD.n18455 0.00089
R18695 DVDD.n18450 DVDD.n18449 0.00089
R18696 DVDD.n18362 DVDD.n18361 0.00089
R18697 DVDD.n14773 DVDD.n14772 0.00089
R18698 DVDD.n20237 DVDD.n20236 0.00089
R18699 DVDD.n7309 DVDD.n7308 0.00089
R18700 DVDD.n380 DVDD.n379 0.000885714
R18701 DVDD.n383 DVDD.n382 0.000885714
R18702 DVDD.n611 DVDD.n610 0.000885714
R18703 DVDD.n614 DVDD.n613 0.000885714
R18704 DVDD.n15255 DVDD.n15254 0.000884205
R18705 DVDD.n15985 DVDD.n15984 0.000876569
R18706 DVDD.n8238 DVDD.n8237 0.000876569
R18707 DVDD.n9427 DVDD.n9426 0.000876569
R18708 DVDD.n8108 DVDD.n8107 0.000876569
R18709 DVDD.n8082 DVDD.n8081 0.000876569
R18710 DVDD.n8086 DVDD.n8085 0.000876569
R18711 DVDD.n13831 DVDD 0.000871429
R18712 DVDD.n3672 DVDD.n3671 0.00086
R18713 DVDD.n2865 DVDD.n2864 0.00086
R18714 DVDD.n2862 DVDD.n2861 0.00086
R18715 DVDD.n2859 DVDD.n2858 0.00086
R18716 DVDD.n2856 DVDD.n2855 0.00086
R18717 DVDD.n2853 DVDD.n2852 0.00086
R18718 DVDD.n2850 DVDD.n2849 0.00086
R18719 DVDD.n2847 DVDD.n2846 0.00086
R18720 DVDD.n2844 DVDD.n2843 0.00086
R18721 DVDD.n2841 DVDD.n2840 0.00086
R18722 DVDD.n2838 DVDD.n2837 0.00086
R18723 DVDD.n2835 DVDD.n2834 0.00086
R18724 DVDD.n3003 DVDD.n3002 0.00086
R18725 DVDD.n2914 DVDD.n2913 0.00086
R18726 DVDD.n7164 DVDD.n7163 0.00086
R18727 DVDD.n7824 DVDD.n7823 0.00086
R18728 DVDD.n9771 DVDD.n9770 0.00086
R18729 DVDD.n9796 DVDD.n9795 0.00086
R18730 DVDD.n9531 DVDD.n9530 0.00086
R18731 DVDD.n9526 DVDD.n9525 0.00086
R18732 DVDD.n9255 DVDD.n9254 0.00086
R18733 DVDD.n9272 DVDD.n9271 0.00086
R18734 DVDD.n9297 DVDD.n9296 0.00086
R18735 DVDD.n6793 DVDD.n6792 0.00086
R18736 DVDD.n6844 DVDD.n6843 0.00086
R18737 DVDD.n6819 DVDD.n6818 0.00086
R18738 DVDD.n6563 DVDD.n6562 0.00086
R18739 DVDD.n6558 DVDD.n6557 0.00086
R18740 DVDD.n3987 DVDD.n3986 0.00086
R18741 DVDD.n3970 DVDD.n3969 0.00086
R18742 DVDD.n3945 DVDD.n3944 0.00086
R18743 DVDD.n4830 DVDD.n4829 0.00086
R18744 DVDD.n4881 DVDD.n4880 0.00086
R18745 DVDD.n4856 DVDD.n4855 0.00086
R18746 DVDD.n5154 DVDD.n5153 0.00086
R18747 DVDD.n5149 DVDD.n5148 0.00086
R18748 DVDD.n5292 DVDD.n5291 0.00086
R18749 DVDD.n5275 DVDD.n5274 0.00086
R18750 DVDD.n5250 DVDD.n5249 0.00086
R18751 DVDD.n1087 DVDD.n1086 0.00086
R18752 DVDD.n1014 DVDD.n1013 0.00086
R18753 DVDD.n1735 DVDD.n1734 0.00086
R18754 DVDD.n1739 DVDD.n1738 0.00086
R18755 DVDD.n1742 DVDD.n1741 0.00086
R18756 DVDD.n1781 DVDD.n1780 0.00086
R18757 DVDD.n1778 DVDD.n1777 0.00086
R18758 DVDD.n1775 DVDD.n1774 0.00086
R18759 DVDD.n1772 DVDD.n1771 0.00086
R18760 DVDD.n1769 DVDD.n1768 0.00086
R18761 DVDD.n1766 DVDD.n1765 0.00086
R18762 DVDD.n1763 DVDD.n1762 0.00086
R18763 DVDD.n1760 DVDD.n1759 0.00086
R18764 DVDD.n1757 DVDD.n1756 0.00086
R18765 DVDD.n11425 DVDD.n11424 0.00086
R18766 DVDD.n1844 DVDD.n1843 0.00086
R18767 DVDD.n1845 DVDD.n1844 0.00086
R18768 DVDD.n19597 DVDD.n19596 0.00086
R18769 DVDD.n18889 DVDD.n18888 0.00086
R18770 DVDD.n18877 DVDD.n18876 0.00086
R18771 DVDD.n18865 DVDD.n18864 0.00086
R18772 DVDD.n18859 DVDD.n18858 0.00086
R18773 DVDD.n18844 DVDD.n18843 0.00086
R18774 DVDD.n7074 DVDD.n3921 0.00086
R18775 DVDD.n19622 DVDD.n19621 0.00086
R18776 DVDD.n19623 DVDD.n19622 0.00086
R18777 DVDD.n20212 DVDD.n20211 0.00086
R18778 DVDD.n19138 DVDD.n19137 0.00086
R18779 DVDD.n19126 DVDD.n19125 0.00086
R18780 DVDD.n19114 DVDD.n19113 0.00086
R18781 DVDD.n19108 DVDD.n19107 0.00086
R18782 DVDD.n19092 DVDD.n19091 0.00086
R18783 DVDD.n4609 DVDD.n4608 0.00086
R18784 DVDD.n8 DVDD.n7 0.00086
R18785 DVDD.n7421 DVDD.n7419 0.00086
R18786 DVDD.n7405 DVDD.n7404 0.00086
R18787 DVDD.n90 DVDD.n89 0.00086
R18788 DVDD.n7469 DVDD.n7467 0.00086
R18789 DVDD.n7453 DVDD.n7452 0.00086
R18790 DVDD.n36 DVDD.n35 0.00086
R18791 DVDD.n7482 DVDD.n7480 0.00086
R18792 DVDD.n7498 DVDD.n7497 0.00086
R18793 DVDD.n1790 DVDD.n1789 0.00086
R18794 DVDD.n250 DVDD.n249 0.00086
R18795 DVDD.n19351 DVDD.n19350 0.00086
R18796 DVDD.n19390 DVDD.n19389 0.00086
R18797 DVDD.n19383 DVDD.n19382 0.00086
R18798 DVDD.n19369 DVDD.n19368 0.00086
R18799 DVDD.n11349 DVDD.n11348 0.00086
R18800 DVDD.n11872 DVDD.n11871 0.00086
R18801 DVDD.n11897 DVDD.n11896 0.00086
R18802 DVDD.n12335 DVDD.n12334 0.00086
R18803 DVDD.n12330 DVDD.n12329 0.00086
R18804 DVDD.n10368 DVDD.n10367 0.00086
R18805 DVDD.n10520 DVDD.n10519 0.00086
R18806 DVDD.n10449 DVDD.n10448 0.00086
R18807 DVDD.n13166 DVDD.n13165 0.00086
R18808 DVDD.n13183 DVDD.n13182 0.00086
R18809 DVDD.n13208 DVDD.n13207 0.00086
R18810 DVDD.n16518 DVDD.n16517 0.00086
R18811 DVDD.n17127 DVDD.n17126 0.00086
R18812 DVDD.n17077 DVDD.n17076 0.00086
R18813 DVDD.n17018 DVDD.n17017 0.00086
R18814 DVDD.n16996 DVDD.n16995 0.00086
R18815 DVDD.n16959 DVDD.n16958 0.00086
R18816 DVDD.n16958 DVDD.n16957 0.00086
R18817 DVDD.n16168 DVDD.n16167 0.00086
R18818 DVDD.n16262 DVDD.n16261 0.00086
R18819 DVDD.n16708 DVDD.n16707 0.00086
R18820 DVDD.n16727 DVDD.n16726 0.00086
R18821 DVDD.n16795 DVDD.n16794 0.00086
R18822 DVDD.n16794 DVDD.n16793 0.00086
R18823 DVDD.n16771 DVDD.n16770 0.00086
R18824 DVDD.n16918 DVDD.n16917 0.00086
R18825 DVDD.n16917 DVDD.n16916 0.00086
R18826 DVDD.n16894 DVDD.n16893 0.00086
R18827 DVDD.n16200 DVDD.n16199 0.00086
R18828 DVDD.n16227 DVDD.n16226 0.00086
R18829 DVDD.n15565 DVDD.n15564 0.00086
R18830 DVDD.n15592 DVDD.n15591 0.00086
R18831 DVDD.n16539 DVDD.n16538 0.00086
R18832 DVDD.n16558 DVDD.n16557 0.00086
R18833 DVDD.n16673 DVDD.n16672 0.00086
R18834 DVDD.n16672 DVDD.n16671 0.00086
R18835 DVDD.n16648 DVDD.n16647 0.00086
R18836 DVDD.n16616 DVDD.n16615 0.00086
R18837 DVDD.n16615 DVDD.n16614 0.00086
R18838 DVDD.n16591 DVDD.n16590 0.00086
R18839 DVDD.n15779 DVDD.n15778 0.00086
R18840 DVDD.n15807 DVDD.n15806 0.00086
R18841 DVDD.n15842 DVDD.n15841 0.00086
R18842 DVDD.n15870 DVDD.n15869 0.00086
R18843 DVDD.n3644 DVDD.n3643 0.00086
R18844 DVDD.n18580 DVDD.n18566 0.00086
R18845 DVDD.n18454 DVDD.n18453 0.00086
R18846 DVDD.n18397 DVDD.n18396 0.00086
R18847 DVDD.n18379 DVDD.n18378 0.00086
R18848 DVDD.n18365 DVDD.n18364 0.00086
R18849 DVDD.n20226 DVDD.n20225 0.00086
R18850 DVDD.n7337 DVDD.n7335 0.00086
R18851 DVDD.n7321 DVDD.n7320 0.00086
R18852 DVDD.n1231 DVDD.n1230 0.000854331
R18853 DVDD.n1568 DVDD.n1567 0.000854331
R18854 DVDD.n1573 DVDD.n1572 0.000854331
R18855 DVDD.n1575 DVDD.n1574 0.000854331
R18856 DVDD.n1583 DVDD.n1582 0.000854331
R18857 DVDD.n1590 DVDD.n1589 0.000854331
R18858 DVDD.n1598 DVDD.n1597 0.000854331
R18859 DVDD.n1605 DVDD.n1604 0.000854331
R18860 DVDD.n1611 DVDD.n1610 0.000854331
R18861 DVDD.n1617 DVDD.n1616 0.000854331
R18862 DVDD.n1618 DVDD.n1617 0.000854331
R18863 DVDD.n1624 DVDD.n1623 0.000854331
R18864 DVDD.n1631 DVDD.n1630 0.000854331
R18865 DVDD.n1639 DVDD.n1638 0.000854331
R18866 DVDD.n1653 DVDD.n1652 0.000854331
R18867 DVDD.n899 DVDD.n898 0.000854331
R18868 DVDD.n896 DVDD.n895 0.000854331
R18869 DVDD.n895 DVDD.n894 0.000854331
R18870 DVDD.n19273 DVDD.n19272 0.000854331
R18871 DVDD.n19278 DVDD.n19277 0.000854331
R18872 DVDD.n19281 DVDD.n19280 0.000854331
R18873 DVDD.n19321 DVDD.n19320 0.000854331
R18874 DVDD.n19312 DVDD.n19311 0.000854331
R18875 DVDD.n10167 DVDD.n10166 0.000854331
R18876 DVDD.n10170 DVDD.n10169 0.000854331
R18877 DVDD.n12140 DVDD.n12139 0.000854331
R18878 DVDD.n12145 DVDD.n12144 0.000854331
R18879 DVDD.n12167 DVDD.n12166 0.000854331
R18880 DVDD.n12232 DVDD.n12231 0.000854331
R18881 DVDD.n13433 DVDD.n13432 0.000854331
R18882 DVDD.n13698 DVDD.n13697 0.000854331
R18883 DVDD.n2719 DVDD.n2718 0.000854331
R18884 DVDD.n2760 DVDD.n2759 0.000854331
R18885 DVDD.n2800 DVDD.n2799 0.000854331
R18886 DVDD.n18674 DVDD.n18673 0.000854331
R18887 DVDD.n10059 DVDD.n10058 0.000854331
R18888 DVDD.n15471 DVDD.n15470 0.000854331
R18889 DVDD.n14732 DVDD.n14731 0.000854331
R18890 DVDD.n14649 DVDD.n14648 0.000854331
R18891 DVDD.n14391 DVDD.n14390 0.000854331
R18892 DVDD.n19693 DVDD.n19692 0.000854331
R18893 DVDD.n19708 DVDD.n19707 0.000854331
R18894 DVDD.n19769 DVDD.n19768 0.000854331
R18895 DVDD.n19839 DVDD.n19838 0.000854331
R18896 DVDD.n19861 DVDD.n19860 0.000854331
R18897 DVDD.n19994 DVDD.n19993 0.000854331
R18898 DVDD.n20008 DVDD.n20007 0.000854331
R18899 DVDD.n20052 DVDD.n20051 0.000854331
R18900 DVDD.n20196 DVDD.n20195 0.000854331
R18901 DVDD.n20183 DVDD.n20182 0.000854331
R18902 DVDD.n20180 DVDD.n20179 0.000854331
R18903 DVDD.n20094 DVDD.n20093 0.000854331
R18904 DVDD.n20108 DVDD.n20107 0.000854331
R18905 DVDD.n20111 DVDD.n20110 0.000854331
R18906 DVDD.n19077 DVDD.n19076 0.000854331
R18907 DVDD.n19054 DVDD.n19018 0.000854331
R18908 DVDD.n3860 DVDD.n3859 0.000854331
R18909 DVDD.n3872 DVDD.n3871 0.000854331
R18910 DVDD.n3874 DVDD.n3873 0.000854331
R18911 DVDD.n4679 DVDD.n4678 0.000854331
R18912 DVDD.n4682 DVDD.n4681 0.000854331
R18913 DVDD.n4705 DVDD.n4704 0.000854331
R18914 DVDD.n4775 DVDD.n4774 0.000854331
R18915 DVDD.n4906 DVDD.n4905 0.000854331
R18916 DVDD.n4909 DVDD.n4908 0.000854331
R18917 DVDD.n4919 DVDD.n4918 0.000854331
R18918 DVDD.n4949 DVDD.n4948 0.000854331
R18919 DVDD.n4955 DVDD.n4954 0.000854331
R18920 DVDD.n4993 DVDD.n4992 0.000854331
R18921 DVDD.n5006 DVDD.n5005 0.000854331
R18922 DVDD.n5024 DVDD.n5023 0.000854331
R18923 DVDD.n5091 DVDD.n5090 0.000854331
R18924 DVDD.n5188 DVDD.n5187 0.000854331
R18925 DVDD.n5338 DVDD.n5337 0.000854331
R18926 DVDD.n5386 DVDD.n5385 0.000854331
R18927 DVDD.n5411 DVDD.n5410 0.000854331
R18928 DVDD.n5428 DVDD.n5427 0.000854331
R18929 DVDD.n5434 DVDD.n5433 0.000854331
R18930 DVDD.n5457 DVDD.n5456 0.000854331
R18931 DVDD.n5581 DVDD.n5580 0.000854331
R18932 DVDD.n5585 DVDD.n5584 0.000854331
R18933 DVDD.n5677 DVDD.n5676 0.000854331
R18934 DVDD.n5679 DVDD.n5678 0.000854331
R18935 DVDD.n5953 DVDD.n5952 0.000854331
R18936 DVDD.n1338 DVDD.n1337 0.000854331
R18937 DVDD.n1353 DVDD.n1352 0.000854331
R18938 DVDD.n1357 DVDD.n1356 0.000854331
R18939 DVDD.n1414 DVDD.n1413 0.000854331
R18940 DVDD.n1537 DVDD.n1536 0.000854331
R18941 DVDD.n1515 DVDD.n1514 0.000854331
R18942 DVDD.n1682 DVDD.n1681 0.000854331
R18943 DVDD.n1696 DVDD.n1695 0.000854331
R18944 DVDD.n1721 DVDD.n1720 0.000854331
R18945 DVDD.n274 DVDD.n273 0.000854331
R18946 DVDD.n261 DVDD.n260 0.000854331
R18947 DVDD.n258 DVDD.n257 0.000854331
R18948 DVDD.n19192 DVDD.n19191 0.000854331
R18949 DVDD.n19206 DVDD.n19205 0.000854331
R18950 DVDD.n19209 DVDD.n19208 0.000854331
R18951 DVDD.n19459 DVDD.n19458 0.000854331
R18952 DVDD.n19436 DVDD.n19227 0.000854331
R18953 DVDD.n10107 DVDD.n10106 0.000854331
R18954 DVDD.n10119 DVDD.n10118 0.000854331
R18955 DVDD.n10121 DVDD.n10120 0.000854331
R18956 DVDD.n11386 DVDD.n11385 0.000854331
R18957 DVDD.n11389 DVDD.n11388 0.000854331
R18958 DVDD.n11412 DVDD.n11411 0.000854331
R18959 DVDD.n11601 DVDD.n11600 0.000854331
R18960 DVDD.n11847 DVDD.n11846 0.000854331
R18961 DVDD.n11844 DVDD.n11843 0.000854331
R18962 DVDD.n11834 DVDD.n11833 0.000854331
R18963 DVDD.n11804 DVDD.n11803 0.000854331
R18964 DVDD.n11798 DVDD.n11797 0.000854331
R18965 DVDD.n11760 DVDD.n11759 0.000854331
R18966 DVDD.n11748 DVDD.n11747 0.000854331
R18967 DVDD.n11730 DVDD.n11729 0.000854331
R18968 DVDD.n11663 DVDD.n11662 0.000854331
R18969 DVDD.n12368 DVDD.n12367 0.000854331
R18970 DVDD.n13121 DVDD.n13120 0.000854331
R18971 DVDD.n13075 DVDD.n13074 0.000854331
R18972 DVDD.n13051 DVDD.n13050 0.000854331
R18973 DVDD.n13035 DVDD.n13034 0.000854331
R18974 DVDD.n13029 DVDD.n13028 0.000854331
R18975 DVDD.n13025 DVDD.n13024 0.000854331
R18976 DVDD.n13006 DVDD.n13005 0.000854331
R18977 DVDD.n12846 DVDD.n12845 0.000854331
R18978 DVDD.n12842 DVDD.n12841 0.000854331
R18979 DVDD.n12764 DVDD.n12763 0.000854331
R18980 DVDD.n12762 DVDD.n12761 0.000854331
R18981 DVDD.n12616 DVDD.n12615 0.000854331
R18982 DVDD.n759 DVDD.n758 0.000854331
R18983 DVDD.n796 DVDD.n795 0.000854331
R18984 DVDD.n832 DVDD.n831 0.000854331
R18985 DVDD.n153 DVDD.n152 0.000854331
R18986 DVDD.n10091 DVDD.n10090 0.000854331
R18987 DVDD.n18138 DVDD.n18137 0.000854331
R18988 DVDD.n18083 DVDD.n18082 0.000854331
R18989 DVDD.n18005 DVDD.n18004 0.000854331
R18990 DVDD.n17769 DVDD.n17768 0.000854331
R18991 DVDD.n1915 DVDD.n1914 0.000854331
R18992 DVDD.n1930 DVDD.n1929 0.000854331
R18993 DVDD.n1934 DVDD.n1933 0.000854331
R18994 DVDD.n1991 DVDD.n1990 0.000854331
R18995 DVDD.n2061 DVDD.n2060 0.000854331
R18996 DVDD.n2083 DVDD.n2082 0.000854331
R18997 DVDD.n2215 DVDD.n2214 0.000854331
R18998 DVDD.n2229 DVDD.n2228 0.000854331
R18999 DVDD.n2273 DVDD.n2272 0.000854331
R19000 DVDD.n19581 DVDD.n19580 0.000854331
R19001 DVDD.n19568 DVDD.n19567 0.000854331
R19002 DVDD.n19565 DVDD.n19564 0.000854331
R19003 DVDD.n19479 DVDD.n19478 0.000854331
R19004 DVDD.n19493 DVDD.n19492 0.000854331
R19005 DVDD.n19496 DVDD.n19495 0.000854331
R19006 DVDD.n18969 DVDD.n18968 0.000854331
R19007 DVDD.n18946 DVDD.n18945 0.000854331
R19008 DVDD.n7081 DVDD.n7080 0.000854331
R19009 DVDD.n7093 DVDD.n7092 0.000854331
R19010 DVDD.n7095 DVDD.n7094 0.000854331
R19011 DVDD.n7005 DVDD.n7004 0.000854331
R19012 DVDD.n7002 DVDD.n7001 0.000854331
R19013 DVDD.n6979 DVDD.n6978 0.000854331
R19014 DVDD.n6909 DVDD.n6908 0.000854331
R19015 DVDD.n6778 DVDD.n6777 0.000854331
R19016 DVDD.n6775 DVDD.n6774 0.000854331
R19017 DVDD.n6765 DVDD.n6764 0.000854331
R19018 DVDD.n6735 DVDD.n6734 0.000854331
R19019 DVDD.n6729 DVDD.n6728 0.000854331
R19020 DVDD.n6691 DVDD.n6690 0.000854331
R19021 DVDD.n6678 DVDD.n6677 0.000854331
R19022 DVDD.n6660 DVDD.n6659 0.000854331
R19023 DVDD.n6591 DVDD.n6590 0.000854331
R19024 DVDD.n6494 DVDD.n6493 0.000854331
R19025 DVDD.n6423 DVDD.n6422 0.000854331
R19026 DVDD.n6375 DVDD.n6374 0.000854331
R19027 DVDD.n6350 DVDD.n6349 0.000854331
R19028 DVDD.n6333 DVDD.n6332 0.000854331
R19029 DVDD.n6327 DVDD.n6326 0.000854331
R19030 DVDD.n6323 DVDD.n6322 0.000854331
R19031 DVDD.n6304 DVDD.n6303 0.000854331
R19032 DVDD.n6226 DVDD.n6225 0.000854331
R19033 DVDD.n6222 DVDD.n6221 0.000854331
R19034 DVDD.n6146 DVDD.n6145 0.000854331
R19035 DVDD.n4412 DVDD.n4411 0.000854331
R19036 DVDD.n3265 DVDD.n3264 0.000854331
R19037 DVDD.n3250 DVDD.n3249 0.000854331
R19038 DVDD.n3246 DVDD.n3245 0.000854331
R19039 DVDD.n3189 DVDD.n3188 0.000854331
R19040 DVDD.n3460 DVDD.n3459 0.000854331
R19041 DVDD.n3482 DVDD.n3481 0.000854331
R19042 DVDD.n3567 DVDD.n3566 0.000854331
R19043 DVDD.n3553 DVDD.n2833 0.000854331
R19044 DVDD.n3717 DVDD.n3716 0.000854331
R19045 DVDD.n3760 DVDD.n3759 0.000854331
R19046 DVDD.n3747 DVDD.n3746 0.000854331
R19047 DVDD.n3744 DVDD.n3743 0.000854331
R19048 DVDD.n18496 DVDD.n18495 0.000854331
R19049 DVDD.n18510 DVDD.n18509 0.000854331
R19050 DVDD.n18513 DVDD.n18512 0.000854331
R19051 DVDD.n18806 DVDD.n18805 0.000854331
R19052 DVDD.n18783 DVDD.n18531 0.000854331
R19053 DVDD.n7139 DVDD.n7138 0.000854331
R19054 DVDD.n7151 DVDD.n7150 0.000854331
R19055 DVDD.n7153 DVDD.n7152 0.000854331
R19056 DVDD.n10022 DVDD.n10021 0.000854331
R19057 DVDD.n10019 DVDD.n10018 0.000854331
R19058 DVDD.n9996 DVDD.n9995 0.000854331
R19059 DVDD.n7857 DVDD.n7856 0.000854331
R19060 DVDD.n9746 DVDD.n9745 0.000854331
R19061 DVDD.n9743 DVDD.n9742 0.000854331
R19062 DVDD.n9733 DVDD.n9732 0.000854331
R19063 DVDD.n9703 DVDD.n9702 0.000854331
R19064 DVDD.n9697 DVDD.n9696 0.000854331
R19065 DVDD.n9659 DVDD.n9658 0.000854331
R19066 DVDD.n9646 DVDD.n9645 0.000854331
R19067 DVDD.n9628 DVDD.n9627 0.000854331
R19068 DVDD.n9559 DVDD.n9558 0.000854331
R19069 DVDD.n8389 DVDD.n8388 0.000854331
R19070 DVDD.n9209 DVDD.n9208 0.000854331
R19071 DVDD.n9161 DVDD.n9160 0.000854331
R19072 DVDD.n9136 DVDD.n9135 0.000854331
R19073 DVDD.n9119 DVDD.n9118 0.000854331
R19074 DVDD.n9113 DVDD.n9112 0.000854331
R19075 DVDD.n9109 DVDD.n9108 0.000854331
R19076 DVDD.n9090 DVDD.n9089 0.000854331
R19077 DVDD.n8928 DVDD.n8927 0.000854331
R19078 DVDD.n8924 DVDD.n8923 0.000854331
R19079 DVDD.n8848 DVDD.n8847 0.000854331
R19080 DVDD.n8686 DVDD.n8685 0.000854331
R19081 DVDD.n10564 DVDD.n10563 0.0008375
R19082 DVDD.n10567 DVDD.n10566 0.0008375
R19083 DVDD.n1824 DVDD.n1823 0.00083
R19084 DVDD.n19551 DVDD.n19550 0.00083
R19085 DVDD.n18858 DVDD.n18856 0.00083
R19086 DVDD.n7566 DVDD.n7565 0.00083
R19087 DVDD.n7573 DVDD.n7572 0.00083
R19088 DVDD.n19602 DVDD.n19601 0.00083
R19089 DVDD.n20166 DVDD.n20165 0.00083
R19090 DVDD.n19107 DVDD.n19106 0.00083
R19091 DVDD.n7522 DVDD.n7521 0.00083
R19092 DVDD.n7529 DVDD.n7528 0.00083
R19093 DVDD.n7359 DVDD.n7358 0.00083
R19094 DVDD.n7409 DVDD.n7407 0.00083
R19095 DVDD.n7590 DVDD.n7589 0.00083
R19096 DVDD.n81 DVDD.n80 0.00083
R19097 DVDD.n7457 DVDD.n7455 0.00083
R19098 DVDD.n7546 DVDD.n7545 0.00083
R19099 DVDD.n7232 DVDD.n7231 0.00083
R19100 DVDD.n7494 DVDD.n7492 0.00083
R19101 DVDD.n7192 DVDD.n7191 0.00083
R19102 DVDD.n847 DVDD.n846 0.00083
R19103 DVDD.n223 DVDD.n222 0.00083
R19104 DVDD.n219 DVDD.n218 0.00083
R19105 DVDD.n215 DVDD.n214 0.00083
R19106 DVDD.n210 DVDD.n209 0.00083
R19107 DVDD.n19382 DVDD.n19381 0.00083
R19108 DVDD.n19356 DVDD.n19355 0.00083
R19109 DVDD.n10184 DVDD.n10086 0.00083
R19110 DVDD.n18253 DVDD.n18252 0.00083
R19111 DVDD.n10519 DVDD.n10518 0.00083
R19112 DVDD.n14954 DVDD.n14953 0.00083
R19113 DVDD.n15056 DVDD.n15055 0.00083
R19114 DVDD.n17126 DVDD.n17125 0.00083
R19115 DVDD.n11012 DVDD.n11011 0.00083
R19116 DVDD.n11034 DVDD.n11033 0.00083
R19117 DVDD.n11089 DVDD.n11088 0.00083
R19118 DVDD.n11187 DVDD.n11186 0.00083
R19119 DVDD.n11138 DVDD.n11137 0.00083
R19120 DVDD.n17017 DVDD.n17016 0.00083
R19121 DVDD.n16143 DVDD.n16142 0.00083
R19122 DVDD.n16169 DVDD.n16168 0.00083
R19123 DVDD.n16288 DVDD.n16287 0.00083
R19124 DVDD.n16333 DVDD.n16332 0.00083
R19125 DVDD.n16348 DVDD.n16347 0.00083
R19126 DVDD.n16228 DVDD.n16227 0.00083
R19127 DVDD.n15593 DVDD.n15592 0.00083
R19128 DVDD.n15909 DVDD.n15908 0.00083
R19129 DVDD.n3611 DVDD.n3610 0.00083
R19130 DVDD.n18606 DVDD.n18605 0.00083
R19131 DVDD.n18617 DVDD.n18616 0.00083
R19132 DVDD.n18621 DVDD.n18620 0.00083
R19133 DVDD.n18633 DVDD.n18632 0.00083
R19134 DVDD.n18378 DVDD.n18377 0.00083
R19135 DVDD.n18335 DVDD.n18334 0.00083
R19136 DVDD.n14742 DVDD.n7134 0.00083
R19137 DVDD.n14778 DVDD.n14777 0.00083
R19138 DVDD.n20271 DVDD.n20270 0.00083
R19139 DVDD.n7325 DVDD.n7323 0.00083
R19140 DVDD.n7683 DVDD.n7682 0.00083
R19141 DVDD.n502 DVDD.n501 0.000821429
R19142 DVDD.n497 DVDD.n496 0.000821429
R19143 DVDD.n732 DVDD.n731 0.000821429
R19144 DVDD.n729 DVDD.n728 0.000821429
R19145 DVDD.n16391 DVDD.n16390 0.00082
R19146 DVDD.n15181 DVDD.n15180 0.00082
R19147 DVDD.n3826 DVDD.n3825 0.000812862
R19148 DVDD.n111 DVDD.n110 0.000812862
R19149 DVDD.n1825 DVDD.n1824 0.0008
R19150 DVDD.n19524 DVDD.n19523 0.0008
R19151 DVDD.n19513 DVDD.n19512 0.0008
R19152 DVDD.n18886 DVDD.n18885 0.0008
R19153 DVDD.n18878 DVDD.n18877 0.0008
R19154 DVDD.n19603 DVDD.n19602 0.0008
R19155 DVDD.n20139 DVDD.n20138 0.0008
R19156 DVDD.n20128 DVDD.n20127 0.0008
R19157 DVDD.n19135 DVDD.n19134 0.0008
R19158 DVDD.n19127 DVDD.n19126 0.0008
R19159 DVDD.n7379 DVDD.n7377 0.0008
R19160 DVDD.n61 DVDD.n59 0.0008
R19161 DVDD.n7252 DVDD.n7250 0.0008
R19162 DVDD.n190 DVDD.n189 0.0008
R19163 DVDD.n19354 DVDD.n19353 0.0008
R19164 DVDD.n19407 DVDD.n19406 0.0008
R19165 DVDD.n19402 DVDD.n19401 0.0008
R19166 DVDD.n18255 DVDD.n18254 0.0008
R19167 DVDD.n14974 DVDD.n14972 0.0008
R19168 DVDD.n15051 DVDD.n15049 0.0008
R19169 DVDD.n15383 DVDD.n15381 0.0008
R19170 DVDD.n15341 DVDD.n14828 0.0008
R19171 DVDD.n10428 DVDD.n10427 0.0008
R19172 DVDD.n14975 DVDD.n14971 0.0008
R19173 DVDD.n15052 DVDD.n15048 0.0008
R19174 DVDD.n15055 DVDD.n15054 0.0008
R19175 DVDD.n15385 DVDD.n15384 0.0008
R19176 DVDD.n15343 DVDD.n15342 0.0008
R19177 DVDD.n17060 DVDD.n17059 0.0008
R19178 DVDD.n11030 DVDD.n11029 0.0008
R19179 DVDD.n11085 DVDD.n11084 0.0008
R19180 DVDD.n11088 DVDD.n11087 0.0008
R19181 DVDD.n11194 DVDD.n11193 0.0008
R19182 DVDD.n11148 DVDD.n11147 0.0008
R19183 DVDD.n16937 DVDD.n16936 0.0008
R19184 DVDD.n16165 DVDD.n16164 0.0008
R19185 DVDD.n16283 DVDD.n16282 0.0008
R19186 DVDD.n16287 DVDD.n16286 0.0008
R19187 DVDD.n16329 DVDD.n16326 0.0008
R19188 DVDD.n16353 DVDD.n16352 0.0008
R19189 DVDD.n16224 DVDD.n16220 0.0008
R19190 DVDD.n15589 DVDD.n15585 0.0008
R19191 DVDD.n15738 DVDD.n15737 0.0008
R19192 DVDD.n15699 DVDD.n15695 0.0008
R19193 DVDD.n15804 DVDD.n15800 0.0008
R19194 DVDD.n15867 DVDD.n15863 0.0008
R19195 DVDD.n16097 DVDD.n16096 0.0008
R19196 DVDD.n15911 DVDD.n15907 0.0008
R19197 DVDD.n15803 DVDD.n15801 0.0008
R19198 DVDD.n15866 DVDD.n15864 0.0008
R19199 DVDD.n16095 DVDD.n16093 0.0008
R19200 DVDD.n15912 DVDD.n15904 0.0008
R19201 DVDD.n16223 DVDD.n16221 0.0008
R19202 DVDD.n15588 DVDD.n15586 0.0008
R19203 DVDD.n15736 DVDD.n15734 0.0008
R19204 DVDD.n15698 DVDD.n15696 0.0008
R19205 DVDD.n16172 DVDD.n16171 0.0008
R19206 DVDD.n16292 DVDD.n16291 0.0008
R19207 DVDD.n16351 DVDD.n16343 0.0008
R19208 DVDD.n11036 DVDD.n11035 0.0008
R19209 DVDD.n11093 DVDD.n11092 0.0008
R19210 DVDD.n11192 DVDD.n11190 0.0008
R19211 DVDD.n11146 DVDD.n11125 0.0008
R19212 DVDD.n18732 DVDD.n18731 0.0008
R19213 DVDD.n18451 DVDD.n18450 0.0008
R19214 DVDD.n18414 DVDD.n18413 0.0008
R19215 DVDD.n18409 DVDD.n18408 0.0008
R19216 DVDD.n14780 DVDD.n14779 0.0008
R19217 DVDD.n20251 DVDD.n20249 0.0008
R19218 DVDD.n15252 DVDD.n15251 0.000788154
R19219 DVDD.n15268 DVDD.n15267 0.000788154
R19220 DVDD.n15289 DVDD.n15288 0.000788154
R19221 DVDD.n10643 DVDD.n10642 0.00078125
R19222 DVDD.n10640 DVDD.n10639 0.00078125
R19223 DVDD.n3678 DVDD.n3677 0.00077
R19224 DVDD.n3707 DVDD.n3706 0.00077
R19225 DVDD.n18553 DVDD.n18552 0.00077
R19226 DVDD.n2997 DVDD.n2996 0.00077
R19227 DVDD.n2920 DVDD.n2919 0.00077
R19228 DVDD.n2933 DVDD.n2932 0.00077
R19229 DVDD.n2937 DVDD.n2936 0.00077
R19230 DVDD.n7158 DVDD.n7157 0.00077
R19231 DVDD.n9386 DVDD.n9385 0.00077
R19232 DVDD.n9383 DVDD.n9382 0.00077
R19233 DVDD.n9380 DVDD.n9379 0.00077
R19234 DVDD.n9377 DVDD.n9376 0.00077
R19235 DVDD.n9374 DVDD.n9373 0.00077
R19236 DVDD.n9371 DVDD.n9370 0.00077
R19237 DVDD.n9368 DVDD.n9367 0.00077
R19238 DVDD.n9365 DVDD.n9364 0.00077
R19239 DVDD.n2026 DVDD.n2025 0.00077
R19240 DVDD.n2158 DVDD.n2157 0.00077
R19241 DVDD.n2171 DVDD.n2170 0.00077
R19242 DVDD.n2175 DVDD.n2174 0.00077
R19243 DVDD.n2234 DVDD.n2233 0.00077
R19244 DVDD.n2263 DVDD.n2262 0.00077
R19245 DVDD.n18922 DVDD.n18921 0.00077
R19246 DVDD.n6940 DVDD.n6939 0.00077
R19247 DVDD.n1887 DVDD.n1886 0.00077
R19248 DVDD.n19804 DVDD.n19803 0.00077
R19249 DVDD.n19937 DVDD.n19936 0.00077
R19250 DVDD.n19950 DVDD.n19949 0.00077
R19251 DVDD.n19954 DVDD.n19953 0.00077
R19252 DVDD.n20013 DVDD.n20012 0.00077
R19253 DVDD.n20042 DVDD.n20041 0.00077
R19254 DVDD.n19040 DVDD.n19039 0.00077
R19255 DVDD.n4714 DVDD.n4713 0.00077
R19256 DVDD.n19665 DVDD.n19664 0.00077
R19257 DVDD.n1093 DVDD.n1092 0.00077
R19258 DVDD.n1008 DVDD.n1007 0.00077
R19259 DVDD.n995 DVDD.n994 0.00077
R19260 DVDD.n991 DVDD.n990 0.00077
R19261 DVDD.n1729 DVDD.n1728 0.00077
R19262 DVDD.n950 DVDD.n949 0.00077
R19263 DVDD.n19249 DVDD.n19248 0.00077
R19264 DVDD.n11419 DVDD.n11417 0.00077
R19265 DVDD.n19540 DVDD.n19539 0.00077
R19266 DVDD.n19520 DVDD.n19519 0.00077
R19267 DVDD.n19505 DVDD.n19504 0.00077
R19268 DVDD.n20155 DVDD.n20154 0.00077
R19269 DVDD.n20135 DVDD.n20134 0.00077
R19270 DVDD.n20120 DVDD.n20119 0.00077
R19271 DVDD.n7383 DVDD.n7382 0.00077
R19272 DVDD.n57 DVDD.n56 0.00077
R19273 DVDD.n7256 DVDD.n7255 0.00077
R19274 DVDD.n251 DVDD.n250 0.00077
R19275 DVDD.n235 DVDD.n234 0.00077
R19276 DVDD.n209 DVDD.n208 0.00077
R19277 DVDD.n185 DVDD.n184 0.00077
R19278 DVDD.n165 DVDD.n164 0.00077
R19279 DVDD.n19344 DVDD.n19343 0.00077
R19280 DVDD.n19348 DVDD.n19347 0.00077
R19281 DVDD.n19405 DVDD.n19404 0.00077
R19282 DVDD.n19362 DVDD.n19361 0.00077
R19283 DVDD.n18333 DVDD.n10086 0.00077
R19284 DVDD.n18239 DVDD.n18238 0.00077
R19285 DVDD.n18262 DVDD.n18261 0.00077
R19286 DVDD.n18259 DVDD.n18258 0.00077
R19287 DVDD.n18258 DVDD.n18257 0.00077
R19288 DVDD.n18250 DVDD.n18249 0.00077
R19289 DVDD.n1310 DVDD.n1309 0.00077
R19290 DVDD.n10350 DVDD.n10349 0.00077
R19291 DVDD.n10355 DVDD.n10354 0.00077
R19292 DVDD.n10654 DVDD.n10540 0.00077
R19293 DVDD.n15364 DVDD.n15363 0.00077
R19294 DVDD.n15355 DVDD.n15354 0.00077
R19295 DVDD.n13297 DVDD.n13296 0.00077
R19296 DVDD.n13294 DVDD.n13293 0.00077
R19297 DVDD.n13291 DVDD.n13290 0.00077
R19298 DVDD.n13288 DVDD.n13287 0.00077
R19299 DVDD.n13285 DVDD.n13284 0.00077
R19300 DVDD.n13282 DVDD.n13281 0.00077
R19301 DVDD.n13279 DVDD.n13278 0.00077
R19302 DVDD.n13276 DVDD.n13275 0.00077
R19303 DVDD.n16505 DVDD.n16504 0.00077
R19304 DVDD.n16509 DVDD.n16508 0.00077
R19305 DVDD.n17152 DVDD.n17151 0.00077
R19306 DVDD.n11169 DVDD.n11168 0.00077
R19307 DVDD.n11162 DVDD.n11161 0.00077
R19308 DVDD.n16847 DVDD.n16846 0.00077
R19309 DVDD.n16851 DVDD.n16850 0.00077
R19310 DVDD.n17043 DVDD.n17042 0.00077
R19311 DVDD.n16372 DVDD.n16371 0.00077
R19312 DVDD.n16366 DVDD.n16365 0.00077
R19313 DVDD.n16816 DVDD.n16815 0.00077
R19314 DVDD.n16694 DVDD.n16693 0.00077
R19315 DVDD.n3293 DVDD.n3292 0.00077
R19316 DVDD.n18566 DVDD.n18565 0.00077
R19317 DVDD.n18587 DVDD.n18586 0.00077
R19318 DVDD.n18634 DVDD.n18633 0.00077
R19319 DVDD.n18727 DVDD.n18726 0.00077
R19320 DVDD.n18686 DVDD.n18685 0.00077
R19321 DVDD.n18461 DVDD.n18460 0.00077
R19322 DVDD.n18457 DVDD.n18456 0.00077
R19323 DVDD.n18412 DVDD.n18411 0.00077
R19324 DVDD.n18358 DVDD.n18357 0.00077
R19325 DVDD.n18333 DVDD.n7134 0.00077
R19326 DVDD.n14799 DVDD.n14798 0.00077
R19327 DVDD.n14787 DVDD.n14786 0.00077
R19328 DVDD.n14784 DVDD.n14783 0.00077
R19329 DVDD.n14783 DVDD.n14782 0.00077
R19330 DVDD.n14775 DVDD.n14774 0.00077
R19331 DVDD.n20247 DVDD.n20246 0.00077
R19332 DVDD.n11262 DVDD.n11261 0.000757143
R19333 DVDD.n11250 DVDD.n11249 0.000757143
R19334 DVDD.n11234 DVDD.n11233 0.000757143
R19335 DVDD.n5768 DVDD.n5767 0.000757143
R19336 DVDD.n300 DVDD.n299 0.000757143
R19337 DVDD.n412 DVDD.n411 0.000757143
R19338 DVDD.n485 DVDD.n484 0.000757143
R19339 DVDD.n439 DVDD.n438 0.000757143
R19340 DVDD.n385 DVDD.n384 0.000757143
R19341 DVDD.n414 DVDD.n413 0.000757143
R19342 DVDD.n486 DVDD.n483 0.000757143
R19343 DVDD.n440 DVDD.n437 0.000757143
R19344 DVDD.n531 DVDD.n530 0.000757143
R19345 DVDD.n643 DVDD.n642 0.000757143
R19346 DVDD.n717 DVDD.n716 0.000757143
R19347 DVDD.n671 DVDD.n670 0.000757143
R19348 DVDD.n616 DVDD.n615 0.000757143
R19349 DVDD.n645 DVDD.n644 0.000757143
R19350 DVDD.n718 DVDD.n715 0.000757143
R19351 DVDD.n672 DVDD.n669 0.000757143
R19352 DVDD.n11296 DVDD.n11295 0.000757143
R19353 DVDD.n11278 DVDD.n11277 0.000757143
R19354 DVDD.n12502 DVDD.n12501 0.000757143
R19355 DVDD.n5769 DVDD.n5765 0.000757143
R19356 DVDD.n8295 DVDD.n8294 0.000743243
R19357 DVDD.n1837 DVDD.n1836 0.00074
R19358 DVDD.n19559 DVDD.n19558 0.00074
R19359 DVDD.n19555 DVDD.n19554 0.00074
R19360 DVDD.n19550 DVDD.n19549 0.00074
R19361 DVDD.n19547 DVDD.n19546 0.00074
R19362 DVDD.n19536 DVDD.n19535 0.00074
R19363 DVDD.n18867 DVDD.n18866 0.00074
R19364 DVDD.n18866 DVDD.n18865 0.00074
R19365 DVDD.n18864 DVDD.n18863 0.00074
R19366 DVDD.n18333 DVDD.n7110 0.00074
R19367 DVDD.n3920 DVDD.n3919 0.00074
R19368 DVDD.n19615 DVDD.n19614 0.00074
R19369 DVDD.n20174 DVDD.n20173 0.00074
R19370 DVDD.n20170 DVDD.n20169 0.00074
R19371 DVDD.n20165 DVDD.n20164 0.00074
R19372 DVDD.n20162 DVDD.n20161 0.00074
R19373 DVDD.n20151 DVDD.n20150 0.00074
R19374 DVDD.n19116 DVDD.n19115 0.00074
R19375 DVDD.n19115 DVDD.n19114 0.00074
R19376 DVDD.n19113 DVDD.n19112 0.00074
R19377 DVDD.n18333 DVDD.n3890 0.00074
R19378 DVDD.n4607 DVDD.n4606 0.00074
R19379 DVDD.n7355 DVDD.n7353 0.00074
R19380 DVDD.n7371 DVDD.n7370 0.00074
R19381 DVDD.n7594 DVDD.n7592 0.00074
R19382 DVDD.n85 DVDD.n83 0.00074
R19383 DVDD.n69 DVDD.n68 0.00074
R19384 DVDD.n7550 DVDD.n7548 0.00074
R19385 DVDD.n7228 DVDD.n7226 0.00074
R19386 DVDD.n7244 DVDD.n7243 0.00074
R19387 DVDD.n7196 DVDD.n7194 0.00074
R19388 DVDD.n863 DVDD.n862 0.00074
R19389 DVDD.n233 DVDD.n232 0.00074
R19390 DVDD.n222 DVDD.n221 0.00074
R19391 DVDD.n218 DVDD.n217 0.00074
R19392 DVDD.n216 DVDD.n215 0.00074
R19393 DVDD.n175 DVDD.n174 0.00074
R19394 DVDD.n19397 DVDD.n19396 0.00074
R19395 DVDD.n19391 DVDD.n19390 0.00074
R19396 DVDD.n18242 DVDD.n18241 0.00074
R19397 DVDD.n3627 DVDD.n3626 0.00074
R19398 DVDD.n18589 DVDD.n18588 0.00074
R19399 DVDD.n18607 DVDD.n18606 0.00074
R19400 DVDD.n18618 DVDD.n18617 0.00074
R19401 DVDD.n18620 DVDD.n18619 0.00074
R19402 DVDD.n18710 DVDD.n18702 0.00074
R19403 DVDD.n18404 DVDD.n18403 0.00074
R19404 DVDD.n18398 DVDD.n18397 0.00074
R19405 DVDD.n18334 DVDD.n18333 0.00074
R19406 DVDD.n14796 DVDD.n14795 0.00074
R19407 DVDD.n20275 DVDD.n20273 0.00074
R19408 DVDD.n20259 DVDD.n20258 0.00074
R19409 DVDD.n7679 DVDD.n7677 0.00074
R19410 DVDD.n3809 DVDD.n3808 0.000725
R19411 DVDD.n18994 DVDD.n18993 0.000725
R19412 DVDD.n7217 DVDD.n7216 0.000725
R19413 DVDD.n10073 DVDD.n10072 0.000725
R19414 DVDD.n7116 DVDD.n7115 0.000725
R19415 DVDD.n1809 DVDD.n1808 0.000725
R19416 DVDD.n2818 DVDD.n2817 0.000725
R19417 DVDD.n14845 DVDD.n14844 0.000725
R19418 DVDD.n15076 DVDD.n15075 0.000725
R19419 DVDD.n10478 DVDD.n10477 0.000725
R19420 DVDD.n10671 DVDD.n10670 0.000725
R19421 DVDD.n10683 DVDD.n10682 0.000725
R19422 DVDD.n10694 DVDD.n10693 0.000725
R19423 DVDD.n10597 DVDD.n10596 0.000725
R19424 DVDD.n10400 DVDD.n10399 0.000725
R19425 DVDD.n10569 DVDD.n10568 0.000725
R19426 DVDD.n10591 DVDD.n10590 0.000725
R19427 DVDD.n7288 DVDD.n7287 0.000725
R19428 DVDD.n1823 DVDD.n1822 0.00071
R19429 DVDD.n1826 DVDD.n1825 0.00071
R19430 DVDD.n1838 DVDD.n1837 0.00071
R19431 DVDD.n1840 DVDD.n1839 0.00071
R19432 DVDD.n19544 DVDD.n19543 0.00071
R19433 DVDD.n19530 DVDD.n19529 0.00071
R19434 DVDD.n19528 DVDD.n19527 0.00071
R19435 DVDD.n19517 DVDD.n19516 0.00071
R19436 DVDD.n19514 DVDD.n19513 0.00071
R19437 DVDD.n18880 DVDD.n18879 0.00071
R19438 DVDD.n18848 DVDD.n18847 0.00071
R19439 DVDD.n19601 DVDD.n19600 0.00071
R19440 DVDD.n19604 DVDD.n19603 0.00071
R19441 DVDD.n19616 DVDD.n19615 0.00071
R19442 DVDD.n19618 DVDD.n19617 0.00071
R19443 DVDD.n20159 DVDD.n20158 0.00071
R19444 DVDD.n20145 DVDD.n20144 0.00071
R19445 DVDD.n20143 DVDD.n20142 0.00071
R19446 DVDD.n20132 DVDD.n20131 0.00071
R19447 DVDD.n20129 DVDD.n20128 0.00071
R19448 DVDD.n19129 DVDD.n19128 0.00071
R19449 DVDD.n19096 DVDD.n19095 0.00071
R19450 DVDD.n7367 DVDD.n7365 0.00071
R19451 DVDD.n7417 DVDD.n7416 0.00071
R19452 DVDD.n73 DVDD.n71 0.00071
R19453 DVDD.n7465 DVDD.n7464 0.00071
R19454 DVDD.n7240 DVDD.n7238 0.00071
R19455 DVDD.n7486 DVDD.n7485 0.00071
R19456 DVDD.n7185 DVDD.n7177 0.00071
R19457 DVDD.n846 DVDD.n845 0.00071
R19458 DVDD.n848 DVDD.n847 0.00071
R19459 DVDD.n850 DVDD.n849 0.00071
R19460 DVDD.n1783 DVDD.n863 0.00071
R19461 DVDD.n1785 DVDD.n1784 0.00071
R19462 DVDD.n1791 DVDD.n1790 0.00071
R19463 DVDD.n20215 DVDD.n254 0.00071
R19464 DVDD.n249 DVDD.n235 0.00071
R19465 DVDD.n228 DVDD.n227 0.00071
R19466 DVDD.n220 DVDD.n219 0.00071
R19467 DVDD.n214 DVDD.n213 0.00071
R19468 DVDD.n211 DVDD.n210 0.00071
R19469 DVDD.n204 DVDD.n203 0.00071
R19470 DVDD.n197 DVDD.n196 0.00071
R19471 DVDD.n195 DVDD.n194 0.00071
R19472 DVDD.n193 DVDD.n192 0.00071
R19473 DVDD.n181 DVDD.n180 0.00071
R19474 DVDD.n177 DVDD.n176 0.00071
R19475 DVDD.n172 DVDD.n171 0.00071
R19476 DVDD.n168 DVDD.n167 0.00071
R19477 DVDD.n144 DVDD.n143 0.00071
R19478 DVDD.n19340 DVDD.n19164 0.00071
R19479 DVDD.n19409 DVDD.n19408 0.00071
R19480 DVDD.n19392 DVDD.n19391 0.00071
R19481 DVDD.n19388 DVDD.n19387 0.00071
R19482 DVDD.n19373 DVDD.n19372 0.00071
R19483 DVDD.n15054 DVDD.n15053 0.00071
R19484 DVDD.n15057 DVDD.n15056 0.00071
R19485 DVDD.n15348 DVDD.n15347 0.00071
R19486 DVDD.n15345 DVDD.n15344 0.00071
R19487 DVDD.n11087 DVDD.n11086 0.00071
R19488 DVDD.n11090 DVDD.n11089 0.00071
R19489 DVDD.n16359 DVDD.n16358 0.00071
R19490 DVDD.n16355 DVDD.n16354 0.00071
R19491 DVDD.n3610 DVDD.n3609 0.00071
R19492 DVDD.n3612 DVDD.n3611 0.00071
R19493 DVDD.n3614 DVDD.n3613 0.00071
R19494 DVDD.n3650 DVDD.n3627 0.00071
R19495 DVDD.n3649 DVDD.n3648 0.00071
R19496 DVDD.n3643 DVDD.n3642 0.00071
R19497 DVDD.n20215 DVDD.n2301 0.00071
R19498 DVDD.n18586 DVDD.n18580 0.00071
R19499 DVDD.n18601 DVDD.n18593 0.00071
R19500 DVDD.n18616 DVDD.n18608 0.00071
R19501 DVDD.n18622 DVDD.n18621 0.00071
R19502 DVDD.n18632 DVDD.n18624 0.00071
R19503 DVDD.n18649 DVDD.n18638 0.00071
R19504 DVDD.n18656 DVDD.n18655 0.00071
R19505 DVDD.n18658 DVDD.n18657 0.00071
R19506 DVDD.n18735 DVDD.n18734 0.00071
R19507 DVDD.n18716 DVDD.n18715 0.00071
R19508 DVDD.n18712 DVDD.n18711 0.00071
R19509 DVDD.n18700 DVDD.n18699 0.00071
R19510 DVDD.n18696 DVDD.n18688 0.00071
R19511 DVDD.n18660 DVDD.n18659 0.00071
R19512 DVDD.n18468 DVDD.n18467 0.00071
R19513 DVDD.n18416 DVDD.n18415 0.00071
R19514 DVDD.n18399 DVDD.n18398 0.00071
R19515 DVDD.n18395 DVDD.n18383 0.00071
R19516 DVDD.n18369 DVDD.n18368 0.00071
R19517 DVDD.n20263 DVDD.n20261 0.00071
R19518 DVDD.n7333 DVDD.n7332 0.00071
R19519 DVDD.n7689 DVDD.n7176 0.00071
R19520 DVDD.n18984 DVDD.n18983 0.000708575
R19521 DVDD.n3835 DVDD.n3834 0.000708575
R19522 DVDD.n120 DVDD.n119 0.000708575
R19523 DVDD.n10551 DVDD.n10550 0.000708575
R19524 DVDD.n3096 DVDD.n3095 0.000700893
R19525 DVDD.n3049 DVDD.n3048 0.000700893
R19526 DVDD.n381 DVDD.n380 0.000692857
R19527 DVDD.n408 DVDD.n407 0.000692857
R19528 DVDD.n489 DVDD.n488 0.000692857
R19529 DVDD.n443 DVDD.n442 0.000692857
R19530 DVDD.n612 DVDD.n611 0.000692857
R19531 DVDD.n639 DVDD.n638 0.000692857
R19532 DVDD.n721 DVDD.n720 0.000692857
R19533 DVDD.n675 DVDD.n674 0.000692857
R19534 DVDD.n13730 DVDD.n13729 0.000692857
R19535 DVDD.n11281 DVDD.n11280 0.000692857
R19536 DVDD.n12504 DVDD.n12492 0.000692857
R19537 DVDD.n5771 DVDD.n5746 0.000692857
R19538 DVDD.n15198 DVDD.n15197 0.000692102
R19539 DVDD.n15269 DVDD.n15268 0.000692102
R19540 DVDD.n15277 DVDD.n15275 0.000692102
R19541 DVDD.n16057 DVDD.n16056 0.000688285
R19542 DVDD.n15994 DVDD.n15993 0.000688285
R19543 DVDD.n15669 DVDD.n15668 0.000688285
R19544 DVDD.n15938 DVDD.n15937 0.000688285
R19545 DVDD.n8287 DVDD.n8286 0.000688285
R19546 DVDD.n8279 DVDD.n8278 0.000688285
R19547 DVDD.n8271 DVDD.n8270 0.000688285
R19548 DVDD.n8265 DVDD.n8264 0.000688285
R19549 DVDD.n8259 DVDD.n8258 0.000688285
R19550 DVDD.n8250 DVDD.n8249 0.000688285
R19551 DVDD.n8241 DVDD.n8240 0.000688285
R19552 DVDD.n8232 DVDD.n8231 0.000688285
R19553 DVDD.n8224 DVDD.n8223 0.000688285
R19554 DVDD.n8216 DVDD.n8215 0.000688285
R19555 DVDD.n8208 DVDD.n8207 0.000688285
R19556 DVDD.n8202 DVDD.n8201 0.000688285
R19557 DVDD.n8196 DVDD.n8195 0.000688285
R19558 DVDD.n8187 DVDD.n8186 0.000688285
R19559 DVDD.n8174 DVDD.n8173 0.000688285
R19560 DVDD.n9395 DVDD.n9394 0.000688285
R19561 DVDD.n9394 DVDD.n9393 0.000688285
R19562 DVDD.n9392 DVDD.n8360 0.000688285
R19563 DVDD.n7963 DVDD.n7962 0.000688285
R19564 DVDD.n8094 DVDD.n8093 0.000688285
R19565 DVDD.n7740 DVDD.n7739 0.00068
R19566 DVDD.n7738 DVDD.n7737 0.00068
R19567 DVDD.n7734 DVDD.n7733 0.00068
R19568 DVDD.n7765 DVDD.n7764 0.00068
R19569 DVDD.n7763 DVDD.n7762 0.00068
R19570 DVDD.n3456 DVDD.n3455 0.00068
R19571 DVDD.n3571 DVDD.n3570 0.00068
R19572 DVDD.n2904 DVDD.n2903 0.00068
R19573 DVDD.n2901 DVDD.n2900 0.00068
R19574 DVDD.n2898 DVDD.n2897 0.00068
R19575 DVDD.n2895 DVDD.n2894 0.00068
R19576 DVDD.n2892 DVDD.n2891 0.00068
R19577 DVDD.n2889 DVDD.n2888 0.00068
R19578 DVDD.n2886 DVDD.n2885 0.00068
R19579 DVDD.n2883 DVDD.n2882 0.00068
R19580 DVDD.n2880 DVDD.n2879 0.00068
R19581 DVDD.n2877 DVDD.n2876 0.00068
R19582 DVDD.n2874 DVDD.n2873 0.00068
R19583 DVDD.n9962 DVDD.n9961 0.00068
R19584 DVDD.n9761 DVDD.n9760 0.00068
R19585 DVDD.n9775 DVDD.n9774 0.00068
R19586 DVDD.n9792 DVDD.n9791 0.00068
R19587 DVDD.n9886 DVDD.n9885 0.00068
R19588 DVDD.n7911 DVDD.n7910 0.00068
R19589 DVDD.n9486 DVDD.n9485 0.00068
R19590 DVDD.n9251 DVDD.n9250 0.00068
R19591 DVDD.n9276 DVDD.n9275 0.00068
R19592 DVDD.n9293 DVDD.n9292 0.00068
R19593 DVDD.n9307 DVDD.n9306 0.00068
R19594 DVDD.n9391 DVDD.n9390 0.00068
R19595 DVDD.n2057 DVDD.n2056 0.00068
R19596 DVDD.n2211 DVDD.n2210 0.00068
R19597 DVDD.n7100 DVDD.n7097 0.00068
R19598 DVDD.n7102 DVDD.n7101 0.00068
R19599 DVDD.n7035 DVDD.n7034 0.00068
R19600 DVDD.n6945 DVDD.n6944 0.00068
R19601 DVDD.n6854 DVDD.n6853 0.00068
R19602 DVDD.n6840 DVDD.n6839 0.00068
R19603 DVDD.n6823 DVDD.n6822 0.00068
R19604 DVDD.n6544 DVDD.n6543 0.00068
R19605 DVDD.n1864 DVDD.n1863 0.00068
R19606 DVDD.n3991 DVDD.n3990 0.00068
R19607 DVDD.n3966 DVDD.n3965 0.00068
R19608 DVDD.n3949 DVDD.n3948 0.00068
R19609 DVDD.n3935 DVDD.n3934 0.00068
R19610 DVDD.n19835 DVDD.n19834 0.00068
R19611 DVDD.n19990 DVDD.n19989 0.00068
R19612 DVDD.n3879 DVDD.n3876 0.00068
R19613 DVDD.n3881 DVDD.n3880 0.00068
R19614 DVDD.n4615 DVDD.n4614 0.00068
R19615 DVDD.n4719 DVDD.n4718 0.00068
R19616 DVDD.n4891 DVDD.n4890 0.00068
R19617 DVDD.n4877 DVDD.n4876 0.00068
R19618 DVDD.n4860 DVDD.n4859 0.00068
R19619 DVDD.n5135 DVDD.n5134 0.00068
R19620 DVDD.n19642 DVDD.n19641 0.00068
R19621 DVDD.n5296 DVDD.n5295 0.00068
R19622 DVDD.n5271 DVDD.n5270 0.00068
R19623 DVDD.n5254 DVDD.n5253 0.00068
R19624 DVDD.n5240 DVDD.n5239 0.00068
R19625 DVDD.n1541 DVDD.n1540 0.00068
R19626 DVDD.n1678 DVDD.n1677 0.00068
R19627 DVDD.n1024 DVDD.n1023 0.00068
R19628 DVDD.n1027 DVDD.n1026 0.00068
R19629 DVDD.n1030 DVDD.n1029 0.00068
R19630 DVDD.n1033 DVDD.n1032 0.00068
R19631 DVDD.n1036 DVDD.n1035 0.00068
R19632 DVDD.n1039 DVDD.n1038 0.00068
R19633 DVDD.n1042 DVDD.n1041 0.00068
R19634 DVDD.n1045 DVDD.n1044 0.00068
R19635 DVDD.n1048 DVDD.n1047 0.00068
R19636 DVDD.n1051 DVDD.n1050 0.00068
R19637 DVDD.n1054 DVDD.n1053 0.00068
R19638 DVDD.n11545 DVDD.n11544 0.00068
R19639 DVDD.n18280 DVDD.n18279 0.00068
R19640 DVDD.n18278 DVDD.n10124 0.00068
R19641 DVDD.n18291 DVDD.n18290 0.00068
R19642 DVDD.n18277 DVDD.n18276 0.00068
R19643 DVDD.n18275 DVDD.n18274 0.00068
R19644 DVDD.n1839 DVDD.n1838 0.00068
R19645 DVDD.n19509 DVDD.n19508 0.00068
R19646 DVDD.n19464 DVDD.n18897 0.00068
R19647 DVDD.n18879 DVDD.n18878 0.00068
R19648 DVDD.n18847 DVDD.n18846 0.00068
R19649 DVDD.n7568 DVDD.n7567 0.00068
R19650 DVDD.n7581 DVDD.n7580 0.00068
R19651 DVDD.n19617 DVDD.n19616 0.00068
R19652 DVDD.n20124 DVDD.n20123 0.00068
R19653 DVDD.n19464 DVDD.n19146 0.00068
R19654 DVDD.n19128 DVDD.n19127 0.00068
R19655 DVDD.n19095 DVDD.n19094 0.00068
R19656 DVDD.n7524 DVDD.n7523 0.00068
R19657 DVDD.n7537 DVDD.n7536 0.00068
R19658 DVDD.n15 DVDD.n13 0.00068
R19659 DVDD.n7397 DVDD.n7395 0.00068
R19660 DVDD.n97 DVDD.n95 0.00068
R19661 DVDD.n7445 DVDD.n7443 0.00068
R19662 DVDD.n43 DVDD.n41 0.00068
R19663 DVDD.n7506 DVDD.n7504 0.00068
R19664 DVDD.n858 DVDD.n857 0.00068
R19665 DVDD.n1784 DVDD.n1783 0.00068
R19666 DVDD.n170 DVDD.n169 0.00068
R19667 DVDD.n19464 DVDD.n19164 0.00068
R19668 DVDD.n19408 DVDD.n19407 0.00068
R19669 DVDD.n19372 DVDD.n19371 0.00068
R19670 DVDD.n18260 DVDD.n18259 0.00068
R19671 DVDD.n7182 DVDD.n7181 0.00068
R19672 DVDD.n11862 DVDD.n11861 0.00068
R19673 DVDD.n11876 DVDD.n11875 0.00068
R19674 DVDD.n11893 DVDD.n11892 0.00068
R19675 DVDD.n11987 DVDD.n11986 0.00068
R19676 DVDD.n1287 DVDD.n1286 0.00068
R19677 DVDD.n11313 DVDD.n11312 0.00068
R19678 DVDD.n12291 DVDD.n12290 0.00068
R19679 DVDD.n10340 DVDD.n10339 0.00068
R19680 DVDD.n10343 DVDD.n10342 0.00068
R19681 DVDD.n13162 DVDD.n13161 0.00068
R19682 DVDD.n13187 DVDD.n13186 0.00068
R19683 DVDD.n13204 DVDD.n13203 0.00068
R19684 DVDD.n13218 DVDD.n13217 0.00068
R19685 DVDD.n13302 DVDD.n13301 0.00068
R19686 DVDD.n16840 DVDD.n16839 0.00068
R19687 DVDD.n16843 DVDD.n16842 0.00068
R19688 DVDD.n3316 DVDD.n3315 0.00068
R19689 DVDD.n3622 DVDD.n3621 0.00068
R19690 DVDD.n3650 DVDD.n3649 0.00068
R19691 DVDD.n18698 DVDD.n18697 0.00068
R19692 DVDD.n19464 DVDD.n18468 0.00068
R19693 DVDD.n18415 DVDD.n18414 0.00068
R19694 DVDD.n18368 DVDD.n18367 0.00068
R19695 DVDD.n14785 DVDD.n14784 0.00068
R19696 DVDD.n7174 DVDD.n7173 0.00068
R19697 DVDD.n20233 DVDD.n20231 0.00068
R19698 DVDD.n7313 DVDD.n7311 0.00068
R19699 DVDD.n1217 DVDD.n1216 0.000677165
R19700 DVDD.n1171 DVDD.n1170 0.000677165
R19701 DVDD.n1629 DVDD.n1628 0.000677165
R19702 DVDD.n1640 DVDD.n1639 0.000677165
R19703 DVDD.n884 DVDD.n883 0.000677165
R19704 DVDD.n878 DVDD.n877 0.000677165
R19705 DVDD.n875 DVDD.n874 0.000677165
R19706 DVDD.n19333 DVDD.n19332 0.000677165
R19707 DVDD.n19323 DVDD.n19322 0.000677165
R19708 DVDD.n19319 DVDD.n19318 0.000677165
R19709 DVDD.n11437 DVDD.n11436 0.000677165
R19710 DVDD.n11443 DVDD.n11442 0.000677165
R19711 DVDD.n11446 DVDD.n11445 0.000677165
R19712 DVDD.n12018 DVDD.n12017 0.000677165
R19713 DVDD.n12153 DVDD.n12152 0.000677165
R19714 DVDD.n12201 DVDD.n12200 0.000677165
R19715 DVDD.n12200 DVDD.n11298 0.000677165
R19716 DVDD.n13304 DVDD.n13303 0.000677165
R19717 DVDD.n13373 DVDD.n13372 0.000677165
R19718 DVDD.n13382 DVDD.n13381 0.000677165
R19719 DVDD.n13391 DVDD.n13390 0.000677165
R19720 DVDD.n13400 DVDD.n13399 0.000677165
R19721 DVDD.n13406 DVDD.n13405 0.000677165
R19722 DVDD.n13412 DVDD.n13411 0.000677165
R19723 DVDD.n13421 DVDD.n13420 0.000677165
R19724 DVDD.n13430 DVDD.n13429 0.000677165
R19725 DVDD.n13439 DVDD.n13438 0.000677165
R19726 DVDD.n13448 DVDD.n13447 0.000677165
R19727 DVDD.n13457 DVDD.n13456 0.000677165
R19728 DVDD.n13466 DVDD.n13465 0.000677165
R19729 DVDD.n13472 DVDD.n13471 0.000677165
R19730 DVDD.n13478 DVDD.n13477 0.000677165
R19731 DVDD.n13487 DVDD.n13486 0.000677165
R19732 DVDD.n13500 DVDD.n13499 0.000677165
R19733 DVDD.n13554 DVDD.n13553 0.000677165
R19734 DVDD.n13610 DVDD.n13609 0.000677165
R19735 DVDD.n13635 DVDD.n13634 0.000677165
R19736 DVDD.n13691 DVDD.n13690 0.000677165
R19737 DVDD.n2747 DVDD.n2746 0.000677165
R19738 DVDD.n2788 DVDD.n2787 0.000677165
R19739 DVDD.n18572 DVDD.n18571 0.000677165
R19740 DVDD.n14808 DVDD.n14807 0.000677165
R19741 DVDD.n15399 DVDD.n15398 0.000677165
R19742 DVDD.n15462 DVDD.n15461 0.000677165
R19743 DVDD.n14704 DVDD.n14703 0.000677165
R19744 DVDD.n14621 DVDD.n14620 0.000677165
R19745 DVDD.n14567 DVDD.n14566 0.000677165
R19746 DVDD.n14504 DVDD.n14503 0.000677165
R19747 DVDD.n14479 DVDD.n14478 0.000677165
R19748 DVDD.n14400 DVDD.n14399 0.000677165
R19749 DVDD.n19695 DVDD.n19694 0.000677165
R19750 DVDD.n19737 DVDD.n19736 0.000677165
R19751 DVDD.n19743 DVDD.n19742 0.000677165
R19752 DVDD.n19750 DVDD.n19749 0.000677165
R19753 DVDD.n19892 DVDD.n19891 0.000677165
R19754 DVDD.n19910 DVDD.n19909 0.000677165
R19755 DVDD.n19917 DVDD.n19916 0.000677165
R19756 DVDD.n20050 DVDD.n20008 0.000677165
R19757 DVDD.n20206 DVDD.n20205 0.000677165
R19758 DVDD.n20203 DVDD.n20202 0.000677165
R19759 DVDD.n20197 DVDD.n20196 0.000677165
R19760 DVDD.n20189 DVDD.n20188 0.000677165
R19761 DVDD.n20085 DVDD.n20084 0.000677165
R19762 DVDD.n20088 DVDD.n20087 0.000677165
R19763 DVDD.n20102 DVDD.n20101 0.000677165
R19764 DVDD.n19057 DVDD.n19056 0.000677165
R19765 DVDD.n19055 DVDD.n19054 0.000677165
R19766 DVDD.n19015 DVDD.n19014 0.000677165
R19767 DVDD.n4659 DVDD.n4658 0.000677165
R19768 DVDD.n4664 DVDD.n4663 0.000677165
R19769 DVDD.n4673 DVDD.n4672 0.000677165
R19770 DVDD.n4806 DVDD.n4805 0.000677165
R19771 DVDD.n4809 DVDD.n4808 0.000677165
R19772 DVDD.n4814 DVDD.n4813 0.000677165
R19773 DVDD.n4900 DVDD.n4899 0.000677165
R19774 DVDD.n4998 DVDD.n4997 0.000677165
R19775 DVDD.n5009 DVDD.n5008 0.000677165
R19776 DVDD.n5020 DVDD.n5019 0.000677165
R19777 DVDD.n5032 DVDD.n5031 0.000677165
R19778 DVDD.n5187 DVDD.n5186 0.000677165
R19779 DVDD.n5190 DVDD.n5189 0.000677165
R19780 DVDD.n5221 DVDD.n5220 0.000677165
R19781 DVDD.n5307 DVDD.n5227 0.000677165
R19782 DVDD.n5310 DVDD.n5309 0.000677165
R19783 DVDD.n5397 DVDD.n5396 0.000677165
R19784 DVDD.n5401 DVDD.n5400 0.000677165
R19785 DVDD.n5463 DVDD.n5462 0.000677165
R19786 DVDD.n5468 DVDD.n5467 0.000677165
R19787 DVDD.n5591 DVDD.n5590 0.000677165
R19788 DVDD.n5610 DVDD.n5609 0.000677165
R19789 DVDD.n5694 DVDD.n5693 0.000677165
R19790 DVDD.n6102 DVDD.n6101 0.000677165
R19791 DVDD.n6075 DVDD.n6074 0.000677165
R19792 DVDD.n5960 DVDD.n5959 0.000677165
R19793 DVDD.n1340 DVDD.n1339 0.000677165
R19794 DVDD.n1378 DVDD.n1377 0.000677165
R19795 DVDD.n1382 DVDD.n1381 0.000677165
R19796 DVDD.n1388 DVDD.n1387 0.000677165
R19797 DVDD.n1395 DVDD.n1394 0.000677165
R19798 DVDD.n1485 DVDD.n1484 0.000677165
R19799 DVDD.n1467 DVDD.n1466 0.000677165
R19800 DVDD.n1460 DVDD.n1459 0.000677165
R19801 DVDD.n1722 DVDD.n1696 0.000677165
R19802 DVDD.n284 DVDD.n283 0.000677165
R19803 DVDD.n281 DVDD.n280 0.000677165
R19804 DVDD.n275 DVDD.n274 0.000677165
R19805 DVDD.n267 DVDD.n266 0.000677165
R19806 DVDD.n19183 DVDD.n19182 0.000677165
R19807 DVDD.n19186 DVDD.n19185 0.000677165
R19808 DVDD.n19200 DVDD.n19199 0.000677165
R19809 DVDD.n19439 DVDD.n19438 0.000677165
R19810 DVDD.n19437 DVDD.n19436 0.000677165
R19811 DVDD.n19224 DVDD.n19223 0.000677165
R19812 DVDD.n11366 DVDD.n11365 0.000677165
R19813 DVDD.n11371 DVDD.n11370 0.000677165
R19814 DVDD.n11380 DVDD.n11379 0.000677165
R19815 DVDD.n11632 DVDD.n11631 0.000677165
R19816 DVDD.n11635 DVDD.n11634 0.000677165
R19817 DVDD.n11640 DVDD.n11639 0.000677165
R19818 DVDD.n11853 DVDD.n11852 0.000677165
R19819 DVDD.n11780 DVDD.n11779 0.000677165
R19820 DVDD.n11755 DVDD.n11754 0.000677165
R19821 DVDD.n11745 DVDD.n11744 0.000677165
R19822 DVDD.n11734 DVDD.n11733 0.000677165
R19823 DVDD.n11722 DVDD.n11721 0.000677165
R19824 DVDD.n12367 DVDD.n12366 0.000677165
R19825 DVDD.n12370 DVDD.n12369 0.000677165
R19826 DVDD.n12401 DVDD.n12400 0.000677165
R19827 DVDD.n13150 DVDD.n12407 0.000677165
R19828 DVDD.n13148 DVDD.n13147 0.000677165
R19829 DVDD.n13142 DVDD.n13141 0.000677165
R19830 DVDD.n13064 DVDD.n13063 0.000677165
R19831 DVDD.n13011 DVDD.n13010 0.000677165
R19832 DVDD.n13004 DVDD.n13003 0.000677165
R19833 DVDD.n13000 DVDD.n12999 0.000677165
R19834 DVDD.n12995 DVDD.n12994 0.000677165
R19835 DVDD.n12836 DVDD.n12835 0.000677165
R19836 DVDD.n12817 DVDD.n12816 0.000677165
R19837 DVDD.n12747 DVDD.n12746 0.000677165
R19838 DVDD.n12734 DVDD.n12733 0.000677165
R19839 DVDD.n12707 DVDD.n12706 0.000677165
R19840 DVDD.n12623 DVDD.n12622 0.000677165
R19841 DVDD.n785 DVDD.n784 0.000677165
R19842 DVDD.n822 DVDD.n821 0.000677165
R19843 DVDD.n241 DVDD.n240 0.000677165
R19844 DVDD.n18230 DVDD.n18229 0.000677165
R19845 DVDD.n18201 DVDD.n18200 0.000677165
R19846 DVDD.n18145 DVDD.n18144 0.000677165
R19847 DVDD.n18057 DVDD.n18056 0.000677165
R19848 DVDD.n17979 DVDD.n17978 0.000677165
R19849 DVDD.n17927 DVDD.n17926 0.000677165
R19850 DVDD.n17871 DVDD.n17870 0.000677165
R19851 DVDD.n17846 DVDD.n17845 0.000677165
R19852 DVDD.n17776 DVDD.n17775 0.000677165
R19853 DVDD.n1917 DVDD.n1916 0.000677165
R19854 DVDD.n1955 DVDD.n1954 0.000677165
R19855 DVDD.n1959 DVDD.n1958 0.000677165
R19856 DVDD.n1965 DVDD.n1964 0.000677165
R19857 DVDD.n1972 DVDD.n1971 0.000677165
R19858 DVDD.n2113 DVDD.n2112 0.000677165
R19859 DVDD.n2131 DVDD.n2130 0.000677165
R19860 DVDD.n2138 DVDD.n2137 0.000677165
R19861 DVDD.n2271 DVDD.n2229 0.000677165
R19862 DVDD.n19591 DVDD.n19590 0.000677165
R19863 DVDD.n19588 DVDD.n19587 0.000677165
R19864 DVDD.n19582 DVDD.n19581 0.000677165
R19865 DVDD.n19574 DVDD.n19573 0.000677165
R19866 DVDD.n19470 DVDD.n19469 0.000677165
R19867 DVDD.n19473 DVDD.n19472 0.000677165
R19868 DVDD.n19487 DVDD.n19486 0.000677165
R19869 DVDD.n18949 DVDD.n18948 0.000677165
R19870 DVDD.n18947 DVDD.n18946 0.000677165
R19871 DVDD.n18942 DVDD.n18941 0.000677165
R19872 DVDD.n7025 DVDD.n7024 0.000677165
R19873 DVDD.n7020 DVDD.n7019 0.000677165
R19874 DVDD.n7011 DVDD.n7010 0.000677165
R19875 DVDD.n6878 DVDD.n6877 0.000677165
R19876 DVDD.n6875 DVDD.n6874 0.000677165
R19877 DVDD.n6870 DVDD.n6869 0.000677165
R19878 DVDD.n6862 DVDD.n6783 0.000677165
R19879 DVDD.n6711 DVDD.n6710 0.000677165
R19880 DVDD.n6686 DVDD.n6685 0.000677165
R19881 DVDD.n6675 DVDD.n6674 0.000677165
R19882 DVDD.n6664 DVDD.n6663 0.000677165
R19883 DVDD.n6652 DVDD.n6651 0.000677165
R19884 DVDD.n6495 DVDD.n6494 0.000677165
R19885 DVDD.n6492 DVDD.n6491 0.000677165
R19886 DVDD.n6461 DVDD.n6460 0.000677165
R19887 DVDD.n6454 DVDD.n6453 0.000677165
R19888 DVDD.n6451 DVDD.n6450 0.000677165
R19889 DVDD.n6445 DVDD.n6444 0.000677165
R19890 DVDD.n6364 DVDD.n6363 0.000677165
R19891 DVDD.n6309 DVDD.n6308 0.000677165
R19892 DVDD.n6302 DVDD.n6301 0.000677165
R19893 DVDD.n6298 DVDD.n6297 0.000677165
R19894 DVDD.n6293 DVDD.n6292 0.000677165
R19895 DVDD.n6216 DVDD.n6215 0.000677165
R19896 DVDD.n6129 DVDD.n6128 0.000677165
R19897 DVDD.n4551 DVDD.n4550 0.000677165
R19898 DVDD.n4525 DVDD.n4524 0.000677165
R19899 DVDD.n4421 DVDD.n4420 0.000677165
R19900 DVDD.n3263 DVDD.n3262 0.000677165
R19901 DVDD.n3225 DVDD.n3224 0.000677165
R19902 DVDD.n3221 DVDD.n3220 0.000677165
R19903 DVDD.n3215 DVDD.n3214 0.000677165
R19904 DVDD.n3208 DVDD.n3207 0.000677165
R19905 DVDD.n3512 DVDD.n3511 0.000677165
R19906 DVDD.n3530 DVDD.n3529 0.000677165
R19907 DVDD.n3537 DVDD.n3536 0.000677165
R19908 DVDD.n3715 DVDD.n2833 0.000677165
R19909 DVDD.n3770 DVDD.n3769 0.000677165
R19910 DVDD.n3767 DVDD.n3766 0.000677165
R19911 DVDD.n3761 DVDD.n3760 0.000677165
R19912 DVDD.n3753 DVDD.n3752 0.000677165
R19913 DVDD.n18487 DVDD.n18486 0.000677165
R19914 DVDD.n18490 DVDD.n18489 0.000677165
R19915 DVDD.n18504 DVDD.n18503 0.000677165
R19916 DVDD.n18786 DVDD.n18785 0.000677165
R19917 DVDD.n18784 DVDD.n18783 0.000677165
R19918 DVDD.n18528 DVDD.n18527 0.000677165
R19919 DVDD.n10042 DVDD.n10041 0.000677165
R19920 DVDD.n10037 DVDD.n10036 0.000677165
R19921 DVDD.n10028 DVDD.n10027 0.000677165
R19922 DVDD.n7888 DVDD.n7887 0.000677165
R19923 DVDD.n7891 DVDD.n7890 0.000677165
R19924 DVDD.n7896 DVDD.n7895 0.000677165
R19925 DVDD.n9752 DVDD.n9751 0.000677165
R19926 DVDD.n9679 DVDD.n9678 0.000677165
R19927 DVDD.n9654 DVDD.n9653 0.000677165
R19928 DVDD.n9643 DVDD.n9642 0.000677165
R19929 DVDD.n9632 DVDD.n9631 0.000677165
R19930 DVDD.n9620 DVDD.n9619 0.000677165
R19931 DVDD.n8388 DVDD.n8387 0.000677165
R19932 DVDD.n8391 DVDD.n8390 0.000677165
R19933 DVDD.n8422 DVDD.n8421 0.000677165
R19934 DVDD.n9239 DVDD.n8428 0.000677165
R19935 DVDD.n9237 DVDD.n9236 0.000677165
R19936 DVDD.n9231 DVDD.n9230 0.000677165
R19937 DVDD.n9150 DVDD.n9149 0.000677165
R19938 DVDD.n9095 DVDD.n9094 0.000677165
R19939 DVDD.n9088 DVDD.n9087 0.000677165
R19940 DVDD.n9084 DVDD.n9083 0.000677165
R19941 DVDD.n9079 DVDD.n9078 0.000677165
R19942 DVDD.n8918 DVDD.n8917 0.000677165
R19943 DVDD.n8831 DVDD.n8830 0.000677165
R19944 DVDD.n8818 DVDD.n8817 0.000677165
R19945 DVDD.n8792 DVDD.n8791 0.000677165
R19946 DVDD.n8695 DVDD.n8694 0.000677165
R19947 DVDD.n10403 DVDD.n10402 0.00066875
R19948 DVDD.n10565 DVDD.n10564 0.00066875
R19949 DVDD.n10588 DVDD.n10587 0.00066875
R19950 DVDD.n10636 DVDD.n10635 0.00066875
R19951 DVDD.n19534 DVDD.n19533 0.00065
R19952 DVDD.n18887 DVDD.n18886 0.00065
R19953 DVDD.n18884 DVDD.n18883 0.00065
R19954 DVDD.n18881 DVDD.n18880 0.00065
R19955 DVDD.n3918 DVDD.n3917 0.00065
R19956 DVDD.n3915 DVDD.n3914 0.00065
R19957 DVDD.n20149 DVDD.n20148 0.00065
R19958 DVDD.n19136 DVDD.n19135 0.00065
R19959 DVDD.n19133 DVDD.n19132 0.00065
R19960 DVDD.n19130 DVDD.n19129 0.00065
R19961 DVDD.n4605 DVDD.n4604 0.00065
R19962 DVDD.n7519 DVDD.n7518 0.00065
R19963 DVDD.n853 DVDD.n852 0.00065
R19964 DVDD.n1788 DVDD.n1787 0.00065
R19965 DVDD.n1792 DVDD.n1791 0.00065
R19966 DVDD.n201 DVDD.n200 0.00065
R19967 DVDD.n19353 DVDD.n19352 0.00065
R19968 DVDD.n19414 DVDD.n19413 0.00065
R19969 DVDD.n18244 DVDD.n18243 0.00065
R19970 DVDD.n18265 DVDD.n18246 0.00065
R19971 DVDD.n18254 DVDD.n18253 0.00065
R19972 DVDD.n18249 DVDD.n18248 0.00065
R19973 DVDD.n10521 DVDD.n10520 0.00065
R19974 DVDD.n10518 DVDD.n10517 0.00065
R19975 DVDD.n17128 DVDD.n17127 0.00065
R19976 DVDD.n17125 DVDD.n17124 0.00065
R19977 DVDD.n16167 DVDD.n16166 0.00065
R19978 DVDD.n16170 DVDD.n16169 0.00065
R19979 DVDD.n16285 DVDD.n16284 0.00065
R19980 DVDD.n16289 DVDD.n16288 0.00065
R19981 DVDD.n16226 DVDD.n16225 0.00065
R19982 DVDD.n16229 DVDD.n16228 0.00065
R19983 DVDD.n15591 DVDD.n15590 0.00065
R19984 DVDD.n15594 DVDD.n15593 0.00065
R19985 DVDD.n15806 DVDD.n15805 0.00065
R19986 DVDD.n15810 DVDD.n15809 0.00065
R19987 DVDD.n15869 DVDD.n15868 0.00065
R19988 DVDD.n15873 DVDD.n15872 0.00065
R19989 DVDD.n3617 DVDD.n3616 0.00065
R19990 DVDD.n3646 DVDD.n3645 0.00065
R19991 DVDD.n3642 DVDD.n3641 0.00065
R19992 DVDD.n18652 DVDD.n18651 0.00065
R19993 DVDD.n18452 DVDD.n18451 0.00065
R19994 DVDD.n18449 DVDD.n18420 0.00065
R19995 DVDD.n14794 DVDD.n14793 0.00065
R19996 DVDD.n14791 DVDD.n14790 0.00065
R19997 DVDD.n14779 DVDD.n14778 0.00065
R19998 DVDD.n14774 DVDD.n14773 0.00065
R19999 DVDD.n4133 DVDD.n4132 0.000628571
R20000 DVDD.n8515 DVDD.n8514 0.000628571
R20001 DVDD.n11217 DVDD.n11216 0.000628571
R20002 DVDD.n13848 DVDD.n13847 0.000628571
R20003 DVDD.n2328 DVDD.n2327 0.000628571
R20004 DVDD.n2337 DVDD.n2336 0.000628571
R20005 DVDD.n2379 DVDD.n2378 0.000628571
R20006 DVDD.n2388 DVDD.n2387 0.000628571
R20007 DVDD.n2426 DVDD.n2425 0.000628571
R20008 DVDD.n2501 DVDD.n2500 0.000628571
R20009 DVDD.n2672 DVDD.n2671 0.000628571
R20010 DVDD.n2526 DVDD.n2525 0.000628571
R20011 DVDD.n2535 DVDD.n2534 0.000628571
R20012 DVDD.n2577 DVDD.n2576 0.000628571
R20013 DVDD.n2586 DVDD.n2585 0.000628571
R20014 DVDD.n2622 DVDD.n2621 0.000628571
R20015 DVDD.n2713 DVDD.n2712 0.000628571
R20016 DVDD.n2674 DVDD.n2673 0.000628571
R20017 DVDD.n2686 DVDD.n2685 0.000628571
R20018 DVDD.n4135 DVDD.n4134 0.000628571
R20019 DVDD.n4159 DVDD.n4158 0.000628571
R20020 DVDD.n8517 DVDD.n8516 0.000628571
R20021 DVDD.n8541 DVDD.n8540 0.000628571
R20022 DVDD.n11219 DVDD.n11218 0.000628571
R20023 DVDD.n13873 DVDD.n13872 0.000628571
R20024 DVDD.n13849 DVDD.n13845 0.000628571
R20025 DVDD.n13838 DVDD.n13837 0.000628571
R20026 DVDD.n1828 DVDD.n1827 0.00062
R20027 DVDD.n1843 DVDD.n1842 0.00062
R20028 DVDD.n1846 DVDD.n1845 0.00062
R20029 DVDD.n1852 DVDD.n1851 0.00062
R20030 DVDD.n1855 DVDD.n1854 0.00062
R20031 DVDD.n20215 DVDD.n1856 0.00062
R20032 DVDD.n19515 DVDD.n19514 0.00062
R20033 DVDD.n18892 DVDD.n18891 0.00062
R20034 DVDD.n18835 DVDD.n18834 0.00062
R20035 DVDD.n3916 DVDD.n3915 0.00062
R20036 DVDD.n7567 DVDD.n7566 0.00062
R20037 DVDD.n7570 DVDD.n7569 0.00062
R20038 DVDD.n19606 DVDD.n19605 0.00062
R20039 DVDD.n19621 DVDD.n19620 0.00062
R20040 DVDD.n19624 DVDD.n19623 0.00062
R20041 DVDD.n19630 DVDD.n19629 0.00062
R20042 DVDD.n19633 DVDD.n19632 0.00062
R20043 DVDD.n20215 DVDD.n19634 0.00062
R20044 DVDD.n20130 DVDD.n20129 0.00062
R20045 DVDD.n19141 DVDD.n19140 0.00062
R20046 DVDD.n19083 DVDD.n19082 0.00062
R20047 DVDD.n7518 DVDD.n7517 0.00062
R20048 DVDD.n7523 DVDD.n7522 0.00062
R20049 DVDD.n7526 DVDD.n7525 0.00062
R20050 DVDD.n23 DVDD.n22 0.00062
R20051 DVDD.n7389 DVDD.n7388 0.00062
R20052 DVDD.n105 DVDD.n104 0.00062
R20053 DVDD.n7437 DVDD.n7436 0.00062
R20054 DVDD.n51 DVDD.n50 0.00062
R20055 DVDD.n7624 DVDD.n7623 0.00062
R20056 DVDD.n852 DVDD.n851 0.00062
R20057 DVDD.n1789 DVDD.n1788 0.00062
R20058 DVDD.n1793 DVDD.n1792 0.00062
R20059 DVDD.n1800 DVDD.n1799 0.00062
R20060 DVDD.n1804 DVDD.n1803 0.00062
R20061 DVDD.n20215 DVDD.n1806 0.00062
R20062 DVDD.n178 DVDD.n177 0.00062
R20063 DVDD.n19347 DVDD.n19346 0.00062
R20064 DVDD.n19358 DVDD.n19357 0.00062
R20065 DVDD.n18246 DVDD.n18245 0.00062
R20066 DVDD.n18261 DVDD.n18260 0.00062
R20067 DVDD.n18257 DVDD.n18256 0.00062
R20068 DVDD.n10346 DVDD.n10345 0.00062
R20069 DVDD.n10380 DVDD.n10379 0.00062
R20070 DVDD.n10506 DVDD.n10505 0.00062
R20071 DVDD.n10435 DVDD.n10434 0.00062
R20072 DVDD.n10348 DVDD.n10347 0.00062
R20073 DVDD.n10382 DVDD.n10381 0.00062
R20074 DVDD.n10507 DVDD.n10503 0.00062
R20075 DVDD.n10436 DVDD.n10431 0.00062
R20076 DVDD.n16503 DVDD.n16502 0.00062
R20077 DVDD.n17164 DVDD.n17160 0.00062
R20078 DVDD.n17117 DVDD.n17114 0.00062
R20079 DVDD.n17067 DVDD.n17064 0.00062
R20080 DVDD.n16845 DVDD.n16844 0.00062
R20081 DVDD.n16870 DVDD.n16869 0.00062
R20082 DVDD.n17019 DVDD.n17018 0.00062
R20083 DVDD.n17015 DVDD.n17014 0.00062
R20084 DVDD.n17009 DVDD.n17008 0.00062
R20085 DVDD.n17006 DVDD.n17002 0.00062
R20086 DVDD.n17001 DVDD.n17000 0.00062
R20087 DVDD.n16960 DVDD.n16959 0.00062
R20088 DVDD.n16957 DVDD.n16956 0.00062
R20089 DVDD.n16951 DVDD.n16950 0.00062
R20090 DVDD.n16948 DVDD.n16944 0.00062
R20091 DVDD.n16943 DVDD.n16942 0.00062
R20092 DVDD.n16153 DVDD.n16152 0.00062
R20093 DVDD.n16161 DVDD.n16160 0.00062
R20094 DVDD.n16271 DVDD.n16270 0.00062
R20095 DVDD.n16279 DVDD.n16278 0.00062
R20096 DVDD.n16716 DVDD.n16715 0.00062
R20097 DVDD.n16740 DVDD.n16739 0.00062
R20098 DVDD.n16796 DVDD.n16795 0.00062
R20099 DVDD.n16793 DVDD.n16792 0.00062
R20100 DVDD.n16784 DVDD.n16783 0.00062
R20101 DVDD.n16781 DVDD.n16777 0.00062
R20102 DVDD.n16776 DVDD.n16775 0.00062
R20103 DVDD.n16919 DVDD.n16918 0.00062
R20104 DVDD.n16916 DVDD.n16915 0.00062
R20105 DVDD.n16907 DVDD.n16906 0.00062
R20106 DVDD.n16904 DVDD.n16900 0.00062
R20107 DVDD.n16899 DVDD.n16898 0.00062
R20108 DVDD.n16209 DVDD.n16208 0.00062
R20109 DVDD.n16217 DVDD.n16216 0.00062
R20110 DVDD.n15574 DVDD.n15573 0.00062
R20111 DVDD.n15582 DVDD.n15581 0.00062
R20112 DVDD.n16547 DVDD.n16546 0.00062
R20113 DVDD.n16572 DVDD.n16571 0.00062
R20114 DVDD.n16674 DVDD.n16673 0.00062
R20115 DVDD.n16671 DVDD.n16670 0.00062
R20116 DVDD.n16661 DVDD.n16660 0.00062
R20117 DVDD.n16658 DVDD.n16654 0.00062
R20118 DVDD.n16653 DVDD.n16652 0.00062
R20119 DVDD.n16617 DVDD.n16616 0.00062
R20120 DVDD.n16614 DVDD.n16613 0.00062
R20121 DVDD.n16604 DVDD.n16603 0.00062
R20122 DVDD.n16601 DVDD.n16597 0.00062
R20123 DVDD.n16596 DVDD.n16595 0.00062
R20124 DVDD.n15788 DVDD.n15787 0.00062
R20125 DVDD.n15796 DVDD.n15795 0.00062
R20126 DVDD.n15851 DVDD.n15850 0.00062
R20127 DVDD.n15859 DVDD.n15858 0.00062
R20128 DVDD.n16532 DVDD.n16531 0.00062
R20129 DVDD.n16657 DVDD.n16656 0.00062
R20130 DVDD.n16600 DVDD.n16599 0.00062
R20131 DVDD.n16701 DVDD.n16700 0.00062
R20132 DVDD.n16780 DVDD.n16779 0.00062
R20133 DVDD.n16903 DVDD.n16902 0.00062
R20134 DVDD.n16827 DVDD.n16826 0.00062
R20135 DVDD.n16877 DVDD.n16876 0.00062
R20136 DVDD.n17005 DVDD.n17004 0.00062
R20137 DVDD.n16947 DVDD.n16946 0.00062
R20138 DVDD.n16483 DVDD.n16482 0.00062
R20139 DVDD.n17163 DVDD.n17162 0.00062
R20140 DVDD.n17116 DVDD.n17115 0.00062
R20141 DVDD.n17066 DVDD.n17065 0.00062
R20142 DVDD.n3616 DVDD.n3615 0.00062
R20143 DVDD.n3645 DVDD.n3644 0.00062
R20144 DVDD.n3641 DVDD.n3640 0.00062
R20145 DVDD.n3634 DVDD.n3633 0.00062
R20146 DVDD.n3630 DVDD.n3629 0.00062
R20147 DVDD.n20215 DVDD.n2812 0.00062
R20148 DVDD.n18713 DVDD.n18712 0.00062
R20149 DVDD.n18458 DVDD.n18457 0.00062
R20150 DVDD.n18337 DVDD.n18336 0.00062
R20151 DVDD.n14792 DVDD.n14791 0.00062
R20152 DVDD.n14786 DVDD.n14785 0.00062
R20153 DVDD.n14782 DVDD.n14781 0.00062
R20154 DVDD.n20241 DVDD.n20240 0.00062
R20155 DVDD.n7305 DVDD.n7304 0.00062
R20156 DVDD.n14918 DVDD.n14917 0.0006125
R20157 DVDD.n14924 DVDD.n14923 0.0006125
R20158 DVDD.n14887 DVDD.n14886 0.0006125
R20159 DVDD.n15216 DVDD.n15215 0.0006125
R20160 DVDD.n15222 DVDD.n15221 0.0006125
R20161 DVDD.n15239 DVDD.n15238 0.0006125
R20162 DVDD.n15248 DVDD.n15247 0.0006125
R20163 DVDD.n15309 DVDD.n15308 0.0006125
R20164 DVDD.n15295 DVDD.n15294 0.0006125
R20165 DVDD.n15000 DVDD.n14999 0.0006125
R20166 DVDD.n18976 DVDD.n18975 0.000604287
R20167 DVDD.n10543 DVDD.n10542 0.000604287
R20168 DVDD.n15199 DVDD.n15198 0.000596051
R20169 DVDD.n15122 DVDD.n15121 0.000596051
R20170 DVDD.n7701 DVDD.n7700 0.00059
R20171 DVDD.n3693 DVDD.n3692 0.00059
R20172 DVDD.n18539 DVDD.n18538 0.00059
R20173 DVDD.n18775 DVDD.n18774 0.00059
R20174 DVDD.n2947 DVDD.n2946 0.00059
R20175 DVDD.n2955 DVDD.n2954 0.00059
R20176 DVDD.n9805 DVDD.n9804 0.00059
R20177 DVDD.n9362 DVDD.n9361 0.00059
R20178 DVDD.n9359 DVDD.n9358 0.00059
R20179 DVDD.n9356 DVDD.n9355 0.00059
R20180 DVDD.n9353 DVDD.n9352 0.00059
R20181 DVDD.n9350 DVDD.n9349 0.00059
R20182 DVDD.n9347 DVDD.n9346 0.00059
R20183 DVDD.n9344 DVDD.n9343 0.00059
R20184 DVDD.n9341 DVDD.n9340 0.00059
R20185 DVDD.n9338 DVDD.n9337 0.00059
R20186 DVDD.n9335 DVDD.n9334 0.00059
R20187 DVDD.n9332 DVDD.n9331 0.00059
R20188 DVDD.n9329 DVDD.n9328 0.00059
R20189 DVDD.n9326 DVDD.n9325 0.00059
R20190 DVDD.n9323 DVDD.n9322 0.00059
R20191 DVDD.n9320 DVDD.n9319 0.00059
R20192 DVDD.n9315 DVDD.n9314 0.00059
R20193 DVDD.n2185 DVDD.n2184 0.00059
R20194 DVDD.n2193 DVDD.n2192 0.00059
R20195 DVDD.n2249 DVDD.n2248 0.00059
R20196 DVDD.n18908 DVDD.n18907 0.00059
R20197 DVDD.n7068 DVDD.n7067 0.00059
R20198 DVDD.n6810 DVDD.n6809 0.00059
R20199 DVDD.n1901 DVDD.n1900 0.00059
R20200 DVDD.n19964 DVDD.n19963 0.00059
R20201 DVDD.n19972 DVDD.n19971 0.00059
R20202 DVDD.n20028 DVDD.n20027 0.00059
R20203 DVDD.n19026 DVDD.n19025 0.00059
R20204 DVDD.n4648 DVDD.n4647 0.00059
R20205 DVDD.n4847 DVDD.n4846 0.00059
R20206 DVDD.n19679 DVDD.n19678 0.00059
R20207 DVDD.n981 DVDD.n980 0.00059
R20208 DVDD.n973 DVDD.n972 0.00059
R20209 DVDD.n936 DVDD.n935 0.00059
R20210 DVDD.n19235 DVDD.n19234 0.00059
R20211 DVDD.n19428 DVDD.n19427 0.00059
R20212 DVDD.n18324 DVDD.n18323 0.00059
R20213 DVDD.n1830 DVDD.n1829 0.00059
R20214 DVDD.n1851 DVDD.n1850 0.00059
R20215 DVDD.n18896 DVDD.n18895 0.00059
R20216 DVDD.n18869 DVDD.n18868 0.00059
R20217 DVDD.n18863 DVDD.n18862 0.00059
R20218 DVDD.n18853 DVDD.n18852 0.00059
R20219 DVDD.n18839 DVDD.n18838 0.00059
R20220 DVDD.n18837 DVDD.n18836 0.00059
R20221 DVDD.n19608 DVDD.n19607 0.00059
R20222 DVDD.n19629 DVDD.n19628 0.00059
R20223 DVDD.n19145 DVDD.n19144 0.00059
R20224 DVDD.n19118 DVDD.n19117 0.00059
R20225 DVDD.n19112 DVDD.n19111 0.00059
R20226 DVDD.n19101 DVDD.n19100 0.00059
R20227 DVDD.n19087 DVDD.n19086 0.00059
R20228 DVDD.n19085 DVDD.n19084 0.00059
R20229 DVDD.n11 DVDD.n10 0.00059
R20230 DVDD.n7425 DVDD.n7423 0.00059
R20231 DVDD.n7401 DVDD.n7400 0.00059
R20232 DVDD.n93 DVDD.n92 0.00059
R20233 DVDD.n7473 DVDD.n7471 0.00059
R20234 DVDD.n7449 DVDD.n7448 0.00059
R20235 DVDD.n39 DVDD.n38 0.00059
R20236 DVDD.n7478 DVDD.n7476 0.00059
R20237 DVDD.n7502 DVDD.n7501 0.00059
R20238 DVDD.n845 DVDD.n844 0.00059
R20239 DVDD.n849 DVDD.n848 0.00059
R20240 DVDD.n855 DVDD.n854 0.00059
R20241 DVDD.n1797 DVDD.n1796 0.00059
R20242 DVDD.n1799 DVDD.n1798 0.00059
R20243 DVDD.n1801 DVDD.n1800 0.00059
R20244 DVDD.n19342 DVDD.n19341 0.00059
R20245 DVDD.n19411 DVDD.n19410 0.00059
R20246 DVDD.n19406 DVDD.n19405 0.00059
R20247 DVDD.n19395 DVDD.n19394 0.00059
R20248 DVDD.n19387 DVDD.n19386 0.00059
R20249 DVDD.n19378 DVDD.n19377 0.00059
R20250 DVDD.n19363 DVDD.n19362 0.00059
R20251 DVDD.n19360 DVDD.n19359 0.00059
R20252 DVDD.n10187 DVDD.n10186 0.00059
R20253 DVDD.n18240 DVDD.n18239 0.00059
R20254 DVDD.n11906 DVDD.n11905 0.00059
R20255 DVDD.n1324 DVDD.n1323 0.00059
R20256 DVDD.n10341 DVDD.n10340 0.00059
R20257 DVDD.n10376 DVDD.n10375 0.00059
R20258 DVDD.n10511 DVDD.n10510 0.00059
R20259 DVDD.n13273 DVDD.n13272 0.00059
R20260 DVDD.n13270 DVDD.n13269 0.00059
R20261 DVDD.n13267 DVDD.n13266 0.00059
R20262 DVDD.n13264 DVDD.n13263 0.00059
R20263 DVDD.n13261 DVDD.n13260 0.00059
R20264 DVDD.n13258 DVDD.n13257 0.00059
R20265 DVDD.n13255 DVDD.n13254 0.00059
R20266 DVDD.n13252 DVDD.n13251 0.00059
R20267 DVDD.n13249 DVDD.n13248 0.00059
R20268 DVDD.n13246 DVDD.n13245 0.00059
R20269 DVDD.n13243 DVDD.n13242 0.00059
R20270 DVDD.n13240 DVDD.n13239 0.00059
R20271 DVDD.n13237 DVDD.n13236 0.00059
R20272 DVDD.n13234 DVDD.n13233 0.00059
R20273 DVDD.n13231 DVDD.n13230 0.00059
R20274 DVDD.n13226 DVDD.n13225 0.00059
R20275 DVDD.n16498 DVDD.n16497 0.00059
R20276 DVDD.n17167 DVDD.n16525 0.00059
R20277 DVDD.n17121 DVDD.n17120 0.00059
R20278 DVDD.n17071 DVDD.n17070 0.00059
R20279 DVDD.n16841 DVDD.n16840 0.00059
R20280 DVDD.n17010 DVDD.n17009 0.00059
R20281 DVDD.n16952 DVDD.n16951 0.00059
R20282 DVDD.n16713 DVDD.n16712 0.00059
R20283 DVDD.n16735 DVDD.n16734 0.00059
R20284 DVDD.n16785 DVDD.n16784 0.00059
R20285 DVDD.n16908 DVDD.n16907 0.00059
R20286 DVDD.n16544 DVDD.n16543 0.00059
R20287 DVDD.n3279 DVDD.n3278 0.00059
R20288 DVDD.n3609 DVDD.n3608 0.00059
R20289 DVDD.n3613 DVDD.n3612 0.00059
R20290 DVDD.n3619 DVDD.n3618 0.00059
R20291 DVDD.n3637 DVDD.n3636 0.00059
R20292 DVDD.n3635 DVDD.n3634 0.00059
R20293 DVDD.n3633 DVDD.n3632 0.00059
R20294 DVDD.n18463 DVDD.n18462 0.00059
R20295 DVDD.n18418 DVDD.n18417 0.00059
R20296 DVDD.n18413 DVDD.n18412 0.00059
R20297 DVDD.n18402 DVDD.n18401 0.00059
R20298 DVDD.n18383 DVDD.n18382 0.00059
R20299 DVDD.n18374 DVDD.n18373 0.00059
R20300 DVDD.n18359 DVDD.n18358 0.00059
R20301 DVDD.n18339 DVDD.n18338 0.00059
R20302 DVDD.n14745 DVDD.n14744 0.00059
R20303 DVDD.n14798 DVDD.n14797 0.00059
R20304 DVDD.n20229 DVDD.n20228 0.00059
R20305 DVDD.n7341 DVDD.n7339 0.00059
R20306 DVDD.n7317 DVDD.n7316 0.00059
R20307 DVDD.n4163 DVDD.n4161 0.000564286
R20308 DVDD.n8545 DVDD.n8543 0.000564286
R20309 DVDD.n13877 DVDD.n13875 0.000564286
R20310 DVDD.n2333 DVDD.n2332 0.000564286
R20311 DVDD.n2384 DVDD.n2383 0.000564286
R20312 DVDD.n2449 DVDD.n2430 0.000564286
R20313 DVDD.n2334 DVDD.n2330 0.000564286
R20314 DVDD.n2374 DVDD.n2373 0.000564286
R20315 DVDD.n2385 DVDD.n2381 0.000564286
R20316 DVDD.n2421 DVDD.n2420 0.000564286
R20317 DVDD.n2450 DVDD.n2428 0.000564286
R20318 DVDD.n2531 DVDD.n2530 0.000564286
R20319 DVDD.n2582 DVDD.n2581 0.000564286
R20320 DVDD.n2645 DVDD.n2626 0.000564286
R20321 DVDD.n2681 DVDD.n2679 0.000564286
R20322 DVDD.n2520 DVDD.n2519 0.000564286
R20323 DVDD.n2532 DVDD.n2528 0.000564286
R20324 DVDD.n2572 DVDD.n2571 0.000564286
R20325 DVDD.n2583 DVDD.n2579 0.000564286
R20326 DVDD.n2617 DVDD.n2616 0.000564286
R20327 DVDD.n2646 DVDD.n2624 0.000564286
R20328 DVDD.n2668 DVDD.n2667 0.000564286
R20329 DVDD.n2682 DVDD.n2678 0.000564286
R20330 DVDD.n4129 DVDD.n4128 0.000564286
R20331 DVDD.n4165 DVDD.n4164 0.000564286
R20332 DVDD.n8511 DVDD.n8510 0.000564286
R20333 DVDD.n8547 DVDD.n8546 0.000564286
R20334 DVDD.n11213 DVDD.n11212 0.000564286
R20335 DVDD.n13879 DVDD.n13878 0.000564286
R20336 DVDD.n13852 DVDD.n13851 0.000564286
R20337 DVDD.n13843 DVDD.n13842 0.000564286
R20338 DVDD.n1831 DVDD.n1830 0.00056
R20339 DVDD.n1834 DVDD.n1833 0.00056
R20340 DVDD.n19549 DVDD.n19548 0.00056
R20341 DVDD.n19543 DVDD.n19542 0.00056
R20342 DVDD.n19538 DVDD.n19537 0.00056
R20343 DVDD.n19535 DVDD.n19534 0.00056
R20344 DVDD.n19522 DVDD.n19521 0.00056
R20345 DVDD.n19510 DVDD.n19509 0.00056
R20346 DVDD.n19507 DVDD.n19506 0.00056
R20347 DVDD.n18893 DVDD.n18892 0.00056
R20348 DVDD.n18872 DVDD.n18871 0.00056
R20349 DVDD.n18871 DVDD.n18870 0.00056
R20350 DVDD.n18852 DVDD.n18851 0.00056
R20351 DVDD.n7574 DVDD.n7573 0.00056
R20352 DVDD.n7579 DVDD.n7578 0.00056
R20353 DVDD.n7582 DVDD.n7581 0.00056
R20354 DVDD.n19609 DVDD.n19608 0.00056
R20355 DVDD.n19612 DVDD.n19611 0.00056
R20356 DVDD.n20164 DVDD.n20163 0.00056
R20357 DVDD.n20158 DVDD.n20157 0.00056
R20358 DVDD.n20153 DVDD.n20152 0.00056
R20359 DVDD.n20150 DVDD.n20149 0.00056
R20360 DVDD.n20137 DVDD.n20136 0.00056
R20361 DVDD.n20125 DVDD.n20124 0.00056
R20362 DVDD.n20122 DVDD.n20121 0.00056
R20363 DVDD.n19142 DVDD.n19141 0.00056
R20364 DVDD.n19121 DVDD.n19120 0.00056
R20365 DVDD.n19120 DVDD.n19119 0.00056
R20366 DVDD.n19100 DVDD.n19099 0.00056
R20367 DVDD.n7530 DVDD.n7529 0.00056
R20368 DVDD.n7535 DVDD.n7534 0.00056
R20369 DVDD.n7538 DVDD.n7537 0.00056
R20370 DVDD.n7363 DVDD.n7362 0.00056
R20371 DVDD.n7413 DVDD.n7411 0.00056
R20372 DVDD.n7586 DVDD.n7585 0.00056
R20373 DVDD.n77 DVDD.n76 0.00056
R20374 DVDD.n7461 DVDD.n7459 0.00056
R20375 DVDD.n7542 DVDD.n7541 0.00056
R20376 DVDD.n7236 DVDD.n7235 0.00056
R20377 DVDD.n7490 DVDD.n7488 0.00056
R20378 DVDD.n7188 DVDD.n7187 0.00056
R20379 DVDD.n856 DVDD.n855 0.00056
R20380 DVDD.n860 DVDD.n859 0.00056
R20381 DVDD.n221 DVDD.n220 0.00056
R20382 DVDD.n213 DVDD.n212 0.00056
R20383 DVDD.n206 DVDD.n205 0.00056
R20384 DVDD.n202 DVDD.n201 0.00056
R20385 DVDD.n187 DVDD.n186 0.00056
R20386 DVDD.n180 DVDD.n179 0.00056
R20387 DVDD.n176 DVDD.n175 0.00056
R20388 DVDD.n171 DVDD.n170 0.00056
R20389 DVDD.n167 DVDD.n166 0.00056
R20390 DVDD.n19346 DVDD.n19345 0.00056
R20391 DVDD.n19410 DVDD.n19409 0.00056
R20392 DVDD.n19399 DVDD.n19398 0.00056
R20393 DVDD.n19398 DVDD.n19397 0.00056
R20394 DVDD.n19377 DVDD.n19376 0.00056
R20395 DVDD.n18263 DVDD.n18262 0.00056
R20396 DVDD.n18252 DVDD.n18251 0.00056
R20397 DVDD.n7179 DVDD.n7178 0.00056
R20398 DVDD.n7183 DVDD.n7182 0.00056
R20399 DVDD.n14962 DVDD.n14961 0.00056
R20400 DVDD.n15360 DVDD.n15359 0.00056
R20401 DVDD.n14957 DVDD.n14956 0.00056
R20402 DVDD.n15036 DVDD.n15035 0.00056
R20403 DVDD.n15047 DVDD.n15046 0.00056
R20404 DVDD.n15321 DVDD.n15320 0.00056
R20405 DVDD.n15387 DVDD.n15386 0.00056
R20406 DVDD.n15361 DVDD.n15357 0.00056
R20407 DVDD.n15346 DVDD.n15345 0.00056
R20408 DVDD.n11017 DVDD.n11016 0.00056
R20409 DVDD.n11028 DVDD.n11027 0.00056
R20410 DVDD.n11073 DVDD.n11072 0.00056
R20411 DVDD.n11083 DVDD.n11082 0.00056
R20412 DVDD.n15530 DVDD.n15527 0.00056
R20413 DVDD.n15518 DVDD.n11195 0.00056
R20414 DVDD.n11165 DVDD.n11164 0.00056
R20415 DVDD.n11152 DVDD.n11151 0.00056
R20416 DVDD.n16938 DVDD.n16937 0.00056
R20417 DVDD.n16935 DVDD.n16934 0.00056
R20418 DVDD.n16150 DVDD.n16149 0.00056
R20419 DVDD.n16162 DVDD.n16161 0.00056
R20420 DVDD.n16268 DVDD.n16267 0.00056
R20421 DVDD.n16280 DVDD.n16279 0.00056
R20422 DVDD.n16286 DVDD.n16285 0.00056
R20423 DVDD.n16290 DVDD.n16289 0.00056
R20424 DVDD.n16318 DVDD.n16317 0.00056
R20425 DVDD.n16325 DVDD.n16324 0.00056
R20426 DVDD.n16369 DVDD.n16368 0.00056
R20427 DVDD.n16206 DVDD.n16205 0.00056
R20428 DVDD.n16218 DVDD.n16217 0.00056
R20429 DVDD.n15571 DVDD.n15570 0.00056
R20430 DVDD.n15583 DVDD.n15582 0.00056
R20431 DVDD.n15752 DVDD.n15747 0.00056
R20432 DVDD.n15740 DVDD.n15739 0.00056
R20433 DVDD.n15716 DVDD.n15711 0.00056
R20434 DVDD.n15694 DVDD.n15693 0.00056
R20435 DVDD.n15785 DVDD.n15784 0.00056
R20436 DVDD.n15848 DVDD.n15847 0.00056
R20437 DVDD.n16112 DVDD.n16107 0.00056
R20438 DVDD.n16074 DVDD.n16069 0.00056
R20439 DVDD.n15906 DVDD.n15905 0.00056
R20440 DVDD.n15783 DVDD.n15782 0.00056
R20441 DVDD.n15846 DVDD.n15845 0.00056
R20442 DVDD.n16111 DVDD.n16110 0.00056
R20443 DVDD.n16073 DVDD.n16072 0.00056
R20444 DVDD.n16204 DVDD.n16203 0.00056
R20445 DVDD.n15569 DVDD.n15568 0.00056
R20446 DVDD.n15751 DVDD.n15750 0.00056
R20447 DVDD.n15715 DVDD.n15714 0.00056
R20448 DVDD.n16148 DVDD.n16147 0.00056
R20449 DVDD.n16266 DVDD.n16265 0.00056
R20450 DVDD.n11118 DVDD.n11117 0.00056
R20451 DVDD.n16378 DVDD.n16377 0.00056
R20452 DVDD.n11174 DVDD.n11173 0.00056
R20453 DVDD.n3620 DVDD.n3619 0.00056
R20454 DVDD.n3624 DVDD.n3623 0.00056
R20455 DVDD.n18608 DVDD.n18607 0.00056
R20456 DVDD.n18623 DVDD.n18622 0.00056
R20457 DVDD.n18637 DVDD.n18636 0.00056
R20458 DVDD.n18651 DVDD.n18650 0.00056
R20459 DVDD.n18729 DVDD.n18728 0.00056
R20460 DVDD.n18715 DVDD.n18714 0.00056
R20461 DVDD.n18711 DVDD.n18710 0.00056
R20462 DVDD.n18699 DVDD.n18698 0.00056
R20463 DVDD.n18688 DVDD.n18687 0.00056
R20464 DVDD.n18459 DVDD.n18458 0.00056
R20465 DVDD.n18417 DVDD.n18416 0.00056
R20466 DVDD.n18406 DVDD.n18405 0.00056
R20467 DVDD.n18405 DVDD.n18404 0.00056
R20468 DVDD.n18373 DVDD.n18372 0.00056
R20469 DVDD.n14788 DVDD.n14787 0.00056
R20470 DVDD.n14777 DVDD.n14776 0.00056
R20471 DVDD.n7171 DVDD.n7170 0.00056
R20472 DVDD.n7175 DVDD.n7174 0.00056
R20473 DVDD.n20267 DVDD.n20266 0.00056
R20474 DVDD.n7329 DVDD.n7327 0.00056
R20475 DVDD.n7687 DVDD.n7686 0.00056
R20476 DVDD.n14914 DVDD.n14913 0.00055625
R20477 DVDD.n14921 DVDD.n14920 0.00055625
R20478 DVDD.n14884 DVDD.n14883 0.00055625
R20479 DVDD.n15213 DVDD.n14904 0.00055625
R20480 DVDD.n15219 DVDD.n15218 0.00055625
R20481 DVDD.n15235 DVDD.n15234 0.00055625
R20482 DVDD.n15244 DVDD.n15243 0.00055625
R20483 DVDD.n15106 DVDD.n15105 0.00055625
R20484 DVDD.n15307 DVDD.n15306 0.00055625
R20485 DVDD.n15293 DVDD.n15292 0.00055625
R20486 DVDD.n15002 DVDD.n15001 0.00055625
R20487 DVDD.n10559 DVDD.n10558 0.00055625
R20488 DVDD.n1832 DVDD.n1831 0.00053
R20489 DVDD.n19557 DVDD.n19556 0.00053
R20490 DVDD.n19554 DVDD.n19553 0.00053
R20491 DVDD.n19542 DVDD.n19541 0.00053
R20492 DVDD.n19529 DVDD.n19528 0.00053
R20493 DVDD.n19526 DVDD.n19525 0.00053
R20494 DVDD.n19521 DVDD.n19520 0.00053
R20495 DVDD.n18875 DVDD.n18874 0.00053
R20496 DVDD.n18873 DVDD.n18872 0.00053
R20497 DVDD.n7575 DVDD.n7574 0.00053
R20498 DVDD.n19610 DVDD.n19609 0.00053
R20499 DVDD.n20172 DVDD.n20171 0.00053
R20500 DVDD.n20169 DVDD.n20168 0.00053
R20501 DVDD.n20157 DVDD.n20156 0.00053
R20502 DVDD.n20144 DVDD.n20143 0.00053
R20503 DVDD.n20141 DVDD.n20140 0.00053
R20504 DVDD.n20136 DVDD.n20135 0.00053
R20505 DVDD.n19124 DVDD.n19123 0.00053
R20506 DVDD.n19122 DVDD.n19121 0.00053
R20507 DVDD.n7531 DVDD.n7530 0.00053
R20508 DVDD.n7375 DVDD.n7373 0.00053
R20509 DVDD.n65 DVDD.n63 0.00053
R20510 DVDD.n7248 DVDD.n7246 0.00053
R20511 DVDD.n857 DVDD.n856 0.00053
R20512 DVDD.n231 DVDD.n230 0.00053
R20513 DVDD.n230 DVDD.n229 0.00053
R20514 DVDD.n227 DVDD.n226 0.00053
R20515 DVDD.n226 DVDD.n225 0.00053
R20516 DVDD.n212 DVDD.n211 0.00053
R20517 DVDD.n207 DVDD.n206 0.00053
R20518 DVDD.n203 DVDD.n202 0.00053
R20519 DVDD.n196 DVDD.n195 0.00053
R20520 DVDD.n192 DVDD.n191 0.00053
R20521 DVDD.n189 DVDD.n188 0.00053
R20522 DVDD.n186 DVDD.n185 0.00053
R20523 DVDD.n184 DVDD.n183 0.00053
R20524 DVDD.n163 DVDD.n162 0.00053
R20525 DVDD.n147 DVDD.n146 0.00053
R20526 DVDD.n19403 DVDD.n19402 0.00053
R20527 DVDD.n19400 DVDD.n19399 0.00053
R20528 DVDD.n19393 DVDD.n19392 0.00053
R20529 DVDD.n19389 DVDD.n19388 0.00053
R20530 DVDD.n18251 DVDD.n18250 0.00053
R20531 DVDD.n7180 DVDD.n7179 0.00053
R20532 DVDD.n7184 DVDD.n7183 0.00053
R20533 DVDD.n14965 DVDD.n14963 0.00053
R20534 DVDD.n15042 DVDD.n15040 0.00053
R20535 DVDD.n15325 DVDD.n14831 0.00053
R20536 DVDD.n15351 DVDD.n15349 0.00053
R20537 DVDD.n14953 DVDD.n14952 0.00053
R20538 DVDD.n14966 DVDD.n14959 0.00053
R20539 DVDD.n15043 DVDD.n15038 0.00053
R20540 DVDD.n15316 DVDD.n15315 0.00053
R20541 DVDD.n15324 DVDD.n15323 0.00053
R20542 DVDD.n15365 DVDD.n15364 0.00053
R20543 DVDD.n15353 DVDD.n15352 0.00053
R20544 DVDD.n11011 DVDD.n11010 0.00053
R20545 DVDD.n11024 DVDD.n11019 0.00053
R20546 DVDD.n11067 DVDD.n11066 0.00053
R20547 DVDD.n11079 DVDD.n11075 0.00053
R20548 DVDD.n15534 DVDD.n15533 0.00053
R20549 DVDD.n15525 DVDD.n15524 0.00053
R20550 DVDD.n11170 DVDD.n11169 0.00053
R20551 DVDD.n11160 DVDD.n11159 0.00053
R20552 DVDD.n17020 DVDD.n17019 0.00053
R20553 DVDD.n17016 DVDD.n17015 0.00053
R20554 DVDD.n16140 DVDD.n16139 0.00053
R20555 DVDD.n16142 DVDD.n16141 0.00053
R20556 DVDD.n16144 DVDD.n16143 0.00053
R20557 DVDD.n16158 DVDD.n16154 0.00053
R20558 DVDD.n16261 DVDD.n16260 0.00053
R20559 DVDD.n16276 DVDD.n16272 0.00053
R20560 DVDD.n16321 DVDD.n16320 0.00053
R20561 DVDD.n16364 DVDD.n16363 0.00053
R20562 DVDD.n16214 DVDD.n16210 0.00053
R20563 DVDD.n15579 DVDD.n15575 0.00053
R20564 DVDD.n15755 DVDD.n15754 0.00053
R20565 DVDD.n15745 DVDD.n15744 0.00053
R20566 DVDD.n15719 DVDD.n15718 0.00053
R20567 DVDD.n15709 DVDD.n15708 0.00053
R20568 DVDD.n15778 DVDD.n15777 0.00053
R20569 DVDD.n15793 DVDD.n15789 0.00053
R20570 DVDD.n15841 DVDD.n15840 0.00053
R20571 DVDD.n15856 DVDD.n15852 0.00053
R20572 DVDD.n16116 DVDD.n16115 0.00053
R20573 DVDD.n16105 DVDD.n16104 0.00053
R20574 DVDD.n16078 DVDD.n16077 0.00053
R20575 DVDD.n15919 DVDD.n15918 0.00053
R20576 DVDD.n15792 DVDD.n15790 0.00053
R20577 DVDD.n15855 DVDD.n15853 0.00053
R20578 DVDD.n16213 DVDD.n16211 0.00053
R20579 DVDD.n15578 DVDD.n15576 0.00053
R20580 DVDD.n16157 DVDD.n16155 0.00053
R20581 DVDD.n16275 DVDD.n16273 0.00053
R20582 DVDD.n11116 DVDD.n11115 0.00053
R20583 DVDD.n16362 DVDD.n16360 0.00053
R20584 DVDD.n11023 DVDD.n11021 0.00053
R20585 DVDD.n11078 DVDD.n11077 0.00053
R20586 DVDD.n15523 DVDD.n15521 0.00053
R20587 DVDD.n11158 DVDD.n11156 0.00053
R20588 DVDD.n3621 DVDD.n3620 0.00053
R20589 DVDD.n18591 DVDD.n18590 0.00053
R20590 DVDD.n18592 DVDD.n18591 0.00053
R20591 DVDD.n18602 DVDD.n18601 0.00053
R20592 DVDD.n18603 DVDD.n18602 0.00053
R20593 DVDD.n18624 DVDD.n18623 0.00053
R20594 DVDD.n18636 DVDD.n18635 0.00053
R20595 DVDD.n18650 DVDD.n18649 0.00053
R20596 DVDD.n18657 DVDD.n18656 0.00053
R20597 DVDD.n18734 DVDD.n18733 0.00053
R20598 DVDD.n18731 DVDD.n18730 0.00053
R20599 DVDD.n18728 DVDD.n18727 0.00053
R20600 DVDD.n18726 DVDD.n18725 0.00053
R20601 DVDD.n18684 DVDD.n18683 0.00053
R20602 DVDD.n18668 DVDD.n18662 0.00053
R20603 DVDD.n18410 DVDD.n18409 0.00053
R20604 DVDD.n18407 DVDD.n18406 0.00053
R20605 DVDD.n18400 DVDD.n18399 0.00053
R20606 DVDD.n18396 DVDD.n18395 0.00053
R20607 DVDD.n14776 DVDD.n14775 0.00053
R20608 DVDD.n7172 DVDD.n7171 0.00053
R20609 DVDD.n7690 DVDD.n7175 0.00053
R20610 DVDD.n20255 DVDD.n20253 0.00053
R20611 DVSS.n349 DVSS.n348 4017.81
R20612 DVSS.n343 DVSS.n342 4017.81
R20613 DVSS.n14893 DVSS.n14892 99.2437
R20614 DVSS.n3402 DVSS.n3401 32.468
R20615 DVSS.n12787 DVSS.n12786 32.468
R20616 DVSS.n2471 DVSS.n1742 11.6508
R20617 DVSS.n2484 DVSS.n2476 11.435
R20618 DVSS.n6729 DVSS.n6728 10.5721
R20619 DVSS.n357 DVSS.n356 7.57947
R20620 DVSS.n13728 DVSS.n13727 6.79968
R20621 DVSS.n7358 DVSS.n7356 6.79968
R20622 DVSS.n13766 DVSS.n13765 6.79968
R20623 DVSS.n7383 DVSS.n7382 6.79968
R20624 DVSS.n2374 DVSS.n2373 5.91395
R20625 DVSS.n11713 DVSS.n11712 5.86071
R20626 DVSS.n8036 DVSS.n8035 5.86071
R20627 DVSS.n1374 DVSS.n1373 5.84304
R20628 DVSS.n6400 DVSS.n6399 5.84304
R20629 DVSS.n2539 DVSS.n2538 5.84304
R20630 DVSS.n6707 DVSS.n6706 5.84304
R20631 DVSS.n6762 DVSS.n6761 5.84304
R20632 DVSS.n6889 DVSS.n6888 5.84304
R20633 DVSS.n4523 DVSS.n4522 5.84304
R20634 DVSS.n5507 DVSS.n5506 5.84304
R20635 DVSS.n5402 DVSS.n5401 5.84304
R20636 DVSS.n4577 DVSS.n4576 5.84304
R20637 DVSS.n1747 DVSS.n1746 5.7217
R20638 DVSS.n1733 DVSS.n1730 5.70148
R20639 DVSS.n1899 DVSS.n1897 5.70148
R20640 DVSS.n14944 DVSS.n14943 5.2293
R20641 DVSS.n7434 DVSS.n7433 5.2293
R20642 DVSS.n13805 DVSS.n13804 5.2005
R20643 DVSS.n7403 DVSS.n7402 5.2005
R20644 DVSS.n13807 DVSS.n13806 5.2005
R20645 DVSS.n7405 DVSS.n7404 5.2005
R20646 DVSS.n13733 DVSS.n13732 5.2005
R20647 DVSS.n7363 DVSS.n7362 5.2005
R20648 DVSS.n7348 DVSS.n7347 5.2005
R20649 DVSS.n7355 DVSS.n7354 5.2005
R20650 DVSS.n7354 DVSS.n7353 5.2005
R20651 DVSS.n7845 DVSS.n7844 5.2005
R20652 DVSS.n13726 DVSS.n13725 5.2005
R20653 DVSS.n13725 DVSS.n13724 5.2005
R20654 DVSS.n351 DVSS.n350 5.2005
R20655 DVSS.n350 DVSS.n349 5.2005
R20656 DVSS.n353 DVSS.n352 5.2005
R20657 DVSS.n11475 DVSS.n11474 5.2005
R20658 DVSS.n11474 DVSS.n11473 5.2005
R20659 DVSS.n11476 DVSS.n11471 5.2005
R20660 DVSS.n11476 DVSS.n11470 5.2005
R20661 DVSS.n6402 DVSS.n6401 5.2005
R20662 DVSS.n6432 DVSS.n6431 5.2005
R20663 DVSS.n6420 DVSS.n6419 5.2005
R20664 DVSS.n6417 DVSS.n6416 5.2005
R20665 DVSS.n6412 DVSS.n6411 5.2005
R20666 DVSS.n6407 DVSS.n6406 5.2005
R20667 DVSS.n4474 DVSS.n4473 5.2005
R20668 DVSS.n16262 DVSS.n16261 5.2005
R20669 DVSS.n16268 DVSS.n16267 5.2005
R20670 DVSS.n16284 DVSS.n16283 5.2005
R20671 DVSS.n16281 DVSS.n16280 5.2005
R20672 DVSS.n16278 DVSS.n16277 5.2005
R20673 DVSS.n7622 DVSS.n7621 5.2005
R20674 DVSS.n17942 DVSS.n17941 5.2005
R20675 DVSS.n7670 DVSS.n7669 5.2005
R20676 DVSS.n15830 DVSS.n15829 5.2005
R20677 DVSS.n15834 DVSS.n15833 5.2005
R20678 DVSS.n15839 DVSS.n15838 5.2005
R20679 DVSS.n15844 DVSS.n15843 5.2005
R20680 DVSS.n15852 DVSS.n15851 5.2005
R20681 DVSS.n8930 DVSS.n8929 5.2005
R20682 DVSS.n8935 DVSS.n8934 5.2005
R20683 DVSS.n9795 DVSS.n9794 5.2005
R20684 DVSS.n9792 DVSS.n9791 5.2005
R20685 DVSS.n9789 DVSS.n9788 5.2005
R20686 DVSS.n9786 DVSS.n9785 5.2005
R20687 DVSS.n9783 DVSS.n9782 5.2005
R20688 DVSS.n8952 DVSS.n8951 5.2005
R20689 DVSS.n8949 DVSS.n8948 5.2005
R20690 DVSS.n11463 DVSS.n11462 5.2005
R20691 DVSS.n11476 DVSS.n11469 5.2005
R20692 DVSS.n11476 DVSS.n11468 5.2005
R20693 DVSS.n11513 DVSS.n11509 5.2005
R20694 DVSS.n11513 DVSS.n11511 5.2005
R20695 DVSS.n2541 DVSS.n2540 5.2005
R20696 DVSS.n6568 DVSS.n6567 5.2005
R20697 DVSS.n6556 DVSS.n6555 5.2005
R20698 DVSS.n6553 DVSS.n6552 5.2005
R20699 DVSS.n6548 DVSS.n6547 5.2005
R20700 DVSS.n6543 DVSS.n6542 5.2005
R20701 DVSS.n6538 DVSS.n6537 5.2005
R20702 DVSS.n16223 DVSS.n16222 5.2005
R20703 DVSS.n16229 DVSS.n16228 5.2005
R20704 DVSS.n16245 DVSS.n16244 5.2005
R20705 DVSS.n16242 DVSS.n16241 5.2005
R20706 DVSS.n16239 DVSS.n16238 5.2005
R20707 DVSS.n7614 DVSS.n7613 5.2005
R20708 DVSS.n18083 DVSS.n18082 5.2005
R20709 DVSS.n7678 DVSS.n7677 5.2005
R20710 DVSS.n15732 DVSS.n15731 5.2005
R20711 DVSS.n15729 DVSS.n15728 5.2005
R20712 DVSS.n15726 DVSS.n15725 5.2005
R20713 DVSS.n15723 DVSS.n15722 5.2005
R20714 DVSS.n7693 DVSS.n7692 5.2005
R20715 DVSS.n8955 DVSS.n8954 5.2005
R20716 DVSS.n8960 DVSS.n8959 5.2005
R20717 DVSS.n9722 DVSS.n9721 5.2005
R20718 DVSS.n9727 DVSS.n9726 5.2005
R20719 DVSS.n9731 DVSS.n9730 5.2005
R20720 DVSS.n9736 DVSS.n9735 5.2005
R20721 DVSS.n9741 DVSS.n9740 5.2005
R20722 DVSS.n9749 DVSS.n9748 5.2005
R20723 DVSS.n9746 DVSS.n9745 5.2005
R20724 DVSS.n11500 DVSS.n11499 5.2005
R20725 DVSS.n11513 DVSS.n11508 5.2005
R20726 DVSS.n11513 DVSS.n11512 5.2005
R20727 DVSS.n11632 DVSS.n11631 5.2005
R20728 DVSS.n11631 DVSS.n11630 5.2005
R20729 DVSS.n11638 DVSS.n11634 5.2005
R20730 DVSS.n11638 DVSS.n11636 5.2005
R20731 DVSS.n6709 DVSS.n6708 5.2005
R20732 DVSS.n6711 DVSS.n6710 5.2005
R20733 DVSS.n2551 DVSS.n2550 5.2005
R20734 DVSS.n2556 DVSS.n2555 5.2005
R20735 DVSS.n4355 DVSS.n4354 5.2005
R20736 DVSS.n4359 DVSS.n4358 5.2005
R20737 DVSS.n4364 DVSS.n4363 5.2005
R20738 DVSS.n4369 DVSS.n4368 5.2005
R20739 DVSS.n4374 DVSS.n4373 5.2005
R20740 DVSS.n7551 DVSS.n7550 5.2005
R20741 DVSS.n7557 DVSS.n7556 5.2005
R20742 DVSS.n18374 DVSS.n18373 5.2005
R20743 DVSS.n18371 DVSS.n18370 5.2005
R20744 DVSS.n18368 DVSS.n18367 5.2005
R20745 DVSS.n18365 DVSS.n18364 5.2005
R20746 DVSS.n18362 DVSS.n18361 5.2005
R20747 DVSS.n7699 DVSS.n7698 5.2005
R20748 DVSS.n15584 DVSS.n15583 5.2005
R20749 DVSS.n15588 DVSS.n15587 5.2005
R20750 DVSS.n15593 DVSS.n15592 5.2005
R20751 DVSS.n15598 DVSS.n15597 5.2005
R20752 DVSS.n15606 DVSS.n15605 5.2005
R20753 DVSS.n8963 DVSS.n8962 5.2005
R20754 DVSS.n8968 DVSS.n8967 5.2005
R20755 DVSS.n9603 DVSS.n9602 5.2005
R20756 DVSS.n9600 DVSS.n9599 5.2005
R20757 DVSS.n9597 DVSS.n9596 5.2005
R20758 DVSS.n9594 DVSS.n9593 5.2005
R20759 DVSS.n9591 DVSS.n9590 5.2005
R20760 DVSS.n8985 DVSS.n8984 5.2005
R20761 DVSS.n8982 DVSS.n8981 5.2005
R20762 DVSS.n11625 DVSS.n11624 5.2005
R20763 DVSS.n11638 DVSS.n11633 5.2005
R20764 DVSS.n11638 DVSS.n11637 5.2005
R20765 DVSS.n11669 DVSS.n11668 5.2005
R20766 DVSS.n11668 DVSS.n11667 5.2005
R20767 DVSS.n11675 DVSS.n11671 5.2005
R20768 DVSS.n11675 DVSS.n11673 5.2005
R20769 DVSS.n6764 DVSS.n6763 5.2005
R20770 DVSS.n6766 DVSS.n6765 5.2005
R20771 DVSS.n2564 DVSS.n2563 5.2005
R20772 DVSS.n2569 DVSS.n2568 5.2005
R20773 DVSS.n4115 DVSS.n4114 5.2005
R20774 DVSS.n4112 DVSS.n4111 5.2005
R20775 DVSS.n4107 DVSS.n4106 5.2005
R20776 DVSS.n4102 DVSS.n4101 5.2005
R20777 DVSS.n4097 DVSS.n4096 5.2005
R20778 DVSS.n7462 DVSS.n7461 5.2005
R20779 DVSS.n7468 DVSS.n7467 5.2005
R20780 DVSS.n18394 DVSS.n18393 5.2005
R20781 DVSS.n18399 DVSS.n18398 5.2005
R20782 DVSS.n18403 DVSS.n18402 5.2005
R20783 DVSS.n18408 DVSS.n18407 5.2005
R20784 DVSS.n18414 DVSS.n18413 5.2005
R20785 DVSS.n15248 DVSS.n15247 5.2005
R20786 DVSS.n7710 DVSS.n7709 5.2005
R20787 DVSS.n14959 DVSS.n14958 5.2005
R20788 DVSS.n14964 DVSS.n14963 5.2005
R20789 DVSS.n14969 DVSS.n14968 5.2005
R20790 DVSS.n14977 DVSS.n14976 5.2005
R20791 DVSS.n9005 DVSS.n9004 5.2005
R20792 DVSS.n9010 DVSS.n9009 5.2005
R20793 DVSS.n9110 DVSS.n9109 5.2005
R20794 DVSS.n9115 DVSS.n9114 5.2005
R20795 DVSS.n9119 DVSS.n9118 5.2005
R20796 DVSS.n9124 DVSS.n9123 5.2005
R20797 DVSS.n9129 DVSS.n9128 5.2005
R20798 DVSS.n9137 DVSS.n9136 5.2005
R20799 DVSS.n9134 DVSS.n9133 5.2005
R20800 DVSS.n11662 DVSS.n11661 5.2005
R20801 DVSS.n11675 DVSS.n11670 5.2005
R20802 DVSS.n11675 DVSS.n11674 5.2005
R20803 DVSS.n11718 DVSS.n11717 5.2005
R20804 DVSS.n11717 DVSS.n11716 5.2005
R20805 DVSS.n8024 DVSS.n8023 5.2005
R20806 DVSS.n6485 DVSS.n6484 5.2005
R20807 DVSS.n6481 DVSS.n6480 5.2005
R20808 DVSS.n11009 DVSS.n11008 5.2005
R20809 DVSS.n4525 DVSS.n4524 5.2005
R20810 DVSS.n6476 DVSS.n6475 5.2005
R20811 DVSS.n11197 DVSS.n11196 5.2005
R20812 DVSS.n11205 DVSS.n11204 5.2005
R20813 DVSS.n11172 DVSS.n11171 5.2005
R20814 DVSS.n11211 DVSS.n11210 5.2005
R20815 DVSS.n11208 DVSS.n11207 5.2005
R20816 DVSS.n11167 DVSS.n11166 5.2005
R20817 DVSS.n9821 DVSS.n9820 5.2005
R20818 DVSS.n9830 DVSS.n9829 5.2005
R20819 DVSS.n9827 DVSS.n9826 5.2005
R20820 DVSS.n9816 DVSS.n9815 5.2005
R20821 DVSS.n17656 DVSS.n17655 5.2005
R20822 DVSS.n7664 DVSS.n7663 5.2005
R20823 DVSS.n7661 DVSS.n7660 5.2005
R20824 DVSS.n17661 DVSS.n17660 5.2005
R20825 DVSS.n16333 DVSS.n16332 5.2005
R20826 DVSS.n7633 DVSS.n7632 5.2005
R20827 DVSS.n7653 DVSS.n7652 5.2005
R20828 DVSS.n7650 DVSS.n7649 5.2005
R20829 DVSS.n11179 DVSS.n11178 5.2005
R20830 DVSS.n11185 DVSS.n11181 5.2005
R20831 DVSS.n11015 DVSS.n11011 5.2005
R20832 DVSS.n4579 DVSS.n4578 5.2005
R20833 DVSS.n11036 DVSS.n11035 5.2005
R20834 DVSS.n11041 DVSS.n11040 5.2005
R20835 DVSS.n11049 DVSS.n11048 5.2005
R20836 DVSS.n11054 DVSS.n11053 5.2005
R20837 DVSS.n11058 DVSS.n11057 5.2005
R20838 DVSS.n11063 DVSS.n11062 5.2005
R20839 DVSS.n11072 DVSS.n11071 5.2005
R20840 DVSS.n11070 DVSS.n11069 5.2005
R20841 DVSS.n16894 DVSS.n16893 5.2005
R20842 DVSS.n16899 DVSS.n16898 5.2005
R20843 DVSS.n17549 DVSS.n17548 5.2005
R20844 DVSS.n17547 DVSS.n17546 5.2005
R20845 DVSS.n17543 DVSS.n17542 5.2005
R20846 DVSS.n17534 DVSS.n17533 5.2005
R20847 DVSS.n17276 DVSS.n17275 5.2005
R20848 DVSS.n5386 DVSS.n5385 5.2005
R20849 DVSS.n5400 DVSS.n5399 5.2005
R20850 DVSS.n10261 DVSS.n10260 5.2005
R20851 DVSS.n10266 DVSS.n10265 5.2005
R20852 DVSS.n10245 DVSS.n10244 5.2005
R20853 DVSS.n10213 DVSS.n10212 5.2005
R20854 DVSS.n16993 DVSS.n16992 5.2005
R20855 DVSS.n17301 DVSS.n17300 5.2005
R20856 DVSS.n17296 DVSS.n17295 5.2005
R20857 DVSS.n17293 DVSS.n17292 5.2005
R20858 DVSS.n17290 DVSS.n17289 5.2005
R20859 DVSS.n10252 DVSS.n10251 5.2005
R20860 DVSS.n10278 DVSS.n10277 5.2005
R20861 DVSS.n10282 DVSS.n10281 5.2005
R20862 DVSS.n10289 DVSS.n10288 5.2005
R20863 DVSS.n10220 DVSS.n10219 5.2005
R20864 DVSS.n10227 DVSS.n10226 5.2005
R20865 DVSS.n10232 DVSS.n10231 5.2005
R20866 DVSS.n10239 DVSS.n10238 5.2005
R20867 DVSS.n17000 DVSS.n16999 5.2005
R20868 DVSS.n17017 DVSS.n17016 5.2005
R20869 DVSS.n17021 DVSS.n17020 5.2005
R20870 DVSS.n17028 DVSS.n17027 5.2005
R20871 DVSS.n16977 DVSS.n16976 5.2005
R20872 DVSS.n16982 DVSS.n16981 5.2005
R20873 DVSS.n16987 DVSS.n16986 5.2005
R20874 DVSS.n5381 DVSS.n5380 5.2005
R20875 DVSS.n5376 DVSS.n5375 5.2005
R20876 DVSS.n5373 DVSS.n5372 5.2005
R20877 DVSS.n5368 DVSS.n5367 5.2005
R20878 DVSS.n5363 DVSS.n5362 5.2005
R20879 DVSS.n10624 DVSS.n10622 5.2005
R20880 DVSS.n10624 DVSS.n10620 5.2005
R20881 DVSS.n10624 DVSS.n10623 5.2005
R20882 DVSS.n10019 DVSS.n10018 5.2005
R20883 DVSS.n10018 DVSS.n10017 5.2005
R20884 DVSS.n5606 DVSS.n5605 5.2005
R20885 DVSS.n5594 DVSS.n5593 5.2005
R20886 DVSS.n17321 DVSS.n17320 5.2005
R20887 DVSS.n17324 DVSS.n17323 5.2005
R20888 DVSS.n17312 DVSS.n17311 5.2005
R20889 DVSS.n17315 DVSS.n17314 5.2005
R20890 DVSS.n5578 DVSS.n5577 5.2005
R20891 DVSS.n5597 DVSS.n5596 5.2005
R20892 DVSS.n11015 DVSS.n11013 5.2005
R20893 DVSS.n17461 DVSS.n17460 5.2005
R20894 DVSS.n17453 DVSS.n17452 5.2005
R20895 DVSS.n17451 DVSS.n17450 5.2005
R20896 DVSS.n16126 DVSS.n16125 5.2005
R20897 DVSS.n17444 DVSS.n17443 5.2005
R20898 DVSS.n17440 DVSS.n17439 5.2005
R20899 DVSS.n17434 DVSS.n17433 5.2005
R20900 DVSS.n5808 DVSS.n5807 5.2005
R20901 DVSS.n4583 DVSS.n4582 5.2005
R20902 DVSS.n5818 DVSS.n5817 5.2005
R20903 DVSS.n5823 DVSS.n5822 5.2005
R20904 DVSS.n5827 DVSS.n5826 5.2005
R20905 DVSS.n5832 DVSS.n5831 5.2005
R20906 DVSS.n11032 DVSS.n11031 5.2005
R20907 DVSS.n11026 DVSS.n11025 5.2005
R20908 DVSS.n11015 DVSS.n11010 5.2005
R20909 DVSS.n11015 DVSS.n11014 5.2005
R20910 DVSS.n16338 DVSS.n16337 5.2005
R20911 DVSS.n6501 DVSS.n6500 5.2005
R20912 DVSS.n6498 DVSS.n6497 5.2005
R20913 DVSS.n6495 DVSS.n6494 5.2005
R20914 DVSS.n16307 DVSS.n16306 5.2005
R20915 DVSS.n16312 DVSS.n16311 5.2005
R20916 DVSS.n16319 DVSS.n16318 5.2005
R20917 DVSS.n16314 DVSS.n16313 5.2005
R20918 DVSS.n11185 DVSS.n11183 5.2005
R20919 DVSS.n11185 DVSS.n11180 5.2005
R20920 DVSS.n11185 DVSS.n11184 5.2005
R20921 DVSS.n1901 DVSS.n1900 5.2005
R20922 DVSS.n1873 DVSS.n1872 5.2005
R20923 DVSS.n1872 DVSS.n1871 5.2005
R20924 DVSS.n1866 DVSS.n1865 5.2005
R20925 DVSS.n1860 DVSS.n1859 5.2005
R20926 DVSS.n1859 DVSS.n1858 5.2005
R20927 DVSS.n1852 DVSS.n1851 5.2005
R20928 DVSS.n1851 DVSS.n1850 5.2005
R20929 DVSS.n1844 DVSS.n1843 5.2005
R20930 DVSS.n1843 DVSS.n1842 5.2005
R20931 DVSS.n1837 DVSS.n1836 5.2005
R20932 DVSS.n1830 DVSS.n1829 5.2005
R20933 DVSS.n1824 DVSS.n1823 5.2005
R20934 DVSS.n1823 DVSS.n1822 5.2005
R20935 DVSS.n1817 DVSS.n1816 5.2005
R20936 DVSS.n1810 DVSS.n1809 5.2005
R20937 DVSS.n1804 DVSS.n1803 5.2005
R20938 DVSS.n1803 DVSS.n1802 5.2005
R20939 DVSS.n1797 DVSS.n1796 5.2005
R20940 DVSS.n1796 DVSS.n1795 5.2005
R20941 DVSS.n1789 DVSS.n1788 5.2005
R20942 DVSS.n1788 DVSS.n1787 5.2005
R20943 DVSS.n1781 DVSS.n1780 5.2005
R20944 DVSS.n1774 DVSS.n1773 5.2005
R20945 DVSS.n1767 DVSS.n1766 5.2005
R20946 DVSS.n1766 DVSS.n1765 5.2005
R20947 DVSS.n1760 DVSS.n1759 5.2005
R20948 DVSS.n1753 DVSS.n1752 5.2005
R20949 DVSS.n1752 DVSS.n1751 5.2005
R20950 DVSS.n1495 DVSS.n1494 5.2005
R20951 DVSS.n1494 DVSS.n1493 5.2005
R20952 DVSS.n1500 DVSS.n1499 5.2005
R20953 DVSS.n1480 DVSS.n1479 5.2005
R20954 DVSS.n1488 DVSS.n1487 5.2005
R20955 DVSS.n1487 DVSS.n1486 5.2005
R20956 DVSS.n10016 DVSS.n10014 5.2005
R20957 DVSS.n1411 DVSS.n1410 5.2005
R20958 DVSS.n1418 DVSS.n1417 5.2005
R20959 DVSS.n1417 DVSS.n1416 5.2005
R20960 DVSS.n1425 DVSS.n1424 5.2005
R20961 DVSS.n1432 DVSS.n1431 5.2005
R20962 DVSS.n1431 DVSS.n1430 5.2005
R20963 DVSS.n1439 DVSS.n1438 5.2005
R20964 DVSS.n1438 DVSS.n1437 5.2005
R20965 DVSS.n1445 DVSS.n1444 5.2005
R20966 DVSS.n1451 DVSS.n1450 5.2005
R20967 DVSS.n1458 DVSS.n1457 5.2005
R20968 DVSS.n1466 DVSS.n1465 5.2005
R20969 DVSS.n1465 DVSS.n1464 5.2005
R20970 DVSS.n1473 DVSS.n1472 5.2005
R20971 DVSS.n1472 DVSS.n1471 5.2005
R20972 DVSS.n1506 DVSS.n1505 5.2005
R20973 DVSS.n1512 DVSS.n1511 5.2005
R20974 DVSS.n1520 DVSS.n1519 5.2005
R20975 DVSS.n1519 DVSS.n1518 5.2005
R20976 DVSS.n1527 DVSS.n1526 5.2005
R20977 DVSS.n1736 DVSS.n1735 5.2005
R20978 DVSS.n1735 DVSS.n1734 5.2005
R20979 DVSS.n10016 DVSS.n10015 5.2005
R20980 DVSS.n6728 DVSS.n6726 5.2005
R20981 DVSS.n6728 DVSS.n6727 5.2005
R20982 DVSS.n345 DVSS.n344 5.2005
R20983 DVSS.n344 DVSS.n343 5.2005
R20984 DVSS.n347 DVSS.n346 5.2005
R20985 DVSS.n21215 DVSS.n21214 5.2005
R20986 DVSS.n12813 DVSS.n12812 5.2005
R20987 DVSS.n12768 DVSS.n12767 5.2005
R20988 DVSS.n12140 DVSS.n12139 5.2005
R20989 DVSS.n12148 DVSS.n12147 5.2005
R20990 DVSS.n12739 DVSS.n12738 5.2005
R20991 DVSS.n12505 DVSS.n12504 5.2005
R20992 DVSS.n12513 DVSS.n12512 5.2005
R20993 DVSS.n12520 DVSS.n12519 5.2005
R20994 DVSS.n12527 DVSS.n12526 5.2005
R20995 DVSS.n12535 DVSS.n12534 5.2005
R20996 DVSS.n12543 DVSS.n12542 5.2005
R20997 DVSS.n12550 DVSS.n12549 5.2005
R20998 DVSS.n12552 DVSS.n12551 5.2005
R20999 DVSS.n12667 DVSS.n12666 5.2005
R21000 DVSS.n12659 DVSS.n12658 5.2005
R21001 DVSS.n12651 DVSS.n12650 5.2005
R21002 DVSS.n12644 DVSS.n12643 5.2005
R21003 DVSS.n12637 DVSS.n12636 5.2005
R21004 DVSS.n12629 DVSS.n12628 5.2005
R21005 DVSS.n12621 DVSS.n12620 5.2005
R21006 DVSS.n12613 DVSS.n12612 5.2005
R21007 DVSS.n12605 DVSS.n12604 5.2005
R21008 DVSS.n12597 DVSS.n12596 5.2005
R21009 DVSS.n12589 DVSS.n12588 5.2005
R21010 DVSS.n12582 DVSS.n12581 5.2005
R21011 DVSS.n12575 DVSS.n12574 5.2005
R21012 DVSS.n12567 DVSS.n12566 5.2005
R21013 DVSS.n12217 DVSS.n12216 5.2005
R21014 DVSS.n12219 DVSS.n12218 5.2005
R21015 DVSS.n12379 DVSS.n12378 5.2005
R21016 DVSS.n12371 DVSS.n12370 5.2005
R21017 DVSS.n12363 DVSS.n12362 5.2005
R21018 DVSS.n12356 DVSS.n12355 5.2005
R21019 DVSS.n12349 DVSS.n12348 5.2005
R21020 DVSS.n12341 DVSS.n12340 5.2005
R21021 DVSS.n12333 DVSS.n12332 5.2005
R21022 DVSS.n12325 DVSS.n12324 5.2005
R21023 DVSS.n12317 DVSS.n12316 5.2005
R21024 DVSS.n12309 DVSS.n12308 5.2005
R21025 DVSS.n12301 DVSS.n12300 5.2005
R21026 DVSS.n12294 DVSS.n12293 5.2005
R21027 DVSS.n12287 DVSS.n12286 5.2005
R21028 DVSS.n12279 DVSS.n12278 5.2005
R21029 DVSS.n12271 DVSS.n12270 5.2005
R21030 DVSS.n12263 DVSS.n12262 5.2005
R21031 DVSS.n12255 DVSS.n12254 5.2005
R21032 DVSS.n12247 DVSS.n12246 5.2005
R21033 DVSS.n12240 DVSS.n12239 5.2005
R21034 DVSS.n12233 DVSS.n12232 5.2005
R21035 DVSS.n12225 DVSS.n12224 5.2005
R21036 DVSS.n21335 DVSS.n21334 5.2005
R21037 DVSS.n21337 DVSS.n21336 5.2005
R21038 DVSS.n21320 DVSS.n21319 5.2005
R21039 DVSS.n21160 DVSS.n21159 5.2005
R21040 DVSS.n19156 DVSS.n19155 5.2005
R21041 DVSS.n19155 DVSS.n19154 5.2005
R21042 DVSS.n20388 DVSS.n20387 5.2005
R21043 DVSS.n20387 DVSS.n20386 5.2005
R21044 DVSS.n1328 DVSS.n1327 5.2005
R21045 DVSS.n13341 DVSS.n13340 5.2005
R21046 DVSS.n13290 DVSS.n13289 5.2005
R21047 DVSS.n7020 DVSS.n7019 5.2005
R21048 DVSS.n8029 DVSS.n8027 5.2005
R21049 DVSS.n8029 DVSS.n8025 5.2005
R21050 DVSS.n8029 DVSS.n8028 5.2005
R21051 DVSS.n11724 DVSS.n11720 5.2005
R21052 DVSS.n11724 DVSS.n11722 5.2005
R21053 DVSS.n6891 DVSS.n6890 5.2005
R21054 DVSS.n6893 DVSS.n6892 5.2005
R21055 DVSS.n2579 DVSS.n2578 5.2005
R21056 DVSS.n4006 DVSS.n4005 5.2005
R21057 DVSS.n4011 DVSS.n4010 5.2005
R21058 DVSS.n4015 DVSS.n4014 5.2005
R21059 DVSS.n4020 DVSS.n4019 5.2005
R21060 DVSS.n4025 DVSS.n4024 5.2005
R21061 DVSS.n4031 DVSS.n4030 5.2005
R21062 DVSS.n7472 DVSS.n7471 5.2005
R21063 DVSS.n7478 DVSS.n7477 5.2005
R21064 DVSS.n7496 DVSS.n7495 5.2005
R21065 DVSS.n7493 DVSS.n7492 5.2005
R21066 DVSS.n7490 DVSS.n7489 5.2005
R21067 DVSS.n7487 DVSS.n7486 5.2005
R21068 DVSS.n7457 DVSS.n7456 5.2005
R21069 DVSS.n15059 DVSS.n15058 5.2005
R21070 DVSS.n15056 DVSS.n15055 5.2005
R21071 DVSS.n15053 DVSS.n15052 5.2005
R21072 DVSS.n15050 DVSS.n15049 5.2005
R21073 DVSS.n15047 DVSS.n15046 5.2005
R21074 DVSS.n7783 DVSS.n7782 5.2005
R21075 DVSS.n7779 DVSS.n7778 5.2005
R21076 DVSS.n9015 DVSS.n9014 5.2005
R21077 DVSS.n9038 DVSS.n9037 5.2005
R21078 DVSS.n9035 DVSS.n9034 5.2005
R21079 DVSS.n9032 DVSS.n9031 5.2005
R21080 DVSS.n9029 DVSS.n9028 5.2005
R21081 DVSS.n9026 DVSS.n9025 5.2005
R21082 DVSS.n8058 DVSS.n8057 5.2005
R21083 DVSS.n8055 DVSS.n8054 5.2005
R21084 DVSS.n11711 DVSS.n11710 5.2005
R21085 DVSS.n11724 DVSS.n11719 5.2005
R21086 DVSS.n11724 DVSS.n11723 5.2005
R21087 DVSS.n1352 DVSS.n1351 5.2005
R21088 DVSS.n1351 DVSS.n1350 5.2005
R21089 DVSS.n6877 DVSS.n6876 5.2005
R21090 DVSS.n6872 DVSS.n6871 5.2005
R21091 DVSS.n6859 DVSS.n6858 5.2005
R21092 DVSS.n6854 DVSS.n6853 5.2005
R21093 DVSS.n6850 DVSS.n6849 5.2005
R21094 DVSS.n6750 DVSS.n6749 5.2005
R21095 DVSS.n6745 DVSS.n6744 5.2005
R21096 DVSS.n6741 DVSS.n6740 5.2005
R21097 DVSS.n6736 DVSS.n6735 5.2005
R21098 DVSS.n6732 DVSS.n6731 5.2005
R21099 DVSS.n6695 DVSS.n6694 5.2005
R21100 DVSS.n6690 DVSS.n6689 5.2005
R21101 DVSS.n6677 DVSS.n6676 5.2005
R21102 DVSS.n6672 DVSS.n6671 5.2005
R21103 DVSS.n6668 DVSS.n6667 5.2005
R21104 DVSS.n2527 DVSS.n2526 5.2005
R21105 DVSS.n2518 DVSS.n2517 5.2005
R21106 DVSS.n2497 DVSS.n2496 5.2005
R21107 DVSS.n2488 DVSS.n2487 5.2005
R21108 DVSS.n6388 DVSS.n6387 5.2005
R21109 DVSS.n6383 DVSS.n6382 5.2005
R21110 DVSS.n6370 DVSS.n6369 5.2005
R21111 DVSS.n6365 DVSS.n6364 5.2005
R21112 DVSS.n6361 DVSS.n6360 5.2005
R21113 DVSS.n4510 DVSS.n4509 5.2005
R21114 DVSS.n4505 DVSS.n4504 5.2005
R21115 DVSS.n4492 DVSS.n4491 5.2005
R21116 DVSS.n4487 DVSS.n4486 5.2005
R21117 DVSS.n4483 DVSS.n4482 5.2005
R21118 DVSS.n4482 DVSS.n4481 5.2005
R21119 DVSS.n4564 DVSS.n4563 5.2005
R21120 DVSS.n4559 DVSS.n4558 5.2005
R21121 DVSS.n4542 DVSS.n4541 5.2005
R21122 DVSS.n4537 DVSS.n4536 5.2005
R21123 DVSS.n4533 DVSS.n4532 5.2005
R21124 DVSS.n4532 DVSS.n4531 5.2005
R21125 DVSS.n4587 DVSS.n4586 5.2005
R21126 DVSS.n5338 DVSS.n5337 5.2005
R21127 DVSS.n5343 DVSS.n5342 5.2005
R21128 DVSS.n5346 DVSS.n5345 5.2005
R21129 DVSS.n4612 DVSS.n4611 5.2005
R21130 DVSS.n4609 DVSS.n4608 5.2005
R21131 DVSS.n4596 DVSS.n4595 5.2005
R21132 DVSS.n4591 DVSS.n4590 5.2005
R21133 DVSS.n5548 DVSS.n5547 5.2005
R21134 DVSS.n5536 DVSS.n5535 5.2005
R21135 DVSS.n5527 DVSS.n5526 5.2005
R21136 DVSS.n5517 DVSS.n5516 5.2005
R21137 DVSS.n5509 DVSS.n5508 5.2005
R21138 DVSS.n5522 DVSS.n5521 5.2005
R21139 DVSS.n5532 DVSS.n5531 5.2005
R21140 DVSS.n5551 DVSS.n5550 5.2005
R21141 DVSS.n5545 DVSS.n5544 5.2005
R21142 DVSS.n16427 DVSS.n16426 5.2005
R21143 DVSS.n10037 DVSS.n10036 5.2005
R21144 DVSS.n10044 DVSS.n10043 5.2005
R21145 DVSS.n10052 DVSS.n10051 5.2005
R21146 DVSS.n10002 DVSS.n10001 5.2005
R21147 DVSS.n9993 DVSS.n9992 5.2005
R21148 DVSS.n9853 DVSS.n9852 5.2005
R21149 DVSS.n16888 DVSS.n16887 5.2005
R21150 DVSS.n17107 DVSS.n17106 5.2005
R21151 DVSS.n16872 DVSS.n16871 5.2005
R21152 DVSS.n17246 DVSS.n17245 5.2005
R21153 DVSS.n17238 DVSS.n17237 5.2005
R21154 DVSS.n10047 DVSS.n10046 5.2005
R21155 DVSS.n10006 DVSS.n10005 5.2005
R21156 DVSS.n9998 DVSS.n9997 5.2005
R21157 DVSS.n9858 DVSS.n9857 5.2005
R21158 DVSS.n16883 DVSS.n16882 5.2005
R21159 DVSS.n17104 DVSS.n17103 5.2005
R21160 DVSS.n17110 DVSS.n17109 5.2005
R21161 DVSS.n17243 DVSS.n17242 5.2005
R21162 DVSS.n16442 DVSS.n16441 5.2005
R21163 DVSS.n16437 DVSS.n16436 5.2005
R21164 DVSS.n10025 DVSS.n10021 5.2005
R21165 DVSS.n10025 DVSS.n10023 5.2005
R21166 DVSS.n10025 DVSS.n10020 5.2005
R21167 DVSS.n10025 DVSS.n10024 5.2005
R21168 DVSS.n16432 DVSS.n16431 5.2005
R21169 DVSS.n925 DVSS.n923 5.2005
R21170 DVSS.n911 DVSS.n910 5.2005
R21171 DVSS.n903 DVSS.n902 5.2005
R21172 DVSS.n895 DVSS.n894 5.2005
R21173 DVSS.n887 DVSS.n886 5.2005
R21174 DVSS.n879 DVSS.n878 5.2005
R21175 DVSS.n2860 DVSS.n2859 5.2005
R21176 DVSS.n2867 DVSS.n2866 5.2005
R21177 DVSS.n2874 DVSS.n2873 5.2005
R21178 DVSS.n2882 DVSS.n2881 5.2005
R21179 DVSS.n2890 DVSS.n2889 5.2005
R21180 DVSS.n2898 DVSS.n2897 5.2005
R21181 DVSS.n2906 DVSS.n2905 5.2005
R21182 DVSS.n2914 DVSS.n2913 5.2005
R21183 DVSS.n2921 DVSS.n2920 5.2005
R21184 DVSS.n2928 DVSS.n2927 5.2005
R21185 DVSS.n2936 DVSS.n2935 5.2005
R21186 DVSS.n2944 DVSS.n2943 5.2005
R21187 DVSS.n2952 DVSS.n2951 5.2005
R21188 DVSS.n2960 DVSS.n2959 5.2005
R21189 DVSS.n2968 DVSS.n2967 5.2005
R21190 DVSS.n2976 DVSS.n2975 5.2005
R21191 DVSS.n2983 DVSS.n2982 5.2005
R21192 DVSS.n2990 DVSS.n2989 5.2005
R21193 DVSS.n2998 DVSS.n2997 5.2005
R21194 DVSS.n3006 DVSS.n3005 5.2005
R21195 DVSS.n2849 DVSS.n2848 5.2005
R21196 DVSS.n2847 DVSS.n2846 5.2005
R21197 DVSS.n3191 DVSS.n3190 5.2005
R21198 DVSS.n3199 DVSS.n3198 5.2005
R21199 DVSS.n3206 DVSS.n3205 5.2005
R21200 DVSS.n3213 DVSS.n3212 5.2005
R21201 DVSS.n3221 DVSS.n3220 5.2005
R21202 DVSS.n3229 DVSS.n3228 5.2005
R21203 DVSS.n3237 DVSS.n3236 5.2005
R21204 DVSS.n3245 DVSS.n3244 5.2005
R21205 DVSS.n3253 DVSS.n3252 5.2005
R21206 DVSS.n3261 DVSS.n3260 5.2005
R21207 DVSS.n3268 DVSS.n3267 5.2005
R21208 DVSS.n3275 DVSS.n3274 5.2005
R21209 DVSS.n3283 DVSS.n3282 5.2005
R21210 DVSS.n3291 DVSS.n3290 5.2005
R21211 DVSS.n3176 DVSS.n3175 5.2005
R21212 DVSS.n3174 DVSS.n3173 5.2005
R21213 DVSS.n3167 DVSS.n3166 5.2005
R21214 DVSS.n3159 DVSS.n3158 5.2005
R21215 DVSS.n3151 DVSS.n3150 5.2005
R21216 DVSS.n3144 DVSS.n3143 5.2005
R21217 DVSS.n3137 DVSS.n3136 5.2005
R21218 DVSS.n3129 DVSS.n3128 5.2005
R21219 DVSS.n2777 DVSS.n2776 5.2005
R21220 DVSS.n2768 DVSS.n2767 5.2005
R21221 DVSS.n2760 DVSS.n2759 5.2005
R21222 DVSS.n3380 DVSS.n3379 5.2005
R21223 DVSS.n3425 DVSS.n3424 5.2005
R21224 DVSS.n925 DVSS.n919 5.2005
R21225 DVSS.n3423 DVSS.n3422 5.2005
R21226 DVSS.n3419 DVSS.n3418 5.2005
R21227 DVSS.n3415 DVSS.n3414 5.2005
R21228 DVSS.n3412 DVSS.n3396 5.2005
R21229 DVSS.n3396 DVSS.n3395 5.2005
R21230 DVSS.n12811 DVSS.n12810 5.2005
R21231 DVSS.n12807 DVSS.n12806 5.2005
R21232 DVSS.n12803 DVSS.n12802 5.2005
R21233 DVSS.n12800 DVSS.n12794 5.2005
R21234 DVSS.n12794 DVSS.n12793 5.2005
R21235 DVSS.n12785 DVSS.n12784 5.2005
R21236 DVSS.n3400 DVSS.n3399 5.2005
R21237 DVSS.n21155 DVSS.n21154 5.2005
R21238 DVSS.n7438 DVSS.n7437 5.2005
R21239 DVSS.n7443 DVSS.n7442 5.2005
R21240 DVSS.n7448 DVSS.n7447 5.2005
R21241 DVSS.n18568 DVSS.n18567 5.2005
R21242 DVSS.n18563 DVSS.n18562 5.2005
R21243 DVSS.n7450 DVSS.n7449 5.2005
R21244 DVSS.n14888 DVSS.n14887 5.2005
R21245 DVSS.n14914 DVSS.n14913 5.2005
R21246 DVSS.n14922 DVSS.n14921 5.2005
R21247 DVSS.n14927 DVSS.n14926 5.2005
R21248 DVSS.n14931 DVSS.n14930 5.2005
R21249 DVSS.n14936 DVSS.n14935 5.2005
R21250 DVSS.n14941 DVSS.n14940 5.2005
R21251 DVSS.n14949 DVSS.n14948 5.2005
R21252 DVSS.n8010 DVSS.n8009 5.2005
R21253 DVSS.n8015 DVSS.n8014 5.2005
R21254 DVSS.n8020 DVSS.n8019 5.2005
R21255 DVSS.n13176 DVSS.n13175 5.2005
R21256 DVSS.n13171 DVSS.n13170 5.2005
R21257 DVSS.n13167 DVSS.n13166 5.2005
R21258 DVSS.n13162 DVSS.n13161 5.2005
R21259 DVSS.n13157 DVSS.n13156 5.2005
R21260 DVSS.n8048 DVSS.n8047 5.2005
R21261 DVSS.n8043 DVSS.n8042 5.2005
R21262 DVSS.n8038 DVSS.n8037 5.2005
R21263 DVSS.n1376 DVSS.n1375 5.2005
R21264 DVSS.n6904 DVSS.n6903 5.2005
R21265 DVSS.n6909 DVSS.n6908 5.2005
R21266 DVSS.n6914 DVSS.n6913 5.2005
R21267 DVSS.n6919 DVSS.n6918 5.2005
R21268 DVSS.n6924 DVSS.n6923 5.2005
R21269 DVSS.n6928 DVSS.n6927 5.2005
R21270 DVSS.n6933 DVSS.n6932 5.2005
R21271 DVSS.n6938 DVSS.n6937 5.2005
R21272 DVSS.n6943 DVSS.n6942 5.2005
R21273 DVSS.n6947 DVSS.n6946 5.2005
R21274 DVSS.n1356 DVSS.n1355 5.2005
R21275 DVSS.n1361 DVSS.n1360 5.2005
R21276 DVSS.n1364 DVSS.n1363 5.2005
R21277 DVSS.n354 DVSS.n353 5.11349
R21278 DVSS.n354 DVSS.n347 5.07814
R21279 DVSS.n1495 DVSS.n1492 4.83394
R21280 DVSS.n1498 DVSS.n1495 4.83394
R21281 DVSS.n1837 DVSS.n1835 4.83394
R21282 DVSS.n1841 DVSS.n1837 4.83394
R21283 DVSS.n6415 DVSS.n6414 4.5005
R21284 DVSS.n6410 DVSS.n6409 4.5005
R21285 DVSS.n4477 DVSS.n4476 4.5005
R21286 DVSS.n4472 DVSS.n4471 4.5005
R21287 DVSS.n6551 DVSS.n6550 4.5005
R21288 DVSS.n6546 DVSS.n6545 4.5005
R21289 DVSS.n6541 DVSS.n6540 4.5005
R21290 DVSS.n6536 DVSS.n2545 4.5005
R21291 DVSS.n4362 DVSS.n4361 4.5005
R21292 DVSS.n4367 DVSS.n4366 4.5005
R21293 DVSS.n4372 DVSS.n4371 4.5005
R21294 DVSS.n4376 DVSS.n4375 4.5005
R21295 DVSS.n4110 DVSS.n4109 4.5005
R21296 DVSS.n4105 DVSS.n4104 4.5005
R21297 DVSS.n4100 DVSS.n4099 4.5005
R21298 DVSS.n4095 DVSS.n2573 4.5005
R21299 DVSS.n6502 DVSS.n6486 4.5005
R21300 DVSS.n5608 DVSS.n5604 4.5005
R21301 DVSS.n5585 DVSS.n5584 4.5005
R21302 DVSS.n5600 DVSS.n5599 4.5005
R21303 DVSS.n5576 DVSS.n5575 4.5005
R21304 DVSS.n5581 DVSS.n5580 4.5005
R21305 DVSS.n5810 DVSS.n5809 4.5005
R21306 DVSS.n5806 DVSS.n5805 4.5005
R21307 DVSS.n5816 DVSS.n5815 4.5005
R21308 DVSS.n5821 DVSS.n5820 4.5005
R21309 DVSS.n6499 DVSS.n6488 4.5005
R21310 DVSS.n6496 DVSS.n6490 4.5005
R21311 DVSS.n6493 DVSS.n6492 4.5005
R21312 DVSS.n9787 DVSS.n8942 4.5005
R21313 DVSS.n9784 DVSS.n8944 4.5005
R21314 DVSS.n9781 DVSS.n8946 4.5005
R21315 DVSS.n8950 DVSS.n8947 4.5005
R21316 DVSS.n9734 DVSS.n9733 4.5005
R21317 DVSS.n9739 DVSS.n9738 4.5005
R21318 DVSS.n9750 DVSS.n9743 4.5005
R21319 DVSS.n9747 DVSS.n9744 4.5005
R21320 DVSS.n9595 DVSS.n8975 4.5005
R21321 DVSS.n9592 DVSS.n8977 4.5005
R21322 DVSS.n9589 DVSS.n8979 4.5005
R21323 DVSS.n8983 DVSS.n8980 4.5005
R21324 DVSS.n9122 DVSS.n9121 4.5005
R21325 DVSS.n9127 DVSS.n9126 4.5005
R21326 DVSS.n9138 DVSS.n9131 4.5005
R21327 DVSS.n9135 DVSS.n9132 4.5005
R21328 DVSS.n11206 DVSS.n11175 4.5005
R21329 DVSS.n11170 DVSS.n11169 4.5005
R21330 DVSS.n11214 DVSS.n11213 4.5005
R21331 DVSS.n11209 DVSS.n11174 4.5005
R21332 DVSS.n11039 DVSS.n11038 4.5005
R21333 DVSS.n11044 DVSS.n11043 4.5005
R21334 DVSS.n11052 DVSS.n11051 4.5005
R21335 DVSS.n10269 DVSS.n10268 4.5005
R21336 DVSS.n10250 DVSS.n10248 4.5005
R21337 DVSS.n10256 DVSS.n10255 4.5005
R21338 DVSS.n10283 DVSS.n10280 4.5005
R21339 DVSS.n10291 DVSS.n10287 4.5005
R21340 DVSS.n11034 DVSS.n11033 4.5005
R21341 DVSS.n16276 DVSS.n16275 4.5005
R21342 DVSS.n17943 DVSS.n7624 4.5005
R21343 DVSS.n17940 DVSS.n7625 4.5005
R21344 DVSS.n16237 DVSS.n16236 4.5005
R21345 DVSS.n18084 DVSS.n7616 4.5005
R21346 DVSS.n18081 DVSS.n7617 4.5005
R21347 DVSS.n18366 DVSS.n7564 4.5005
R21348 DVSS.n18363 DVSS.n7610 4.5005
R21349 DVSS.n18360 DVSS.n7611 4.5005
R21350 DVSS.n18406 DVSS.n18405 4.5005
R21351 DVSS.n18415 DVSS.n18410 4.5005
R21352 DVSS.n18412 DVSS.n18411 4.5005
R21353 DVSS.n16336 DVSS.n16335 4.5005
R21354 DVSS.n7634 DVSS.n7629 4.5005
R21355 DVSS.n7631 DVSS.n7630 4.5005
R21356 DVSS.n17459 DVSS.n17458 4.5005
R21357 DVSS.n17298 DVSS.n17280 4.5005
R21358 DVSS.n17294 DVSS.n17282 4.5005
R21359 DVSS.n17291 DVSS.n17284 4.5005
R21360 DVSS.n17287 DVSS.n17286 4.5005
R21361 DVSS.n17463 DVSS.n17462 4.5005
R21362 DVSS.n17455 DVSS.n17454 4.5005
R21363 DVSS.n15837 DVSS.n15836 4.5005
R21364 DVSS.n15842 DVSS.n15841 4.5005
R21365 DVSS.n15853 DVSS.n15846 4.5005
R21366 DVSS.n15850 DVSS.n15847 4.5005
R21367 DVSS.n15727 DVSS.n7683 4.5005
R21368 DVSS.n15724 DVSS.n7685 4.5005
R21369 DVSS.n15721 DVSS.n7687 4.5005
R21370 DVSS.n7691 DVSS.n7688 4.5005
R21371 DVSS.n15591 DVSS.n15590 4.5005
R21372 DVSS.n15596 DVSS.n15595 4.5005
R21373 DVSS.n15607 DVSS.n15600 4.5005
R21374 DVSS.n15604 DVSS.n15601 4.5005
R21375 DVSS.n14962 DVSS.n14961 4.5005
R21376 DVSS.n14967 DVSS.n14966 4.5005
R21377 DVSS.n14978 DVSS.n14971 4.5005
R21378 DVSS.n14975 DVSS.n14972 4.5005
R21379 DVSS.n17644 DVSS.n17641 4.5005
R21380 DVSS.n17659 DVSS.n17658 4.5005
R21381 DVSS.n17654 DVSS.n7657 4.5005
R21382 DVSS.n7662 DVSS.n7659 4.5005
R21383 DVSS.n16892 DVSS.n16891 4.5005
R21384 DVSS.n16897 DVSS.n16896 4.5005
R21385 DVSS.n16902 DVSS.n16901 4.5005
R21386 DVSS.n17552 DVSS.n17551 4.5005
R21387 DVSS.n17008 DVSS.n17007 4.5005
R21388 DVSS.n16998 DVSS.n16996 4.5005
R21389 DVSS.n17004 DVSS.n17003 4.5005
R21390 DVSS.n17022 DVSS.n17019 4.5005
R21391 DVSS.n17030 DVSS.n17026 4.5005
R21392 DVSS.n7668 DVSS.n7667 4.5005
R21393 DVSS.n15828 DVSS.n7672 4.5005
R21394 DVSS.n15832 DVSS.n15831 4.5005
R21395 DVSS.n7676 DVSS.n7675 4.5005
R21396 DVSS.n15733 DVSS.n7680 4.5005
R21397 DVSS.n15730 DVSS.n7681 4.5005
R21398 DVSS.n7697 DVSS.n7696 4.5005
R21399 DVSS.n15582 DVSS.n7701 4.5005
R21400 DVSS.n15586 DVSS.n15585 4.5005
R21401 DVSS.n15249 DVSS.n7706 4.5005
R21402 DVSS.n15246 DVSS.n7708 4.5005
R21403 DVSS.n14957 DVSS.n14956 4.5005
R21404 DVSS.n17663 DVSS.n17662 4.5005
R21405 DVSS.n17675 DVSS.n17674 4.5005
R21406 DVSS.n17545 DVSS.n17544 4.5005
R21407 DVSS.n17541 DVSS.n17540 4.5005
R21408 DVSS.n17536 DVSS.n17535 4.5005
R21409 DVSS.n16990 DVSS.n16989 4.5005
R21410 DVSS.n16974 DVSS.n16973 4.5005
R21411 DVSS.n16980 DVSS.n16979 4.5005
R21412 DVSS.n16985 DVSS.n16984 4.5005
R21413 DVSS.n7651 DVSS.n7648 4.5005
R21414 DVSS.n8031 DVSS.n8030 4.5005
R21415 DVSS.n11480 DVSS.n11477 4.5005
R21416 DVSS.n11480 DVSS.n11467 4.5005
R21417 DVSS.n11461 DVSS.n11460 4.5005
R21418 DVSS.n11465 DVSS.n11464 4.5005
R21419 DVSS.n11480 DVSS.n11478 4.5005
R21420 DVSS.n11480 DVSS.n11466 4.5005
R21421 DVSS.n11480 DVSS.n11479 4.5005
R21422 DVSS.n11517 DVSS.n11514 4.5005
R21423 DVSS.n11517 DVSS.n11504 4.5005
R21424 DVSS.n11498 DVSS.n11497 4.5005
R21425 DVSS.n11502 DVSS.n11501 4.5005
R21426 DVSS.n11517 DVSS.n11515 4.5005
R21427 DVSS.n11517 DVSS.n11503 4.5005
R21428 DVSS.n11517 DVSS.n11516 4.5005
R21429 DVSS.n11642 DVSS.n11639 4.5005
R21430 DVSS.n11642 DVSS.n11629 4.5005
R21431 DVSS.n11623 DVSS.n11622 4.5005
R21432 DVSS.n11627 DVSS.n11626 4.5005
R21433 DVSS.n11642 DVSS.n11640 4.5005
R21434 DVSS.n11642 DVSS.n11628 4.5005
R21435 DVSS.n11642 DVSS.n11641 4.5005
R21436 DVSS.n11679 DVSS.n11676 4.5005
R21437 DVSS.n11679 DVSS.n11666 4.5005
R21438 DVSS.n11660 DVSS.n11659 4.5005
R21439 DVSS.n11664 DVSS.n11663 4.5005
R21440 DVSS.n11679 DVSS.n11677 4.5005
R21441 DVSS.n11679 DVSS.n11665 4.5005
R21442 DVSS.n11679 DVSS.n11678 4.5005
R21443 DVSS.n8031 DVSS.n8022 4.5005
R21444 DVSS.n8031 DVSS.n8021 4.5005
R21445 DVSS.n11189 DVSS.n11186 4.5005
R21446 DVSS.n11189 DVSS.n11177 4.5005
R21447 DVSS.n11201 DVSS.n11200 4.5005
R21448 DVSS.n11019 DVSS.n11016 4.5005
R21449 DVSS.n11019 DVSS.n11007 4.5005
R21450 DVSS.n10263 DVSS.n10259 4.5005
R21451 DVSS.n10627 DVSS.n10625 4.5005
R21452 DVSS.n10627 DVSS.n10619 4.5005
R21453 DVSS.n10627 DVSS.n10626 4.5005
R21454 DVSS.n10640 DVSS.n10639 4.5005
R21455 DVSS.n11019 DVSS.n11017 4.5005
R21456 DVSS.n11028 DVSS.n11004 4.5005
R21457 DVSS.n11024 DVSS.n11005 4.5005
R21458 DVSS.n11019 DVSS.n11006 4.5005
R21459 DVSS.n11019 DVSS.n11018 4.5005
R21460 DVSS.n11189 DVSS.n11187 4.5005
R21461 DVSS.n11195 DVSS.n11194 4.5005
R21462 DVSS.n11189 DVSS.n11176 4.5005
R21463 DVSS.n11189 DVSS.n11188 4.5005
R21464 DVSS.n11728 DVSS.n11725 4.5005
R21465 DVSS.n11728 DVSS.n11715 4.5005
R21466 DVSS.n4018 DVSS.n4017 4.5005
R21467 DVSS.n4023 DVSS.n4022 4.5005
R21468 DVSS.n4032 DVSS.n4027 4.5005
R21469 DVSS.n4029 DVSS.n4028 4.5005
R21470 DVSS.n7488 DVSS.n7485 4.5005
R21471 DVSS.n7458 DVSS.n7453 4.5005
R21472 DVSS.n7455 DVSS.n7454 4.5005
R21473 DVSS.n15060 DVSS.n7726 4.5005
R21474 DVSS.n15057 DVSS.n7767 4.5005
R21475 DVSS.n15054 DVSS.n7769 4.5005
R21476 DVSS.n15051 DVSS.n7770 4.5005
R21477 DVSS.n15048 DVSS.n7772 4.5005
R21478 DVSS.n15045 DVSS.n7774 4.5005
R21479 DVSS.n7781 DVSS.n7776 4.5005
R21480 DVSS.n9030 DVSS.n9022 4.5005
R21481 DVSS.n9027 DVSS.n9024 4.5005
R21482 DVSS.n8059 DVSS.n8051 4.5005
R21483 DVSS.n8056 DVSS.n8053 4.5005
R21484 DVSS.n11709 DVSS.n11708 4.5005
R21485 DVSS.n11728 DVSS.n11726 4.5005
R21486 DVSS.n11728 DVSS.n11714 4.5005
R21487 DVSS.n11728 DVSS.n11727 4.5005
R21488 DVSS.n5546 DVSS.n5540 4.5005
R21489 DVSS.n5549 DVSS.n5538 4.5005
R21490 DVSS.n5553 DVSS.n5552 4.5005
R21491 DVSS.n5543 DVSS.n5542 4.5005
R21492 DVSS.n10039 DVSS.n10011 4.5005
R21493 DVSS.n10045 DVSS.n10009 4.5005
R21494 DVSS.n10050 DVSS.n10049 4.5005
R21495 DVSS.n10053 DVSS.n10008 4.5005
R21496 DVSS.n10004 DVSS.n10003 4.5005
R21497 DVSS.n16881 DVSS.n16878 4.5005
R21498 DVSS.n16886 DVSS.n16885 4.5005
R21499 DVSS.n17102 DVSS.n16877 4.5005
R21500 DVSS.n17105 DVSS.n16875 4.5005
R21501 DVSS.n17108 DVSS.n16874 4.5005
R21502 DVSS.n17113 DVSS.n17112 4.5005
R21503 DVSS.n16870 DVSS.n16869 4.5005
R21504 DVSS.n17244 DVSS.n16443 4.5005
R21505 DVSS.n17236 DVSS.n16444 4.5005
R21506 DVSS.n17241 DVSS.n17240 4.5005
R21507 DVSS.n10029 DVSS.n10026 4.5005
R21508 DVSS.n10029 DVSS.n10013 4.5005
R21509 DVSS.n10029 DVSS.n10027 4.5005
R21510 DVSS.n10029 DVSS.n10012 4.5005
R21511 DVSS.n10029 DVSS.n10028 4.5005
R21512 DVSS.n10035 DVSS.n10034 4.5005
R21513 DVSS.n5534 DVSS.n5533 4.5005
R21514 DVSS.n5530 DVSS.n5529 4.5005
R21515 DVSS.n5525 DVSS.n5524 4.5005
R21516 DVSS.n5520 DVSS.n5519 4.5005
R21517 DVSS.n5383 DVSS.n5354 4.5005
R21518 DVSS.n5378 DVSS.n5356 4.5005
R21519 DVSS.n5374 DVSS.n5358 4.5005
R21520 DVSS.n5370 DVSS.n5360 4.5005
R21521 DVSS.n5365 DVSS.n5361 4.5005
R21522 DVSS.n6430 DVSS.n6404 4.5005
R21523 DVSS.n6418 DVSS.n6405 4.5005
R21524 DVSS.n6566 DVSS.n2543 4.5005
R21525 DVSS.n6554 DVSS.n2544 4.5005
R21526 DVSS.n6483 DVSS.n6482 4.5005
R21527 DVSS.n6479 DVSS.n6478 4.5005
R21528 DVSS.n5825 DVSS.n5824 4.5005
R21529 DVSS.n5830 DVSS.n5829 4.5005
R21530 DVSS.n2549 DVSS.n2548 4.5005
R21531 DVSS.n2554 DVSS.n2553 4.5005
R21532 DVSS.n4353 DVSS.n2558 4.5005
R21533 DVSS.n4357 DVSS.n4356 4.5005
R21534 DVSS.n2562 DVSS.n2561 4.5005
R21535 DVSS.n2567 DVSS.n2566 4.5005
R21536 DVSS.n4116 DVSS.n2571 4.5005
R21537 DVSS.n4113 DVSS.n2572 4.5005
R21538 DVSS.n2577 DVSS.n2576 4.5005
R21539 DVSS.n4004 DVSS.n4003 4.5005
R21540 DVSS.n4009 DVSS.n4008 4.5005
R21541 DVSS.n4013 DVSS.n4012 4.5005
R21542 DVSS.n925 DVSS.n924 4.5005
R21543 DVSS.n3410 DVSS.n3403 4.5005
R21544 DVSS.n3410 DVSS.n3398 4.5005
R21545 DVSS.n12791 DVSS.n12788 4.5005
R21546 DVSS.n12791 DVSS.n12790 4.5005
R21547 DVSS.n8933 DVSS.n8932 4.5005
R21548 DVSS.n9796 DVSS.n8937 4.5005
R21549 DVSS.n9793 DVSS.n8939 4.5005
R21550 DVSS.n9790 DVSS.n8940 4.5005
R21551 DVSS.n8958 DVSS.n8957 4.5005
R21552 DVSS.n9720 DVSS.n9719 4.5005
R21553 DVSS.n9725 DVSS.n9724 4.5005
R21554 DVSS.n9729 DVSS.n9728 4.5005
R21555 DVSS.n8966 DVSS.n8965 4.5005
R21556 DVSS.n9604 DVSS.n8970 4.5005
R21557 DVSS.n9601 DVSS.n8972 4.5005
R21558 DVSS.n9598 DVSS.n8973 4.5005
R21559 DVSS.n9008 DVSS.n9007 4.5005
R21560 DVSS.n9108 DVSS.n9107 4.5005
R21561 DVSS.n9113 DVSS.n9112 4.5005
R21562 DVSS.n9117 DVSS.n9116 4.5005
R21563 DVSS.n9013 DVSS.n9012 4.5005
R21564 DVSS.n9039 DVSS.n9017 4.5005
R21565 DVSS.n9036 DVSS.n9019 4.5005
R21566 DVSS.n9033 DVSS.n9021 4.5005
R21567 DVSS.n11165 DVSS.n8927 4.5005
R21568 DVSS.n9819 DVSS.n9818 4.5005
R21569 DVSS.n9831 DVSS.n9823 4.5005
R21570 DVSS.n9828 DVSS.n9825 4.5005
R21571 DVSS.n11056 DVSS.n11055 4.5005
R21572 DVSS.n11061 DVSS.n11060 4.5005
R21573 DVSS.n11066 DVSS.n11065 4.5005
R21574 DVSS.n11075 DVSS.n11074 4.5005
R21575 DVSS.n10000 DVSS.n9999 4.5005
R21576 DVSS.n9996 DVSS.n9995 4.5005
R21577 DVSS.n9991 DVSS.n9860 4.5005
R21578 DVSS.n9856 DVSS.n9855 4.5005
R21579 DVSS.n10242 DVSS.n10241 4.5005
R21580 DVSS.n10217 DVSS.n10216 4.5005
R21581 DVSS.n10224 DVSS.n10223 4.5005
R21582 DVSS.n10230 DVSS.n10229 4.5005
R21583 DVSS.n10236 DVSS.n10235 4.5005
R21584 DVSS.n16266 DVSS.n16265 4.5005
R21585 DVSS.n16285 DVSS.n16270 4.5005
R21586 DVSS.n16282 DVSS.n16272 4.5005
R21587 DVSS.n16279 DVSS.n16273 4.5005
R21588 DVSS.n16227 DVSS.n16226 4.5005
R21589 DVSS.n16246 DVSS.n16231 4.5005
R21590 DVSS.n16243 DVSS.n16233 4.5005
R21591 DVSS.n16240 DVSS.n16234 4.5005
R21592 DVSS.n7555 DVSS.n7554 4.5005
R21593 DVSS.n18375 DVSS.n7559 4.5005
R21594 DVSS.n18372 DVSS.n7561 4.5005
R21595 DVSS.n18369 DVSS.n7562 4.5005
R21596 DVSS.n7466 DVSS.n7465 4.5005
R21597 DVSS.n18392 DVSS.n18391 4.5005
R21598 DVSS.n18397 DVSS.n18396 4.5005
R21599 DVSS.n18401 DVSS.n18400 4.5005
R21600 DVSS.n7476 DVSS.n7475 4.5005
R21601 DVSS.n7497 DVSS.n7480 4.5005
R21602 DVSS.n7494 DVSS.n7482 4.5005
R21603 DVSS.n7491 DVSS.n7483 4.5005
R21604 DVSS.n16430 DVSS.n16429 4.5005
R21605 DVSS.n16435 DVSS.n16434 4.5005
R21606 DVSS.n17248 DVSS.n17247 4.5005
R21607 DVSS.n16440 DVSS.n16439 4.5005
R21608 DVSS.n17303 DVSS.n17278 4.5005
R21609 DVSS.n17274 DVSS.n17272 4.5005
R21610 DVSS.n17327 DVSS.n17326 4.5005
R21611 DVSS.n17270 DVSS.n17269 4.5005
R21612 DVSS.n17318 DVSS.n17317 4.5005
R21613 DVSS.n17449 DVSS.n16127 4.5005
R21614 DVSS.n16124 DVSS.n16123 4.5005
R21615 DVSS.n17445 DVSS.n17442 4.5005
R21616 DVSS.n17438 DVSS.n17437 4.5005
R21617 DVSS.n16340 DVSS.n16339 4.5005
R21618 DVSS.n16310 DVSS.n16309 4.5005
R21619 DVSS.n16322 DVSS.n16321 4.5005
R21620 DVSS.n16317 DVSS.n16316 4.5005
R21621 DVSS.n7436 DVSS.n7435 4.5005
R21622 DVSS.n7441 DVSS.n7440 4.5005
R21623 DVSS.n7446 DVSS.n7445 4.5005
R21624 DVSS.n18571 DVSS.n18570 4.5005
R21625 DVSS.n18566 DVSS.n18565 4.5005
R21626 DVSS.n18561 DVSS.n18560 4.5005
R21627 DVSS.n14886 DVSS.n14885 4.5005
R21628 DVSS.n14910 DVSS.n14909 4.5005
R21629 DVSS.n14920 DVSS.n14919 4.5005
R21630 DVSS.n14925 DVSS.n14924 4.5005
R21631 DVSS.n14929 DVSS.n14928 4.5005
R21632 DVSS.n14934 DVSS.n14933 4.5005
R21633 DVSS.n14939 DVSS.n14938 4.5005
R21634 DVSS.n14952 DVSS.n14951 4.5005
R21635 DVSS.n14947 DVSS.n14946 4.5005
R21636 DVSS.n8008 DVSS.n8007 4.5005
R21637 DVSS.n8013 DVSS.n8012 4.5005
R21638 DVSS.n8018 DVSS.n8017 4.5005
R21639 DVSS.n13179 DVSS.n13178 4.5005
R21640 DVSS.n13174 DVSS.n13173 4.5005
R21641 DVSS.n13169 DVSS.n13168 4.5005
R21642 DVSS.n13165 DVSS.n13164 4.5005
R21643 DVSS.n13160 DVSS.n13159 4.5005
R21644 DVSS.n13155 DVSS.n13154 4.5005
R21645 DVSS.n8046 DVSS.n8045 4.5005
R21646 DVSS.n8040 DVSS.n8039 4.5005
R21647 DVSS.n6907 DVSS.n6906 4.5005
R21648 DVSS.n6912 DVSS.n6911 4.5005
R21649 DVSS.n6917 DVSS.n6916 4.5005
R21650 DVSS.n6922 DVSS.n6921 4.5005
R21651 DVSS.n6926 DVSS.n6925 4.5005
R21652 DVSS.n6931 DVSS.n6930 4.5005
R21653 DVSS.n6936 DVSS.n6935 4.5005
R21654 DVSS.n6941 DVSS.n6940 4.5005
R21655 DVSS.n6950 DVSS.n6949 4.5005
R21656 DVSS.n6945 DVSS.n6944 4.5005
R21657 DVSS.n6901 DVSS.n1377 4.5005
R21658 DVSS.n6435 DVSS.n6434 4.5005
R21659 DVSS.n6571 DVSS.n6570 4.5005
R21660 DVSS.n6714 DVSS.n6713 4.5005
R21661 DVSS.n6769 DVSS.n6768 4.5005
R21662 DVSS.n6896 DVSS.n6895 4.5005
R21663 DVSS.n5512 DVSS.n5511 4.5005
R21664 DVSS.n5388 DVSS.n5352 4.5005
R21665 DVSS.n5835 DVSS.n4581 4.5005
R21666 DVSS.n6472 DVSS.n4527 4.5005
R21667 DVSS.n2482 DVSS.n2480 4.06502
R21668 DVSS.n2482 DVSS.n2481 4.06502
R21669 DVSS.n2505 DVSS.n2503 4.06502
R21670 DVSS.n2505 DVSS.n2504 4.06502
R21671 DVSS.n2470 DVSS.n1743 4.06502
R21672 DVSS.n2470 DVSS.n1744 4.06502
R21673 DVSS.n2479 DVSS.n2477 4.06502
R21674 DVSS.n2479 DVSS.n2478 4.06502
R21675 DVSS.n2502 DVSS.n2500 4.06502
R21676 DVSS.n2502 DVSS.n2501 4.06502
R21677 DVSS.n1741 DVSS.n1403 4.06502
R21678 DVSS.n1741 DVSS.n1404 4.06502
R21679 DVSS.n7158 DVSS.n7157 3.71156
R21680 DVSS.n7968 DVSS.n7967 3.71156
R21681 DVSS.n7026 DVSS.n7025 3.71156
R21682 DVSS.n13323 DVSS.n13322 3.71156
R21683 DVSS.n14906 DVSS.n14891 3.62347
R21684 DVSS.n21148 DVSS.n21147 3.58891
R21685 DVSS DVSS.t31 3.33845
R21686 DVSS DVSS.t24 3.33845
R21687 DVSS DVSS.t20 3.33845
R21688 DVSS DVSS.t18 3.33845
R21689 DVSS DVSS.t0 3.33845
R21690 DVSS DVSS.t27 3.33845
R21691 DVSS DVSS.t26 3.33845
R21692 DVSS DVSS.t19 3.33845
R21693 DVSS DVSS.t8 3.33845
R21694 DVSS DVSS.t2 3.33845
R21695 DVSS DVSS.t7 3.33845
R21696 DVSS DVSS.t33 3.33845
R21697 DVSS DVSS.t22 3.33845
R21698 DVSS DVSS.t11 3.33845
R21699 DVSS DVSS.t5 3.33845
R21700 DVSS DVSS.t36 3.33845
R21701 DVSS DVSS.t29 3.33845
R21702 DVSS DVSS.t32 3.33845
R21703 DVSS.n7432 DVSS.t25 3.2597
R21704 DVSS.n7432 DVSS.t32 3.2597
R21705 DVSS.n17432 DVSS.t23 3.2597
R21706 DVSS.n17432 DVSS.t31 3.2597
R21707 DVSS.n16889 DVSS.t24 3.2597
R21708 DVSS.n16889 DVSS.t10 3.2597
R21709 DVSS.n7460 DVSS.t17 3.2597
R21710 DVSS.n7460 DVSS.t20 3.2597
R21711 DVSS.n14973 DVSS.t18 3.2597
R21712 DVSS.n14973 DVSS.t34 3.2597
R21713 DVSS.n7549 DVSS.t30 3.2597
R21714 DVSS.n7549 DVSS.t0 3.2597
R21715 DVSS.n15602 DVSS.t27 3.2597
R21716 DVSS.n15602 DVSS.t12 3.2597
R21717 DVSS.n16221 DVSS.t21 3.2597
R21718 DVSS.n16221 DVSS.t26 3.2597
R21719 DVSS.n7689 DVSS.t19 3.2597
R21720 DVSS.n7689 DVSS.t6 3.2597
R21721 DVSS.n16305 DVSS.t1 3.2597
R21722 DVSS.n16305 DVSS.t8 3.2597
R21723 DVSS.n17642 DVSS.t2 3.2597
R21724 DVSS.n17642 DVSS.t15 3.2597
R21725 DVSS.n16260 DVSS.t35 3.2597
R21726 DVSS.n16260 DVSS.t7 3.2597
R21727 DVSS.n15848 DVSS.t33 3.2597
R21728 DVSS.n15848 DVSS.t14 3.2597
R21729 DVSS.n14942 DVSS.t22 3.2597
R21730 DVSS.n14942 DVSS.t9 3.2597
R21731 DVSS.n7470 DVSS.t4 3.2597
R21732 DVSS.n7470 DVSS.t11 3.2597
R21733 DVSS.n7777 DVSS.t5 3.2597
R21734 DVSS.n7777 DVSS.t16 3.2597
R21735 DVSS.n16425 DVSS.t28 3.2597
R21736 DVSS.n16425 DVSS.t36 3.2597
R21737 DVSS.n16879 DVSS.t29 3.2597
R21738 DVSS.n16879 DVSS.t13 3.2597
R21739 DVSS.n16800 DVSS.n16799 3.1505
R21740 DVSS.n15115 DVSS.n15114 3.1505
R21741 DVSS.n7638 DVSS.n7637 3.1505
R21742 DVSS.n16012 DVSS.n16007 3.1505
R21743 DVSS.n15309 DVSS.n15304 3.1505
R21744 DVSS.n18298 DVSS.n18297 3.1505
R21745 DVSS.n18011 DVSS.n18006 3.1505
R21746 DVSS.n17870 DVSS.n17865 3.1505
R21747 DVSS.n13916 DVSS.n13915 3.1505
R21748 DVSS.n18353 DVSS.n18352 3.14853
R21749 DVSS.n15072 DVSS.n15071 3.14797
R21750 DVSS.n13969 DVSS.n13968 3.14797
R21751 DVSS.n14908 DVSS.n14907 3.14395
R21752 DVSS.n21148 DVSS.n21146 3.10592
R21753 DVSS.n915 DVSS.n913 2.91885
R21754 DVSS.n918 DVSS.n916 2.91885
R21755 DVSS.n21158 DVSS.n21156 2.91885
R21756 DVSS.n21151 DVSS.n21149 2.73983
R21757 DVSS.n14890 DVSS.n14889 2.72092
R21758 DVSS.n7387 DVSS.n7386 2.61893
R21759 DVSS.n13770 DVSS.n13769 2.61893
R21760 DVSS.n1325 DVSS.n1319 2.61893
R21761 DVSS.n13338 DVSS.n13332 2.61893
R21762 DVSS.n13809 DVSS.n13808 2.6005
R21763 DVSS.n7790 DVSS.n7789 2.6005
R21764 DVSS.n7785 DVSS.n7784 2.6005
R21765 DVSS.n7798 DVSS.n7797 2.6005
R21766 DVSS.n7793 DVSS.n7792 2.6005
R21767 DVSS.n13837 DVSS.n13836 2.6005
R21768 DVSS.n13988 DVSS.n13987 2.6005
R21769 DVSS.n13985 DVSS.n13984 2.6005
R21770 DVSS.n13982 DVSS.n13981 2.6005
R21771 DVSS.n14234 DVSS.n14233 2.6005
R21772 DVSS.n14229 DVSS.n14228 2.6005
R21773 DVSS.n14211 DVSS.n14210 2.6005
R21774 DVSS.n18587 DVSS.n18586 2.6005
R21775 DVSS.n7429 DVSS.n7428 2.6005
R21776 DVSS.n7426 DVSS.n7425 2.6005
R21777 DVSS.n18597 DVSS.n18596 2.6005
R21778 DVSS.n18594 DVSS.n18593 2.6005
R21779 DVSS.n7407 DVSS.n7406 2.6005
R21780 DVSS.n7384 DVSS.n7383 2.6005
R21781 DVSS.n13814 DVSS.n13813 2.6005
R21782 DVSS.n7412 DVSS.n7411 2.6005
R21783 DVSS.n13767 DVSS.n13766 2.6005
R21784 DVSS.n13722 DVSS.n13721 2.6005
R21785 DVSS.n13723 DVSS.n13722 2.6005
R21786 DVSS.n13774 DVSS.n13773 2.6005
R21787 DVSS.n7391 DVSS.n7390 2.6005
R21788 DVSS.n7352 DVSS.n7351 2.6005
R21789 DVSS.n7359 DVSS.n7358 2.6005
R21790 DVSS.n7358 DVSS.n7357 2.6005
R21791 DVSS.n13736 DVSS.n13735 2.6005
R21792 DVSS.n13735 DVSS.n13734 2.6005
R21793 DVSS.n7366 DVSS.n7365 2.6005
R21794 DVSS.n7365 DVSS.n7364 2.6005
R21795 DVSS.n13729 DVSS.n13728 2.6005
R21796 DVSS.n18697 DVSS.n18696 2.6005
R21797 DVSS.n18699 DVSS.n18698 2.6005
R21798 DVSS.n7338 DVSS.n7337 2.6005
R21799 DVSS.n7344 DVSS.n7343 2.6005
R21800 DVSS.n7340 DVSS.n7339 2.6005
R21801 DVSS.n14340 DVSS.n14339 2.6005
R21802 DVSS.n14327 DVSS.n14326 2.6005
R21803 DVSS.n14331 DVSS.n14330 2.6005
R21804 DVSS.n14801 DVSS.n14800 2.6005
R21805 DVSS.n7849 DVSS.n7848 2.6005
R21806 DVSS.n7837 DVSS.n7836 2.6005
R21807 DVSS.n14803 DVSS.n14802 2.6005
R21808 DVSS.n14043 DVSS.n14042 2.6005
R21809 DVSS.n13691 DVSS.n13690 2.6005
R21810 DVSS.n13693 DVSS.n13692 2.6005
R21811 DVSS.n7842 DVSS.n7841 2.6005
R21812 DVSS.n17939 DVSS.n17938 2.6005
R21813 DVSS.n18080 DVSS.n18079 2.6005
R21814 DVSS.n18359 DVSS.n18358 2.6005
R21815 DVSS.n15261 DVSS.n15260 2.6005
R21816 DVSS.n17532 DVSS.n17531 2.6005
R21817 DVSS.n17678 DVSS.n17677 2.6005
R21818 DVSS.n11507 DVSS.n11506 2.6005
R21819 DVSS.n11506 DVSS.n11505 2.6005
R21820 DVSS.n1746 DVSS.n1745 2.6005
R21821 DVSS.n355 DVSS.n354 2.6005
R21822 DVSS.n356 DVSS.n355 2.6005
R21823 DVSS.n12560 DVSS.n12559 2.6005
R21824 DVSS.n20396 DVSS.n20395 2.6005
R21825 DVSS.n20421 DVSS.n20420 2.6005
R21826 DVSS.n20437 DVSS.n20436 2.6005
R21827 DVSS.n20151 DVSS.n20150 2.6005
R21828 DVSS.n20173 DVSS.n20172 2.6005
R21829 DVSS.n19877 DVSS.n19876 2.6005
R21830 DVSS.n19898 DVSS.n19897 2.6005
R21831 DVSS.n19677 DVSS.n19676 2.6005
R21832 DVSS.n19661 DVSS.n19660 2.6005
R21833 DVSS.n19640 DVSS.n19639 2.6005
R21834 DVSS.n19388 DVSS.n19387 2.6005
R21835 DVSS.n19413 DVSS.n19412 2.6005
R21836 DVSS.n19429 DVSS.n19428 2.6005
R21837 DVSS.n19106 DVSS.n19105 2.6005
R21838 DVSS.n19165 DVSS.n19164 2.6005
R21839 DVSS.n19139 DVSS.n19138 2.6005
R21840 DVSS.n19113 DVSS.n19112 2.6005
R21841 DVSS.n19435 DVSS.n19434 2.6005
R21842 DVSS.n19378 DVSS.n19377 2.6005
R21843 DVSS.n19382 DVSS.n19381 2.6005
R21844 DVSS.n19870 DVSS.n19869 2.6005
R21845 DVSS.n20166 DVSS.n20165 2.6005
R21846 DVSS.n20138 DVSS.n20137 2.6005
R21847 DVSS.n20145 DVSS.n20144 2.6005
R21848 DVSS.n20443 DVSS.n20442 2.6005
R21849 DVSS.n20383 DVSS.n20382 2.6005
R21850 DVSS.n13334 DVSS.n13333 2.6005
R21851 DVSS.n1324 DVSS.n1323 2.6005
R21852 DVSS.n1321 DVSS.n1320 2.6005
R21853 DVSS.n7160 DVSS.n7159 2.6005
R21854 DVSS.n7970 DVSS.n7969 2.6005
R21855 DVSS.n13337 DVSS.n13336 2.6005
R21856 DVSS.n1331 DVSS.n1330 2.6005
R21857 DVSS.n1330 DVSS.n1329 2.6005
R21858 DVSS.n13344 DVSS.n13343 2.6005
R21859 DVSS.n13343 DVSS.n13342 2.6005
R21860 DVSS.n1317 DVSS.n1316 2.6005
R21861 DVSS.n1316 DVSS.n1315 2.6005
R21862 DVSS.n13292 DVSS.n13291 2.6005
R21863 DVSS.n13330 DVSS.n13329 2.6005
R21864 DVSS.n13329 DVSS.n13328 2.6005
R21865 DVSS.n7028 DVSS.n7027 2.6005
R21866 DVSS.n13325 DVSS.n13324 2.6005
R21867 DVSS.n7022 DVSS.n7021 2.6005
R21868 DVSS.n13675 DVSS.n13674 2.6005
R21869 DVSS.n7860 DVSS.n7859 2.6005
R21870 DVSS.n7852 DVSS.n7851 2.6005
R21871 DVSS.n13682 DVSS.n13681 2.6005
R21872 DVSS.n14053 DVSS.n14052 2.6005
R21873 DVSS.n14360 DVSS.n14359 2.6005
R21874 DVSS.n18713 DVSS.n18712 2.6005
R21875 DVSS.n18733 DVSS.n18732 2.6005
R21876 DVSS.n18730 DVSS.n18729 2.6005
R21877 DVSS.n18723 DVSS.n18722 2.6005
R21878 DVSS.n18720 DVSS.n18719 2.6005
R21879 DVSS.n7004 DVSS.n7003 2.6005
R21880 DVSS.n7007 DVSS.n7006 2.6005
R21881 DVSS.n7010 DVSS.n7009 2.6005
R21882 DVSS.n7013 DVSS.n7012 2.6005
R21883 DVSS.n7016 DVSS.n7015 2.6005
R21884 DVSS.n7862 DVSS.n7861 2.6005
R21885 DVSS.n7854 DVSS.n7853 2.6005
R21886 DVSS.n14057 DVSS.n14056 2.6005
R21887 DVSS.n14788 DVSS.n14787 2.6005
R21888 DVSS.n14362 DVSS.n14361 2.6005
R21889 DVSS.n14352 DVSS.n14351 2.6005
R21890 DVSS.n13196 DVSS.n13195 2.6005
R21891 DVSS.n13276 DVSS.n13275 2.6005
R21892 DVSS.n13280 DVSS.n13279 2.6005
R21893 DVSS.n13284 DVSS.n13283 2.6005
R21894 DVSS.n15064 DVSS.n15063 2.6005
R21895 DVSS.n2475 DVSS.n2474 2.6005
R21896 DVSS.n17235 DVSS.n17234 2.6005
R21897 DVSS.n3184 DVSS.n3183 2.6005
R21898 DVSS.n15063 DVSS.n15061 2.54004
R21899 DVSS.n15063 DVSS.n15062 2.54004
R21900 DVSS.n17234 DVSS.n17232 2.54004
R21901 DVSS.n17234 DVSS.n17233 2.54004
R21902 DVSS.n21158 DVSS.n21157 2.52606
R21903 DVSS.n918 DVSS.n917 2.52606
R21904 DVSS.n915 DVSS.n914 2.52606
R21905 DVSS.n1733 DVSS.n1732 2.41287
R21906 DVSS.n1732 DVSS.n1731 2.41287
R21907 DVSS.n1899 DVSS.n1896 2.41287
R21908 DVSS.n1841 DVSS.n1840 2.41287
R21909 DVSS.n1840 DVSS.n1839 2.41287
R21910 DVSS.n1492 DVSS.n1491 2.41287
R21911 DVSS.n1463 DVSS.n1462 2.41287
R21912 DVSS.n1462 DVSS.n1461 2.41287
R21913 DVSS.n1449 DVSS.n1448 2.41287
R21914 DVSS.n1436 DVSS.n1435 2.41287
R21915 DVSS.n1423 DVSS.n1422 2.41287
R21916 DVSS.n1422 DVSS.n1421 2.41287
R21917 DVSS.n1409 DVSS.n1408 2.41287
R21918 DVSS.n1408 DVSS.n1407 2.41287
R21919 DVSS.n1415 DVSS.n1414 2.41287
R21920 DVSS.n1429 DVSS.n1428 2.41287
R21921 DVSS.n1443 DVSS.n1442 2.41287
R21922 DVSS.n1456 DVSS.n1455 2.41287
R21923 DVSS.n1455 DVSS.n1454 2.41287
R21924 DVSS.n1470 DVSS.n1469 2.41287
R21925 DVSS.n1478 DVSS.n1477 2.41287
R21926 DVSS.n1477 DVSS.n1476 2.41287
R21927 DVSS.n1485 DVSS.n1484 2.41287
R21928 DVSS.n1484 DVSS.n1483 2.41287
R21929 DVSS.n1504 DVSS.n1503 2.41287
R21930 DVSS.n1510 DVSS.n1509 2.41287
R21931 DVSS.n1517 DVSS.n1516 2.41287
R21932 DVSS.n1516 DVSS.n1515 2.41287
R21933 DVSS.n1525 DVSS.n1524 2.41287
R21934 DVSS.n1524 DVSS.n1523 2.41287
R21935 DVSS.n1531 DVSS.n1530 2.41287
R21936 DVSS.n2483 DVSS.n2479 2.41287
R21937 DVSS.n2492 DVSS.n2490 2.41287
R21938 DVSS.n2506 DVSS.n2502 2.41287
R21939 DVSS.n2522 DVSS.n2520 2.41287
R21940 DVSS.n1741 DVSS.n1740 2.41287
R21941 DVSS.n2471 DVSS.n1741 2.41287
R21942 DVSS.n1738 DVSS.n1737 2.41287
R21943 DVSS.n1498 DVSS.n1497 2.41287
R21944 DVSS.n2464 DVSS.n2463 2.41287
R21945 DVSS.n2463 DVSS.n2462 2.41287
R21946 DVSS.n2470 DVSS.n2469 2.41287
R21947 DVSS.n2471 DVSS.n2470 2.41287
R21948 DVSS.n2522 DVSS.n2521 2.41287
R21949 DVSS.n2506 DVSS.n2505 2.41287
R21950 DVSS.n2492 DVSS.n2491 2.41287
R21951 DVSS.n2483 DVSS.n2482 2.41287
R21952 DVSS.n1878 DVSS.n1877 2.41287
R21953 DVSS.n1877 DVSS.n1876 2.41287
R21954 DVSS.n1870 DVSS.n1869 2.41287
R21955 DVSS.n1864 DVSS.n1863 2.41287
R21956 DVSS.n1857 DVSS.n1856 2.41287
R21957 DVSS.n1856 DVSS.n1855 2.41287
R21958 DVSS.n1849 DVSS.n1848 2.41287
R21959 DVSS.n1848 DVSS.n1847 2.41287
R21960 DVSS.n1835 DVSS.n1834 2.41287
R21961 DVSS.n1834 DVSS.n1833 2.41287
R21962 DVSS.n1828 DVSS.n1827 2.41287
R21963 DVSS.n1821 DVSS.n1820 2.41287
R21964 DVSS.n1815 DVSS.n1814 2.41287
R21965 DVSS.n1814 DVSS.n1813 2.41287
R21966 DVSS.n1808 DVSS.n1807 2.41287
R21967 DVSS.n1801 DVSS.n1800 2.41287
R21968 DVSS.n1794 DVSS.n1793 2.41287
R21969 DVSS.n1793 DVSS.n1792 2.41287
R21970 DVSS.n1786 DVSS.n1785 2.41287
R21971 DVSS.n1785 DVSS.n1784 2.41287
R21972 DVSS.n1779 DVSS.n1778 2.41287
R21973 DVSS.n1778 DVSS.n1777 2.41287
R21974 DVSS.n1772 DVSS.n1771 2.41287
R21975 DVSS.n1771 DVSS.n1770 2.41287
R21976 DVSS.n1764 DVSS.n1763 2.41287
R21977 DVSS.n1758 DVSS.n1757 2.41287
R21978 DVSS.n1757 DVSS.n1756 2.41287
R21979 DVSS.n1750 DVSS.n1749 2.41287
R21980 DVSS.n4614 DVSS.n4613 2.41287
R21981 DVSS.n1349 DVSS.n1348 2.41287
R21982 DVSS.n4508 DVSS.n4507 2.41287
R21983 DVSS.n4485 DVSS.n4484 2.41287
R21984 DVSS.n4535 DVSS.n4534 2.41287
R21985 DVSS.n4490 DVSS.n4489 2.41287
R21986 DVSS.n4503 DVSS.n4502 2.41287
R21987 DVSS.n4530 DVSS.n4529 2.41287
R21988 DVSS.n4540 DVSS.n4539 2.41287
R21989 DVSS.n4594 DVSS.n4593 2.41287
R21990 DVSS.n5336 DVSS.n5335 2.41287
R21991 DVSS.n5334 DVSS.n5333 2.41287
R21992 DVSS.n4589 DVSS.n4588 2.41287
R21993 DVSS.n4607 DVSS.n4606 2.41287
R21994 DVSS.n4585 DVSS.n4584 2.41287
R21995 DVSS.n4557 DVSS.n4556 2.41287
R21996 DVSS.n4562 DVSS.n4561 2.41287
R21997 DVSS.n1354 DVSS.n1353 2.41287
R21998 DVSS.n1359 DVSS.n1358 2.41287
R21999 DVSS.n6848 DVSS.n6847 2.41287
R22000 DVSS.n6875 DVSS.n6874 2.41287
R22001 DVSS.n6870 DVSS.n6869 2.41287
R22002 DVSS.n6857 DVSS.n6856 2.41287
R22003 DVSS.n6852 DVSS.n6851 2.41287
R22004 DVSS.n6730 DVSS.n6729 2.41287
R22005 DVSS.n6748 DVSS.n6747 2.41287
R22006 DVSS.n6739 DVSS.n6738 2.41287
R22007 DVSS.n6734 DVSS.n6733 2.41287
R22008 DVSS.n6666 DVSS.n6665 2.41287
R22009 DVSS.n6693 DVSS.n6692 2.41287
R22010 DVSS.n6688 DVSS.n6687 2.41287
R22011 DVSS.n6675 DVSS.n6674 2.41287
R22012 DVSS.n6670 DVSS.n6669 2.41287
R22013 DVSS.n2473 DVSS.n2472 2.41287
R22014 DVSS.n2524 DVSS.n2523 2.41287
R22015 DVSS.n2515 DVSS.n2514 2.41287
R22016 DVSS.n2494 DVSS.n2493 2.41287
R22017 DVSS.n2485 DVSS.n2484 2.41287
R22018 DVSS.n6359 DVSS.n6358 2.41287
R22019 DVSS.n6386 DVSS.n6385 2.41287
R22020 DVSS.n6381 DVSS.n6380 2.41287
R22021 DVSS.n6368 DVSS.n6367 2.41287
R22022 DVSS.n6363 DVSS.n6362 2.41287
R22023 DVSS.n4480 DVSS.n4479 2.41287
R22024 DVSS.n5341 DVSS.n5340 2.41287
R22025 DVSS.n6753 DVSS.n6730 2.41258
R22026 DVSS.n6698 DVSS.n6666 2.41258
R22027 DVSS.n2530 DVSS.n2473 2.41258
R22028 DVSS.n6391 DVSS.n6359 2.41258
R22029 DVSS.n4513 DVSS.n4480 2.41258
R22030 DVSS.n4567 DVSS.n4530 2.41258
R22031 DVSS.n4617 DVSS.n4585 2.41258
R22032 DVSS.n6880 DVSS.n6848 2.41258
R22033 DVSS.n1365 DVSS.n1349 2.41193
R22034 DVSS.n5347 DVSS.n5334 2.41193
R22035 DVSS.n948 DVSS.n947 2.41108
R22036 DVSS.n940 DVSS.n939 2.41079
R22037 DVSS.n21180 DVSS.n21179 2.41079
R22038 DVSS.n930 DVSS.n928 2.40893
R22039 DVSS.n21172 DVSS.n21170 2.40888
R22040 DVSS.n21151 DVSS.n21150 2.37114
R22041 DVSS.n20392 DVSS.n20391 2.35296
R22042 DVSS.n13286 DVSS.n13285 2.35296
R22043 DVSS.n19160 DVSS.n19159 2.32427
R22044 DVSS.n6998 DVSS.n6997 2.32427
R22045 DVSS.n16969 DVSS.n16968 2.3132
R22046 DVSS.n14905 DVSS.n14894 2.3132
R22047 DVSS.n5609 DVSS.n5608 2.25096
R22048 DVSS.n10292 DVSS.n10291 2.25096
R22049 DVSS.n17031 DVSS.n17030 2.25096
R22050 DVSS.n17328 DVSS.n17327 2.25096
R22051 DVSS.n7196 DVSS.n7195 2.25096
R22052 DVSS.n13523 DVSS.n7890 2.25096
R22053 DVSS.n10641 DVSS.n10640 2.25096
R22054 DVSS.n13400 DVSS.n13399 2.25096
R22055 DVSS.n18856 DVSS.n18855 2.25096
R22056 DVSS.n5404 DVSS.n5403 2.25096
R22057 DVSS.n21345 DVSS.n21299 2.25096
R22058 DVSS.n21345 DVSS.n21293 2.25096
R22059 DVSS.n14497 DVSS.n14496 2.25095
R22060 DVSS.n14630 DVSS.n14629 2.25095
R22061 DVSS.n5389 DVSS.n5351 2.25094
R22062 DVSS.n791 DVSS.n768 2.25091
R22063 DVSS.n21253 DVSS.n21237 2.25091
R22064 DVSS.n21345 DVSS.n21344 2.25091
R22065 DVSS.n7170 DVSS.n7169 2.25087
R22066 DVSS.n13536 DVSS.n7873 2.25087
R22067 DVSS.n14473 DVSS.n14472 2.25084
R22068 DVSS.n19144 DVSS.n19116 2.25082
R22069 DVSS.n20426 DVSS.n20398 2.25082
R22070 DVSS.n19418 DVSS.n19390 2.25082
R22071 DVSS.n19666 DVSS.n19643 2.25079
R22072 DVSS.n718 DVSS.n713 2.25078
R22073 DVSS.n21190 DVSS.n21134 2.25078
R22074 DVSS.n718 DVSS.n703 2.25073
R22075 DVSS.n21190 DVSS.n21189 2.25073
R22076 DVSS.n21253 DVSS.n21199 2.25073
R22077 DVSS.n791 DVSS.n784 2.25073
R22078 DVSS.n718 DVSS.n711 2.25069
R22079 DVSS.n21269 DVSS.n21268 2.25069
R22080 DVSS.n791 DVSS.n758 2.25065
R22081 DVSS.n21253 DVSS.n21228 2.25065
R22082 DVSS.n791 DVSS.n772 2.25056
R22083 DVSS.n21253 DVSS.n21241 2.25056
R22084 DVSS.n21190 DVSS.n21128 2.25056
R22085 DVSS.n679 DVSS.n672 2.25051
R22086 DVSS.n718 DVSS.n717 2.25051
R22087 DVSS.n21345 DVSS.n21308 2.25051
R22088 DVSS.n21190 DVSS.n21125 2.25051
R22089 DVSS.n21345 DVSS.n21328 2.25051
R22090 DVSS.n679 DVSS.n678 2.25051
R22091 DVSS.n5586 DVSS.n5576 2.2505
R22092 DVSS.n5586 DVSS.n5581 2.2505
R22093 DVSS.n5586 DVSS.n5585 2.2505
R22094 DVSS.n5601 DVSS.n5600 2.2505
R22095 DVSS.n10270 DVSS.n10250 2.2505
R22096 DVSS.n10270 DVSS.n10256 2.2505
R22097 DVSS.n10270 DVSS.n10269 2.2505
R22098 DVSS.n10284 DVSS.n10283 2.2505
R22099 DVSS.n14341 DVSS.n14336 2.2505
R22100 DVSS.n14338 DVSS.n14337 2.2505
R22101 DVSS.n14333 DVSS.n14332 2.2505
R22102 DVSS.n14329 DVSS.n14328 2.2505
R22103 DVSS.n14232 DVSS.n14231 2.2505
R22104 DVSS.n14235 DVSS.n14230 2.2505
R22105 DVSS.n14225 DVSS.n14224 2.2505
R22106 DVSS.n14212 DVSS.n14209 2.2505
R22107 DVSS.n19663 DVSS.n19662 2.2505
R22108 DVSS.n19638 DVSS.n19637 2.2505
R22109 DVSS.n19167 DVSS.n19160 2.2505
R22110 DVSS.n19162 DVSS.n19161 2.2505
R22111 DVSS.n19141 DVSS.n19140 2.2505
R22112 DVSS.n19116 DVSS.n19115 2.2505
R22113 DVSS.n19110 DVSS.n19109 2.2505
R22114 DVSS.n19643 DVSS.n19642 2.2505
R22115 DVSS.n19681 DVSS.n19680 2.2505
R22116 DVSS.n20175 DVSS.n20168 2.2505
R22117 DVSS.n7788 DVSS.n7787 2.2505
R22118 DVSS.n7791 DVSS.n7786 2.2505
R22119 DVSS.n7796 DVSS.n7795 2.2505
R22120 DVSS.n7799 DVSS.n7794 2.2505
R22121 DVSS.n13839 DVSS.n13838 2.2505
R22122 DVSS.n13695 DVSS.n13694 2.2505
R22123 DVSS.n7838 DVSS.n7835 2.2505
R22124 DVSS.n7840 DVSS.n7839 2.2505
R22125 DVSS.n7850 DVSS.n7843 2.2505
R22126 DVSS.n7847 DVSS.n7846 2.2505
R22127 DVSS.n17009 DVSS.n16998 2.2505
R22128 DVSS.n17009 DVSS.n17004 2.2505
R22129 DVSS.n17009 DVSS.n17008 2.2505
R22130 DVSS.n17023 DVSS.n17022 2.2505
R22131 DVSS.n20170 DVSS.n20169 2.2505
R22132 DVSS.n20152 DVSS.n20139 2.2505
R22133 DVSS.n20148 DVSS.n20147 2.2505
R22134 DVSS.n20142 DVSS.n20141 2.2505
R22135 DVSS.n14475 DVSS.n14139 2.2505
R22136 DVSS.n13676 DVSS.n13673 2.2505
R22137 DVSS.n7864 DVSS.n7863 2.2505
R22138 DVSS.n7858 DVSS.n7857 2.2505
R22139 DVSS.n7856 DVSS.n7855 2.2505
R22140 DVSS.n13684 DVSS.n13683 2.2505
R22141 DVSS.n14180 DVSS.n14179 2.2505
R22142 DVSS.n14364 DVSS.n14363 2.2505
R22143 DVSS.n14354 DVSS.n14353 2.2505
R22144 DVSS.n14348 DVSS.n14347 2.2505
R22145 DVSS.n7005 DVSS.n7002 2.2505
R22146 DVSS.n7008 DVSS.n7001 2.2505
R22147 DVSS.n7011 DVSS.n7000 2.2505
R22148 DVSS.n7014 DVSS.n6999 2.2505
R22149 DVSS.n7017 DVSS.n6998 2.2505
R22150 DVSS.n14790 DVSS.n14789 2.2505
R22151 DVSS.n14644 DVSS.n14643 2.2505
R22152 DVSS.n14055 DVSS.n14054 2.2505
R22153 DVSS.n14059 DVSS.n14058 2.2505
R22154 DVSS.n14051 DVSS.n14050 2.2505
R22155 DVSS.n13990 DVSS.n13989 2.2505
R22156 DVSS.n13977 DVSS.n13976 2.2505
R22157 DVSS.n13986 DVSS.n13983 2.2505
R22158 DVSS.n13980 DVSS.n13979 2.2505
R22159 DVSS.n14805 DVSS.n14804 2.2505
R22160 DVSS.n14045 DVSS.n14044 2.2505
R22161 DVSS.n14041 DVSS.n14040 2.2505
R22162 DVSS.n14049 DVSS.n14048 2.2505
R22163 DVSS.n19900 DVSS.n19894 2.2505
R22164 DVSS.n19896 DVSS.n19895 2.2505
R22165 DVSS.n19878 DVSS.n19871 2.2505
R22166 DVSS.n19874 DVSS.n19873 2.2505
R22167 DVSS.n10630 DVSS.n10629 2.2505
R22168 DVSS.n13194 DVSS.n13193 2.2505
R22169 DVSS.n13198 DVSS.n13197 2.2505
R22170 DVSS.n13278 DVSS.n13277 2.2505
R22171 DVSS.n13282 DVSS.n13281 2.2505
R22172 DVSS.n13287 DVSS.n13286 2.2505
R22173 DVSS.n20446 DVSS.n20445 2.2505
R22174 DVSS.n20440 DVSS.n20439 2.2505
R22175 DVSS.n20423 DVSS.n20422 2.2505
R22176 DVSS.n20398 DVSS.n20385 2.2505
R22177 DVSS.n20393 DVSS.n20392 2.2505
R22178 DVSS.n7350 DVSS.n7349 2.2505
R22179 DVSS.n18701 DVSS.n18700 2.2505
R22180 DVSS.n7336 DVSS.n7335 2.2505
R22181 DVSS.n7346 DVSS.n7345 2.2505
R22182 DVSS.n7342 DVSS.n7341 2.2505
R22183 DVSS.n18588 DVSS.n18585 2.2505
R22184 DVSS.n7430 DVSS.n7427 2.2505
R22185 DVSS.n7424 DVSS.n7423 2.2505
R22186 DVSS.n18598 DVSS.n18595 2.2505
R22187 DVSS.n18592 DVSS.n18591 2.2505
R22188 DVSS.n18714 DVSS.n18711 2.2505
R22189 DVSS.n18734 DVSS.n18731 2.2505
R22190 DVSS.n18728 DVSS.n18727 2.2505
R22191 DVSS.n18724 DVSS.n18721 2.2505
R22192 DVSS.n18718 DVSS.n18717 2.2505
R22193 DVSS.n17304 DVSS.n17270 2.2505
R22194 DVSS.n17304 DVSS.n17274 2.2505
R22195 DVSS.n17304 DVSS.n17303 2.2505
R22196 DVSS.n17319 DVSS.n17318 2.2505
R22197 DVSS.n19438 DVSS.n19437 2.2505
R22198 DVSS.n19432 DVSS.n19431 2.2505
R22199 DVSS.n19415 DVSS.n19414 2.2505
R22200 DVSS.n19390 DVSS.n19380 2.2505
R22201 DVSS.n19385 DVSS.n19384 2.2505
R22202 DVSS.n5389 DVSS.n5388 2.2505
R22203 DVSS.n805 DVSS.n804 2.2505
R22204 DVSS.n21345 DVSS.n21312 2.2505
R22205 DVSS.n21253 DVSS.n21197 2.2505
R22206 DVSS.n19168 DVSS.n19167 2.25047
R22207 DVSS.n20176 DVSS.n20175 2.25047
R22208 DVSS.n13525 DVSS.n7883 2.25047
R22209 DVSS.n7187 DVSS.n7186 2.25047
R22210 DVSS.n13391 DVSS.n7962 2.25047
R22211 DVSS.n20447 DVSS.n20446 2.25047
R22212 DVSS.n18849 DVSS.n7307 2.25047
R22213 DVSS.n19439 DVSS.n19438 2.25047
R22214 DVSS.n718 DVSS.n715 2.25047
R22215 DVSS.n21190 DVSS.n21131 2.25047
R22216 DVSS.n19142 DVSS.n19141 2.25042
R22217 DVSS.n20153 DVSS.n20152 2.25042
R22218 DVSS.n13832 DVSS.n7791 2.25042
R22219 DVSS.n13840 DVSS.n13839 2.25042
R22220 DVSS.n13830 DVSS.n7799 2.25042
R22221 DVSS.n13696 DVSS.n13695 2.25042
R22222 DVSS.n13698 DVSS.n7850 2.25042
R22223 DVSS.n13671 DVSS.n7864 2.25042
R22224 DVSS.n13677 DVSS.n13676 2.25042
R22225 DVSS.n13685 DVSS.n13684 2.25042
R22226 DVSS.n20424 DVSS.n20423 2.25042
R22227 DVSS.n18735 DVSS.n18734 2.25042
R22228 DVSS.n19416 DVSS.n19415 2.25042
R22229 DVSS.n18599 DVSS.n18598 2.25042
R22230 DVSS.n18702 DVSS.n18701 2.25042
R22231 DVSS.n18725 DVSS.n18724 2.25042
R22232 DVSS.n18704 DVSS.n7346 2.25042
R22233 DVSS.n18601 DVSS.n7430 2.25042
R22234 DVSS.n791 DVSS.n754 2.25038
R22235 DVSS.n21253 DVSS.n21225 2.25038
R22236 DVSS.n791 DVSS.n747 2.25038
R22237 DVSS.n21253 DVSS.n21249 2.25038
R22238 DVSS.n19682 DVSS.n19681 2.25037
R22239 DVSS.n14491 DVSS.n14490 2.25037
R22240 DVSS.n14632 DVSS.n14081 2.25037
R22241 DVSS.n19901 DVSS.n19900 2.25037
R22242 DVSS.n14334 DVSS.n14333 2.25031
R22243 DVSS.n14236 DVSS.n14235 2.25031
R22244 DVSS.n14342 DVSS.n14341 2.25031
R22245 DVSS.n14238 DVSS.n14212 2.25031
R22246 DVSS.n19664 DVSS.n19663 2.25031
R22247 DVSS.n14365 DVSS.n14364 2.25031
R22248 DVSS.n14357 DVSS.n14180 2.25031
R22249 DVSS.n14349 DVSS.n14348 2.25031
R22250 DVSS.n14784 DVSS.n14059 2.25031
R22251 DVSS.n19879 DVSS.n19878 2.25031
R22252 DVSS.n14791 DVSS.n14790 2.25031
R22253 DVSS.n14870 DVSS.n13986 2.25031
R22254 DVSS.n14806 DVSS.n14805 2.25031
R22255 DVSS.n14812 DVSS.n14041 2.25031
R22256 DVSS.n14868 DVSS.n13990 2.25031
R22257 DVSS.n14808 DVSS.n14049 2.25031
R22258 DVSS.n791 DVSS.n778 2.25029
R22259 DVSS.n21253 DVSS.n21246 2.25029
R22260 DVSS.n21253 DVSS.n21210 2.25029
R22261 DVSS.n791 DVSS.n790 2.25029
R22262 DVSS.n5505 DVSS.n5504 2.2502
R22263 DVSS.n679 DVSS.n667 2.25016
R22264 DVSS.n21345 DVSS.n21304 2.25016
R22265 DVSS.n679 DVSS.n662 2.25016
R22266 DVSS.n21345 DVSS.n21285 2.25016
R22267 DVSS.n7172 DVSS.n1314 2.25007
R22268 DVSS.n13382 DVSS.n7973 2.25007
R22269 DVSS.n18840 DVSS.n7313 2.25007
R22270 DVSS.n21253 DVSS.n21252 2.24994
R22271 DVSS.n791 DVSS.n735 2.24994
R22272 DVSS.n14651 DVSS.n14650 2.24989
R22273 DVSS.n13378 DVSS.n13377 2.24839
R22274 DVSS.n18836 DVSS.n7316 2.24839
R22275 DVSS.n13700 DVSS.n7838 2.24737
R22276 DVSS.n13679 DVSS.n7856 2.24737
R22277 DVSS.n13199 DVSS.n13198 2.24737
R22278 DVSS.n18715 DVSS.n18714 2.24737
R22279 DVSS.n18694 DVSS.n7350 2.24737
R22280 DVSS.n18589 DVSS.n18588 2.24737
R22281 DVSS.n14226 DVSS.n14225 2.24668
R22282 DVSS.n14355 DVSS.n14354 2.24668
R22283 DVSS.n14793 DVSS.n14051 2.24668
R22284 DVSS.n14810 DVSS.n14045 2.24668
R22285 DVSS.n14872 DVSS.n13977 2.24668
R22286 DVSS.n8029 DVSS.n8024 2.20815
R22287 DVSS.n1364 DVSS.n1352 2.20815
R22288 DVSS.n4566 DVSS.n4533 2.18432
R22289 DVSS.n4512 DVSS.n4483 2.18432
R22290 DVSS.n6390 DVSS.n6361 2.18432
R22291 DVSS.n2529 DVSS.n2475 2.18432
R22292 DVSS.n6697 DVSS.n6668 2.18432
R22293 DVSS.n6752 DVSS.n6732 2.18432
R22294 DVSS.n6879 DVSS.n6850 2.18432
R22295 DVSS.n11185 DVSS.n11179 2.18432
R22296 DVSS.n11015 DVSS.n11009 2.18432
R22297 DVSS.n11724 DVSS.n11718 2.18432
R22298 DVSS.n11675 DVSS.n11669 2.18432
R22299 DVSS.n11638 DVSS.n11632 2.18432
R22300 DVSS.n11513 DVSS.n11507 2.18432
R22301 DVSS.n11476 DVSS.n11475 2.18432
R22302 DVSS.n4616 DVSS.n4587 2.15918
R22303 DVSS.n10025 DVSS.n10019 2.15918
R22304 DVSS.n16804 DVSS.n16803 2.0983
R22305 DVSS.n7642 DVSS.n7641 2.0983
R22306 DVSS.n16011 DVSS.n16010 2.0983
R22307 DVSS.n15308 DVSS.n15307 2.0983
R22308 DVSS.n18010 DVSS.n18009 2.0983
R22309 DVSS.n17869 DVSS.n17868 2.0983
R22310 DVSS.n16969 DVSS.n16966 2.0485
R22311 DVSS.n14905 DVSS.n14904 2.0485
R22312 DVSS.n6879 DVSS.n6878 1.85305
R22313 DVSS.n6879 DVSS.n6873 1.85305
R22314 DVSS.n6879 DVSS.n6860 1.85305
R22315 DVSS.n6879 DVSS.n6855 1.85305
R22316 DVSS.n6752 DVSS.n6751 1.85305
R22317 DVSS.n6752 DVSS.n6746 1.85305
R22318 DVSS.n6752 DVSS.n6742 1.85305
R22319 DVSS.n6752 DVSS.n6737 1.85305
R22320 DVSS.n6697 DVSS.n6696 1.85305
R22321 DVSS.n6697 DVSS.n6691 1.85305
R22322 DVSS.n6697 DVSS.n6678 1.85305
R22323 DVSS.n6697 DVSS.n6673 1.85305
R22324 DVSS.n2529 DVSS.n2528 1.85305
R22325 DVSS.n2529 DVSS.n2519 1.85305
R22326 DVSS.n2529 DVSS.n2498 1.85305
R22327 DVSS.n2529 DVSS.n2489 1.85305
R22328 DVSS.n6390 DVSS.n6389 1.85305
R22329 DVSS.n6390 DVSS.n6384 1.85305
R22330 DVSS.n6390 DVSS.n6371 1.85305
R22331 DVSS.n6390 DVSS.n6366 1.85305
R22332 DVSS.n4512 DVSS.n4511 1.85305
R22333 DVSS.n4512 DVSS.n4506 1.85305
R22334 DVSS.n4512 DVSS.n4493 1.85305
R22335 DVSS.n4512 DVSS.n4488 1.85305
R22336 DVSS.n4566 DVSS.n4565 1.85305
R22337 DVSS.n4566 DVSS.n4560 1.85305
R22338 DVSS.n4566 DVSS.n4543 1.85305
R22339 DVSS.n4566 DVSS.n4538 1.85305
R22340 DVSS.n5346 DVSS.n5339 1.85305
R22341 DVSS.n5346 DVSS.n5344 1.85305
R22342 DVSS.n4616 DVSS.n4615 1.85305
R22343 DVSS.n4616 DVSS.n4610 1.85305
R22344 DVSS.n4616 DVSS.n4597 1.85305
R22345 DVSS.n4616 DVSS.n4592 1.85305
R22346 DVSS.n1364 DVSS.n1357 1.85305
R22347 DVSS.n1364 DVSS.n1362 1.85305
R22348 DVSS.n913 DVSS.n912 1.83783
R22349 DVSS.n1409 DVSS.n1405 1.83517
R22350 DVSS.n1750 DVSS.n1747 1.83517
R22351 DVSS.n13817 DVSS.n13816 1.73383
R22352 DVSS.n13801 DVSS.n13800 1.73383
R22353 DVSS.n7808 DVSS.n7807 1.73383
R22354 DVSS.n7805 DVSS.n7804 1.73383
R22355 DVSS.n7801 DVSS.n7800 1.73383
R22356 DVSS.n14002 DVSS.n14001 1.73383
R22357 DVSS.n13997 DVSS.n13996 1.73383
R22358 DVSS.n13994 DVSS.n13993 1.73383
R22359 DVSS.n14204 DVSS.n14203 1.73383
R22360 DVSS.n14253 DVSS.n14252 1.73383
R22361 DVSS.n14250 DVSS.n14249 1.73383
R22362 DVSS.n18615 DVSS.n18614 1.73383
R22363 DVSS.n18618 DVSS.n18617 1.73383
R22364 DVSS.n18611 DVSS.n18610 1.73383
R22365 DVSS.n7421 DVSS.n7420 1.73383
R22366 DVSS.n7416 DVSS.n7415 1.73383
R22367 DVSS.n13778 DVSS.n13777 1.73383
R22368 DVSS.n13764 DVSS.n13763 1.73383
R22369 DVSS.n7817 DVSS.n7816 1.73383
R22370 DVSS.n7815 DVSS.n7814 1.73383
R22371 DVSS.n7811 DVSS.n7810 1.73383
R22372 DVSS.n14016 DVSS.n14015 1.73383
R22373 DVSS.n14010 DVSS.n14009 1.73383
R22374 DVSS.n14008 DVSS.n14007 1.73383
R22375 DVSS.n14196 DVSS.n14195 1.73383
R22376 DVSS.n14277 DVSS.n14276 1.73383
R22377 DVSS.n14275 DVSS.n14274 1.73383
R22378 DVSS.n18640 DVSS.n18639 1.73383
R22379 DVSS.n18644 DVSS.n18643 1.73383
R22380 DVSS.n18638 DVSS.n18637 1.73383
R22381 DVSS.n7399 DVSS.n7398 1.73383
R22382 DVSS.n7395 DVSS.n7394 1.73383
R22383 DVSS.n13741 DVSS.n13740 1.73383
R22384 DVSS.n13717 DVSS.n13716 1.73383
R22385 DVSS.n7832 DVSS.n7831 1.73383
R22386 DVSS.n7827 DVSS.n7826 1.73383
R22387 DVSS.n7821 DVSS.n7820 1.73383
R22388 DVSS.n14035 DVSS.n14034 1.73383
R22389 DVSS.n14028 DVSS.n14027 1.73383
R22390 DVSS.n14023 DVSS.n14022 1.73383
R22391 DVSS.n14185 DVSS.n14184 1.73383
R22392 DVSS.n14306 DVSS.n14305 1.73383
R22393 DVSS.n14301 DVSS.n14300 1.73383
R22394 DVSS.n18672 DVSS.n18671 1.73383
R22395 DVSS.n18676 DVSS.n18675 1.73383
R22396 DVSS.n18665 DVSS.n18664 1.73383
R22397 DVSS.n7379 DVSS.n7378 1.73383
R22398 DVSS.n7371 DVSS.n7370 1.73383
R22399 DVSS.n7372 DVSS.n7371 1.73383
R22400 DVSS.n7380 DVSS.n7379 1.73383
R22401 DVSS.n18666 DVSS.n18665 1.73383
R22402 DVSS.n18677 DVSS.n18676 1.73383
R22403 DVSS.n18673 DVSS.n18672 1.73383
R22404 DVSS.n14302 DVSS.n14301 1.73383
R22405 DVSS.n14307 DVSS.n14306 1.73383
R22406 DVSS.n14186 DVSS.n14185 1.73383
R22407 DVSS.n14024 DVSS.n14023 1.73383
R22408 DVSS.n14029 DVSS.n14028 1.73383
R22409 DVSS.n14036 DVSS.n14035 1.73383
R22410 DVSS.n7822 DVSS.n7821 1.73383
R22411 DVSS.n7828 DVSS.n7827 1.73383
R22412 DVSS.n7833 DVSS.n7832 1.73383
R22413 DVSS.n13718 DVSS.n13717 1.73383
R22414 DVSS.n13742 DVSS.n13741 1.73383
R22415 DVSS.n16970 DVSS.n16969 1.73383
R22416 DVSS.n7958 DVSS.n7957 1.73383
R22417 DVSS.n14494 DVSS.n14493 1.73383
R22418 DVSS.n14484 DVSS.n14483 1.73383
R22419 DVSS.n7309 DVSS.n7308 1.73383
R22420 DVSS.n18853 DVSS.n18852 1.73383
R22421 DVSS.n7304 DVSS.n7303 1.73383
R22422 DVSS.n7301 DVSS.n7300 1.73383
R22423 DVSS.n7295 DVSS.n7294 1.73383
R22424 DVSS.n7183 DVSS.n7182 1.73383
R22425 DVSS.n7193 DVSS.n7192 1.73383
R22426 DVSS.n7191 DVSS.n7190 1.73383
R22427 DVSS.n7166 DVSS.n7165 1.73383
R22428 DVSS.n7964 DVSS.n7963 1.73383
R22429 DVSS.n7870 DVSS.n7869 1.73383
R22430 DVSS.n14137 DVSS.n14136 1.73383
R22431 DVSS.n14487 DVSS.n14486 1.73383
R22432 DVSS.n13397 DVSS.n13396 1.73383
R22433 DVSS.n13394 DVSS.n13393 1.73383
R22434 DVSS.n7952 DVSS.n7951 1.73383
R22435 DVSS.n7886 DVSS.n7885 1.73383
R22436 DVSS.n7888 DVSS.n7887 1.73383
R22437 DVSS.n7880 DVSS.n7879 1.73383
R22438 DVSS.n14647 DVSS.n14646 1.73383
R22439 DVSS.n14641 DVSS.n14640 1.73383
R22440 DVSS.n14628 DVSS.n14627 1.73383
R22441 DVSS.n14625 DVSS.n14624 1.73383
R22442 DVSS.n13350 DVSS.n13349 1.73383
R22443 DVSS.n13349 DVSS.n13348 1.73383
R22444 DVSS.n13272 DVSS.n13271 1.73383
R22445 DVSS.n13271 DVSS.n13270 1.73383
R22446 DVSS.n8004 DVSS.n8003 1.73383
R22447 DVSS.n8003 DVSS.n8002 1.73383
R22448 DVSS.n7996 DVSS.n7995 1.73383
R22449 DVSS.n7995 DVSS.n7994 1.73383
R22450 DVSS.n7990 DVSS.n7989 1.73383
R22451 DVSS.n7989 DVSS.n7988 1.73383
R22452 DVSS.n7985 DVSS.n7984 1.73383
R22453 DVSS.n7981 DVSS.n7980 1.73383
R22454 DVSS.n7977 DVSS.n7976 1.73383
R22455 DVSS.n14067 DVSS.n14066 1.73383
R22456 DVSS.n14072 DVSS.n14071 1.73383
R22457 DVSS.n14071 DVSS.n14070 1.73383
R22458 DVSS.n14685 DVSS.n14684 1.73383
R22459 DVSS.n14684 DVSS.n14683 1.73383
R22460 DVSS.n14142 DVSS.n14141 1.73383
R22461 DVSS.n14141 DVSS.n14140 1.73383
R22462 DVSS.n18807 DVSS.n18806 1.73383
R22463 DVSS.n18806 DVSS.n18805 1.73383
R22464 DVSS.n18811 DVSS.n18810 1.73383
R22465 DVSS.n18810 DVSS.n18809 1.73383
R22466 DVSS.n18800 DVSS.n18799 1.73383
R22467 DVSS.n18799 DVSS.n18798 1.73383
R22468 DVSS.n7333 DVSS.n7332 1.73383
R22469 DVSS.n7332 DVSS.n7331 1.73383
R22470 DVSS.n7325 DVSS.n7324 1.73383
R22471 DVSS.n7324 DVSS.n7323 1.73383
R22472 DVSS.n7319 DVSS.n7318 1.73383
R22473 DVSS.n7318 DVSS.n7317 1.73383
R22474 DVSS.n14065 DVSS.n14064 1.73383
R22475 DVSS.n14064 DVSS.n14063 1.73383
R22476 DVSS.n14689 DVSS.n14688 1.73383
R22477 DVSS.n14688 DVSS.n14687 1.73383
R22478 DVSS.n14439 DVSS.n14438 1.73383
R22479 DVSS.n14438 DVSS.n14437 1.73383
R22480 DVSS.n14148 DVSS.n14147 1.73383
R22481 DVSS.n14147 DVSS.n14146 1.73383
R22482 DVSS.n7127 DVSS.n7126 1.73383
R22483 DVSS.n7126 DVSS.n7125 1.73383
R22484 DVSS.n7121 DVSS.n7120 1.73383
R22485 DVSS.n7120 DVSS.n7119 1.73383
R22486 DVSS.n1343 DVSS.n1342 1.73383
R22487 DVSS.n1342 DVSS.n1341 1.73383
R22488 DVSS.n1337 DVSS.n1336 1.73383
R22489 DVSS.n1336 DVSS.n1335 1.73383
R22490 DVSS.n13627 DVSS.n13626 1.73383
R22491 DVSS.n13626 DVSS.n13625 1.73383
R22492 DVSS.n13636 DVSS.n13635 1.73383
R22493 DVSS.n13635 DVSS.n13634 1.73383
R22494 DVSS.n13616 DVSS.n13615 1.73383
R22495 DVSS.n13615 DVSS.n13614 1.73383
R22496 DVSS.n13607 DVSS.n13606 1.73383
R22497 DVSS.n13606 DVSS.n13605 1.73383
R22498 DVSS.n13598 DVSS.n13597 1.73383
R22499 DVSS.n14749 DVSS.n14748 1.73383
R22500 DVSS.n14169 DVSS.n14168 1.73383
R22501 DVSS.n14158 DVSS.n14157 1.73383
R22502 DVSS.n7049 DVSS.n7048 1.73383
R22503 DVSS.n7054 DVSS.n7053 1.73383
R22504 DVSS.n7057 DVSS.n7056 1.73383
R22505 DVSS.n7063 DVSS.n7062 1.73383
R22506 DVSS.n7069 DVSS.n7068 1.73383
R22507 DVSS.n7076 DVSS.n7075 1.73383
R22508 DVSS.n7082 DVSS.n7081 1.73383
R22509 DVSS.n7042 DVSS.n7041 1.73383
R22510 DVSS.n7035 DVSS.n7034 1.73383
R22511 DVSS.n14745 DVSS.n14744 1.73383
R22512 DVSS.n14738 DVSS.n14737 1.73383
R22513 DVSS.n14176 DVSS.n14175 1.73383
R22514 DVSS.n13305 DVSS.n13304 1.73383
R22515 DVSS.n13316 DVSS.n13315 1.73383
R22516 DVSS.n13309 DVSS.n13308 1.73383
R22517 DVSS.n13299 DVSS.n13298 1.73383
R22518 DVSS.n13620 DVSS.n13619 1.73383
R22519 DVSS.n14165 DVSS.n14164 1.73383
R22520 DVSS.n14910 DVSS.n14890 1.68445
R22521 DVSS.n14910 DVSS.n14908 1.68445
R22522 DVSS.n4556 DVSS.n4553 1.61232
R22523 DVSS.n4556 DVSS.n4549 1.61232
R22524 DVSS.n4556 DVSS.n4548 1.61232
R22525 DVSS.n4556 DVSS.n4554 1.61232
R22526 DVSS.n1456 DVSS.n1453 1.5005
R22527 DVSS.n1899 DVSS.n1898 1.5005
R22528 DVSS.n1733 DVSS.n1729 1.5005
R22529 DVSS.n1841 DVSS.n1838 1.5005
R22530 DVSS.n1492 DVSS.n1490 1.5005
R22531 DVSS.n1470 DVSS.n1468 1.5005
R22532 DVSS.n1463 DVSS.n1460 1.5005
R22533 DVSS.n1449 DVSS.n1447 1.5005
R22534 DVSS.n1443 DVSS.n1441 1.5005
R22535 DVSS.n1436 DVSS.n1434 1.5005
R22536 DVSS.n1429 DVSS.n1427 1.5005
R22537 DVSS.n1423 DVSS.n1420 1.5005
R22538 DVSS.n1415 DVSS.n1413 1.5005
R22539 DVSS.n1409 DVSS.n1406 1.5005
R22540 DVSS.n1478 DVSS.n1475 1.5005
R22541 DVSS.n1485 DVSS.n1482 1.5005
R22542 DVSS.n1504 DVSS.n1502 1.5005
R22543 DVSS.n1510 DVSS.n1508 1.5005
R22544 DVSS.n1517 DVSS.n1514 1.5005
R22545 DVSS.n1525 DVSS.n1522 1.5005
R22546 DVSS.n1531 DVSS.n1529 1.5005
R22547 DVSS.n1535 DVSS.n1534 1.5005
R22548 DVSS.n1539 DVSS.n1538 1.5005
R22549 DVSS.n1543 DVSS.n1542 1.5005
R22550 DVSS.n1547 DVSS.n1546 1.5005
R22551 DVSS.n1740 DVSS.n1551 1.5005
R22552 DVSS.n1738 DVSS.n1728 1.5005
R22553 DVSS.n1498 DVSS.n1496 1.5005
R22554 DVSS.n2464 DVSS.n2461 1.5005
R22555 DVSS.n2469 DVSS.n2468 1.5005
R22556 DVSS.n1894 DVSS.n1893 1.5005
R22557 DVSS.n1890 DVSS.n1889 1.5005
R22558 DVSS.n1886 DVSS.n1885 1.5005
R22559 DVSS.n1882 DVSS.n1881 1.5005
R22560 DVSS.n1878 DVSS.n1875 1.5005
R22561 DVSS.n1870 DVSS.n1868 1.5005
R22562 DVSS.n1864 DVSS.n1862 1.5005
R22563 DVSS.n1857 DVSS.n1854 1.5005
R22564 DVSS.n1849 DVSS.n1846 1.5005
R22565 DVSS.n1835 DVSS.n1832 1.5005
R22566 DVSS.n1828 DVSS.n1826 1.5005
R22567 DVSS.n1821 DVSS.n1819 1.5005
R22568 DVSS.n1815 DVSS.n1812 1.5005
R22569 DVSS.n1808 DVSS.n1806 1.5005
R22570 DVSS.n1801 DVSS.n1799 1.5005
R22571 DVSS.n1794 DVSS.n1791 1.5005
R22572 DVSS.n1786 DVSS.n1783 1.5005
R22573 DVSS.n1779 DVSS.n1776 1.5005
R22574 DVSS.n1772 DVSS.n1769 1.5005
R22575 DVSS.n1764 DVSS.n1762 1.5005
R22576 DVSS.n1758 DVSS.n1755 1.5005
R22577 DVSS.n1750 DVSS.n1748 1.5005
R22578 DVSS.n18290 DVSS.n18275 1.5005
R22579 DVSS.n18096 DVSS.n18095 1.5005
R22580 DVSS.n17872 DVSS.n17871 1.5005
R22581 DVSS.n17858 DVSS.n17857 1.5005
R22582 DVSS.n17850 DVSS.n17849 1.5005
R22583 DVSS.n17842 DVSS.n17841 1.5005
R22584 DVSS.n17834 DVSS.n17833 1.5005
R22585 DVSS.n17826 DVSS.n17825 1.5005
R22586 DVSS.n17818 DVSS.n17817 1.5005
R22587 DVSS.n17814 DVSS.n17813 1.5005
R22588 DVSS.n17822 DVSS.n17821 1.5005
R22589 DVSS.n17830 DVSS.n17829 1.5005
R22590 DVSS.n17838 DVSS.n17837 1.5005
R22591 DVSS.n17846 DVSS.n17845 1.5005
R22592 DVSS.n17854 DVSS.n17853 1.5005
R22593 DVSS.n17862 DVSS.n17861 1.5005
R22594 DVSS.n17898 DVSS.n17897 1.5005
R22595 DVSS.n18013 DVSS.n18012 1.5005
R22596 DVSS.n17999 DVSS.n17998 1.5005
R22597 DVSS.n17991 DVSS.n17990 1.5005
R22598 DVSS.n17983 DVSS.n17982 1.5005
R22599 DVSS.n17975 DVSS.n17974 1.5005
R22600 DVSS.n17967 DVSS.n17966 1.5005
R22601 DVSS.n17959 DVSS.n17958 1.5005
R22602 DVSS.n17955 DVSS.n17954 1.5005
R22603 DVSS.n17963 DVSS.n17962 1.5005
R22604 DVSS.n17971 DVSS.n17970 1.5005
R22605 DVSS.n17979 DVSS.n17978 1.5005
R22606 DVSS.n17987 DVSS.n17986 1.5005
R22607 DVSS.n17995 DVSS.n17994 1.5005
R22608 DVSS.n18003 DVSS.n18002 1.5005
R22609 DVSS.n18039 DVSS.n18038 1.5005
R22610 DVSS.n14208 DVSS.n14205 1.5005
R22611 DVSS.n14202 DVSS.n14201 1.5005
R22612 DVSS.n14254 DVSS.n14251 1.5005
R22613 DVSS.n14248 DVSS.n14247 1.5005
R22614 DVSS.n14200 DVSS.n14199 1.5005
R22615 DVSS.n14194 DVSS.n14193 1.5005
R22616 DVSS.n14279 DVSS.n14278 1.5005
R22617 DVSS.n14273 DVSS.n14272 1.5005
R22618 DVSS.n14299 DVSS.n14298 1.5005
R22619 DVSS.n14298 DVSS.n14297 1.5005
R22620 DVSS.n14308 DVSS.n14304 1.5005
R22621 DVSS.n14304 DVSS.n14303 1.5005
R22622 DVSS.n14183 DVSS.n14182 1.5005
R22623 DVSS.n14182 DVSS.n14181 1.5005
R22624 DVSS.n14192 DVSS.n14188 1.5005
R22625 DVSS.n14188 DVSS.n14187 1.5005
R22626 DVSS.n17491 DVSS.n17490 1.5005
R22627 DVSS.n16448 DVSS.n16447 1.5005
R22628 DVSS.n16456 DVSS.n16455 1.5005
R22629 DVSS.n16464 DVSS.n16463 1.5005
R22630 DVSS.n16472 DVSS.n16471 1.5005
R22631 DVSS.n16480 DVSS.n16479 1.5005
R22632 DVSS.n16488 DVSS.n16487 1.5005
R22633 DVSS.n16499 DVSS.n16498 1.5005
R22634 DVSS.n16492 DVSS.n16491 1.5005
R22635 DVSS.n16484 DVSS.n16483 1.5005
R22636 DVSS.n16476 DVSS.n16475 1.5005
R22637 DVSS.n16468 DVSS.n16467 1.5005
R22638 DVSS.n16460 DVSS.n16459 1.5005
R22639 DVSS.n16452 DVSS.n16451 1.5005
R22640 DVSS.n16014 DVSS.n16013 1.5005
R22641 DVSS.n16630 DVSS.n16629 1.5005
R22642 DVSS.n16624 DVSS.n16623 1.5005
R22643 DVSS.n16620 DVSS.n16619 1.5005
R22644 DVSS.n16616 DVSS.n16615 1.5005
R22645 DVSS.n16612 DVSS.n16611 1.5005
R22646 DVSS.n17721 DVSS.n17720 1.5005
R22647 DVSS.n7644 DVSS.n7643 1.5005
R22648 DVSS.n16018 DVSS.n16017 1.5005
R22649 DVSS.n16022 DVSS.n16021 1.5005
R22650 DVSS.n16026 DVSS.n16025 1.5005
R22651 DVSS.n16030 DVSS.n16029 1.5005
R22652 DVSS.n16034 DVSS.n16033 1.5005
R22653 DVSS.n16038 DVSS.n16037 1.5005
R22654 DVSS.n16042 DVSS.n16041 1.5005
R22655 DVSS.n16058 DVSS.n16057 1.5005
R22656 DVSS.n16085 DVSS.n16084 1.5005
R22657 DVSS.n16098 DVSS.n16097 1.5005
R22658 DVSS.n13815 DVSS.n13803 1.5005
R22659 DVSS.n13818 DVSS.n13802 1.5005
R22660 DVSS.n13799 DVSS.n13798 1.5005
R22661 DVSS.n7809 DVSS.n7806 1.5005
R22662 DVSS.n7803 DVSS.n7802 1.5005
R22663 DVSS.n13738 DVSS.n13737 1.5005
R22664 DVSS.n13776 DVSS.n13775 1.5005
R22665 DVSS.n13780 DVSS.n13779 1.5005
R22666 DVSS.n13762 DVSS.n13761 1.5005
R22667 DVSS.n7819 DVSS.n7818 1.5005
R22668 DVSS.n7813 DVSS.n7812 1.5005
R22669 DVSS.n7825 DVSS.n7824 1.5005
R22670 DVSS.n7824 DVSS.n7823 1.5005
R22671 DVSS.n7834 DVSS.n7830 1.5005
R22672 DVSS.n7830 DVSS.n7829 1.5005
R22673 DVSS.n13715 DVSS.n13714 1.5005
R22674 DVSS.n13714 DVSS.n13713 1.5005
R22675 DVSS.n13743 DVSS.n13720 1.5005
R22676 DVSS.n13720 DVSS.n13719 1.5005
R22677 DVSS.n13739 DVSS.n13738 1.5005
R22678 DVSS.n14472 DVSS.n14471 1.5005
R22679 DVSS.n14139 DVSS.n14138 1.5005
R22680 DVSS.n14490 DVSS.n14489 1.5005
R22681 DVSS.n1314 DVSS.n1313 1.5005
R22682 DVSS.n7186 DVSS.n7185 1.5005
R22683 DVSS.n7195 DVSS.n7194 1.5005
R22684 DVSS.n7169 DVSS.n7168 1.5005
R22685 DVSS.n7873 DVSS.n7872 1.5005
R22686 DVSS.n7890 DVSS.n7889 1.5005
R22687 DVSS.n7883 DVSS.n7882 1.5005
R22688 DVSS.n7877 DVSS.n7876 1.5005
R22689 DVSS.n7867 DVSS.n7866 1.5005
R22690 DVSS.n7163 DVSS.n7162 1.5005
R22691 DVSS.n14496 DVSS.n14495 1.5005
R22692 DVSS.n7987 DVSS.n7986 1.5005
R22693 DVSS.n7983 DVSS.n7982 1.5005
R22694 DVSS.n7979 DVSS.n7978 1.5005
R22695 DVSS.n7975 DVSS.n7974 1.5005
R22696 DVSS.n14069 DVSS.n14068 1.5005
R22697 DVSS.n14442 DVSS.n14441 1.5005
R22698 DVSS.n14441 DVSS.n14440 1.5005
R22699 DVSS.n14436 DVSS.n14435 1.5005
R22700 DVSS.n14435 DVSS.n14434 1.5005
R22701 DVSS.n14145 DVSS.n14144 1.5005
R22702 DVSS.n14144 DVSS.n14143 1.5005
R22703 DVSS.n14151 DVSS.n14150 1.5005
R22704 DVSS.n14150 DVSS.n14149 1.5005
R22705 DVSS.n7124 DVSS.n7123 1.5005
R22706 DVSS.n7123 DVSS.n7122 1.5005
R22707 DVSS.n7130 DVSS.n7129 1.5005
R22708 DVSS.n7129 DVSS.n7128 1.5005
R22709 DVSS.n1340 DVSS.n1339 1.5005
R22710 DVSS.n1339 DVSS.n1338 1.5005
R22711 DVSS.n1346 DVSS.n1345 1.5005
R22712 DVSS.n1345 DVSS.n1344 1.5005
R22713 DVSS.n1334 DVSS.n1333 1.5005
R22714 DVSS.n1333 DVSS.n1332 1.5005
R22715 DVSS.n13623 DVSS.n13618 1.5005
R22716 DVSS.n13618 DVSS.n13617 1.5005
R22717 DVSS.n13632 DVSS.n13631 1.5005
R22718 DVSS.n13631 DVSS.n13630 1.5005
R22719 DVSS.n13639 DVSS.n13638 1.5005
R22720 DVSS.n13638 DVSS.n13637 1.5005
R22721 DVSS.n13612 DVSS.n13611 1.5005
R22722 DVSS.n13611 DVSS.n13610 1.5005
R22723 DVSS.n13603 DVSS.n13602 1.5005
R22724 DVSS.n13602 DVSS.n13601 1.5005
R22725 DVSS.n14172 DVSS.n14170 1.5005
R22726 DVSS.n14178 DVSS.n14177 1.5005
R22727 DVSS.n7073 DVSS.n7072 1.5005
R22728 DVSS.n7079 DVSS.n7043 1.5005
R22729 DVSS.n7039 DVSS.n7038 1.5005
R22730 DVSS.n7032 DVSS.n7031 1.5005
R22731 DVSS.n7084 DVSS.n7083 1.5005
R22732 DVSS.n14162 DVSS.n14161 1.5005
R22733 DVSS.n14167 DVSS.n14166 1.5005
R22734 DVSS.n14742 DVSS.n14739 1.5005
R22735 DVSS.n14747 DVSS.n14746 1.5005
R22736 DVSS.n14751 DVSS.n14750 1.5005
R22737 DVSS.n15402 DVSS.n15401 1.5005
R22738 DVSS.n15438 DVSS.n15437 1.5005
R22739 DVSS.n14004 DVSS.n14003 1.5005
R22740 DVSS.n14000 DVSS.n13999 1.5005
R22741 DVSS.n13998 DVSS.n13995 1.5005
R22742 DVSS.n13992 DVSS.n13991 1.5005
R22743 DVSS.n14018 DVSS.n14017 1.5005
R22744 DVSS.n14014 DVSS.n14013 1.5005
R22745 DVSS.n14012 DVSS.n14011 1.5005
R22746 DVSS.n14006 DVSS.n14005 1.5005
R22747 DVSS.n14021 DVSS.n14020 1.5005
R22748 DVSS.n14020 DVSS.n14019 1.5005
R22749 DVSS.n14030 DVSS.n14026 1.5005
R22750 DVSS.n14026 DVSS.n14025 1.5005
R22751 DVSS.n14033 DVSS.n14032 1.5005
R22752 DVSS.n14032 DVSS.n14031 1.5005
R22753 DVSS.n14039 DVSS.n14038 1.5005
R22754 DVSS.n14038 DVSS.n14037 1.5005
R22755 DVSS.n15191 DVSS.n15190 1.5005
R22756 DVSS.n15209 DVSS.n15208 1.5005
R22757 DVSS.n15216 DVSS.n15215 1.5005
R22758 DVSS.n15301 DVSS.n15300 1.5005
R22759 DVSS.n15311 DVSS.n15310 1.5005
R22760 DVSS.n15315 DVSS.n15314 1.5005
R22761 DVSS.n15319 DVSS.n15318 1.5005
R22762 DVSS.n15323 DVSS.n15322 1.5005
R22763 DVSS.n15327 DVSS.n15326 1.5005
R22764 DVSS.n15331 DVSS.n15330 1.5005
R22765 DVSS.n15335 DVSS.n15334 1.5005
R22766 DVSS.n15339 DVSS.n15338 1.5005
R22767 DVSS.n15343 DVSS.n15342 1.5005
R22768 DVSS.n15347 DVSS.n15346 1.5005
R22769 DVSS.n15351 DVSS.n15350 1.5005
R22770 DVSS.n15355 DVSS.n15354 1.5005
R22771 DVSS.n15359 DVSS.n15358 1.5005
R22772 DVSS.n15366 DVSS.n15365 1.5005
R22773 DVSS.n15157 DVSS.n15156 1.5005
R22774 DVSS.n15117 DVSS.n15116 1.5005
R22775 DVSS.n16783 DVSS.n16782 1.5005
R22776 DVSS.n16787 DVSS.n16786 1.5005
R22777 DVSS.n16792 DVSS.n16791 1.5005
R22778 DVSS.n16796 DVSS.n16795 1.5005
R22779 DVSS.n16806 DVSS.n16805 1.5005
R22780 DVSS.n17189 DVSS.n17188 1.5005
R22781 DVSS.n14075 DVSS.n14074 1.5005
R22782 DVSS.n14074 DVSS.n14073 1.5005
R22783 DVSS.n14062 DVSS.n14061 1.5005
R22784 DVSS.n14061 DVSS.n14060 1.5005
R22785 DVSS.n14686 DVSS.n14682 1.5005
R22786 DVSS.n14682 DVSS.n14681 1.5005
R22787 DVSS.n14690 DVSS.n14680 1.5005
R22788 DVSS.n14680 DVSS.n14679 1.5005
R22789 DVSS.n14734 DVSS.n14733 1.5005
R22790 DVSS.n14650 DVSS.n14649 1.5005
R22791 DVSS.n14643 DVSS.n14642 1.5005
R22792 DVSS.n14081 DVSS.n14079 1.5005
R22793 DVSS.n14629 DVSS.n14626 1.5005
R22794 DVSS.n13918 DVSS.n13917 1.5005
R22795 DVSS.n13908 DVSS.n13907 1.5005
R22796 DVSS.n13900 DVSS.n13899 1.5005
R22797 DVSS.n13892 DVSS.n13891 1.5005
R22798 DVSS.n13884 DVSS.n13883 1.5005
R22799 DVSS.n13876 DVSS.n13875 1.5005
R22800 DVSS.n13868 DVSS.n13867 1.5005
R22801 DVSS.n13864 DVSS.n13863 1.5005
R22802 DVSS.n13872 DVSS.n13871 1.5005
R22803 DVSS.n13880 DVSS.n13879 1.5005
R22804 DVSS.n13888 DVSS.n13887 1.5005
R22805 DVSS.n13896 DVSS.n13895 1.5005
R22806 DVSS.n13904 DVSS.n13903 1.5005
R22807 DVSS.n13912 DVSS.n13911 1.5005
R22808 DVSS.n13933 DVSS.n13932 1.5005
R22809 DVSS.n13319 DVSS.n13318 1.5005
R22810 DVSS.n13313 DVSS.n13312 1.5005
R22811 DVSS.n13307 DVSS.n13306 1.5005
R22812 DVSS.n13302 DVSS.n13301 1.5005
R22813 DVSS.n13295 DVSS.n13294 1.5005
R22814 DVSS.n13346 DVSS.n13345 1.5005
R22815 DVSS.n13351 DVSS.n13274 1.5005
R22816 DVSS.n13274 DVSS.n13273 1.5005
R22817 DVSS.n8001 DVSS.n8000 1.5005
R22818 DVSS.n8000 DVSS.n7999 1.5005
R22819 DVSS.n8005 DVSS.n7998 1.5005
R22820 DVSS.n7998 DVSS.n7997 1.5005
R22821 DVSS.n7993 DVSS.n7992 1.5005
R22822 DVSS.n7992 DVSS.n7991 1.5005
R22823 DVSS.n13347 DVSS.n13346 1.5005
R22824 DVSS.n13377 DVSS.n13375 1.5005
R22825 DVSS.n13399 DVSS.n13398 1.5005
R22826 DVSS.n7962 DVSS.n7960 1.5005
R22827 DVSS.n7955 DVSS.n7954 1.5005
R22828 DVSS.n7973 DVSS.n7972 1.5005
R22829 DVSS.n7313 DVSS.n7312 1.5005
R22830 DVSS.n7316 DVSS.n7315 1.5005
R22831 DVSS.n18855 DVSS.n18854 1.5005
R22832 DVSS.n7307 DVSS.n7306 1.5005
R22833 DVSS.n7298 DVSS.n7297 1.5005
R22834 DVSS.n14154 DVSS.n14153 1.5005
R22835 DVSS.n7051 DVSS.n7047 1.5005
R22836 DVSS.n7055 DVSS.n7046 1.5005
R22837 DVSS.n7060 DVSS.n7045 1.5005
R22838 DVSS.n7065 DVSS.n7044 1.5005
R22839 DVSS.n18616 DVSS.n18613 1.5005
R22840 DVSS.n18619 DVSS.n18612 1.5005
R22841 DVSS.n7419 DVSS.n7418 1.5005
R22842 DVSS.n7422 DVSS.n7417 1.5005
R22843 DVSS.n18642 DVSS.n18641 1.5005
R22844 DVSS.n18646 DVSS.n18645 1.5005
R22845 DVSS.n7397 DVSS.n7396 1.5005
R22846 DVSS.n7401 DVSS.n7400 1.5005
R22847 DVSS.n7393 DVSS.n7392 1.5005
R22848 DVSS.n7369 DVSS.n7368 1.5005
R22849 DVSS.n7368 DVSS.n7367 1.5005
R22850 DVSS.n7381 DVSS.n7374 1.5005
R22851 DVSS.n7374 DVSS.n7373 1.5005
R22852 DVSS.n7377 DVSS.n7376 1.5005
R22853 DVSS.n7376 DVSS.n7375 1.5005
R22854 DVSS.n18678 DVSS.n18668 1.5005
R22855 DVSS.n18668 DVSS.n18667 1.5005
R22856 DVSS.n18674 DVSS.n18670 1.5005
R22857 DVSS.n18670 DVSS.n18669 1.5005
R22858 DVSS.n7414 DVSS.n7413 1.5005
R22859 DVSS.n18808 DVSS.n18804 1.5005
R22860 DVSS.n18804 DVSS.n18803 1.5005
R22861 DVSS.n18812 DVSS.n18802 1.5005
R22862 DVSS.n18802 DVSS.n18801 1.5005
R22863 DVSS.n7330 DVSS.n7329 1.5005
R22864 DVSS.n7329 DVSS.n7328 1.5005
R22865 DVSS.n7334 DVSS.n7327 1.5005
R22866 DVSS.n7327 DVSS.n7326 1.5005
R22867 DVSS.n7322 DVSS.n7321 1.5005
R22868 DVSS.n7321 DVSS.n7320 1.5005
R22869 DVSS.n5816 DVSS.n5813 1.50017
R22870 DVSS.n11045 DVSS.n11044 1.50017
R22871 DVSS.n16903 DVSS.n16902 1.50017
R22872 DVSS.n7131 DVSS.n7130 1.50017
R22873 DVSS.n10968 DVSS.n10053 1.50017
R22874 DVSS.n17102 DVSS.n17101 1.50017
R22875 DVSS.n5677 DVSS.n5553 1.50017
R22876 DVSS.n9991 DVSS.n9990 1.50017
R22877 DVSS.n11067 DVSS.n11066 1.50017
R22878 DVSS.n13352 DVSS.n13351 1.50017
R22879 DVSS.n18620 DVSS.n18619 1.50017
R22880 DVSS.n18647 DVSS.n18646 1.50017
R22881 DVSS.n18679 DVSS.n18678 1.50017
R22882 DVSS.n17446 DVSS.n17445 1.50017
R22883 DVSS.n17396 DVSS.n17248 1.50017
R22884 DVSS.n5836 DVSS.n5835 1.50017
R22885 DVSS.n6472 DVSS.n6471 1.50017
R22886 DVSS.n7133 DVSS.n1346 1.50013
R22887 DVSS.n13354 DVSS.n8005 1.50013
R22888 DVSS.n13746 DVSS.n7834 1.50006
R22889 DVSS.n13783 DVSS.n7819 1.50006
R22890 DVSS.n13821 DVSS.n7809 1.50006
R22891 DVSS.n18813 DVSS.n18812 1.50006
R22892 DVSS.n5811 DVSS.n5810 1.50002
R22893 DVSS.n11052 DVSS.n11047 1.50002
R22894 DVSS.n13744 DVSS.n13743 1.50002
R22895 DVSS.n13781 DVSS.n13780 1.50002
R22896 DVSS.n13819 DVSS.n13818 1.50002
R22897 DVSS.n17553 DVSS.n17552 1.50002
R22898 DVSS.n13640 DVSS.n13639 1.50002
R22899 DVSS.n7085 DVSS.n7084 1.50002
R22900 DVSS.n11076 DVSS.n11075 1.50002
R22901 DVSS.n18622 DVSS.n7422 1.50002
R22902 DVSS.n18649 DVSS.n7401 1.50002
R22903 DVSS.n18681 DVSS.n7381 1.50002
R22904 DVSS.n18815 DVSS.n7334 1.50002
R22905 DVSS.n17449 DVSS.n17448 1.50002
R22906 DVSS.n14693 DVSS.n14075 1.49999
R22907 DVSS.n17114 DVSS.n17113 1.49999
R22908 DVSS.n17236 DVSS.n16708 1.49999
R22909 DVSS.n17464 DVSS.n17463 1.49999
R22910 DVSS.n14443 DVSS.n14442 1.49999
R22911 DVSS.n17541 DVSS.n17539 1.49999
R22912 DVSS.n11215 DVSS.n11214 1.49998
R22913 DVSS.n6503 DVSS.n6502 1.49998
R22914 DVSS.n17654 DVSS.n17653 1.49998
R22915 DVSS.n17645 DVSS.n17644 1.49998
R22916 DVSS.n9832 DVSS.n9831 1.49998
R22917 DVSS.n11165 DVSS.n11164 1.49998
R22918 DVSS.n16323 DVSS.n16322 1.49998
R22919 DVSS.n16341 DVSS.n16340 1.49998
R22920 DVSS.n14445 DVSS.n14151 1.49994
R22921 DVSS.n17798 DVSS.n7634 1.49989
R22922 DVSS.n14309 DVSS.n14308 1.49987
R22923 DVSS.n14280 DVSS.n14279 1.49987
R22924 DVSS.n14255 DVSS.n14254 1.49987
R22925 DVSS.n14859 DVSS.n13998 1.49987
R22926 DVSS.n14842 DVSS.n14012 1.49987
R22927 DVSS.n14825 DVSS.n14030 1.49987
R22928 DVSS.n14311 DVSS.n14192 1.49983
R22929 DVSS.n14282 DVSS.n14200 1.49983
R22930 DVSS.n14257 DVSS.n14208 1.49983
R22931 DVSS.n17456 DVSS.n17455 1.49983
R22932 DVSS.n14397 DVSS.n14178 1.49983
R22933 DVSS.n14752 DVSS.n14751 1.49983
R22934 DVSS.n14857 DVSS.n14004 1.49983
R22935 DVSS.n14840 DVSS.n14018 1.49983
R22936 DVSS.n14823 DVSS.n14039 1.49983
R22937 DVSS.n17537 DVSS.n17536 1.49983
R22938 DVSS.n14691 DVSS.n14690 1.49983
R22939 DVSS.n17675 DVSS.n17672 1.49978
R22940 DVSS.n17664 DVSS.n17663 1.49978
R22941 DVSS.n5344 DVSS.n5343 1.49689
R22942 DVSS.n5339 DVSS.n5338 1.49689
R22943 DVSS.n4592 DVSS.n4591 1.49689
R22944 DVSS.n4597 DVSS.n4596 1.49689
R22945 DVSS.n4610 DVSS.n4609 1.49689
R22946 DVSS.n4615 DVSS.n4614 1.49689
R22947 DVSS.n4538 DVSS.n4537 1.49689
R22948 DVSS.n4543 DVSS.n4542 1.49689
R22949 DVSS.n4560 DVSS.n4559 1.49689
R22950 DVSS.n4565 DVSS.n4564 1.49689
R22951 DVSS.n4488 DVSS.n4487 1.49689
R22952 DVSS.n4493 DVSS.n4492 1.49689
R22953 DVSS.n4506 DVSS.n4505 1.49689
R22954 DVSS.n4511 DVSS.n4510 1.49689
R22955 DVSS.n6366 DVSS.n6365 1.49689
R22956 DVSS.n6371 DVSS.n6370 1.49689
R22957 DVSS.n6384 DVSS.n6383 1.49689
R22958 DVSS.n6389 DVSS.n6388 1.49689
R22959 DVSS.n2489 DVSS.n2488 1.49689
R22960 DVSS.n2498 DVSS.n2497 1.49689
R22961 DVSS.n2519 DVSS.n2518 1.49689
R22962 DVSS.n2528 DVSS.n2527 1.49689
R22963 DVSS.n6673 DVSS.n6672 1.49689
R22964 DVSS.n6678 DVSS.n6677 1.49689
R22965 DVSS.n6691 DVSS.n6690 1.49689
R22966 DVSS.n6696 DVSS.n6695 1.49689
R22967 DVSS.n6737 DVSS.n6736 1.49689
R22968 DVSS.n6742 DVSS.n6741 1.49689
R22969 DVSS.n6746 DVSS.n6745 1.49689
R22970 DVSS.n6751 DVSS.n6750 1.49689
R22971 DVSS.n6855 DVSS.n6852 1.49689
R22972 DVSS.n6860 DVSS.n6857 1.49689
R22973 DVSS.n6873 DVSS.n6870 1.49689
R22974 DVSS.n6878 DVSS.n6875 1.49689
R22975 DVSS.n1362 DVSS.n1361 1.49689
R22976 DVSS.n1357 DVSS.n1356 1.49689
R22977 DVSS.n6878 DVSS.n6877 1.49689
R22978 DVSS.n6873 DVSS.n6872 1.49689
R22979 DVSS.n6860 DVSS.n6859 1.49689
R22980 DVSS.n6855 DVSS.n6854 1.49689
R22981 DVSS.n6751 DVSS.n6748 1.49689
R22982 DVSS.n6746 DVSS.n6743 1.49689
R22983 DVSS.n6742 DVSS.n6739 1.49689
R22984 DVSS.n6737 DVSS.n6734 1.49689
R22985 DVSS.n6696 DVSS.n6693 1.49689
R22986 DVSS.n6691 DVSS.n6688 1.49689
R22987 DVSS.n6678 DVSS.n6675 1.49689
R22988 DVSS.n6673 DVSS.n6670 1.49689
R22989 DVSS.n2528 DVSS.n2524 1.49689
R22990 DVSS.n2519 DVSS.n2515 1.49689
R22991 DVSS.n2498 DVSS.n2494 1.49689
R22992 DVSS.n2489 DVSS.n2485 1.49689
R22993 DVSS.n6389 DVSS.n6386 1.49689
R22994 DVSS.n6384 DVSS.n6381 1.49689
R22995 DVSS.n6371 DVSS.n6368 1.49689
R22996 DVSS.n6366 DVSS.n6363 1.49689
R22997 DVSS.n4511 DVSS.n4508 1.49689
R22998 DVSS.n4506 DVSS.n4503 1.49689
R22999 DVSS.n4493 DVSS.n4490 1.49689
R23000 DVSS.n4488 DVSS.n4485 1.49689
R23001 DVSS.n4565 DVSS.n4562 1.49689
R23002 DVSS.n4560 DVSS.n4557 1.49689
R23003 DVSS.n4543 DVSS.n4540 1.49689
R23004 DVSS.n4538 DVSS.n4535 1.49689
R23005 DVSS.n5339 DVSS.n5336 1.49689
R23006 DVSS.n5344 DVSS.n5341 1.49689
R23007 DVSS.n4615 DVSS.n4612 1.49689
R23008 DVSS.n4610 DVSS.n4607 1.49689
R23009 DVSS.n4597 DVSS.n4594 1.49689
R23010 DVSS.n4592 DVSS.n4589 1.49689
R23011 DVSS.n1357 DVSS.n1354 1.49689
R23012 DVSS.n1362 DVSS.n1359 1.49689
R23013 DVSS.n13420 DVSS.n13419 1.49675
R23014 DVSS.n13517 DVSS.n13503 1.49675
R23015 DVSS.n18875 DVSS.n18874 1.49675
R23016 DVSS.n7215 DVSS.n7214 1.49675
R23017 DVSS.n20967 DVSS.n20952 1.49632
R23018 DVSS.n10942 DVSS.n10192 1.49617
R23019 DVSS.n4974 DVSS.n4719 1.49617
R23020 DVSS.n20965 DVSS.n20964 1.49613
R23021 DVSS.n14527 DVSS.n14521 1.49592
R23022 DVSS.n14618 DVSS.n14599 1.49581
R23023 DVSS.n5538 DVSS.n5537 1.49526
R23024 DVSS.n5540 DVSS.n5539 1.49526
R23025 DVSS.n17112 DVSS.n17111 1.49526
R23026 DVSS.n16874 DVSS.n16873 1.49526
R23027 DVSS.n16877 DVSS.n16876 1.49526
R23028 DVSS.n16885 DVSS.n16884 1.49526
R23029 DVSS.n10008 DVSS.n10007 1.49526
R23030 DVSS.n10049 DVSS.n10048 1.49526
R23031 DVSS.n4017 DVSS.n4016 1.49526
R23032 DVSS.n4022 DVSS.n4021 1.49526
R23033 DVSS.n4027 DVSS.n4026 1.49526
R23034 DVSS.n7485 DVSS.n7484 1.49526
R23035 DVSS.n7453 DVSS.n7452 1.49526
R23036 DVSS.n4109 DVSS.n4108 1.49526
R23037 DVSS.n4104 DVSS.n4103 1.49526
R23038 DVSS.n4099 DVSS.n4098 1.49526
R23039 DVSS.n4361 DVSS.n4360 1.49526
R23040 DVSS.n4366 DVSS.n4365 1.49526
R23041 DVSS.n4371 DVSS.n4370 1.49526
R23042 DVSS.n6550 DVSS.n6549 1.49526
R23043 DVSS.n6545 DVSS.n6544 1.49526
R23044 DVSS.n6540 DVSS.n6539 1.49526
R23045 DVSS.n6414 DVSS.n6413 1.49526
R23046 DVSS.n6409 DVSS.n6408 1.49526
R23047 DVSS.n4476 DVSS.n4475 1.49526
R23048 DVSS.n5805 DVSS.n5804 1.49526
R23049 DVSS.n5815 DVSS.n5814 1.49526
R23050 DVSS.n5820 DVSS.n5819 1.49526
R23051 DVSS.n6488 DVSS.n6487 1.49526
R23052 DVSS.n6490 DVSS.n6489 1.49526
R23053 DVSS.n6492 DVSS.n6491 1.49526
R23054 DVSS.n8942 DVSS.n8941 1.49526
R23055 DVSS.n8944 DVSS.n8943 1.49526
R23056 DVSS.n8946 DVSS.n8945 1.49526
R23057 DVSS.n9733 DVSS.n9732 1.49526
R23058 DVSS.n9738 DVSS.n9737 1.49526
R23059 DVSS.n9743 DVSS.n9742 1.49526
R23060 DVSS.n8975 DVSS.n8974 1.49526
R23061 DVSS.n8977 DVSS.n8976 1.49526
R23062 DVSS.n8979 DVSS.n8978 1.49526
R23063 DVSS.n9121 DVSS.n9120 1.49526
R23064 DVSS.n9126 DVSS.n9125 1.49526
R23065 DVSS.n9131 DVSS.n9130 1.49526
R23066 DVSS.n11169 DVSS.n11168 1.49526
R23067 DVSS.n11213 DVSS.n11212 1.49526
R23068 DVSS.n11174 DVSS.n11173 1.49526
R23069 DVSS.n11038 DVSS.n11037 1.49526
R23070 DVSS.n11043 DVSS.n11042 1.49526
R23071 DVSS.n11051 DVSS.n11050 1.49526
R23072 DVSS.n16275 DVSS.n16274 1.49526
R23073 DVSS.n7624 DVSS.n7623 1.49526
R23074 DVSS.n16236 DVSS.n16235 1.49526
R23075 DVSS.n7616 DVSS.n7615 1.49526
R23076 DVSS.n7564 DVSS.n7563 1.49526
R23077 DVSS.n7610 DVSS.n7609 1.49526
R23078 DVSS.n18405 DVSS.n18404 1.49526
R23079 DVSS.n18410 DVSS.n18409 1.49526
R23080 DVSS.n16335 DVSS.n16334 1.49526
R23081 DVSS.n7629 DVSS.n7628 1.49526
R23082 DVSS.n15836 DVSS.n15835 1.49526
R23083 DVSS.n15841 DVSS.n15840 1.49526
R23084 DVSS.n15846 DVSS.n15845 1.49526
R23085 DVSS.n7683 DVSS.n7682 1.49526
R23086 DVSS.n7685 DVSS.n7684 1.49526
R23087 DVSS.n7687 DVSS.n7686 1.49526
R23088 DVSS.n15590 DVSS.n15589 1.49526
R23089 DVSS.n15595 DVSS.n15594 1.49526
R23090 DVSS.n15600 DVSS.n15599 1.49526
R23091 DVSS.n14961 DVSS.n14960 1.49526
R23092 DVSS.n14966 DVSS.n14965 1.49526
R23093 DVSS.n14971 DVSS.n14970 1.49526
R23094 DVSS.n17658 DVSS.n17657 1.49526
R23095 DVSS.n7657 DVSS.n7656 1.49526
R23096 DVSS.n7659 DVSS.n7658 1.49526
R23097 DVSS.n16896 DVSS.n16895 1.49526
R23098 DVSS.n16901 DVSS.n16900 1.49526
R23099 DVSS.n17551 DVSS.n17550 1.49526
R23100 DVSS.n7667 DVSS.n7666 1.49526
R23101 DVSS.n7672 DVSS.n7671 1.49526
R23102 DVSS.n7675 DVSS.n7674 1.49526
R23103 DVSS.n7680 DVSS.n7679 1.49526
R23104 DVSS.n7696 DVSS.n7695 1.49526
R23105 DVSS.n7701 DVSS.n7700 1.49526
R23106 DVSS.n7706 DVSS.n7705 1.49526
R23107 DVSS.n7708 DVSS.n7707 1.49526
R23108 DVSS.n17674 DVSS.n17673 1.49526
R23109 DVSS.n7648 DVSS.n7647 1.49526
R23110 DVSS.n7767 DVSS.n7766 1.49526
R23111 DVSS.n7769 DVSS.n7768 1.49526
R23112 DVSS.n7772 DVSS.n7771 1.49526
R23113 DVSS.n7774 DVSS.n7773 1.49526
R23114 DVSS.n7776 DVSS.n7775 1.49526
R23115 DVSS.n9024 DVSS.n9023 1.49526
R23116 DVSS.n8051 DVSS.n8050 1.49526
R23117 DVSS.n8053 DVSS.n8052 1.49526
R23118 DVSS.n5542 DVSS.n5541 1.49526
R23119 DVSS.n17240 DVSS.n17239 1.49526
R23120 DVSS.n5529 DVSS.n5528 1.49526
R23121 DVSS.n5524 DVSS.n5523 1.49526
R23122 DVSS.n5519 DVSS.n5518 1.49526
R23123 DVSS.n6404 DVSS.n6403 1.49526
R23124 DVSS.n2543 DVSS.n2542 1.49526
R23125 DVSS.n6478 DVSS.n6477 1.49526
R23126 DVSS.n5829 DVSS.n5828 1.49526
R23127 DVSS.n2548 DVSS.n2547 1.49526
R23128 DVSS.n2553 DVSS.n2552 1.49526
R23129 DVSS.n2558 DVSS.n2557 1.49526
R23130 DVSS.n2561 DVSS.n2560 1.49526
R23131 DVSS.n2566 DVSS.n2565 1.49526
R23132 DVSS.n2571 DVSS.n2570 1.49526
R23133 DVSS.n2576 DVSS.n2575 1.49526
R23134 DVSS.n4003 DVSS.n4002 1.49526
R23135 DVSS.n4008 DVSS.n4007 1.49526
R23136 DVSS.n8932 DVSS.n8931 1.49526
R23137 DVSS.n8937 DVSS.n8936 1.49526
R23138 DVSS.n8939 DVSS.n8938 1.49526
R23139 DVSS.n8957 DVSS.n8956 1.49526
R23140 DVSS.n9719 DVSS.n9718 1.49526
R23141 DVSS.n9724 DVSS.n9723 1.49526
R23142 DVSS.n8965 DVSS.n8964 1.49526
R23143 DVSS.n8970 DVSS.n8969 1.49526
R23144 DVSS.n8972 DVSS.n8971 1.49526
R23145 DVSS.n9007 DVSS.n9006 1.49526
R23146 DVSS.n9107 DVSS.n9106 1.49526
R23147 DVSS.n9112 DVSS.n9111 1.49526
R23148 DVSS.n9017 DVSS.n9016 1.49526
R23149 DVSS.n9019 DVSS.n9018 1.49526
R23150 DVSS.n9021 DVSS.n9020 1.49526
R23151 DVSS.n9818 DVSS.n9817 1.49526
R23152 DVSS.n9823 DVSS.n9822 1.49526
R23153 DVSS.n9825 DVSS.n9824 1.49526
R23154 DVSS.n11060 DVSS.n11059 1.49526
R23155 DVSS.n11065 DVSS.n11064 1.49526
R23156 DVSS.n11074 DVSS.n11073 1.49526
R23157 DVSS.n9995 DVSS.n9994 1.49526
R23158 DVSS.n9860 DVSS.n9859 1.49526
R23159 DVSS.n9855 DVSS.n9854 1.49526
R23160 DVSS.n16265 DVSS.n16264 1.49526
R23161 DVSS.n16270 DVSS.n16269 1.49526
R23162 DVSS.n16272 DVSS.n16271 1.49526
R23163 DVSS.n16226 DVSS.n16225 1.49526
R23164 DVSS.n16231 DVSS.n16230 1.49526
R23165 DVSS.n16233 DVSS.n16232 1.49526
R23166 DVSS.n7554 DVSS.n7553 1.49526
R23167 DVSS.n7559 DVSS.n7558 1.49526
R23168 DVSS.n7561 DVSS.n7560 1.49526
R23169 DVSS.n7465 DVSS.n7464 1.49526
R23170 DVSS.n18391 DVSS.n18390 1.49526
R23171 DVSS.n18396 DVSS.n18395 1.49526
R23172 DVSS.n7475 DVSS.n7474 1.49526
R23173 DVSS.n7480 DVSS.n7479 1.49526
R23174 DVSS.n7482 DVSS.n7481 1.49526
R23175 DVSS.n16434 DVSS.n16433 1.49526
R23176 DVSS.n16439 DVSS.n16438 1.49526
R23177 DVSS.n16123 DVSS.n16122 1.49526
R23178 DVSS.n17442 DVSS.n17441 1.49526
R23179 DVSS.n17437 DVSS.n17436 1.49526
R23180 DVSS.n16321 DVSS.n16320 1.49526
R23181 DVSS.n16316 DVSS.n16315 1.49526
R23182 DVSS.n2460 DVSS.n2459 1.47742
R23183 DVSS.n17531 DVSS.n17530 1.47233
R23184 DVSS.n17677 DVSS.n17676 1.47233
R23185 DVSS.n15260 DVSS.n15259 1.47233
R23186 DVSS.n18358 DVSS.n18357 1.47233
R23187 DVSS.n18079 DVSS.n18078 1.47233
R23188 DVSS.n17938 DVSS.n17937 1.47233
R23189 DVSS.n16966 DVSS.n16965 1.4635
R23190 DVSS.n14904 DVSS.n14903 1.4635
R23191 DVSS.n5604 DVSS.n5603 1.36071
R23192 DVSS.n5584 DVSS.n5583 1.36071
R23193 DVSS.n5599 DVSS.n5598 1.36071
R23194 DVSS.n5575 DVSS.n5574 1.36071
R23195 DVSS.n10248 DVSS.n10247 1.36071
R23196 DVSS.n10255 DVSS.n10254 1.36071
R23197 DVSS.n10280 DVSS.n10279 1.36071
R23198 DVSS.n10287 DVSS.n10286 1.36071
R23199 DVSS.n17280 DVSS.n17279 1.36071
R23200 DVSS.n17282 DVSS.n17281 1.36071
R23201 DVSS.n17284 DVSS.n17283 1.36071
R23202 DVSS.n16996 DVSS.n16995 1.36071
R23203 DVSS.n17003 DVSS.n17002 1.36071
R23204 DVSS.n17019 DVSS.n17018 1.36071
R23205 DVSS.n17026 DVSS.n17025 1.36071
R23206 DVSS.n16973 DVSS.n16972 1.36071
R23207 DVSS.n16979 DVSS.n16978 1.36071
R23208 DVSS.n16984 DVSS.n16983 1.36071
R23209 DVSS.n11460 DVSS.n11459 1.36071
R23210 DVSS.n11497 DVSS.n11496 1.36071
R23211 DVSS.n11622 DVSS.n11621 1.36071
R23212 DVSS.n11659 DVSS.n11658 1.36071
R23213 DVSS.n11200 DVSS.n11199 1.36071
R23214 DVSS.n10259 DVSS.n10258 1.36071
R23215 DVSS.n11004 DVSS.n11003 1.36071
R23216 DVSS.n10011 DVSS.n10010 1.36071
R23217 DVSS.n5354 DVSS.n5353 1.36071
R23218 DVSS.n5356 DVSS.n5355 1.36071
R23219 DVSS.n5358 DVSS.n5357 1.36071
R23220 DVSS.n5360 DVSS.n5359 1.36071
R23221 DVSS.n10216 DVSS.n10215 1.36071
R23222 DVSS.n10223 DVSS.n10222 1.36071
R23223 DVSS.n10229 DVSS.n10228 1.36071
R23224 DVSS.n10235 DVSS.n10234 1.36071
R23225 DVSS.n17272 DVSS.n17271 1.36071
R23226 DVSS.n17269 DVSS.n17268 1.36071
R23227 DVSS.n17317 DVSS.n17316 1.36071
R23228 DVSS.n6906 DVSS.n6905 1.36071
R23229 DVSS.n6911 DVSS.n6910 1.36071
R23230 DVSS.n6916 DVSS.n6915 1.36071
R23231 DVSS.n6921 DVSS.n6920 1.36071
R23232 DVSS.n6930 DVSS.n6929 1.36071
R23233 DVSS.n6935 DVSS.n6934 1.36071
R23234 DVSS.n6940 DVSS.n6939 1.36071
R23235 DVSS.n6949 DVSS.n6948 1.36071
R23236 DVSS.n7440 DVSS.n7439 1.36071
R23237 DVSS.n7445 DVSS.n7444 1.36071
R23238 DVSS.n18570 DVSS.n18569 1.36071
R23239 DVSS.n18565 DVSS.n18564 1.36071
R23240 DVSS.n14885 DVSS.n14884 1.36071
R23241 DVSS.n14919 DVSS.n14918 1.36071
R23242 DVSS.n14924 DVSS.n14923 1.36071
R23243 DVSS.n14933 DVSS.n14932 1.36071
R23244 DVSS.n14938 DVSS.n14937 1.36071
R23245 DVSS.n14951 DVSS.n14950 1.36071
R23246 DVSS.n14946 DVSS.n14945 1.36071
R23247 DVSS.n8012 DVSS.n8011 1.36071
R23248 DVSS.n8017 DVSS.n8016 1.36071
R23249 DVSS.n13178 DVSS.n13177 1.36071
R23250 DVSS.n13173 DVSS.n13172 1.36071
R23251 DVSS.n13164 DVSS.n13163 1.36071
R23252 DVSS.n13159 DVSS.n13158 1.36071
R23253 DVSS.n13154 DVSS.n13153 1.36071
R23254 DVSS.n8045 DVSS.n8044 1.36071
R23255 DVSS.n7386 DVSS.n7385 1.35477
R23256 DVSS.n13769 DVSS.n13768 1.35477
R23257 DVSS.n1319 DVSS.n1318 1.35477
R23258 DVSS.n13332 DVSS.n13331 1.35477
R23259 DVSS.n12948 DVSS.n12947 1.30851
R23260 DVSS.n13044 DVSS.n13043 1.30851
R23261 DVSS.n3781 DVSS.n3780 1.30851
R23262 DVSS.n3580 DVSS.n3579 1.30851
R23263 DVSS.n20516 DVSS.n20515 1.3005
R23264 DVSS.n20515 DVSS.n20514 1.3005
R23265 DVSS.n20506 DVSS.n20505 1.3005
R23266 DVSS.n20505 DVSS.n20504 1.3005
R23267 DVSS.n20244 DVSS.n20243 1.3005
R23268 DVSS.n20243 DVSS.n20242 1.3005
R23269 DVSS.n20230 DVSS.n20229 1.3005
R23270 DVSS.n20229 DVSS.n20228 1.3005
R23271 DVSS.n19959 DVSS.n19958 1.3005
R23272 DVSS.n19958 DVSS.n19957 1.3005
R23273 DVSS.n19734 DVSS.n19733 1.3005
R23274 DVSS.n19733 DVSS.n19732 1.3005
R23275 DVSS.n19495 DVSS.n19494 1.3005
R23276 DVSS.n19494 DVSS.n19493 1.3005
R23277 DVSS.n19505 DVSS.n19504 1.3005
R23278 DVSS.n19504 DVSS.n19503 1.3005
R23279 DVSS.n19234 DVSS.n19233 1.3005
R23280 DVSS.n19233 DVSS.n19232 1.3005
R23281 DVSS.n19220 DVSS.n19219 1.3005
R23282 DVSS.n19219 DVSS.n19218 1.3005
R23283 DVSS.n19226 DVSS.n19225 1.3005
R23284 DVSS.n19225 DVSS.n19224 1.3005
R23285 DVSS.n19485 DVSS.n19484 1.3005
R23286 DVSS.n19484 DVSS.n19483 1.3005
R23287 DVSS.n19499 DVSS.n19498 1.3005
R23288 DVSS.n19498 DVSS.n19497 1.3005
R23289 DVSS.n19729 DVSS.n19728 1.3005
R23290 DVSS.n19728 DVSS.n19727 1.3005
R23291 DVSS.n19738 DVSS.n19737 1.3005
R23292 DVSS.n19737 DVSS.n19736 1.3005
R23293 DVSS.n19963 DVSS.n19962 1.3005
R23294 DVSS.n19962 DVSS.n19961 1.3005
R23295 DVSS.n20224 DVSS.n20223 1.3005
R23296 DVSS.n20223 DVSS.n20222 1.3005
R23297 DVSS.n20236 DVSS.n20235 1.3005
R23298 DVSS.n20235 DVSS.n20234 1.3005
R23299 DVSS.n20495 DVSS.n20494 1.3005
R23300 DVSS.n20494 DVSS.n20493 1.3005
R23301 DVSS.n20510 DVSS.n20509 1.3005
R23302 DVSS.n20509 DVSS.n20508 1.3005
R23303 DVSS.n20500 DVSS.n20499 1.3005
R23304 DVSS.n20499 DVSS.n20498 1.3005
R23305 DVSS.n19214 DVSS.n19213 1.3005
R23306 DVSS.n19213 DVSS.n19212 1.3005
R23307 DVSS.n952 DVSS.n951 1.3005
R23308 DVSS.n951 DVSS.n950 1.3005
R23309 DVSS.n365 DVSS.n364 1.3005
R23310 DVSS.n364 DVSS.n363 1.3005
R23311 DVSS.n20961 DVSS.n20960 1.3005
R23312 DVSS.n20960 DVSS.n20959 1.3005
R23313 DVSS.n1189 DVSS.n1188 1.3005
R23314 DVSS.n1188 DVSS.n1187 1.3005
R23315 DVSS.n332 DVSS.n331 1.3005
R23316 DVSS.n331 DVSS.n330 1.3005
R23317 DVSS.n20733 DVSS.n20732 1.3005
R23318 DVSS.n20732 DVSS.n20731 1.3005
R23319 DVSS.n20945 DVSS.n20944 1.3005
R23320 DVSS.n20944 DVSS.n20943 1.3005
R23321 DVSS.n20940 DVSS.n20939 1.3005
R23322 DVSS.n20939 DVSS.n20938 1.3005
R23323 DVSS.n20949 DVSS.n20948 1.3005
R23324 DVSS.n20948 DVSS.n20947 1.3005
R23325 DVSS.n20716 DVSS.n20715 1.3005
R23326 DVSS.n20715 DVSS.n20714 1.3005
R23327 DVSS.n20711 DVSS.n20710 1.3005
R23328 DVSS.n20710 DVSS.n20709 1.3005
R23329 DVSS.n20720 DVSS.n20719 1.3005
R23330 DVSS.n20719 DVSS.n20718 1.3005
R23331 DVSS.n20727 DVSS.n20726 1.3005
R23332 DVSS.n20726 DVSS.n20725 1.3005
R23333 DVSS.n371 DVSS.n370 1.3005
R23334 DVSS.n370 DVSS.n369 1.3005
R23335 DVSS.n338 DVSS.n337 1.3005
R23336 DVSS.n337 DVSS.n336 1.3005
R23337 DVSS.n1168 DVSS.n1167 1.3005
R23338 DVSS.n1167 DVSS.n1166 1.3005
R23339 DVSS.n1178 DVSS.n1177 1.3005
R23340 DVSS.n1177 DVSS.n1176 1.3005
R23341 DVSS.n1172 DVSS.n1171 1.3005
R23342 DVSS.n1171 DVSS.n1170 1.3005
R23343 DVSS.n1186 DVSS.n1185 1.3005
R23344 DVSS.n1185 DVSS.n1184 1.3005
R23345 DVSS.n970 DVSS.n969 1.3005
R23346 DVSS.n969 DVSS.n968 1.3005
R23347 DVSS.n964 DVSS.n963 1.3005
R23348 DVSS.n963 DVSS.n962 1.3005
R23349 DVSS.n958 DVSS.n957 1.3005
R23350 DVSS.n957 DVSS.n956 1.3005
R23351 DVSS.n7365 DVSS.n7363 1.24924
R23352 DVSS.n7390 DVSS.n7389 1.24924
R23353 DVSS.n7411 DVSS.n7410 1.24924
R23354 DVSS.n7159 DVSS.n7158 1.24924
R23355 DVSS.n1330 DVSS.n1328 1.24924
R23356 DVSS.n7027 DVSS.n7026 1.24924
R23357 DVSS.n13735 DVSS.n13733 1.23166
R23358 DVSS.n13773 DVSS.n13772 1.23166
R23359 DVSS.n13813 DVSS.n13812 1.23166
R23360 DVSS.n7969 DVSS.n7968 1.23166
R23361 DVSS.n13343 DVSS.n13341 1.23166
R23362 DVSS.n13324 DVSS.n13323 1.23166
R23363 DVSS.n6959 DVSS.n6958 1.17298
R23364 DVSS.n13188 DVSS.n13187 1.17298
R23365 DVSS.n21160 DVSS.n21151 1.14278
R23366 DVSS.n947 DVSS.n946 1.13013
R23367 DVSS.n13975 DVSS.n13974 1.1255
R23368 DVSS.n14916 DVSS.n14915 1.1255
R23369 DVSS.n19223 DVSS.n19222 1.1255
R23370 DVSS.n19222 DVSS.n19221 1.1255
R23371 DVSS.n19235 DVSS.n19228 1.1255
R23372 DVSS.n19228 DVSS.n19227 1.1255
R23373 DVSS.n19231 DVSS.n19230 1.1255
R23374 DVSS.n19230 DVSS.n19229 1.1255
R23375 DVSS.n19741 DVSS.n19740 1.1255
R23376 DVSS.n19740 DVSS.n19739 1.1255
R23377 DVSS.n19735 DVSS.n19731 1.1255
R23378 DVSS.n19731 DVSS.n19730 1.1255
R23379 DVSS.n19948 DVSS.n19947 1.1255
R23380 DVSS.n19947 DVSS.n19946 1.1255
R23381 DVSS.n19966 DVSS.n19965 1.1255
R23382 DVSS.n19965 DVSS.n19964 1.1255
R23383 DVSS.n19960 DVSS.n19953 1.1255
R23384 DVSS.n19953 DVSS.n19952 1.1255
R23385 DVSS.n19956 DVSS.n19955 1.1255
R23386 DVSS.n19955 DVSS.n19954 1.1255
R23387 DVSS.n20227 DVSS.n20226 1.1255
R23388 DVSS.n20226 DVSS.n20225 1.1255
R23389 DVSS.n20233 DVSS.n20232 1.1255
R23390 DVSS.n20232 DVSS.n20231 1.1255
R23391 DVSS.n20245 DVSS.n20238 1.1255
R23392 DVSS.n20238 DVSS.n20237 1.1255
R23393 DVSS.n20241 DVSS.n20240 1.1255
R23394 DVSS.n20240 DVSS.n20239 1.1255
R23395 DVSS.n19217 DVSS.n19216 1.1255
R23396 DVSS.n19216 DVSS.n19215 1.1255
R23397 DVSS.n20519 DVSS.n20518 1.1255
R23398 DVSS.n20518 DVSS.n20517 1.1255
R23399 DVSS.n20513 DVSS.n20512 1.1255
R23400 DVSS.n20512 DVSS.n20511 1.1255
R23401 DVSS.n20507 DVSS.n20497 1.1255
R23402 DVSS.n20497 DVSS.n20496 1.1255
R23403 DVSS.n20503 DVSS.n20502 1.1255
R23404 DVSS.n20502 DVSS.n20501 1.1255
R23405 DVSS.n20952 DVSS.n20951 1.1255
R23406 DVSS.n20951 DVSS.n20950 1.1255
R23407 DVSS.n20946 DVSS.n20942 1.1255
R23408 DVSS.n20942 DVSS.n20941 1.1255
R23409 DVSS.n20958 DVSS.n20957 1.1255
R23410 DVSS.n20957 DVSS.n20956 1.1255
R23411 DVSS.n20736 DVSS.n20735 1.1255
R23412 DVSS.n20735 DVSS.n20734 1.1255
R23413 DVSS.n20723 DVSS.n20722 1.1255
R23414 DVSS.n20722 DVSS.n20721 1.1255
R23415 DVSS.n20717 DVSS.n20713 1.1255
R23416 DVSS.n20713 DVSS.n20712 1.1255
R23417 DVSS.n20730 DVSS.n20729 1.1255
R23418 DVSS.n20729 DVSS.n20728 1.1255
R23419 DVSS.n368 DVSS.n367 1.1255
R23420 DVSS.n367 DVSS.n366 1.1255
R23421 DVSS.n374 DVSS.n373 1.1255
R23422 DVSS.n373 DVSS.n372 1.1255
R23423 DVSS.n362 DVSS.n361 1.1255
R23424 DVSS.n361 DVSS.n360 1.1255
R23425 DVSS.n335 DVSS.n334 1.1255
R23426 DVSS.n334 DVSS.n333 1.1255
R23427 DVSS.n341 DVSS.n340 1.1255
R23428 DVSS.n340 DVSS.n339 1.1255
R23429 DVSS.n329 DVSS.n328 1.1255
R23430 DVSS.n328 DVSS.n327 1.1255
R23431 DVSS.n967 DVSS.n966 1.1255
R23432 DVSS.n966 DVSS.n965 1.1255
R23433 DVSS.n973 DVSS.n972 1.1255
R23434 DVSS.n972 DVSS.n971 1.1255
R23435 DVSS.n961 DVSS.n960 1.1255
R23436 DVSS.n960 DVSS.n959 1.1255
R23437 DVSS.n955 DVSS.n954 1.1255
R23438 DVSS.n954 DVSS.n953 1.1255
R23439 DVSS.n20964 DVSS.n20963 1.1255
R23440 DVSS.n20963 DVSS.n20962 1.1255
R23441 DVSS.n1192 DVSS.n1191 1.1255
R23442 DVSS.n19506 DVSS.n19487 1.1255
R23443 DVSS.n19487 DVSS.n19486 1.1255
R23444 DVSS.n19502 DVSS.n19501 1.1255
R23445 DVSS.n19501 DVSS.n19500 1.1255
R23446 DVSS.n19496 DVSS.n19489 1.1255
R23447 DVSS.n19489 DVSS.n19488 1.1255
R23448 DVSS.n19492 DVSS.n19491 1.1255
R23449 DVSS.n19491 DVSS.n19490 1.1255
R23450 DVSS.n1181 DVSS.n1180 1.1255
R23451 DVSS.n1180 DVSS.n1179 1.1255
R23452 DVSS.n1175 DVSS.n1174 1.1255
R23453 DVSS.n1174 DVSS.n1173 1.1255
R23454 DVSS.n1169 DVSS.n1165 1.1255
R23455 DVSS.n1165 DVSS.n1164 1.1255
R23456 DVSS.n1191 DVSS.n1190 1.1255
R23457 DVSS.n14953 DVSS.n14952 1.12142
R23458 DVSS.n13155 DVSS.n13152 1.12142
R23459 DVSS.n13180 DVSS.n13179 1.12142
R23460 DVSS.n18572 DVSS.n18571 1.12142
R23461 DVSS.n6951 DVSS.n6950 1.12142
R23462 DVSS.n6436 DVSS.n6435 1.12124
R23463 DVSS.n6572 DVSS.n6571 1.12124
R23464 DVSS.n6715 DVSS.n6714 1.12124
R23465 DVSS.n6770 DVSS.n6769 1.12124
R23466 DVSS.n6897 DVSS.n6896 1.12124
R23467 DVSS.n6901 DVSS.n6900 1.12124
R23468 DVSS.n6522 DVSS.n4477 1.12072
R23469 DVSS.n9781 DVSS.n9780 1.12072
R23470 DVSS.n9751 DVSS.n9750 1.12072
R23471 DVSS.n9589 DVSS.n9588 1.12072
R23472 DVSS.n9139 DVSS.n9138 1.12072
R23473 DVSS.n13115 DVSS.n13114 1.12072
R23474 DVSS.n9502 DVSS.n9488 1.12072
R23475 DVSS.n11299 DVSS.n11298 1.12072
R23476 DVSS.n12967 DVSS.n12966 1.12072
R23477 DVSS.n10901 DVSS.n10900 1.12072
R23478 DVSS.n11257 DVSS.n8925 1.12072
R23479 DVSS.n15854 DVSS.n15853 1.12072
R23480 DVSS.n15721 DVSS.n15720 1.12072
R23481 DVSS.n15608 DVSS.n15607 1.12072
R23482 DVSS.n14990 DVSS.n14978 1.12072
R23483 DVSS.n13086 DVSS.n13085 1.12072
R23484 DVSS.n11540 DVSS.n8323 1.12072
R23485 DVSS.n11363 DVSS.n11362 1.12072
R23486 DVSS.n13025 DVSS.n13024 1.12072
R23487 DVSS.n10883 DVSS.n10860 1.12072
R23488 DVSS.n10819 DVSS.n10733 1.12072
R23489 DVSS.n11404 DVSS.n8336 1.12072
R23490 DVSS.n4033 DVSS.n4032 1.12072
R23491 DVSS.n15045 DVSS.n15044 1.12072
R23492 DVSS.n13149 DVSS.n8059 1.12072
R23493 DVSS.n5236 DVSS.n5235 1.12072
R23494 DVSS.n4353 DVSS.n4352 1.12072
R23495 DVSS.n4117 DVSS.n4116 1.12072
R23496 DVSS.n4004 DVSS.n4001 1.12072
R23497 DVSS.n3764 DVSS.n2756 1.12072
R23498 DVSS.n3969 DVSS.n3968 1.12072
R23499 DVSS.n4273 DVSS.n4259 1.12072
R23500 DVSS.n19236 DVSS.n19235 1.12072
R23501 DVSS.n20246 DVSS.n20245 1.12072
R23502 DVSS.n9797 DVSS.n9796 1.12072
R23503 DVSS.n9720 DVSS.n9717 1.12072
R23504 DVSS.n9605 DVSS.n9604 1.12072
R23505 DVSS.n9108 DVSS.n9105 1.12072
R23506 DVSS.n9040 DVSS.n9039 1.12072
R23507 DVSS.n977 DVSS.n973 1.12072
R23508 DVSS.n20737 DVSS.n20736 1.12072
R23509 DVSS.n20739 DVSS.n20723 1.12072
R23510 DVSS.n1182 DVSS.n1181 1.12072
R23511 DVSS.n16286 DVSS.n16285 1.12072
R23512 DVSS.n16247 DVSS.n16246 1.12072
R23513 DVSS.n18376 DVSS.n18375 1.12072
R23514 DVSS.n18392 DVSS.n18389 1.12072
R23515 DVSS.n7498 DVSS.n7497 1.12072
R23516 DVSS.n19507 DVSS.n19506 1.12072
R23517 DVSS.n5444 DVSS.n5058 1.12072
R23518 DVSS.n6050 DVSS.n6049 1.12072
R23519 DVSS.n6327 DVSS.n6326 1.12072
R23520 DVSS.n3626 DVSS.n3625 1.12072
R23521 DVSS.n6587 DVSS.n1401 1.12072
R23522 DVSS.n6817 DVSS.n6816 1.12072
R23523 DVSS.n5407 DVSS.n5311 1.12072
R23524 DVSS.n12092 DVSS.n12091 1.12072
R23525 DVSS.n12906 DVSS.n12136 1.12072
R23526 DVSS.n3661 DVSS.n3660 1.12072
R23527 DVSS.n3730 DVSS.n3729 1.12072
R23528 DVSS.n19020 DVSS.n19019 1.12072
R23529 DVSS.n19572 DVSS.n19571 1.12072
R23530 DVSS.n21557 DVSS.n21555 1.12072
R23531 DVSS.n20317 DVSS.n20316 1.12072
R23532 DVSS.n20591 DVSS.n20590 1.12072
R23533 DVSS.n19301 DVSS.n19300 1.12072
R23534 DVSS.n622 DVSS.n621 1.12072
R23535 DVSS.n1271 DVSS.n1270 1.12072
R23536 DVSS.n21467 DVSS.n21392 1.12072
R23537 DVSS.n1056 DVSS.n1055 1.12072
R23538 DVSS.n21088 DVSS.n21087 1.12072
R23539 DVSS.n20862 DVSS.n20861 1.12072
R23540 DVSS.n6536 DVSS.n6535 1.12053
R23541 DVSS.n4377 DVSS.n4376 1.12053
R23542 DVSS.n4095 DVSS.n4094 1.12053
R23543 DVSS.n20520 DVSS.n20519 1.12053
R23544 DVSS.n1193 DVSS.n1192 1.12053
R23545 DVSS.n18561 DVSS.n18559 1.12051
R23546 DVSS.n14920 DVSS.n14917 1.12051
R23547 DVSS.n17944 DVSS.n17943 1.11968
R23548 DVSS.n18085 DVSS.n18084 1.11968
R23549 DVSS.n18363 DVSS.n7608 1.11968
R23550 DVSS.n18416 DVSS.n18415 1.11968
R23551 DVSS.n15828 DVSS.n15827 1.11968
R23552 DVSS.n15734 DVSS.n15733 1.11968
R23553 DVSS.n15582 DVSS.n15581 1.11968
R23554 DVSS.n15246 DVSS.n15245 1.11968
R23555 DVSS.n18524 DVSS.n7458 1.11968
R23556 DVSS.n15057 DVSS.n7765 1.11968
R23557 DVSS.n19742 DVSS.n19741 1.11968
R23558 DVSS.n19967 DVSS.n19966 1.11968
R23559 DVSS.n378 DVSS.n374 1.11968
R23560 DVSS.n19812 DVSS.n19811 1.11968
R23561 DVSS.n20037 DVSS.n20036 1.11968
R23562 DVSS.n253 DVSS.n252 1.11968
R23563 DVSS.n461 DVSS.n460 1.11968
R23564 DVSS.n2353 DVSS.n2336 1.11241
R23565 DVSS.n2413 DVSS.n2412 1.11241
R23566 DVSS.n6430 DVSS.n6425 1.11241
R23567 DVSS.n6430 DVSS.n6429 1.11241
R23568 DVSS.n6566 DVSS.n6561 1.11241
R23569 DVSS.n6566 DVSS.n6565 1.11241
R23570 DVSS.n6271 DVSS.n6269 1.11241
R23571 DVSS.n6271 DVSS.n6270 1.11241
R23572 DVSS.n6264 DVSS.n6144 1.11241
R23573 DVSS.n6022 DVSS.n6007 1.11241
R23574 DVSS.n6026 DVSS.n5913 1.11241
R23575 DVSS.n6022 DVSS.n6021 1.11241
R23576 DVSS.n6022 DVSS.n5914 1.11241
R23577 DVSS.n6026 DVSS.n6025 1.11241
R23578 DVSS.n6026 DVSS.n5912 1.11241
R23579 DVSS.n6264 DVSS.n6145 1.11241
R23580 DVSS.n6264 DVSS.n6142 1.11241
R23581 DVSS.n1727 DVSS.n1726 1.10465
R23582 DVSS.n21160 DVSS.n21158 1.05973
R23583 DVSS.n925 DVSS.n918 1.05973
R23584 DVSS.n925 DVSS.n915 1.05973
R23585 DVSS.n939 DVSS.n936 1.05973
R23586 DVSS.n21179 DVSS.n21177 1.05973
R23587 DVSS.n21179 DVSS.n21176 1.05973
R23588 DVSS.n11683 DVSS.n11682 0.897595
R23589 DVSS.n11646 DVSS.n11645 0.897595
R23590 DVSS.n11521 DVSS.n11520 0.897595
R23591 DVSS.n11484 DVSS.n11483 0.897595
R23592 DVSS.n13057 DVSS.n11731 0.897595
R23593 DVSS.n14906 DVSS.n14905 0.87334
R23594 DVSS.t3 DVSS.n14189 0.867167
R23595 DVSS.n14047 DVSS.n14046 0.867167
R23596 DVSS.n19892 DVSS.n19891 0.867167
R23597 DVSS.t37 DVSS.n14676 0.867167
R23598 DVSS.n12805 DVSS.n12803 0.771929
R23599 DVSS.n12807 DVSS.n12805 0.771929
R23600 DVSS.n12809 DVSS.n12807 0.771929
R23601 DVSS.n12811 DVSS.n12809 0.771929
R23602 DVSS.n12815 DVSS.n12811 0.771929
R23603 DVSS.n12815 DVSS.n12813 0.771929
R23604 DVSS.n12770 DVSS.n12768 0.771929
R23605 DVSS.n12142 DVSS.n12140 0.771929
R23606 DVSS.n12150 DVSS.n12148 0.771929
R23607 DVSS.n12741 DVSS.n12739 0.771929
R23608 DVSS.n12507 DVSS.n12505 0.771929
R23609 DVSS.n12515 DVSS.n12513 0.771929
R23610 DVSS.n12522 DVSS.n12520 0.771929
R23611 DVSS.n12529 DVSS.n12527 0.771929
R23612 DVSS.n12537 DVSS.n12535 0.771929
R23613 DVSS.n12545 DVSS.n12543 0.771929
R23614 DVSS.n12554 DVSS.n12550 0.771929
R23615 DVSS.n12554 DVSS.n12552 0.771929
R23616 DVSS.n12669 DVSS.n12667 0.771929
R23617 DVSS.n12661 DVSS.n12659 0.771929
R23618 DVSS.n12653 DVSS.n12651 0.771929
R23619 DVSS.n12646 DVSS.n12644 0.771929
R23620 DVSS.n12639 DVSS.n12637 0.771929
R23621 DVSS.n12631 DVSS.n12629 0.771929
R23622 DVSS.n12623 DVSS.n12621 0.771929
R23623 DVSS.n12615 DVSS.n12613 0.771929
R23624 DVSS.n12607 DVSS.n12605 0.771929
R23625 DVSS.n12599 DVSS.n12597 0.771929
R23626 DVSS.n12591 DVSS.n12589 0.771929
R23627 DVSS.n12584 DVSS.n12582 0.771929
R23628 DVSS.n12577 DVSS.n12575 0.771929
R23629 DVSS.n12569 DVSS.n12567 0.771929
R23630 DVSS.n12562 DVSS.n12560 0.771929
R23631 DVSS.n12221 DVSS.n12217 0.771929
R23632 DVSS.n12221 DVSS.n12219 0.771929
R23633 DVSS.n12381 DVSS.n12379 0.771929
R23634 DVSS.n12373 DVSS.n12371 0.771929
R23635 DVSS.n12365 DVSS.n12363 0.771929
R23636 DVSS.n12358 DVSS.n12356 0.771929
R23637 DVSS.n12351 DVSS.n12349 0.771929
R23638 DVSS.n12343 DVSS.n12341 0.771929
R23639 DVSS.n12335 DVSS.n12333 0.771929
R23640 DVSS.n12327 DVSS.n12325 0.771929
R23641 DVSS.n12319 DVSS.n12317 0.771929
R23642 DVSS.n12311 DVSS.n12309 0.771929
R23643 DVSS.n12303 DVSS.n12301 0.771929
R23644 DVSS.n12296 DVSS.n12294 0.771929
R23645 DVSS.n12289 DVSS.n12287 0.771929
R23646 DVSS.n12281 DVSS.n12279 0.771929
R23647 DVSS.n12273 DVSS.n12271 0.771929
R23648 DVSS.n12265 DVSS.n12263 0.771929
R23649 DVSS.n12257 DVSS.n12255 0.771929
R23650 DVSS.n12249 DVSS.n12247 0.771929
R23651 DVSS.n12242 DVSS.n12240 0.771929
R23652 DVSS.n12235 DVSS.n12233 0.771929
R23653 DVSS.n12227 DVSS.n12225 0.771929
R23654 DVSS.n21339 DVSS.n21335 0.771929
R23655 DVSS.n21339 DVSS.n21337 0.771929
R23656 DVSS.n21322 DVSS.n21320 0.771929
R23657 DVSS.n21217 DVSS.n21215 0.771929
R23658 DVSS.n21160 DVSS.n21155 0.771929
R23659 DVSS.n21155 DVSS.n21153 0.771929
R23660 DVSS.n21153 DVSS.n21152 0.771929
R23661 DVSS.n21170 DVSS.n21169 0.771929
R23662 DVSS.n21175 DVSS.n21174 0.771929
R23663 DVSS.n21179 DVSS.n21175 0.771929
R23664 DVSS.n3417 DVSS.n3415 0.771929
R23665 DVSS.n3419 DVSS.n3417 0.771929
R23666 DVSS.n3421 DVSS.n3419 0.771929
R23667 DVSS.n3423 DVSS.n3421 0.771929
R23668 DVSS.n3427 DVSS.n3423 0.771929
R23669 DVSS.n3427 DVSS.n3425 0.771929
R23670 DVSS.n3382 DVSS.n3380 0.771929
R23671 DVSS.n2762 DVSS.n2760 0.771929
R23672 DVSS.n2770 DVSS.n2768 0.771929
R23673 DVSS.n2779 DVSS.n2777 0.771929
R23674 DVSS.n3131 DVSS.n3129 0.771929
R23675 DVSS.n3139 DVSS.n3137 0.771929
R23676 DVSS.n3146 DVSS.n3144 0.771929
R23677 DVSS.n3153 DVSS.n3151 0.771929
R23678 DVSS.n3161 DVSS.n3159 0.771929
R23679 DVSS.n3169 DVSS.n3167 0.771929
R23680 DVSS.n3178 DVSS.n3174 0.771929
R23681 DVSS.n3178 DVSS.n3176 0.771929
R23682 DVSS.n3293 DVSS.n3291 0.771929
R23683 DVSS.n3285 DVSS.n3283 0.771929
R23684 DVSS.n3277 DVSS.n3275 0.771929
R23685 DVSS.n3270 DVSS.n3268 0.771929
R23686 DVSS.n3263 DVSS.n3261 0.771929
R23687 DVSS.n3255 DVSS.n3253 0.771929
R23688 DVSS.n3247 DVSS.n3245 0.771929
R23689 DVSS.n3239 DVSS.n3237 0.771929
R23690 DVSS.n3231 DVSS.n3229 0.771929
R23691 DVSS.n3223 DVSS.n3221 0.771929
R23692 DVSS.n3215 DVSS.n3213 0.771929
R23693 DVSS.n3208 DVSS.n3206 0.771929
R23694 DVSS.n3201 DVSS.n3199 0.771929
R23695 DVSS.n3193 DVSS.n3191 0.771929
R23696 DVSS.n3186 DVSS.n3184 0.771929
R23697 DVSS.n2851 DVSS.n2847 0.771929
R23698 DVSS.n2851 DVSS.n2849 0.771929
R23699 DVSS.n3008 DVSS.n3006 0.771929
R23700 DVSS.n3000 DVSS.n2998 0.771929
R23701 DVSS.n2992 DVSS.n2990 0.771929
R23702 DVSS.n2985 DVSS.n2983 0.771929
R23703 DVSS.n2978 DVSS.n2976 0.771929
R23704 DVSS.n2970 DVSS.n2968 0.771929
R23705 DVSS.n2962 DVSS.n2960 0.771929
R23706 DVSS.n2954 DVSS.n2952 0.771929
R23707 DVSS.n2946 DVSS.n2944 0.771929
R23708 DVSS.n2938 DVSS.n2936 0.771929
R23709 DVSS.n2930 DVSS.n2928 0.771929
R23710 DVSS.n2923 DVSS.n2921 0.771929
R23711 DVSS.n2916 DVSS.n2914 0.771929
R23712 DVSS.n2908 DVSS.n2906 0.771929
R23713 DVSS.n2900 DVSS.n2898 0.771929
R23714 DVSS.n2892 DVSS.n2890 0.771929
R23715 DVSS.n2884 DVSS.n2882 0.771929
R23716 DVSS.n2876 DVSS.n2874 0.771929
R23717 DVSS.n2869 DVSS.n2867 0.771929
R23718 DVSS.n2862 DVSS.n2860 0.771929
R23719 DVSS.n881 DVSS.n879 0.771929
R23720 DVSS.n889 DVSS.n887 0.771929
R23721 DVSS.n897 DVSS.n895 0.771929
R23722 DVSS.n905 DVSS.n903 0.771929
R23723 DVSS.n925 DVSS.n911 0.771929
R23724 DVSS.n925 DVSS.n922 0.771929
R23725 DVSS.n922 DVSS.n921 0.771929
R23726 DVSS.n921 DVSS.n920 0.771929
R23727 DVSS.n947 DVSS.n944 0.771929
R23728 DVSS.n947 DVSS.n945 0.771929
R23729 DVSS.n939 DVSS.n937 0.754407
R23730 DVSS.n21184 DVSS.n21183 0.7505
R23731 DVSS.n12817 DVSS.n12816 0.7505
R23732 DVSS.n3429 DVSS.n3428 0.7505
R23733 DVSS.n3363 DVSS.n2772 0.7505
R23734 DVSS.n12750 DVSS.n12152 0.7505
R23735 DVSS.n12773 DVSS.n12772 0.7505
R23736 DVSS.n12744 DVSS.n12743 0.7505
R23737 DVSS.n3370 DVSS.n2764 0.7505
R23738 DVSS.n12757 DVSS.n12144 0.7505
R23739 DVSS.n3385 DVSS.n3384 0.7505
R23740 DVSS.n3357 DVSS.n2781 0.7505
R23741 DVSS.n21207 DVSS.n21206 0.7505
R23742 DVSS.n21342 DVSS.n21341 0.7505
R23743 DVSS.n21326 DVSS.n21325 0.7505
R23744 DVSS.n21221 DVSS.n21220 0.7505
R23745 DVSS.n21160 DVSS.n21148 0.748877
R23746 DVSS.n15259 DVSS.n15258 0.716353
R23747 DVSS.n21179 DVSS.n21178 0.7005
R23748 DVSS.n939 DVSS.n938 0.7005
R23749 DVSS.n12243 DVSS.n12242 0.696929
R23750 DVSS.n12242 DVSS.n12241 0.696929
R23751 DVSS.n12250 DVSS.n12249 0.696929
R23752 DVSS.n12249 DVSS.n12248 0.696929
R23753 DVSS.n12258 DVSS.n12257 0.696929
R23754 DVSS.n12257 DVSS.n12256 0.696929
R23755 DVSS.n12297 DVSS.n12296 0.696929
R23756 DVSS.n12296 DVSS.n12295 0.696929
R23757 DVSS.n12304 DVSS.n12303 0.696929
R23758 DVSS.n12303 DVSS.n12302 0.696929
R23759 DVSS.n12312 DVSS.n12311 0.696929
R23760 DVSS.n12311 DVSS.n12310 0.696929
R23761 DVSS.n12328 DVSS.n12327 0.696929
R23762 DVSS.n12327 DVSS.n12326 0.696929
R23763 DVSS.n12359 DVSS.n12358 0.696929
R23764 DVSS.n12358 DVSS.n12357 0.696929
R23765 DVSS.n12366 DVSS.n12365 0.696929
R23766 DVSS.n12365 DVSS.n12364 0.696929
R23767 DVSS.n12374 DVSS.n12373 0.696929
R23768 DVSS.n12373 DVSS.n12372 0.696929
R23769 DVSS.n12557 DVSS.n12556 0.696929
R23770 DVSS.n12556 DVSS.n12555 0.696929
R23771 DVSS.n12563 DVSS.n12562 0.696929
R23772 DVSS.n12562 DVSS.n12561 0.696929
R23773 DVSS.n12585 DVSS.n12584 0.696929
R23774 DVSS.n12584 DVSS.n12583 0.696929
R23775 DVSS.n12592 DVSS.n12591 0.696929
R23776 DVSS.n12591 DVSS.n12590 0.696929
R23777 DVSS.n12608 DVSS.n12607 0.696929
R23778 DVSS.n12607 DVSS.n12606 0.696929
R23779 DVSS.n12616 DVSS.n12615 0.696929
R23780 DVSS.n12615 DVSS.n12614 0.696929
R23781 DVSS.n12647 DVSS.n12646 0.696929
R23782 DVSS.n12646 DVSS.n12645 0.696929
R23783 DVSS.n12654 DVSS.n12653 0.696929
R23784 DVSS.n12653 DVSS.n12652 0.696929
R23785 DVSS.n12673 DVSS.n12554 0.696929
R23786 DVSS.n12554 DVSS.n12553 0.696929
R23787 DVSS.n12523 DVSS.n12522 0.696929
R23788 DVSS.n12522 DVSS.n12521 0.696929
R23789 DVSS.n12516 DVSS.n12515 0.696929
R23790 DVSS.n12515 DVSS.n12514 0.696929
R23791 DVSS.n12508 DVSS.n12507 0.696929
R23792 DVSS.n12507 DVSS.n12506 0.696929
R23793 DVSS.n21205 DVSS.n21204 0.696929
R23794 DVSS.n21204 DVSS.n21203 0.696929
R23795 DVSS.n12530 DVSS.n12529 0.696929
R23796 DVSS.n12529 DVSS.n12528 0.696929
R23797 DVSS.n12538 DVSS.n12537 0.696929
R23798 DVSS.n12537 DVSS.n12536 0.696929
R23799 DVSS.n12546 DVSS.n12545 0.696929
R23800 DVSS.n12545 DVSS.n12544 0.696929
R23801 DVSS.n12670 DVSS.n12669 0.696929
R23802 DVSS.n12669 DVSS.n12668 0.696929
R23803 DVSS.n12662 DVSS.n12661 0.696929
R23804 DVSS.n12661 DVSS.n12660 0.696929
R23805 DVSS.n12640 DVSS.n12639 0.696929
R23806 DVSS.n12639 DVSS.n12638 0.696929
R23807 DVSS.n12632 DVSS.n12631 0.696929
R23808 DVSS.n12631 DVSS.n12630 0.696929
R23809 DVSS.n12624 DVSS.n12623 0.696929
R23810 DVSS.n12623 DVSS.n12622 0.696929
R23811 DVSS.n12600 DVSS.n12599 0.696929
R23812 DVSS.n12599 DVSS.n12598 0.696929
R23813 DVSS.n12578 DVSS.n12577 0.696929
R23814 DVSS.n12577 DVSS.n12576 0.696929
R23815 DVSS.n12570 DVSS.n12569 0.696929
R23816 DVSS.n12569 DVSS.n12568 0.696929
R23817 DVSS.n12385 DVSS.n12221 0.696929
R23818 DVSS.n12221 DVSS.n12220 0.696929
R23819 DVSS.n12382 DVSS.n12381 0.696929
R23820 DVSS.n12381 DVSS.n12380 0.696929
R23821 DVSS.n12352 DVSS.n12351 0.696929
R23822 DVSS.n12351 DVSS.n12350 0.696929
R23823 DVSS.n12344 DVSS.n12343 0.696929
R23824 DVSS.n12343 DVSS.n12342 0.696929
R23825 DVSS.n12336 DVSS.n12335 0.696929
R23826 DVSS.n12335 DVSS.n12334 0.696929
R23827 DVSS.n12320 DVSS.n12319 0.696929
R23828 DVSS.n12319 DVSS.n12318 0.696929
R23829 DVSS.n12290 DVSS.n12289 0.696929
R23830 DVSS.n12289 DVSS.n12288 0.696929
R23831 DVSS.n12282 DVSS.n12281 0.696929
R23832 DVSS.n12281 DVSS.n12280 0.696929
R23833 DVSS.n12274 DVSS.n12273 0.696929
R23834 DVSS.n12273 DVSS.n12272 0.696929
R23835 DVSS.n12266 DVSS.n12265 0.696929
R23836 DVSS.n12265 DVSS.n12264 0.696929
R23837 DVSS.n12236 DVSS.n12235 0.696929
R23838 DVSS.n12235 DVSS.n12234 0.696929
R23839 DVSS.n12228 DVSS.n12227 0.696929
R23840 DVSS.n12227 DVSS.n12226 0.696929
R23841 DVSS.n21340 DVSS.n21339 0.696929
R23842 DVSS.n21339 DVSS.n21338 0.696929
R23843 DVSS.n12500 DVSS.n12499 0.696929
R23844 DVSS.n12499 DVSS.n12498 0.696929
R23845 DVSS.n12742 DVSS.n12741 0.696929
R23846 DVSS.n12741 DVSS.n12740 0.696929
R23847 DVSS.n12151 DVSS.n12150 0.696929
R23848 DVSS.n12150 DVSS.n12149 0.696929
R23849 DVSS.n12143 DVSS.n12142 0.696929
R23850 DVSS.n12142 DVSS.n12141 0.696929
R23851 DVSS.n12771 DVSS.n12770 0.696929
R23852 DVSS.n12770 DVSS.n12769 0.696929
R23853 DVSS.n12816 DVSS.n12815 0.696929
R23854 DVSS.n12815 DVSS.n12814 0.696929
R23855 DVSS.n21323 DVSS.n21322 0.696929
R23856 DVSS.n21322 DVSS.n21321 0.696929
R23857 DVSS.n21218 DVSS.n21217 0.696929
R23858 DVSS.n21217 DVSS.n21216 0.696929
R23859 DVSS.n21161 DVSS.n21160 0.696929
R23860 DVSS.n926 DVSS.n925 0.696929
R23861 DVSS.n3132 DVSS.n3131 0.696929
R23862 DVSS.n3131 DVSS.n3130 0.696929
R23863 DVSS.n3140 DVSS.n3139 0.696929
R23864 DVSS.n3139 DVSS.n3138 0.696929
R23865 DVSS.n3278 DVSS.n3277 0.696929
R23866 DVSS.n3277 DVSS.n3276 0.696929
R23867 DVSS.n3240 DVSS.n3239 0.696929
R23868 DVSS.n3239 DVSS.n3238 0.696929
R23869 DVSS.n3232 DVSS.n3231 0.696929
R23870 DVSS.n3231 DVSS.n3230 0.696929
R23871 DVSS.n3216 DVSS.n3215 0.696929
R23872 DVSS.n3215 DVSS.n3214 0.696929
R23873 DVSS.n3001 DVSS.n3000 0.696929
R23874 DVSS.n3000 DVSS.n2999 0.696929
R23875 DVSS.n2993 DVSS.n2992 0.696929
R23876 DVSS.n2992 DVSS.n2991 0.696929
R23877 DVSS.n2955 DVSS.n2954 0.696929
R23878 DVSS.n2954 DVSS.n2953 0.696929
R23879 DVSS.n2939 DVSS.n2938 0.696929
R23880 DVSS.n2938 DVSS.n2937 0.696929
R23881 DVSS.n2931 DVSS.n2930 0.696929
R23882 DVSS.n2930 DVSS.n2929 0.696929
R23883 DVSS.n2885 DVSS.n2884 0.696929
R23884 DVSS.n2884 DVSS.n2883 0.696929
R23885 DVSS.n2877 DVSS.n2876 0.696929
R23886 DVSS.n2876 DVSS.n2875 0.696929
R23887 DVSS.n898 DVSS.n897 0.696929
R23888 DVSS.n897 DVSS.n896 0.696929
R23889 DVSS.n3124 DVSS.n3123 0.696929
R23890 DVSS.n3123 DVSS.n3122 0.696929
R23891 DVSS.n3154 DVSS.n3153 0.696929
R23892 DVSS.n3153 DVSS.n3152 0.696929
R23893 DVSS.n3162 DVSS.n3161 0.696929
R23894 DVSS.n3161 DVSS.n3160 0.696929
R23895 DVSS.n3170 DVSS.n3169 0.696929
R23896 DVSS.n3169 DVSS.n3168 0.696929
R23897 DVSS.n3294 DVSS.n3293 0.696929
R23898 DVSS.n3293 DVSS.n3292 0.696929
R23899 DVSS.n3286 DVSS.n3285 0.696929
R23900 DVSS.n3285 DVSS.n3284 0.696929
R23901 DVSS.n3264 DVSS.n3263 0.696929
R23902 DVSS.n3263 DVSS.n3262 0.696929
R23903 DVSS.n3256 DVSS.n3255 0.696929
R23904 DVSS.n3255 DVSS.n3254 0.696929
R23905 DVSS.n3248 DVSS.n3247 0.696929
R23906 DVSS.n3247 DVSS.n3246 0.696929
R23907 DVSS.n3224 DVSS.n3223 0.696929
R23908 DVSS.n3223 DVSS.n3222 0.696929
R23909 DVSS.n3202 DVSS.n3201 0.696929
R23910 DVSS.n3201 DVSS.n3200 0.696929
R23911 DVSS.n3194 DVSS.n3193 0.696929
R23912 DVSS.n3193 DVSS.n3192 0.696929
R23913 DVSS.n3012 DVSS.n2851 0.696929
R23914 DVSS.n2851 DVSS.n2850 0.696929
R23915 DVSS.n3009 DVSS.n3008 0.696929
R23916 DVSS.n3008 DVSS.n3007 0.696929
R23917 DVSS.n2979 DVSS.n2978 0.696929
R23918 DVSS.n2978 DVSS.n2977 0.696929
R23919 DVSS.n2971 DVSS.n2970 0.696929
R23920 DVSS.n2970 DVSS.n2969 0.696929
R23921 DVSS.n2963 DVSS.n2962 0.696929
R23922 DVSS.n2962 DVSS.n2961 0.696929
R23923 DVSS.n2947 DVSS.n2946 0.696929
R23924 DVSS.n2946 DVSS.n2945 0.696929
R23925 DVSS.n2917 DVSS.n2916 0.696929
R23926 DVSS.n2916 DVSS.n2915 0.696929
R23927 DVSS.n2909 DVSS.n2908 0.696929
R23928 DVSS.n2908 DVSS.n2907 0.696929
R23929 DVSS.n2901 DVSS.n2900 0.696929
R23930 DVSS.n2900 DVSS.n2899 0.696929
R23931 DVSS.n2893 DVSS.n2892 0.696929
R23932 DVSS.n2892 DVSS.n2891 0.696929
R23933 DVSS.n2863 DVSS.n2862 0.696929
R23934 DVSS.n2862 DVSS.n2861 0.696929
R23935 DVSS.n2855 DVSS.n2854 0.696929
R23936 DVSS.n2854 DVSS.n2853 0.696929
R23937 DVSS.n882 DVSS.n881 0.696929
R23938 DVSS.n881 DVSS.n880 0.696929
R23939 DVSS.n2771 DVSS.n2770 0.696929
R23940 DVSS.n2770 DVSS.n2769 0.696929
R23941 DVSS.n2763 DVSS.n2762 0.696929
R23942 DVSS.n2762 DVSS.n2761 0.696929
R23943 DVSS.n3383 DVSS.n3382 0.696929
R23944 DVSS.n3382 DVSS.n3381 0.696929
R23945 DVSS.n2780 DVSS.n2779 0.696929
R23946 DVSS.n2779 DVSS.n2778 0.696929
R23947 DVSS.n890 DVSS.n889 0.696929
R23948 DVSS.n889 DVSS.n888 0.696929
R23949 DVSS.n906 DVSS.n905 0.696929
R23950 DVSS.n905 DVSS.n904 0.696929
R23951 DVSS.n3398 DVSS.n3397 0.696929
R23952 DVSS.n3417 DVSS.n3416 0.696929
R23953 DVSS.n12809 DVSS.n12808 0.696929
R23954 DVSS.n3421 DVSS.n3420 0.696929
R23955 DVSS.n3403 DVSS.n3402 0.696929
R23956 DVSS.n3428 DVSS.n3427 0.696929
R23957 DVSS.n3427 DVSS.n3426 0.696929
R23958 DVSS.n3147 DVSS.n3146 0.696929
R23959 DVSS.n3146 DVSS.n3145 0.696929
R23960 DVSS.n3297 DVSS.n3178 0.696929
R23961 DVSS.n3178 DVSS.n3177 0.696929
R23962 DVSS.n3271 DVSS.n3270 0.696929
R23963 DVSS.n3270 DVSS.n3269 0.696929
R23964 DVSS.n3209 DVSS.n3208 0.696929
R23965 DVSS.n3208 DVSS.n3207 0.696929
R23966 DVSS.n3187 DVSS.n3186 0.696929
R23967 DVSS.n3186 DVSS.n3185 0.696929
R23968 DVSS.n3181 DVSS.n3180 0.696929
R23969 DVSS.n3180 DVSS.n3179 0.696929
R23970 DVSS.n2986 DVSS.n2985 0.696929
R23971 DVSS.n2985 DVSS.n2984 0.696929
R23972 DVSS.n2924 DVSS.n2923 0.696929
R23973 DVSS.n2923 DVSS.n2922 0.696929
R23974 DVSS.n2870 DVSS.n2869 0.696929
R23975 DVSS.n2869 DVSS.n2868 0.696929
R23976 DVSS.n12788 DVSS.n12787 0.696929
R23977 DVSS.n12790 DVSS.n12789 0.696929
R23978 DVSS.n12805 DVSS.n12804 0.696929
R23979 DVSS.n12788 DVSS.n12785 0.686214
R23980 DVSS.n3403 DVSS.n3400 0.686214
R23981 DVSS.n353 DVSS.n351 0.685697
R23982 DVSS.n347 DVSS.n345 0.685697
R23983 DVSS.n5833 DVSS 0.66425
R23984 DVSS.n11030 DVSS 0.66425
R23985 DVSS.n6767 DVSS 0.66425
R23986 DVSS.n11657 DVSS 0.66425
R23987 DVSS.n6712 DVSS 0.66425
R23988 DVSS.n11620 DVSS 0.66425
R23989 DVSS.n6569 DVSS 0.66425
R23990 DVSS.n11495 DVSS 0.66425
R23991 DVSS.n6474 DVSS 0.66425
R23992 DVSS.n11203 DVSS 0.66425
R23993 DVSS.n6433 DVSS 0.66425
R23994 DVSS.n11458 DVSS 0.66425
R23995 DVSS.n8041 DVSS 0.66425
R23996 DVSS.n6894 DVSS 0.66425
R23997 DVSS.n11707 DVSS 0.66425
R23998 DVSS.n5515 DVSS 0.66425
R23999 DVSS.n10042 DVSS 0.66425
R24000 DVSS.n6902 DVSS 0.66425
R24001 DVSS.n14207 DVSS.n14206 0.6505
R24002 DVSS.n14198 DVSS.n14197 0.6505
R24003 DVSS.n14190 DVSS.t3 0.6505
R24004 DVSS.n14191 DVSS.n14190 0.6505
R24005 DVSS.n14077 DVSS.n14076 0.6505
R24006 DVSS.n14677 DVSS.t37 0.6505
R24007 DVSS.n14678 DVSS.n14677 0.6505
R24008 DVSS.n14731 DVSS.n14730 0.6505
R24009 DVSS.n10017 DVSS.n10016 0.647738
R24010 DVSS.n16965 DVSS.n16959 0.632106
R24011 DVSS.n16965 DVSS.n16964 0.632106
R24012 DVSS.n14903 DVSS.n14897 0.632106
R24013 DVSS.n14903 DVSS.n14902 0.632106
R24014 DVSS.n14910 DVSS.n14906 0.624161
R24015 DVSS.n11490 DVSS.n11489 0.623413
R24016 DVSS.n11652 DVSS.n11651 0.623413
R24017 DVSS.n6357 DVSS.n6356 0.623413
R24018 DVSS.n6717 DVSS.n6716 0.623413
R24019 DVSS.n10777 DVSS.n10776 0.617744
R24020 DVSS.n5503 DVSS.n5502 0.617744
R24021 DVSS.n13052 DVSS.n13051 0.616858
R24022 DVSS.n6899 DVSS.n6898 0.616858
R24023 DVSS.n6524 DVSS.n6523 0.612075
R24024 DVSS.n4083 DVSS.n2546 0.612075
R24025 DVSS.n9763 DVSS.n9762 0.612075
R24026 DVSS.n9151 DVSS.n9150 0.612075
R24027 DVSS.n15709 DVSS.n7665 0.612075
R24028 DVSS.n14979 DVSS.n7694 0.612075
R24029 DVSS.n4129 DVSS.n4128 0.612075
R24030 DVSS.n9706 DVSS.n8928 0.612075
R24031 DVSS.n9094 DVSS.n8961 0.612075
R24032 DVSS.n16259 DVSS.n16258 0.612075
R24033 DVSS.n18378 DVSS.n18377 0.612075
R24034 DVSS.n5702 DVSS.n5701 0.61172
R24035 DVSS.n10992 DVSS.n10991 0.61172
R24036 DVSS.n16915 DVSS.n16914 0.61172
R24037 DVSS.n9871 DVSS.n9870 0.61172
R24038 DVSS.n17421 DVSS.n17420 0.61172
R24039 DVSS.n2574 DVSS.n1347 0.611189
R24040 DVSS.n13151 DVSS.n13150 0.611189
R24041 DVSS.n14955 DVSS.n14954 0.611189
R24042 DVSS.n3790 DVSS.n3789 0.611189
R24043 DVSS.n9011 DVSS.n8006 0.611189
R24044 DVSS.n7469 DVSS.n7431 0.611189
R24045 DVSS.n11453 DVSS.n11452 0.606228
R24046 DVSS.n6446 DVSS.n6445 0.606228
R24047 DVSS.n6380 DVSS.n6373 0.604265
R24048 DVSS.n2514 DVSS.n2507 0.604265
R24049 DVSS.n4502 DVSS.n4499 0.604265
R24050 DVSS.n16965 DVSS.n16960 0.604265
R24051 DVSS.n16965 DVSS.n16961 0.604265
R24052 DVSS.n4556 DVSS.n4544 0.604265
R24053 DVSS.n14903 DVSS.n14896 0.604265
R24054 DVSS.n14903 DVSS.n14895 0.604265
R24055 DVSS.n6511 DVSS.n6510 0.600559
R24056 DVSS.n9769 DVSS.n9768 0.600559
R24057 DVSS.n15866 DVSS.n15865 0.600559
R24058 DVSS.n9809 DVSS.n9808 0.600559
R24059 DVSS.n16298 DVSS.n16297 0.600559
R24060 DVSS.n6380 DVSS.n6378 0.594741
R24061 DVSS.n2514 DVSS.n2512 0.594741
R24062 DVSS.n6687 DVSS.n6681 0.594741
R24063 DVSS.n6687 DVSS.n6685 0.594741
R24064 DVSS.n15258 DVSS.n15252 0.594741
R24065 DVSS.n15258 DVSS.n15256 0.594741
R24066 DVSS.n4502 DVSS.n4497 0.594741
R24067 DVSS.n4556 DVSS.n4552 0.594741
R24068 DVSS.n6869 DVSS.n6863 0.594741
R24069 DVSS.n6869 DVSS.n6867 0.594741
R24070 DVSS.n4606 DVSS.n4602 0.594741
R24071 DVSS.n4606 DVSS.n4600 0.594741
R24072 DVSS.n6380 DVSS.n6379 0.586651
R24073 DVSS.n2514 DVSS.n2513 0.586651
R24074 DVSS.n6687 DVSS.n6680 0.586651
R24075 DVSS.n6687 DVSS.n6686 0.586651
R24076 DVSS.n15258 DVSS.n15251 0.586651
R24077 DVSS.n15258 DVSS.n15257 0.586651
R24078 DVSS.n4502 DVSS.n4498 0.586651
R24079 DVSS.n4556 DVSS.n4555 0.586651
R24080 DVSS.n6869 DVSS.n6862 0.586651
R24081 DVSS.n6869 DVSS.n6868 0.586651
R24082 DVSS.n4606 DVSS.n4603 0.586651
R24083 DVSS.n4606 DVSS.n4604 0.586651
R24084 DVSS.n16968 DVSS.n16967 0.576595
R24085 DVSS.n14894 DVSS.n14893 0.576595
R24086 DVSS.n19951 DVSS.n19950 0.5205
R24087 DVSS.n19950 DVSS.n19949 0.5205
R24088 DVSS.n359 DVSS.n358 0.5205
R24089 DVSS.n358 DVSS.n357 0.5205
R24090 DVSS.n3298 DVSS.n3297 0.5005
R24091 DVSS.n12674 DVSS.n12673 0.5005
R24092 DVSS.n12386 DVSS.n12385 0.5005
R24093 DVSS.n3013 DVSS.n3012 0.5005
R24094 DVSS.n6380 DVSS.n6374 0.466929
R24095 DVSS.n2514 DVSS.n2508 0.466929
R24096 DVSS.n4502 DVSS.n4500 0.466929
R24097 DVSS.n4556 DVSS.n4545 0.466929
R24098 DVSS.n13809 DVSS.n13807 0.403878
R24099 DVSS.n7407 DVSS.n7405 0.403878
R24100 DVSS.n7359 DVSS.n7355 0.403878
R24101 DVSS.n13729 DVSS.n13726 0.403878
R24102 DVSS.n14344 DVSS.n14343 0.394514
R24103 DVSS.n14799 DVSS.n14798 0.394514
R24104 DVSS.n18588 DVSS.n18587 0.376311
R24105 DVSS.n7342 DVSS.n7340 0.376311
R24106 DVSS.n18714 DVSS.n18713 0.376311
R24107 DVSS.n13839 DVSS.n13837 0.375905
R24108 DVSS.n13695 DVSS.n13691 0.375905
R24109 DVSS.n13684 DVSS.n13682 0.375905
R24110 DVSS.n7005 DVSS.n7004 0.373473
R24111 DVSS.n13676 DVSS.n13675 0.373473
R24112 DVSS.n14944 DVSS 0.37265
R24113 DVSS.n7434 DVSS 0.37265
R24114 DVSS.n19383 DVSS.n19382 0.371446
R24115 DVSS.n20167 DVSS.n20166 0.371041
R24116 DVSS.n19430 DVSS.n19429 0.368608
R24117 DVSS.n20438 DVSS.n20437 0.368608
R24118 DVSS.n5629 DVSS.n5628 0.345264
R24119 DVSS.n10920 DVSS.n10919 0.345264
R24120 DVSS.n17053 DVSS.n17052 0.345264
R24121 DVSS.n10842 DVSS.n10841 0.345264
R24122 DVSS.n9942 DVSS.n9941 0.345264
R24123 DVSS.n17348 DVSS.n17347 0.345264
R24124 DVSS.n5424 DVSS.n5423 0.345264
R24125 DVSS.n5771 DVSS.n5770 0.344378
R24126 DVSS.n11276 DVSS.n11275 0.344378
R24127 DVSS.n17589 DVSS.n17588 0.344378
R24128 DVSS.n11386 DVSS.n11385 0.344378
R24129 DVSS.n11112 DVSS.n11111 0.344378
R24130 DVSS.n16392 DVSS.n16391 0.344378
R24131 DVSS.n6071 DVSS.n6070 0.344378
R24132 DVSS.n12920 DVSS.n12919 0.340835
R24133 DVSS.n12052 DVSS.n12051 0.340835
R24134 DVSS.n3744 DVSS.n3743 0.340835
R24135 DVSS.n3647 DVSS.n3646 0.340835
R24136 DVSS.n17435 DVSS 0.332375
R24137 DVSS.n16890 DVSS 0.332375
R24138 DVSS.n7463 DVSS 0.332375
R24139 DVSS.n14974 DVSS 0.332375
R24140 DVSS.n7552 DVSS 0.332375
R24141 DVSS.n15603 DVSS 0.332375
R24142 DVSS.n16224 DVSS 0.332375
R24143 DVSS.n7690 DVSS 0.332375
R24144 DVSS.n16308 DVSS 0.332375
R24145 DVSS.n17643 DVSS 0.332375
R24146 DVSS.n16263 DVSS 0.332375
R24147 DVSS.n15849 DVSS 0.332375
R24148 DVSS.n7473 DVSS 0.332375
R24149 DVSS.n7780 DVSS 0.332375
R24150 DVSS.n16428 DVSS 0.332375
R24151 DVSS.n16880 DVSS 0.332375
R24152 DVSS.n13689 DVSS.n13688 0.330913
R24153 DVSS.n18706 DVSS.n18705 0.330913
R24154 DVSS.n16965 DVSS.n16962 0.28898
R24155 DVSS.n16965 DVSS.n16957 0.28898
R24156 DVSS.n14903 DVSS.n14901 0.28898
R24157 DVSS.n14903 DVSS.n14898 0.28898
R24158 DVSS.n14903 DVSS.n14900 0.287336
R24159 DVSS.n14903 DVSS.n14899 0.287336
R24160 DVSS.n16965 DVSS.n16958 0.287064
R24161 DVSS.n16965 DVSS.n16963 0.287064
R24162 DVSS.n13063 DVSS.n13062 0.285913
R24163 DVSS.n6838 DVSS.n6837 0.285913
R24164 DVSS.n7847 DVSS.n7845 0.284689
R24165 DVSS.n7350 DVSS.n7348 0.284284
R24166 DVSS.n6380 DVSS.n6372 0.280941
R24167 DVSS.n6380 DVSS.n6377 0.280941
R24168 DVSS.n2514 DVSS.n2499 0.280941
R24169 DVSS.n2514 DVSS.n2511 0.280941
R24170 DVSS.n6687 DVSS.n6679 0.280941
R24171 DVSS.n6687 DVSS.n6684 0.280941
R24172 DVSS.n15258 DVSS.n15250 0.280941
R24173 DVSS.n15258 DVSS.n15255 0.280941
R24174 DVSS.n4502 DVSS.n4496 0.280941
R24175 DVSS.n4556 DVSS.n4551 0.280941
R24176 DVSS.n4556 DVSS.n4546 0.280941
R24177 DVSS.n4502 DVSS.n4501 0.280941
R24178 DVSS.n6869 DVSS.n6861 0.280941
R24179 DVSS.n6869 DVSS.n6866 0.280941
R24180 DVSS.n4606 DVSS.n4601 0.280941
R24181 DVSS.n4606 DVSS.n4605 0.280941
R24182 DVSS.n4045 DVSS.n4044 0.280244
R24183 DVSS.n13138 DVSS.n13137 0.280244
R24184 DVSS.n15033 DVSS.n15032 0.280244
R24185 DVSS.n3990 DVSS.n3989 0.280244
R24186 DVSS.n9052 DVSS.n9051 0.280244
R24187 DVSS.n7510 DVSS.n7509 0.280244
R24188 DVSS.n6869 DVSS.n6865 0.278361
R24189 DVSS.n4606 DVSS.n4599 0.278361
R24190 DVSS.n4606 DVSS.n4598 0.278361
R24191 DVSS.n6380 DVSS.n6375 0.278105
R24192 DVSS.n6380 DVSS.n6376 0.278105
R24193 DVSS.n2514 DVSS.n2509 0.278105
R24194 DVSS.n2514 DVSS.n2510 0.278105
R24195 DVSS.n6687 DVSS.n6682 0.278105
R24196 DVSS.n6687 DVSS.n6683 0.278105
R24197 DVSS.n15258 DVSS.n15253 0.278105
R24198 DVSS.n15258 DVSS.n15254 0.278105
R24199 DVSS.n4502 DVSS.n4495 0.278105
R24200 DVSS.n4556 DVSS.n4550 0.278105
R24201 DVSS.n4556 DVSS.n4547 0.278105
R24202 DVSS.n4502 DVSS.n4494 0.278105
R24203 DVSS.n6869 DVSS.n6864 0.278105
R24204 DVSS.n14219 DVSS.n14218 0.268599
R24205 DVSS.n14878 DVSS.n14877 0.268599
R24206 DVSS.n7022 DVSS.n7020 0.266041
R24207 DVSS.n13292 DVSS.n13290 0.265635
R24208 DVSS.n5060 DVSS.n5059 0.257472
R24209 DVSS.n10862 DVSS.n10861 0.257261
R24210 DVSS.n10868 DVSS.n10867 0.2505
R24211 DVSS.n10879 DVSS.n10878 0.2505
R24212 DVSS.n10880 DVSS.n10879 0.2505
R24213 DVSS.n10888 DVSS.n10887 0.2505
R24214 DVSS.n10887 DVSS.n10886 0.2505
R24215 DVSS.n10591 DVSS.n10590 0.2505
R24216 DVSS.n10587 DVSS.n10586 0.2505
R24217 DVSS.n10583 DVSS.n10582 0.2505
R24218 DVSS.n10576 DVSS.n10575 0.2505
R24219 DVSS.n10896 DVSS.n10895 0.2505
R24220 DVSS.n10897 DVSS.n10896 0.2505
R24221 DVSS.n10559 DVSS.n10558 0.2505
R24222 DVSS.n10560 DVSS.n10559 0.2505
R24223 DVSS.n10496 DVSS.n10495 0.2505
R24224 DVSS.n10480 DVSS.n10479 0.2505
R24225 DVSS.n10470 DVSS.n10469 0.2505
R24226 DVSS.n10462 DVSS.n10461 0.2505
R24227 DVSS.n10453 DVSS.n10452 0.2505
R24228 DVSS.n10441 DVSS.n10440 0.2505
R24229 DVSS.n10435 DVSS.n10434 0.2505
R24230 DVSS.n10433 DVSS.n10432 0.2505
R24231 DVSS.n10431 DVSS.n10430 0.2505
R24232 DVSS.n10421 DVSS.n10420 0.2505
R24233 DVSS.n10411 DVSS.n10410 0.2505
R24234 DVSS.n10403 DVSS.n10402 0.2505
R24235 DVSS.n10394 DVSS.n10393 0.2505
R24236 DVSS.n10388 DVSS.n10387 0.2505
R24237 DVSS.n10386 DVSS.n10385 0.2505
R24238 DVSS.n10384 DVSS.n10383 0.2505
R24239 DVSS.n10380 DVSS.n10379 0.2505
R24240 DVSS.n10378 DVSS.n10377 0.2505
R24241 DVSS.n10372 DVSS.n10371 0.2505
R24242 DVSS.n10363 DVSS.n10362 0.2505
R24243 DVSS.n10354 DVSS.n10353 0.2505
R24244 DVSS.n10341 DVSS.n10340 0.2505
R24245 DVSS.n10335 DVSS.n10334 0.2505
R24246 DVSS.n10323 DVSS.n10322 0.2505
R24247 DVSS.n10314 DVSS.n10313 0.2505
R24248 DVSS.n10306 DVSS.n10305 0.2505
R24249 DVSS.n10302 DVSS.n10301 0.2505
R24250 DVSS.n5084 DVSS.n5083 0.2505
R24251 DVSS.n5089 DVSS.n5088 0.2505
R24252 DVSS.n5096 DVSS.n5095 0.2505
R24253 DVSS.n5106 DVSS.n5105 0.2505
R24254 DVSS.n5114 DVSS.n5113 0.2505
R24255 DVSS.n5120 DVSS.n5119 0.2505
R24256 DVSS.n5126 DVSS.n5125 0.2505
R24257 DVSS.n5132 DVSS.n5131 0.2505
R24258 DVSS.n5134 DVSS.n5133 0.2505
R24259 DVSS.n5138 DVSS.n5137 0.2505
R24260 DVSS.n5143 DVSS.n5142 0.2505
R24261 DVSS.n5150 DVSS.n5149 0.2505
R24262 DVSS.n5160 DVSS.n5159 0.2505
R24263 DVSS.n5170 DVSS.n5169 0.2505
R24264 DVSS.n5172 DVSS.n5171 0.2505
R24265 DVSS.n5174 DVSS.n5173 0.2505
R24266 DVSS.n5176 DVSS.n5175 0.2505
R24267 DVSS.n5181 DVSS.n5180 0.2505
R24268 DVSS.n5188 DVSS.n5187 0.2505
R24269 DVSS.n5066 DVSS.n5064 0.2505
R24270 DVSS.n5067 DVSS.n5066 0.2505
R24271 DVSS.n5307 DVSS.n5306 0.2505
R24272 DVSS.n5308 DVSS.n5307 0.2505
R24273 DVSS.n5264 DVSS.n5263 0.2505
R24274 DVSS.n5259 DVSS.n5258 0.2505
R24275 DVSS.n5243 DVSS.n5242 0.2505
R24276 DVSS.n2457 DVSS.n2456 0.242431
R24277 DVSS.n14927 DVSS.n14925 0.233545
R24278 DVSS.n18563 DVSS.n18561 0.233293
R24279 DVSS.n4626 DVSS.n4625 0.231864
R24280 DVSS.n6789 DVSS.n6788 0.231864
R24281 DVSS.n3597 DVSS.n3596 0.231864
R24282 DVSS.n5861 DVSS.n5860 0.231864
R24283 DVSS.n6088 DVSS.n6087 0.231864
R24284 DVSS.n13089 DVSS.n13088 0.231671
R24285 DVSS.n13006 DVSS.n13005 0.231671
R24286 DVSS.n11341 DVSS.n11340 0.231671
R24287 DVSS.n16993 DVSS.n16991 0.231534
R24288 DVSS.n17301 DVSS.n17299 0.231282
R24289 DVSS.n17302 DVSS.n17301 0.230528
R24290 DVSS.n1722 DVSS.n1721 0.230514
R24291 DVSS.n2052 DVSS.n2051 0.230514
R24292 DVSS.n16994 DVSS.n16993 0.230277
R24293 DVSS.n17322 DVSS.n17321 0.228768
R24294 DVSS.n10214 DVSS.n10213 0.228768
R24295 DVSS.n2021 DVSS.n2020 0.2255
R24296 DVSS.n2023 DVSS.n2022 0.2255
R24297 DVSS.n2025 DVSS.n2024 0.2255
R24298 DVSS.n2027 DVSS.n2026 0.2255
R24299 DVSS.n2029 DVSS.n2028 0.2255
R24300 DVSS.n2031 DVSS.n2030 0.2255
R24301 DVSS.n2033 DVSS.n2032 0.2255
R24302 DVSS.n2035 DVSS.n2034 0.2255
R24303 DVSS.n2037 DVSS.n2036 0.2255
R24304 DVSS.n2041 DVSS.n2040 0.2255
R24305 DVSS.n2042 DVSS.n2041 0.2255
R24306 DVSS.n2333 DVSS.n2330 0.2255
R24307 DVSS.n2334 DVSS.n2333 0.2255
R24308 DVSS.n2066 DVSS.n2065 0.2255
R24309 DVSS.n2069 DVSS.n2068 0.2255
R24310 DVSS.n2071 DVSS.n2070 0.2255
R24311 DVSS.n2073 DVSS.n2072 0.2255
R24312 DVSS.n2075 DVSS.n2074 0.2255
R24313 DVSS.n2077 DVSS.n2076 0.2255
R24314 DVSS.n2079 DVSS.n2078 0.2255
R24315 DVSS.n2081 DVSS.n2080 0.2255
R24316 DVSS.n2083 DVSS.n2082 0.2255
R24317 DVSS.n2085 DVSS.n2084 0.2255
R24318 DVSS.n2087 DVSS.n2086 0.2255
R24319 DVSS.n2089 DVSS.n2088 0.2255
R24320 DVSS.n2091 DVSS.n2090 0.2255
R24321 DVSS.n2093 DVSS.n2092 0.2255
R24322 DVSS.n2095 DVSS.n2094 0.2255
R24323 DVSS.n2097 DVSS.n2096 0.2255
R24324 DVSS.n2099 DVSS.n2098 0.2255
R24325 DVSS.n2101 DVSS.n2100 0.2255
R24326 DVSS.n2103 DVSS.n2102 0.2255
R24327 DVSS.n2105 DVSS.n2104 0.2255
R24328 DVSS.n2107 DVSS.n2106 0.2255
R24329 DVSS.n2109 DVSS.n2108 0.2255
R24330 DVSS.n2111 DVSS.n2110 0.2255
R24331 DVSS.n2113 DVSS.n2112 0.2255
R24332 DVSS.n2115 DVSS.n2114 0.2255
R24333 DVSS.n2117 DVSS.n2116 0.2255
R24334 DVSS.n2119 DVSS.n2118 0.2255
R24335 DVSS.n2121 DVSS.n2120 0.2255
R24336 DVSS.n2123 DVSS.n2122 0.2255
R24337 DVSS.n2125 DVSS.n2124 0.2255
R24338 DVSS.n2127 DVSS.n2126 0.2255
R24339 DVSS.n2129 DVSS.n2128 0.2255
R24340 DVSS.n2131 DVSS.n2130 0.2255
R24341 DVSS.n2133 DVSS.n2132 0.2255
R24342 DVSS.n2135 DVSS.n2134 0.2255
R24343 DVSS.n2137 DVSS.n2136 0.2255
R24344 DVSS.n2139 DVSS.n2138 0.2255
R24345 DVSS.n2141 DVSS.n2140 0.2255
R24346 DVSS.n2144 DVSS.n2143 0.2255
R24347 DVSS.n2148 DVSS.n2147 0.2255
R24348 DVSS.n2151 DVSS.n2150 0.2255
R24349 DVSS.n2153 DVSS.n2152 0.2255
R24350 DVSS.n2155 DVSS.n2154 0.2255
R24351 DVSS.n2157 DVSS.n2156 0.2255
R24352 DVSS.n2159 DVSS.n2158 0.2255
R24353 DVSS.n2161 DVSS.n2160 0.2255
R24354 DVSS.n2163 DVSS.n2162 0.2255
R24355 DVSS.n2165 DVSS.n2164 0.2255
R24356 DVSS.n2167 DVSS.n2166 0.2255
R24357 DVSS.n2169 DVSS.n2168 0.2255
R24358 DVSS.n2171 DVSS.n2170 0.2255
R24359 DVSS.n2173 DVSS.n2172 0.2255
R24360 DVSS.n2175 DVSS.n2174 0.2255
R24361 DVSS.n2177 DVSS.n2176 0.2255
R24362 DVSS.n2179 DVSS.n2178 0.2255
R24363 DVSS.n2181 DVSS.n2180 0.2255
R24364 DVSS.n2183 DVSS.n2182 0.2255
R24365 DVSS.n2185 DVSS.n2184 0.2255
R24366 DVSS.n2187 DVSS.n2186 0.2255
R24367 DVSS.n2189 DVSS.n2188 0.2255
R24368 DVSS.n2191 DVSS.n2190 0.2255
R24369 DVSS.n2193 DVSS.n2192 0.2255
R24370 DVSS.n2195 DVSS.n2194 0.2255
R24371 DVSS.n2197 DVSS.n2196 0.2255
R24372 DVSS.n2199 DVSS.n2198 0.2255
R24373 DVSS.n2201 DVSS.n2200 0.2255
R24374 DVSS.n2203 DVSS.n2202 0.2255
R24375 DVSS.n2205 DVSS.n2204 0.2255
R24376 DVSS.n2207 DVSS.n2206 0.2255
R24377 DVSS.n2209 DVSS.n2208 0.2255
R24378 DVSS.n2211 DVSS.n2210 0.2255
R24379 DVSS.n2213 DVSS.n2212 0.2255
R24380 DVSS.n2215 DVSS.n2214 0.2255
R24381 DVSS.n2218 DVSS.n2217 0.2255
R24382 DVSS.n2221 DVSS.n2220 0.2255
R24383 DVSS.n2223 DVSS.n2222 0.2255
R24384 DVSS.n2225 DVSS.n2224 0.2255
R24385 DVSS.n2227 DVSS.n2226 0.2255
R24386 DVSS.n2229 DVSS.n2228 0.2255
R24387 DVSS.n2232 DVSS.n2231 0.2255
R24388 DVSS.n2236 DVSS.n2235 0.2255
R24389 DVSS.n2239 DVSS.n2238 0.2255
R24390 DVSS.n2242 DVSS.n2241 0.2255
R24391 DVSS.n2241 DVSS.n2240 0.2255
R24392 DVSS.n2060 DVSS.n2059 0.2255
R24393 DVSS.n2059 DVSS.n2058 0.2255
R24394 DVSS.n2057 DVSS.n2056 0.2255
R24395 DVSS.n2056 DVSS.n2055 0.2255
R24396 DVSS.n2054 DVSS.n2053 0.2255
R24397 DVSS.n1998 DVSS.n1997 0.2255
R24398 DVSS.n1994 DVSS.n1993 0.2255
R24399 DVSS.n1992 DVSS.n1991 0.2255
R24400 DVSS.n1990 DVSS.n1989 0.2255
R24401 DVSS.n1988 DVSS.n1987 0.2255
R24402 DVSS.n1986 DVSS.n1985 0.2255
R24403 DVSS.n1984 DVSS.n1983 0.2255
R24404 DVSS.n1982 DVSS.n1981 0.2255
R24405 DVSS.n1980 DVSS.n1979 0.2255
R24406 DVSS.n1978 DVSS.n1977 0.2255
R24407 DVSS.n1976 DVSS.n1975 0.2255
R24408 DVSS.n1974 DVSS.n1973 0.2255
R24409 DVSS.n1972 DVSS.n1971 0.2255
R24410 DVSS.n1966 DVSS.n1965 0.2255
R24411 DVSS.n1964 DVSS.n1963 0.2255
R24412 DVSS.n1962 DVSS.n1961 0.2255
R24413 DVSS.n1958 DVSS.n1957 0.2255
R24414 DVSS.n1956 DVSS.n1955 0.2255
R24415 DVSS.n1954 DVSS.n1953 0.2255
R24416 DVSS.n1952 DVSS.n1951 0.2255
R24417 DVSS.n1950 DVSS.n1949 0.2255
R24418 DVSS.n1948 DVSS.n1947 0.2255
R24419 DVSS.n1942 DVSS.n1941 0.2255
R24420 DVSS.n1940 DVSS.n1939 0.2255
R24421 DVSS.n1574 DVSS.n1573 0.2255
R24422 DVSS.n1576 DVSS.n1575 0.2255
R24423 DVSS.n1578 DVSS.n1577 0.2255
R24424 DVSS.n1580 DVSS.n1579 0.2255
R24425 DVSS.n1582 DVSS.n1581 0.2255
R24426 DVSS.n1584 DVSS.n1583 0.2255
R24427 DVSS.n1586 DVSS.n1585 0.2255
R24428 DVSS.n1588 DVSS.n1587 0.2255
R24429 DVSS.n1590 DVSS.n1589 0.2255
R24430 DVSS.n1592 DVSS.n1591 0.2255
R24431 DVSS.n1594 DVSS.n1593 0.2255
R24432 DVSS.n1596 DVSS.n1595 0.2255
R24433 DVSS.n1598 DVSS.n1597 0.2255
R24434 DVSS.n1600 DVSS.n1599 0.2255
R24435 DVSS.n1602 DVSS.n1601 0.2255
R24436 DVSS.n1604 DVSS.n1603 0.2255
R24437 DVSS.n1606 DVSS.n1605 0.2255
R24438 DVSS.n1608 DVSS.n1607 0.2255
R24439 DVSS.n1610 DVSS.n1609 0.2255
R24440 DVSS.n1612 DVSS.n1611 0.2255
R24441 DVSS.n1614 DVSS.n1613 0.2255
R24442 DVSS.n1616 DVSS.n1615 0.2255
R24443 DVSS.n1618 DVSS.n1617 0.2255
R24444 DVSS.n1620 DVSS.n1619 0.2255
R24445 DVSS.n1622 DVSS.n1621 0.2255
R24446 DVSS.n1624 DVSS.n1623 0.2255
R24447 DVSS.n1626 DVSS.n1625 0.2255
R24448 DVSS.n1628 DVSS.n1627 0.2255
R24449 DVSS.n1630 DVSS.n1629 0.2255
R24450 DVSS.n1632 DVSS.n1631 0.2255
R24451 DVSS.n1634 DVSS.n1633 0.2255
R24452 DVSS.n1636 DVSS.n1635 0.2255
R24453 DVSS.n1638 DVSS.n1637 0.2255
R24454 DVSS.n1640 DVSS.n1639 0.2255
R24455 DVSS.n1642 DVSS.n1641 0.2255
R24456 DVSS.n1645 DVSS.n1644 0.2255
R24457 DVSS.n1644 DVSS.n1643 0.2255
R24458 DVSS.n1648 DVSS.n1647 0.2255
R24459 DVSS.n1647 DVSS.n1646 0.2255
R24460 DVSS.n1651 DVSS.n1650 0.2255
R24461 DVSS.n1650 DVSS.n1649 0.2255
R24462 DVSS.n1654 DVSS.n1653 0.2255
R24463 DVSS.n1653 DVSS.n1652 0.2255
R24464 DVSS.n1657 DVSS.n1656 0.2255
R24465 DVSS.n1656 DVSS.n1655 0.2255
R24466 DVSS.n1660 DVSS.n1659 0.2255
R24467 DVSS.n1659 DVSS.n1658 0.2255
R24468 DVSS.n1663 DVSS.n1662 0.2255
R24469 DVSS.n1662 DVSS.n1661 0.2255
R24470 DVSS.n1666 DVSS.n1665 0.2255
R24471 DVSS.n1665 DVSS.n1664 0.2255
R24472 DVSS.n1669 DVSS.n1668 0.2255
R24473 DVSS.n1668 DVSS.n1667 0.2255
R24474 DVSS.n1672 DVSS.n1671 0.2255
R24475 DVSS.n1671 DVSS.n1670 0.2255
R24476 DVSS.n1675 DVSS.n1674 0.2255
R24477 DVSS.n1674 DVSS.n1673 0.2255
R24478 DVSS.n1678 DVSS.n1677 0.2255
R24479 DVSS.n1677 DVSS.n1676 0.2255
R24480 DVSS.n1681 DVSS.n1680 0.2255
R24481 DVSS.n1680 DVSS.n1679 0.2255
R24482 DVSS.n1684 DVSS.n1683 0.2255
R24483 DVSS.n1683 DVSS.n1682 0.2255
R24484 DVSS.n1687 DVSS.n1686 0.2255
R24485 DVSS.n1686 DVSS.n1685 0.2255
R24486 DVSS.n1690 DVSS.n1689 0.2255
R24487 DVSS.n1689 DVSS.n1688 0.2255
R24488 DVSS.n1693 DVSS.n1692 0.2255
R24489 DVSS.n1692 DVSS.n1691 0.2255
R24490 DVSS.n1696 DVSS.n1695 0.2255
R24491 DVSS.n1695 DVSS.n1694 0.2255
R24492 DVSS.n1699 DVSS.n1698 0.2255
R24493 DVSS.n1698 DVSS.n1697 0.2255
R24494 DVSS.n1702 DVSS.n1701 0.2255
R24495 DVSS.n1701 DVSS.n1700 0.2255
R24496 DVSS.n1705 DVSS.n1704 0.2255
R24497 DVSS.n1704 DVSS.n1703 0.2255
R24498 DVSS.n1708 DVSS.n1707 0.2255
R24499 DVSS.n1707 DVSS.n1706 0.2255
R24500 DVSS.n1710 DVSS.n1709 0.2255
R24501 DVSS.n1711 DVSS.n1710 0.2255
R24502 DVSS.n1718 DVSS.n1717 0.2255
R24503 DVSS.n1717 DVSS.n1716 0.2255
R24504 DVSS.n1715 DVSS.n1714 0.2255
R24505 DVSS.n1713 DVSS.n1712 0.2255
R24506 DVSS.n1553 DVSS.n1552 0.2255
R24507 DVSS.n2435 DVSS.n2434 0.2255
R24508 DVSS.n2006 DVSS.n2005 0.2255
R24509 DVSS.n10652 DVSS.n10651 0.2255
R24510 DVSS.n10729 DVSS.n10728 0.2255
R24511 DVSS.n10730 DVSS.n10729 0.2255
R24512 DVSS.n10726 DVSS.n10725 0.2255
R24513 DVSS.n10725 DVSS.n10724 0.2255
R24514 DVSS.n4764 DVSS.n4763 0.2255
R24515 DVSS.n4752 DVSS.n4751 0.2255
R24516 DVSS.n4743 DVSS.n4742 0.2255
R24517 DVSS.n4731 DVSS.n4730 0.2255
R24518 DVSS.n10064 DVSS.n10063 0.2255
R24519 DVSS.n10075 DVSS.n10074 0.2255
R24520 DVSS.n10119 DVSS.n10118 0.2255
R24521 DVSS.n10128 DVSS.n10127 0.2255
R24522 DVSS.n10150 DVSS.n10149 0.2255
R24523 DVSS.n10163 DVSS.n10162 0.2255
R24524 DVSS.n10165 DVSS.n10164 0.2255
R24525 DVSS.n10167 DVSS.n10166 0.2255
R24526 DVSS.n10176 DVSS.n10175 0.2255
R24527 DVSS.n10188 DVSS.n10187 0.2255
R24528 DVSS.n10701 DVSS.n10700 0.2255
R24529 DVSS.n10710 DVSS.n10709 0.2255
R24530 DVSS.n10713 DVSS.n10712 0.2255
R24531 DVSS.n10715 DVSS.n10714 0.2255
R24532 DVSS.n10717 DVSS.n10716 0.2255
R24533 DVSS.n4838 DVSS.n4837 0.2255
R24534 DVSS.n4836 DVSS.n4835 0.2255
R24535 DVSS.n4834 DVSS.n4833 0.2255
R24536 DVSS.n4830 DVSS.n4829 0.2255
R24537 DVSS.n4828 DVSS.n4827 0.2255
R24538 DVSS.n4826 DVSS.n4825 0.2255
R24539 DVSS.n4824 DVSS.n4823 0.2255
R24540 DVSS.n4807 DVSS.n4806 0.2255
R24541 DVSS.n4796 DVSS.n4795 0.2255
R24542 DVSS.n4781 DVSS.n4780 0.2255
R24543 DVSS.n4942 DVSS.n4941 0.2255
R24544 DVSS.n4926 DVSS.n4925 0.2255
R24545 DVSS.n4914 DVSS.n4913 0.2255
R24546 DVSS.n4898 DVSS.n4897 0.2255
R24547 DVSS.n4882 DVSS.n4881 0.2255
R24548 DVSS.n4876 DVSS.n4875 0.2255
R24549 DVSS.n4866 DVSS.n4865 0.2255
R24550 DVSS.n4854 DVSS.n4853 0.2255
R24551 DVSS.n4845 DVSS.n4844 0.2255
R24552 DVSS.n4632 DVSS.n4631 0.2255
R24553 DVSS.n4643 DVSS.n4642 0.2255
R24554 DVSS.n4644 DVSS.n4643 0.2255
R24555 DVSS.n5055 DVSS.n5054 0.2255
R24556 DVSS.n5056 DVSS.n5055 0.2255
R24557 DVSS.n4986 DVSS.n4985 0.2255
R24558 DVSS.n4970 DVSS.n4969 0.2255
R24559 DVSS.n4958 DVSS.n4957 0.2255
R24560 DVSS.n13095 DVSS.n13094 0.2255
R24561 DVSS.n13102 DVSS.n13101 0.2255
R24562 DVSS.n13101 DVSS.n13100 0.2255
R24563 DVSS.n8321 DVSS.n8320 0.2255
R24564 DVSS.n8314 DVSS.n8313 0.2255
R24565 DVSS.n8312 DVSS.n8311 0.2255
R24566 DVSS.n8310 DVSS.n8309 0.2255
R24567 DVSS.n8308 DVSS.n8307 0.2255
R24568 DVSS.n8306 DVSS.n8305 0.2255
R24569 DVSS.n8301 DVSS.n8300 0.2255
R24570 DVSS.n13111 DVSS.n13110 0.2255
R24571 DVSS.n13112 DVSS.n13111 0.2255
R24572 DVSS.n8286 DVSS.n8285 0.2255
R24573 DVSS.n8287 DVSS.n8286 0.2255
R24574 DVSS.n8230 DVSS.n8229 0.2255
R24575 DVSS.n8228 DVSS.n8227 0.2255
R24576 DVSS.n8226 DVSS.n8225 0.2255
R24577 DVSS.n8224 DVSS.n8223 0.2255
R24578 DVSS.n8222 DVSS.n8221 0.2255
R24579 DVSS.n8216 DVSS.n8215 0.2255
R24580 DVSS.n8208 DVSS.n8207 0.2255
R24581 DVSS.n8201 DVSS.n8200 0.2255
R24582 DVSS.n8195 DVSS.n8194 0.2255
R24583 DVSS.n8193 DVSS.n8192 0.2255
R24584 DVSS.n8191 DVSS.n8190 0.2255
R24585 DVSS.n8189 DVSS.n8188 0.2255
R24586 DVSS.n8187 DVSS.n8186 0.2255
R24587 DVSS.n8185 DVSS.n8184 0.2255
R24588 DVSS.n8183 DVSS.n8182 0.2255
R24589 DVSS.n8181 DVSS.n8180 0.2255
R24590 DVSS.n8179 DVSS.n8178 0.2255
R24591 DVSS.n8177 DVSS.n8176 0.2255
R24592 DVSS.n8175 DVSS.n8174 0.2255
R24593 DVSS.n8173 DVSS.n8172 0.2255
R24594 DVSS.n8171 DVSS.n8170 0.2255
R24595 DVSS.n8165 DVSS.n8164 0.2255
R24596 DVSS.n8157 DVSS.n8156 0.2255
R24597 DVSS.n8150 DVSS.n8149 0.2255
R24598 DVSS.n8144 DVSS.n8143 0.2255
R24599 DVSS.n8142 DVSS.n8141 0.2255
R24600 DVSS.n8140 DVSS.n8139 0.2255
R24601 DVSS.n8138 DVSS.n8137 0.2255
R24602 DVSS.n8136 DVSS.n8135 0.2255
R24603 DVSS.n8134 DVSS.n8133 0.2255
R24604 DVSS.n8132 DVSS.n8131 0.2255
R24605 DVSS.n8130 DVSS.n8129 0.2255
R24606 DVSS.n8128 DVSS.n8127 0.2255
R24607 DVSS.n8126 DVSS.n8125 0.2255
R24608 DVSS.n8124 DVSS.n8123 0.2255
R24609 DVSS.n8122 DVSS.n8121 0.2255
R24610 DVSS.n8120 DVSS.n8119 0.2255
R24611 DVSS.n8115 DVSS.n8114 0.2255
R24612 DVSS.n8106 DVSS.n8105 0.2255
R24613 DVSS.n8095 DVSS.n8094 0.2255
R24614 DVSS.n6795 DVSS.n6793 0.2255
R24615 DVSS.n6796 DVSS.n6795 0.2255
R24616 DVSS.n6813 DVSS.n6812 0.2255
R24617 DVSS.n6814 DVSS.n6813 0.2255
R24618 DVSS.n6805 DVSS.n6804 0.2255
R24619 DVSS.n6802 DVSS.n6801 0.2255
R24620 DVSS.n6800 DVSS.n6799 0.2255
R24621 DVSS.n3808 DVSS.n3807 0.2255
R24622 DVSS.n3810 DVSS.n3809 0.2255
R24623 DVSS.n3812 DVSS.n3811 0.2255
R24624 DVSS.n3823 DVSS.n3821 0.2255
R24625 DVSS.n3824 DVSS.n3823 0.2255
R24626 DVSS.n3965 DVSS.n3964 0.2255
R24627 DVSS.n3966 DVSS.n3965 0.2255
R24628 DVSS.n3927 DVSS.n3926 0.2255
R24629 DVSS.n3924 DVSS.n3923 0.2255
R24630 DVSS.n3922 DVSS.n3921 0.2255
R24631 DVSS.n3920 DVSS.n3919 0.2255
R24632 DVSS.n3918 DVSS.n3917 0.2255
R24633 DVSS.n3916 DVSS.n3915 0.2255
R24634 DVSS.n3911 DVSS.n3910 0.2255
R24635 DVSS.n3902 DVSS.n3901 0.2255
R24636 DVSS.n3897 DVSS.n3896 0.2255
R24637 DVSS.n3894 DVSS.n3893 0.2255
R24638 DVSS.n3892 DVSS.n3891 0.2255
R24639 DVSS.n3890 DVSS.n3889 0.2255
R24640 DVSS.n3888 DVSS.n3887 0.2255
R24641 DVSS.n3886 DVSS.n3885 0.2255
R24642 DVSS.n3884 DVSS.n3883 0.2255
R24643 DVSS.n3882 DVSS.n3881 0.2255
R24644 DVSS.n3880 DVSS.n3879 0.2255
R24645 DVSS.n3878 DVSS.n3877 0.2255
R24646 DVSS.n3876 DVSS.n3875 0.2255
R24647 DVSS.n3874 DVSS.n3873 0.2255
R24648 DVSS.n3872 DVSS.n3871 0.2255
R24649 DVSS.n3870 DVSS.n3869 0.2255
R24650 DVSS.n3865 DVSS.n3864 0.2255
R24651 DVSS.n3856 DVSS.n3855 0.2255
R24652 DVSS.n3851 DVSS.n3850 0.2255
R24653 DVSS.n3848 DVSS.n3847 0.2255
R24654 DVSS.n3846 DVSS.n3845 0.2255
R24655 DVSS.n3844 DVSS.n3843 0.2255
R24656 DVSS.n3842 DVSS.n3841 0.2255
R24657 DVSS.n3840 DVSS.n3839 0.2255
R24658 DVSS.n3838 DVSS.n3837 0.2255
R24659 DVSS.n3836 DVSS.n3835 0.2255
R24660 DVSS.n3834 DVSS.n3833 0.2255
R24661 DVSS.n3828 DVSS.n3827 0.2255
R24662 DVSS.n8062 DVSS.n8061 0.2255
R24663 DVSS.n8064 DVSS.n8063 0.2255
R24664 DVSS.n8070 DVSS.n8069 0.2255
R24665 DVSS.n8079 DVSS.n8078 0.2255
R24666 DVSS.n8089 DVSS.n8088 0.2255
R24667 DVSS.n3612 DVSS.n3610 0.2255
R24668 DVSS.n13012 DVSS.n13011 0.2255
R24669 DVSS.n13021 DVSS.n13020 0.2255
R24670 DVSS.n13022 DVSS.n13021 0.2255
R24671 DVSS.n3613 DVSS.n3612 0.2255
R24672 DVSS.n3623 DVSS.n3622 0.2255
R24673 DVSS.n3624 DVSS.n3623 0.2255
R24674 DVSS.n3618 DVSS.n3617 0.2255
R24675 DVSS.n3616 DVSS.n3615 0.2255
R24676 DVSS.n2581 DVSS.n2580 0.2255
R24677 DVSS.n2583 DVSS.n2582 0.2255
R24678 DVSS.n2585 DVSS.n2584 0.2255
R24679 DVSS.n2592 DVSS.n2591 0.2255
R24680 DVSS.n2604 DVSS.n2603 0.2255
R24681 DVSS.n2605 DVSS.n2604 0.2255
R24682 DVSS.n2754 DVSS.n2753 0.2255
R24683 DVSS.n2755 DVSS.n2754 0.2255
R24684 DVSS.n2720 DVSS.n2719 0.2255
R24685 DVSS.n2718 DVSS.n2717 0.2255
R24686 DVSS.n2716 DVSS.n2715 0.2255
R24687 DVSS.n2714 DVSS.n2713 0.2255
R24688 DVSS.n2712 DVSS.n2711 0.2255
R24689 DVSS.n2705 DVSS.n2704 0.2255
R24690 DVSS.n2694 DVSS.n2693 0.2255
R24691 DVSS.n2687 DVSS.n2686 0.2255
R24692 DVSS.n2682 DVSS.n2681 0.2255
R24693 DVSS.n2680 DVSS.n2679 0.2255
R24694 DVSS.n2678 DVSS.n2677 0.2255
R24695 DVSS.n2676 DVSS.n2675 0.2255
R24696 DVSS.n2674 DVSS.n2673 0.2255
R24697 DVSS.n2672 DVSS.n2671 0.2255
R24698 DVSS.n2670 DVSS.n2669 0.2255
R24699 DVSS.n2668 DVSS.n2667 0.2255
R24700 DVSS.n2666 DVSS.n2665 0.2255
R24701 DVSS.n2664 DVSS.n2663 0.2255
R24702 DVSS.n2662 DVSS.n2661 0.2255
R24703 DVSS.n2660 DVSS.n2659 0.2255
R24704 DVSS.n2658 DVSS.n2657 0.2255
R24705 DVSS.n2651 DVSS.n2650 0.2255
R24706 DVSS.n2640 DVSS.n2639 0.2255
R24707 DVSS.n2633 DVSS.n2632 0.2255
R24708 DVSS.n2628 DVSS.n2627 0.2255
R24709 DVSS.n2626 DVSS.n2625 0.2255
R24710 DVSS.n2624 DVSS.n2623 0.2255
R24711 DVSS.n2622 DVSS.n2621 0.2255
R24712 DVSS.n2620 DVSS.n2619 0.2255
R24713 DVSS.n2618 DVSS.n2617 0.2255
R24714 DVSS.n2616 DVSS.n2615 0.2255
R24715 DVSS.n2614 DVSS.n2613 0.2255
R24716 DVSS.n2612 DVSS.n2611 0.2255
R24717 DVSS.n2610 DVSS.n2609 0.2255
R24718 DVSS.n2608 DVSS.n2607 0.2255
R24719 DVSS.n11739 DVSS.n11738 0.2255
R24720 DVSS.n11741 DVSS.n11740 0.2255
R24721 DVSS.n11749 DVSS.n11748 0.2255
R24722 DVSS.n11758 DVSS.n11757 0.2255
R24723 DVSS.n11767 DVSS.n11766 0.2255
R24724 DVSS.n11773 DVSS.n11772 0.2255
R24725 DVSS.n11783 DVSS.n11782 0.2255
R24726 DVSS.n11792 DVSS.n11791 0.2255
R24727 DVSS.n11799 DVSS.n11798 0.2255
R24728 DVSS.n11801 DVSS.n11800 0.2255
R24729 DVSS.n11803 DVSS.n11802 0.2255
R24730 DVSS.n11805 DVSS.n11804 0.2255
R24731 DVSS.n11807 DVSS.n11806 0.2255
R24732 DVSS.n11809 DVSS.n11808 0.2255
R24733 DVSS.n11811 DVSS.n11810 0.2255
R24734 DVSS.n11813 DVSS.n11812 0.2255
R24735 DVSS.n11815 DVSS.n11814 0.2255
R24736 DVSS.n11817 DVSS.n11816 0.2255
R24737 DVSS.n11819 DVSS.n11818 0.2255
R24738 DVSS.n11821 DVSS.n11820 0.2255
R24739 DVSS.n11823 DVSS.n11822 0.2255
R24740 DVSS.n11832 DVSS.n11831 0.2255
R24741 DVSS.n11840 DVSS.n11839 0.2255
R24742 DVSS.n11850 DVSS.n11849 0.2255
R24743 DVSS.n11858 DVSS.n11857 0.2255
R24744 DVSS.n11860 DVSS.n11859 0.2255
R24745 DVSS.n11862 DVSS.n11861 0.2255
R24746 DVSS.n11864 DVSS.n11863 0.2255
R24747 DVSS.n11866 DVSS.n11865 0.2255
R24748 DVSS.n11868 DVSS.n11867 0.2255
R24749 DVSS.n11870 DVSS.n11869 0.2255
R24750 DVSS.n11872 DVSS.n11871 0.2255
R24751 DVSS.n11874 DVSS.n11873 0.2255
R24752 DVSS.n11876 DVSS.n11875 0.2255
R24753 DVSS.n11878 DVSS.n11877 0.2255
R24754 DVSS.n11880 DVSS.n11879 0.2255
R24755 DVSS.n11882 DVSS.n11881 0.2255
R24756 DVSS.n11891 DVSS.n11890 0.2255
R24757 DVSS.n11899 DVSS.n11898 0.2255
R24758 DVSS.n11909 DVSS.n11908 0.2255
R24759 DVSS.n11917 DVSS.n11916 0.2255
R24760 DVSS.n11919 DVSS.n11918 0.2255
R24761 DVSS.n11921 DVSS.n11920 0.2255
R24762 DVSS.n11923 DVSS.n11922 0.2255
R24763 DVSS.n11925 DVSS.n11924 0.2255
R24764 DVSS.n11981 DVSS.n11980 0.2255
R24765 DVSS.n11982 DVSS.n11981 0.2255
R24766 DVSS.n12994 DVSS.n12993 0.2255
R24767 DVSS.n12993 DVSS.n12992 0.2255
R24768 DVSS.n12987 DVSS.n12986 0.2255
R24769 DVSS.n12980 DVSS.n12979 0.2255
R24770 DVSS.n12978 DVSS.n12977 0.2255
R24771 DVSS.n12976 DVSS.n12975 0.2255
R24772 DVSS.n12974 DVSS.n12973 0.2255
R24773 DVSS.n12972 DVSS.n12971 0.2255
R24774 DVSS.n13002 DVSS.n13001 0.2255
R24775 DVSS.n13003 DVSS.n13002 0.2255
R24776 DVSS.n3603 DVSS.n3602 0.2255
R24777 DVSS.n5910 DVSS.n5909 0.2255
R24778 DVSS.n6046 DVSS.n5910 0.2255
R24779 DVSS.n6041 DVSS.n6040 0.2255
R24780 DVSS.n6036 DVSS.n6035 0.2255
R24781 DVSS.n6034 DVSS.n6033 0.2255
R24782 DVSS.n6030 DVSS.n6029 0.2255
R24783 DVSS.n6028 DVSS.n6027 0.2255
R24784 DVSS.n6024 DVSS.n6023 0.2255
R24785 DVSS.n6006 DVSS.n6005 0.2255
R24786 DVSS.n6004 DVSS.n6003 0.2255
R24787 DVSS.n6002 DVSS.n6001 0.2255
R24788 DVSS.n6000 DVSS.n5999 0.2255
R24789 DVSS.n5998 DVSS.n5997 0.2255
R24790 DVSS.n5996 DVSS.n5995 0.2255
R24791 DVSS.n5994 DVSS.n5993 0.2255
R24792 DVSS.n5989 DVSS.n5988 0.2255
R24793 DVSS.n5980 DVSS.n5979 0.2255
R24794 DVSS.n5975 DVSS.n5974 0.2255
R24795 DVSS.n5972 DVSS.n5971 0.2255
R24796 DVSS.n5970 DVSS.n5969 0.2255
R24797 DVSS.n5966 DVSS.n5965 0.2255
R24798 DVSS.n5964 DVSS.n5963 0.2255
R24799 DVSS.n5962 DVSS.n5961 0.2255
R24800 DVSS.n5960 DVSS.n5959 0.2255
R24801 DVSS.n5958 DVSS.n5957 0.2255
R24802 DVSS.n5956 DVSS.n5955 0.2255
R24803 DVSS.n5954 DVSS.n5953 0.2255
R24804 DVSS.n5952 DVSS.n5951 0.2255
R24805 DVSS.n5950 DVSS.n5949 0.2255
R24806 DVSS.n5948 DVSS.n5947 0.2255
R24807 DVSS.n5943 DVSS.n5942 0.2255
R24808 DVSS.n5934 DVSS.n5933 0.2255
R24809 DVSS.n5929 DVSS.n5928 0.2255
R24810 DVSS.n5926 DVSS.n5925 0.2255
R24811 DVSS.n5922 DVSS.n5921 0.2255
R24812 DVSS.n5920 DVSS.n5919 0.2255
R24813 DVSS.n5918 DVSS.n5917 0.2255
R24814 DVSS.n5916 DVSS.n5915 0.2255
R24815 DVSS.n8344 DVSS.n8343 0.2255
R24816 DVSS.n8346 DVSS.n8345 0.2255
R24817 DVSS.n8348 DVSS.n8347 0.2255
R24818 DVSS.n8350 DVSS.n8349 0.2255
R24819 DVSS.n8352 DVSS.n8351 0.2255
R24820 DVSS.n8354 DVSS.n8353 0.2255
R24821 DVSS.n8356 DVSS.n8355 0.2255
R24822 DVSS.n8362 DVSS.n8361 0.2255
R24823 DVSS.n8371 DVSS.n8370 0.2255
R24824 DVSS.n8381 DVSS.n8380 0.2255
R24825 DVSS.n8387 DVSS.n8386 0.2255
R24826 DVSS.n8398 DVSS.n8397 0.2255
R24827 DVSS.n8407 DVSS.n8406 0.2255
R24828 DVSS.n8412 DVSS.n8411 0.2255
R24829 DVSS.n8414 DVSS.n8413 0.2255
R24830 DVSS.n8416 DVSS.n8415 0.2255
R24831 DVSS.n8418 DVSS.n8417 0.2255
R24832 DVSS.n8420 DVSS.n8419 0.2255
R24833 DVSS.n8422 DVSS.n8421 0.2255
R24834 DVSS.n8424 DVSS.n8423 0.2255
R24835 DVSS.n8426 DVSS.n8425 0.2255
R24836 DVSS.n8430 DVSS.n8429 0.2255
R24837 DVSS.n8432 DVSS.n8431 0.2255
R24838 DVSS.n8434 DVSS.n8433 0.2255
R24839 DVSS.n8436 DVSS.n8435 0.2255
R24840 DVSS.n8442 DVSS.n8441 0.2255
R24841 DVSS.n8449 DVSS.n8448 0.2255
R24842 DVSS.n8457 DVSS.n8456 0.2255
R24843 DVSS.n8463 DVSS.n8462 0.2255
R24844 DVSS.n8465 DVSS.n8464 0.2255
R24845 DVSS.n8467 DVSS.n8466 0.2255
R24846 DVSS.n8469 DVSS.n8468 0.2255
R24847 DVSS.n8471 DVSS.n8470 0.2255
R24848 DVSS.n8473 DVSS.n8472 0.2255
R24849 DVSS.n8475 DVSS.n8474 0.2255
R24850 DVSS.n8479 DVSS.n8478 0.2255
R24851 DVSS.n8481 DVSS.n8480 0.2255
R24852 DVSS.n8483 DVSS.n8482 0.2255
R24853 DVSS.n8487 DVSS.n8486 0.2255
R24854 DVSS.n8493 DVSS.n8492 0.2255
R24855 DVSS.n8500 DVSS.n8499 0.2255
R24856 DVSS.n8508 DVSS.n8507 0.2255
R24857 DVSS.n8514 DVSS.n8513 0.2255
R24858 DVSS.n8516 DVSS.n8515 0.2255
R24859 DVSS.n8518 DVSS.n8517 0.2255
R24860 DVSS.n8520 DVSS.n8519 0.2255
R24861 DVSS.n8522 DVSS.n8521 0.2255
R24862 DVSS.n8583 DVSS.n8582 0.2255
R24863 DVSS.n8584 DVSS.n8583 0.2255
R24864 DVSS.n11328 DVSS.n11327 0.2255
R24865 DVSS.n11327 DVSS.n11326 0.2255
R24866 DVSS.n11321 DVSS.n11320 0.2255
R24867 DVSS.n11314 DVSS.n11313 0.2255
R24868 DVSS.n11312 DVSS.n11311 0.2255
R24869 DVSS.n11308 DVSS.n11307 0.2255
R24870 DVSS.n11306 DVSS.n11305 0.2255
R24871 DVSS.n11336 DVSS.n11335 0.2255
R24872 DVSS.n11337 DVSS.n11336 0.2255
R24873 DVSS.n11358 DVSS.n11357 0.2255
R24874 DVSS.n11359 DVSS.n11358 0.2255
R24875 DVSS.n11347 DVSS.n11346 0.2255
R24876 DVSS.n5867 DVSS.n5866 0.2255
R24877 DVSS.n5868 DVSS.n5867 0.2255
R24878 DVSS.n8331 DVSS.n8330 0.2255
R24879 DVSS.n8332 DVSS.n8331 0.2255
R24880 DVSS.n8909 DVSS.n8907 0.2255
R24881 DVSS.n8910 DVSS.n8909 0.2255
R24882 DVSS.n8899 DVSS.n8898 0.2255
R24883 DVSS.n6094 DVSS.n6092 0.2255
R24884 DVSS.n6095 DVSS.n6094 0.2255
R24885 DVSS.n6106 DVSS.n6105 0.2255
R24886 DVSS.n6105 DVSS.n6104 0.2255
R24887 DVSS.n6323 DVSS.n6322 0.2255
R24888 DVSS.n6324 DVSS.n6323 0.2255
R24889 DVSS.n6284 DVSS.n6283 0.2255
R24890 DVSS.n6261 DVSS.n6260 0.2255
R24891 DVSS.n6242 DVSS.n6241 0.2255
R24892 DVSS.n6231 DVSS.n6230 0.2255
R24893 DVSS.n6215 DVSS.n6214 0.2255
R24894 DVSS.n6207 DVSS.n6206 0.2255
R24895 DVSS.n6203 DVSS.n6202 0.2255
R24896 DVSS.n6201 DVSS.n6200 0.2255
R24897 DVSS.n6199 DVSS.n6198 0.2255
R24898 DVSS.n6197 DVSS.n6196 0.2255
R24899 DVSS.n6195 DVSS.n6194 0.2255
R24900 DVSS.n6191 DVSS.n6190 0.2255
R24901 DVSS.n6184 DVSS.n6183 0.2255
R24902 DVSS.n6173 DVSS.n6172 0.2255
R24903 DVSS.n6157 DVSS.n6156 0.2255
R24904 DVSS.n6151 DVSS.n6150 0.2255
R24905 DVSS.n6147 DVSS.n6146 0.2255
R24906 DVSS.n8590 DVSS.n8589 0.2255
R24907 DVSS.n8594 DVSS.n8593 0.2255
R24908 DVSS.n8596 DVSS.n8595 0.2255
R24909 DVSS.n8598 DVSS.n8597 0.2255
R24910 DVSS.n8600 DVSS.n8599 0.2255
R24911 DVSS.n8607 DVSS.n8606 0.2255
R24912 DVSS.n8619 DVSS.n8618 0.2255
R24913 DVSS.n8631 DVSS.n8630 0.2255
R24914 DVSS.n8637 DVSS.n8636 0.2255
R24915 DVSS.n8649 DVSS.n8648 0.2255
R24916 DVSS.n8660 DVSS.n8659 0.2255
R24917 DVSS.n8666 DVSS.n8665 0.2255
R24918 DVSS.n8668 DVSS.n8667 0.2255
R24919 DVSS.n8672 DVSS.n8671 0.2255
R24920 DVSS.n8674 DVSS.n8673 0.2255
R24921 DVSS.n8676 DVSS.n8675 0.2255
R24922 DVSS.n8678 DVSS.n8677 0.2255
R24923 DVSS.n8686 DVSS.n8685 0.2255
R24924 DVSS.n8690 DVSS.n8689 0.2255
R24925 DVSS.n8709 DVSS.n8708 0.2255
R24926 DVSS.n8719 DVSS.n8718 0.2255
R24927 DVSS.n8749 DVSS.n8748 0.2255
R24928 DVSS.n8751 DVSS.n8750 0.2255
R24929 DVSS.n8759 DVSS.n8758 0.2255
R24930 DVSS.n8770 DVSS.n8769 0.2255
R24931 DVSS.n8780 DVSS.n8779 0.2255
R24932 DVSS.n8790 DVSS.n8789 0.2255
R24933 DVSS.n8792 DVSS.n8791 0.2255
R24934 DVSS.n8794 DVSS.n8793 0.2255
R24935 DVSS.n8796 DVSS.n8795 0.2255
R24936 DVSS.n8860 DVSS.n8859 0.2255
R24937 DVSS.n8859 DVSS.n8858 0.2255
R24938 DVSS.n8920 DVSS.n8918 0.2255
R24939 DVSS.n8921 DVSS.n8920 0.2255
R24940 DVSS.n8875 DVSS.n8874 0.2255
R24941 DVSS.n8882 DVSS.n8881 0.2255
R24942 DVSS.n8884 DVSS.n8883 0.2255
R24943 DVSS.n8886 DVSS.n8885 0.2255
R24944 DVSS.n8888 DVSS.n8887 0.2255
R24945 DVSS.n8890 DVSS.n8889 0.2255
R24946 DVSS.n13844 DVSS.n13843 0.225323
R24947 DVSS.n18580 DVSS.n18579 0.225323
R24948 DVSS.n18616 DVSS.n18615 0.222388
R24949 DVSS.n18642 DVSS.n18640 0.222388
R24950 DVSS.n18674 DVSS.n18673 0.222388
R24951 DVSS.n18808 DVSS.n18807 0.222388
R24952 DVSS.n14075 DVSS.n14072 0.222388
R24953 DVSS.n7803 DVSS.n7801 0.222149
R24954 DVSS.n7813 DVSS.n7811 0.222149
R24955 DVSS.n7825 DVSS.n7822 0.222149
R24956 DVSS.n14072 DVSS.n14069 0.222149
R24957 DVSS.n7322 DVSS.n7319 0.220713
R24958 DVSS.n7990 DVSS.n7987 0.220713
R24959 DVSS.n7993 DVSS.n7990 0.220713
R24960 DVSS.n14648 DVSS.n14647 0.220473
R24961 DVSS.n14485 DVSS.n14484 0.220234
R24962 DVSS.n14159 DVSS.n14158 0.220234
R24963 DVSS.n14158 DVSS.n14156 0.219516
R24964 DVSS.n13599 DVSS.n13598 0.219277
R24965 DVSS.n7296 DVSS.n7295 0.21784
R24966 DVSS.n7953 DVSS.n7952 0.21784
R24967 DVSS.n7070 DVSS.n7069 0.21784
R24968 DVSS.n7069 DVSS.n7067 0.21784
R24969 DVSS.n13621 DVSS.n13620 0.21784
R24970 DVSS.n2484 DVSS.n2483 0.216246
R24971 DVSS.n2487 DVSS.n2486 0.216246
R24972 DVSS.n2493 DVSS.n2492 0.216246
R24973 DVSS.n2496 DVSS.n2495 0.216246
R24974 DVSS.n2514 DVSS.n2506 0.216246
R24975 DVSS.n2517 DVSS.n2516 0.216246
R24976 DVSS.n2523 DVSS.n2522 0.216246
R24977 DVSS.n2526 DVSS.n2525 0.216246
R24978 DVSS.n2472 DVSS.n2471 0.216246
R24979 DVSS.n14453 DVSS.n14452 0.214725
R24980 DVSS.n14669 DVSS.n14668 0.214725
R24981 DVSS.n1325 DVSS.n1317 0.208878
R24982 DVSS.n1322 DVSS.n1321 0.208878
R24983 DVSS.n13338 DVSS.n13337 0.208878
R24984 DVSS.n13337 DVSS.n13335 0.208878
R24985 DVSS.n13335 DVSS.n13334 0.208878
R24986 DVSS.n1325 DVSS.n1324 0.208878
R24987 DVSS.n1324 DVSS.n1322 0.208878
R24988 DVSS.n13327 DVSS.n13292 0.208878
R24989 DVSS.n13330 DVSS.n13327 0.208878
R24990 DVSS.n13338 DVSS.n13330 0.208878
R24991 DVSS.n7023 DVSS.n7022 0.208878
R24992 DVSS.n7409 DVSS.n7408 0.199888
R24993 DVSS.n13811 DVSS.n13810 0.199888
R24994 DVSS.n7388 DVSS.n7387 0.199888
R24995 DVSS.n13771 DVSS.n13770 0.199888
R24996 DVSS.n7361 DVSS.n7360 0.199888
R24997 DVSS.n13731 DVSS.n13730 0.199888
R24998 DVSS.n1169 DVSS.n1168 0.185308
R24999 DVSS.n19741 DVSS.n19729 0.185115
R25000 DVSS.n20227 DVSS.n20224 0.185115
R25001 DVSS.n20730 DVSS.n20727 0.185115
R25002 DVSS.n19506 DVSS.n19485 0.183192
R25003 DVSS.n20519 DVSS.n20495 0.183192
R25004 DVSS.n1192 DVSS.n1186 0.183192
R25005 DVSS.n20717 DVSS.n20716 0.183192
R25006 DVSS.n7141 DVSS.n7140 0.180146
R25007 DVSS.n13552 DVSS.n13551 0.180146
R25008 DVSS.n13362 DVSS.n13361 0.180146
R25009 DVSS.n18823 DVSS.n18822 0.180146
R25010 DVSS.n13815 DVSS.n13814 0.168293
R25011 DVSS.n13776 DVSS.n13774 0.168293
R25012 DVSS.n13739 DVSS.n13736 0.168293
R25013 DVSS.n7414 DVSS.n7412 0.168053
R25014 DVSS.n7393 DVSS.n7391 0.168053
R25015 DVSS.n7369 DVSS.n7366 0.168053
R25016 DVSS.n7436 DVSS.n7434 0.137763
R25017 DVSS.n14947 DVSS.n14944 0.137763
R25018 DVSS.n18566 DVSS 0.136254
R25019 DVSS.n14929 DVSS 0.136254
R25020 DVSS.n14427 DVSS.n14426 0.136134
R25021 DVSS.n14701 DVSS.n14700 0.136134
R25022 DVSS.n17547 DVSS.n17545 0.133972
R25023 DVSS.n14959 DVSS.n14957 0.133972
R25024 DVSS.n15588 DVSS.n15586 0.133972
R25025 DVSS.n15730 DVSS.n15729 0.133972
R25026 DVSS.n17663 DVSS.n17661 0.133972
R25027 DVSS.n15834 DVSS.n15832 0.133972
R25028 DVSS.n15054 DVSS.n15053 0.133972
R25029 DVSS.n17108 DVSS.n17107 0.133972
R25030 DVSS.n17455 DVSS.n17451 0.133833
R25031 DVSS.n18406 DVSS.n18403 0.133833
R25032 DVSS.n18368 DVSS.n18366 0.133833
R25033 DVSS.n16239 DVSS.n16237 0.133833
R25034 DVSS.n16338 DVSS.n16336 0.133833
R25035 DVSS.n16278 DVSS.n16276 0.133833
R25036 DVSS.n7490 DVSS.n7488 0.133833
R25037 DVSS.n17246 DVSS.n17244 0.133833
R25038 DVSS.n14367 DVSS.n14366 0.13381
R25039 DVSS.n14783 DVSS.n14782 0.13381
R25040 DVSS.n11075 DVSS.n11070 0.132444
R25041 DVSS.n9008 DVSS.n9005 0.132444
R25042 DVSS.n8966 DVSS.n8963 0.132444
R25043 DVSS.n8958 DVSS.n8955 0.132444
R25044 DVSS.n9819 DVSS.n9816 0.132444
R25045 DVSS.n8933 DVSS.n8930 0.132444
R25046 DVSS.n9856 DVSS.n9853 0.132444
R25047 DVSS.n14265 DVSS.n14264 0.128739
R25048 DVSS.n14290 DVSS.n14289 0.128739
R25049 DVSS.n14850 DVSS.n14849 0.128739
R25050 DVSS.n14833 DVSS.n14832 0.128739
R25051 DVSS.n14240 DVSS.n14239 0.128106
R25052 DVSS.n14867 DVSS.n14866 0.128106
R25053 DVSS.n14319 DVSS.n14318 0.127894
R25054 DVSS.n14816 DVSS.n14815 0.127894
R25055 DVSS.n2456 DVSS.n2455 0.120204
R25056 DVSS.n2019 DVSS.n2018 0.120204
R25057 DVSS.n1721 DVSS.n1720 0.116325
R25058 DVSS.n2052 VSS 0.115811
R25059 DVSS.n11689 DVSS.n11688 0.114949
R25060 DVSS.n6772 DVSS.n6771 0.114949
R25061 DVSS.n7112 DVSS.n7111 0.11424
R25062 DVSS.n13569 DVSS.n13568 0.11424
R25063 DVSS.n13263 DVSS.n13262 0.11424
R25064 DVSS.n18791 DVSS.n18790 0.11424
R25065 DVSS.n6970 DVSS.n6969 0.112291
R25066 DVSS.n13670 DVSS.n13669 0.112291
R25067 DVSS.n13205 DVSS.n13204 0.112291
R25068 DVSS.n18737 DVSS.n18736 0.112291
R25069 DVSS.n1380 DVSS.n1379 0.110613
R25070 DVSS.n21373 DVSS.n21372 0.110523
R25071 DVSS.n13968 DVSS.t25 0.1097
R25072 DVSS.n16803 DVSS.t28 0.1097
R25073 DVSS.n15071 DVSS.t4 0.1097
R25074 DVSS.n7641 DVSS.t1 0.1097
R25075 DVSS.n16010 DVSS.t23 0.1097
R25076 DVSS.n15307 DVSS.t17 0.1097
R25077 DVSS.n18352 DVSS.t30 0.1097
R25078 DVSS.n18009 DVSS.t21 0.1097
R25079 DVSS.n17868 DVSS.t35 0.1097
R25080 DVSS.n3528 DVSS.n3518 0.109536
R25081 DVSS.n12026 DVSS.n12017 0.109536
R25082 DVSS.n18929 DVSS.n18920 0.109536
R25083 DVSS.n13 DVSS.n3 0.109536
R25084 DVSS.n514 DVSS.n505 0.109536
R25085 DVSS.n4082 DVSS.n4081 0.10928
R25086 DVSS.n9003 DVSS.n9002 0.10928
R25087 DVSS.n14992 DVSS.n14991 0.10928
R25088 DVSS.n3791 DVSS.n2559 0.10928
R25089 DVSS.n9093 DVSS.n9092 0.10928
R25090 DVSS.n7547 DVSS.n7546 0.10928
R25091 DVSS.n17438 DVSS.n17435 0.108278
R25092 DVSS.n16892 DVSS.n16890 0.108278
R25093 DVSS.n7466 DVSS.n7463 0.108278
R25094 DVSS.n14975 DVSS.n14974 0.108278
R25095 DVSS.n7555 DVSS.n7552 0.108278
R25096 DVSS.n15604 DVSS.n15603 0.108278
R25097 DVSS.n16227 DVSS.n16224 0.108278
R25098 DVSS.n7691 DVSS.n7690 0.108278
R25099 DVSS.n16310 DVSS.n16308 0.108278
R25100 DVSS.n17644 DVSS.n17643 0.108278
R25101 DVSS.n16266 DVSS.n16263 0.108278
R25102 DVSS.n15850 DVSS.n15849 0.108278
R25103 DVSS.n7476 DVSS.n7473 0.108278
R25104 DVSS.n7781 DVSS.n7780 0.108278
R25105 DVSS.n16430 DVSS.n16428 0.108278
R25106 DVSS.n16881 DVSS.n16880 0.108278
R25107 DVSS.n13791 DVSS.n13790 0.108039
R25108 DVSS.n13754 DVSS.n13753 0.108039
R25109 DVSS.n18630 DVSS.n18629 0.108039
R25110 DVSS.n18657 DVSS.n18656 0.108039
R25111 DVSS.n1386 DVSS.n1385 0.107643
R25112 DVSS.n9440 DVSS.n9439 0.107643
R25113 DVSS.n9447 DVSS.n9446 0.107643
R25114 DVSS.n9446 DVSS.n9445 0.107643
R25115 DVSS.n4233 DVSS.n4232 0.107643
R25116 DVSS.n4231 DVSS.n4230 0.107643
R25117 DVSS.n4229 DVSS.n4228 0.107643
R25118 DVSS.n4227 DVSS.n4226 0.107643
R25119 DVSS.n4225 DVSS.n4224 0.107643
R25120 DVSS.n4219 DVSS.n4218 0.107643
R25121 DVSS.n4211 DVSS.n4210 0.107643
R25122 DVSS.n4205 DVSS.n4204 0.107643
R25123 DVSS.n4202 DVSS.n4201 0.107643
R25124 DVSS.n4200 DVSS.n4199 0.107643
R25125 DVSS.n4198 DVSS.n4197 0.107643
R25126 DVSS.n4194 DVSS.n4193 0.107643
R25127 DVSS.n4190 DVSS.n4189 0.107643
R25128 DVSS.n4186 DVSS.n4185 0.107643
R25129 DVSS.n4184 DVSS.n4183 0.107643
R25130 DVSS.n4180 DVSS.n4179 0.107643
R25131 DVSS.n4178 DVSS.n4177 0.107643
R25132 DVSS.n4173 DVSS.n4172 0.107643
R25133 DVSS.n4165 DVSS.n4164 0.107643
R25134 DVSS.n4156 DVSS.n4155 0.107643
R25135 DVSS.n4154 DVSS.n4153 0.107643
R25136 DVSS.n4152 DVSS.n4151 0.107643
R25137 DVSS.n4150 DVSS.n4149 0.107643
R25138 DVSS.n4148 DVSS.n4147 0.107643
R25139 DVSS.n9153 DVSS.n9152 0.107643
R25140 DVSS.n9155 DVSS.n9154 0.107643
R25141 DVSS.n9157 DVSS.n9156 0.107643
R25142 DVSS.n9159 DVSS.n9158 0.107643
R25143 DVSS.n9161 DVSS.n9160 0.107643
R25144 DVSS.n9163 DVSS.n9162 0.107643
R25145 DVSS.n9165 DVSS.n9164 0.107643
R25146 DVSS.n9167 DVSS.n9166 0.107643
R25147 DVSS.n9175 DVSS.n9174 0.107643
R25148 DVSS.n9184 DVSS.n9183 0.107643
R25149 DVSS.n9194 DVSS.n9193 0.107643
R25150 DVSS.n9201 DVSS.n9200 0.107643
R25151 DVSS.n9212 DVSS.n9211 0.107643
R25152 DVSS.n9221 DVSS.n9220 0.107643
R25153 DVSS.n9227 DVSS.n9226 0.107643
R25154 DVSS.n9229 DVSS.n9228 0.107643
R25155 DVSS.n9231 DVSS.n9230 0.107643
R25156 DVSS.n9233 DVSS.n9232 0.107643
R25157 DVSS.n9237 DVSS.n9236 0.107643
R25158 DVSS.n9239 DVSS.n9238 0.107643
R25159 DVSS.n9241 DVSS.n9240 0.107643
R25160 DVSS.n9243 DVSS.n9242 0.107643
R25161 DVSS.n9245 DVSS.n9244 0.107643
R25162 DVSS.n9247 DVSS.n9246 0.107643
R25163 DVSS.n9249 DVSS.n9248 0.107643
R25164 DVSS.n9251 DVSS.n9250 0.107643
R25165 DVSS.n9257 DVSS.n9256 0.107643
R25166 DVSS.n9265 DVSS.n9264 0.107643
R25167 DVSS.n9273 DVSS.n9272 0.107643
R25168 DVSS.n9279 DVSS.n9278 0.107643
R25169 DVSS.n9281 DVSS.n9280 0.107643
R25170 DVSS.n9283 DVSS.n9282 0.107643
R25171 DVSS.n9285 DVSS.n9284 0.107643
R25172 DVSS.n9287 DVSS.n9286 0.107643
R25173 DVSS.n9289 DVSS.n9288 0.107643
R25174 DVSS.n9291 DVSS.n9290 0.107643
R25175 DVSS.n9293 DVSS.n9292 0.107643
R25176 DVSS.n9295 DVSS.n9294 0.107643
R25177 DVSS.n9301 DVSS.n9300 0.107643
R25178 DVSS.n9303 DVSS.n9302 0.107643
R25179 DVSS.n9310 DVSS.n9309 0.107643
R25180 DVSS.n9318 DVSS.n9317 0.107643
R25181 DVSS.n9326 DVSS.n9325 0.107643
R25182 DVSS.n9331 DVSS.n9330 0.107643
R25183 DVSS.n9333 DVSS.n9332 0.107643
R25184 DVSS.n9335 DVSS.n9334 0.107643
R25185 DVSS.n9337 DVSS.n9336 0.107643
R25186 DVSS.n9339 DVSS.n9338 0.107643
R25187 DVSS.n9422 DVSS.n9421 0.107643
R25188 DVSS.n9423 DVSS.n9422 0.107643
R25189 DVSS.n9485 DVSS.n9484 0.107643
R25190 DVSS.n9486 DVSS.n9485 0.107643
R25191 DVSS.n9455 DVSS.n9454 0.107643
R25192 DVSS.n9461 DVSS.n9460 0.107643
R25193 DVSS.n9463 DVSS.n9462 0.107643
R25194 DVSS.n9465 DVSS.n9464 0.107643
R25195 DVSS.n9476 DVSS.n9475 0.107643
R25196 DVSS.n9478 DVSS.n9477 0.107643
R25197 DVSS.n9470 DVSS.n9469 0.107643
R25198 DVSS.n1399 DVSS.n1398 0.107643
R25199 DVSS.n1393 DVSS.n1392 0.107643
R25200 DVSS.n1390 DVSS.n1389 0.107643
R25201 DVSS.n4131 DVSS.n4130 0.107643
R25202 DVSS.n4133 DVSS.n4132 0.107643
R25203 DVSS.n4137 DVSS.n4136 0.107643
R25204 DVSS.n4144 DVSS.n4143 0.107643
R25205 DVSS.n4256 DVSS.n4255 0.107643
R25206 DVSS.n4257 DVSS.n4256 0.107643
R25207 DVSS.n4236 DVSS.n4235 0.107643
R25208 DVSS.n18890 DVSS.n18889 0.107643
R25209 DVSS.n18891 DVSS.n18890 0.107643
R25210 DVSS.n12025 DVSS.n12023 0.107643
R25211 DVSS.n12026 DVSS.n12025 0.107643
R25212 DVSS.n12118 DVSS.n12117 0.107643
R25213 DVSS.n12117 DVSS.n12116 0.107643
R25214 DVSS.n12114 DVSS.n12013 0.107643
R25215 DVSS.n12115 DVSS.n12114 0.107643
R25216 DVSS.n12113 DVSS.n12015 0.107643
R25217 DVSS.n12113 DVSS.n12112 0.107643
R25218 DVSS.n12109 DVSS.n12108 0.107643
R25219 DVSS.n12110 DVSS.n12109 0.107643
R25220 DVSS.n12106 DVSS.n12104 0.107643
R25221 DVSS.n12107 DVSS.n12106 0.107643
R25222 DVSS.n12097 DVSS.n12096 0.107643
R25223 DVSS.n12096 DVSS.n12095 0.107643
R25224 DVSS.n12122 DVSS.n12121 0.107643
R25225 DVSS.n12124 DVSS.n12123 0.107643
R25226 DVSS.n12125 DVSS.n12124 0.107643
R25227 DVSS.n12011 DVSS.n12009 0.107643
R25228 DVSS.n12012 DVSS.n12011 0.107643
R25229 DVSS.n12001 DVSS.n12000 0.107643
R25230 DVSS.n12000 DVSS.n11999 0.107643
R25231 DVSS.n11995 DVSS.n11994 0.107643
R25232 DVSS.n11994 DVSS.n11993 0.107643
R25233 DVSS.n11992 DVSS.n11991 0.107643
R25234 DVSS.n11991 DVSS.n11990 0.107643
R25235 DVSS.n11989 DVSS.n11988 0.107643
R25236 DVSS.n11988 DVSS.n11987 0.107643
R25237 DVSS.n7913 DVSS.n7912 0.107643
R25238 DVSS.n7912 DVSS.n7911 0.107643
R25239 DVSS.n13499 DVSS.n13498 0.107643
R25240 DVSS.n13500 DVSS.n13499 0.107643
R25241 DVSS.n13496 DVSS.n13494 0.107643
R25242 DVSS.n13497 DVSS.n13496 0.107643
R25243 DVSS.n13484 DVSS.n13483 0.107643
R25244 DVSS.n13483 DVSS.n13482 0.107643
R25245 DVSS.n7944 DVSS.n7942 0.107643
R25246 DVSS.n7945 DVSS.n7944 0.107643
R25247 DVSS.n7930 DVSS.n7929 0.107643
R25248 DVSS.n7929 DVSS.n7928 0.107643
R25249 DVSS.n7908 DVSS.n7907 0.107643
R25250 DVSS.n7907 DVSS.n7906 0.107643
R25251 DVSS.n7905 DVSS.n7904 0.107643
R25252 DVSS.n7904 DVSS.n7903 0.107643
R25253 DVSS.n7902 DVSS.n7901 0.107643
R25254 DVSS.n7901 DVSS.n7900 0.107643
R25255 DVSS.n7899 DVSS.n7898 0.107643
R25256 DVSS.n7898 DVSS.n7897 0.107643
R25257 DVSS.n14540 DVSS.n14539 0.107643
R25258 DVSS.n14539 DVSS.n14538 0.107643
R25259 DVSS.n14543 DVSS.n14542 0.107643
R25260 DVSS.n14542 DVSS.n14541 0.107643
R25261 DVSS.n14546 DVSS.n14545 0.107643
R25262 DVSS.n14545 DVSS.n14544 0.107643
R25263 DVSS.n14549 DVSS.n14548 0.107643
R25264 DVSS.n14548 DVSS.n14547 0.107643
R25265 DVSS.n14552 DVSS.n14551 0.107643
R25266 DVSS.n14551 DVSS.n14550 0.107643
R25267 DVSS.n14555 DVSS.n14554 0.107643
R25268 DVSS.n14554 DVSS.n14553 0.107643
R25269 DVSS.n14558 DVSS.n14557 0.107643
R25270 DVSS.n14557 DVSS.n14556 0.107643
R25271 DVSS.n14561 DVSS.n14560 0.107643
R25272 DVSS.n14560 DVSS.n14559 0.107643
R25273 DVSS.n14564 DVSS.n14563 0.107643
R25274 DVSS.n14563 DVSS.n14562 0.107643
R25275 DVSS.n14581 DVSS.n14580 0.107643
R25276 DVSS.n14580 DVSS.n14579 0.107643
R25277 DVSS.n13464 DVSS.n13463 0.107643
R25278 DVSS.n13465 DVSS.n13464 0.107643
R25279 DVSS.n13462 DVSS.n13461 0.107643
R25280 DVSS.n13461 DVSS.n13460 0.107643
R25281 DVSS.n13458 DVSS.n13457 0.107643
R25282 DVSS.n13459 DVSS.n13458 0.107643
R25283 DVSS.n13456 DVSS.n13455 0.107643
R25284 DVSS.n13455 DVSS.n13454 0.107643
R25285 DVSS.n13452 DVSS.n13451 0.107643
R25286 DVSS.n13453 DVSS.n13452 0.107643
R25287 DVSS.n13450 DVSS.n13449 0.107643
R25288 DVSS.n13449 DVSS.n13448 0.107643
R25289 DVSS.n13446 DVSS.n13445 0.107643
R25290 DVSS.n13447 DVSS.n13446 0.107643
R25291 DVSS.n13444 DVSS.n13443 0.107643
R25292 DVSS.n13443 DVSS.n13442 0.107643
R25293 DVSS.n13440 DVSS.n13439 0.107643
R25294 DVSS.n13441 DVSS.n13440 0.107643
R25295 DVSS.n13438 DVSS.n13437 0.107643
R25296 DVSS.n13437 DVSS.n13436 0.107643
R25297 DVSS.n13434 DVSS.n13433 0.107643
R25298 DVSS.n13435 DVSS.n13434 0.107643
R25299 DVSS.n13432 DVSS.n13431 0.107643
R25300 DVSS.n13431 DVSS.n13430 0.107643
R25301 DVSS.n13428 DVSS.n13427 0.107643
R25302 DVSS.n13429 DVSS.n13428 0.107643
R25303 DVSS.n13426 DVSS.n13425 0.107643
R25304 DVSS.n13425 DVSS.n13424 0.107643
R25305 DVSS.n14591 DVSS.n14589 0.107643
R25306 DVSS.n14592 DVSS.n14591 0.107643
R25307 DVSS.n14594 DVSS.n14593 0.107643
R25308 DVSS.n14595 DVSS.n14594 0.107643
R25309 DVSS.n14534 DVSS.n14532 0.107643
R25310 DVSS.n14535 DVSS.n14534 0.107643
R25311 DVSS.n14134 DVSS.n14133 0.107643
R25312 DVSS.n14133 DVSS.n14132 0.107643
R25313 DVSS.n14115 DVSS.n14114 0.107643
R25314 DVSS.n14111 DVSS.n14110 0.107643
R25315 DVSS.n14110 DVSS.n14109 0.107643
R25316 DVSS.n14107 DVSS.n14106 0.107643
R25317 DVSS.n14108 DVSS.n14107 0.107643
R25318 DVSS.n14105 DVSS.n14104 0.107643
R25319 DVSS.n14104 DVSS.n14103 0.107643
R25320 DVSS.n14101 DVSS.n14100 0.107643
R25321 DVSS.n14102 DVSS.n14101 0.107643
R25322 DVSS.n14099 DVSS.n14098 0.107643
R25323 DVSS.n14098 DVSS.n14097 0.107643
R25324 DVSS.n14095 DVSS.n14094 0.107643
R25325 DVSS.n14096 DVSS.n14095 0.107643
R25326 DVSS.n14093 DVSS.n14092 0.107643
R25327 DVSS.n14092 DVSS.n14091 0.107643
R25328 DVSS.n14089 DVSS.n14088 0.107643
R25329 DVSS.n14090 DVSS.n14089 0.107643
R25330 DVSS.n14087 DVSS.n14086 0.107643
R25331 DVSS.n14086 DVSS.n14085 0.107643
R25332 DVSS.n18917 DVSS.n18915 0.107643
R25333 DVSS.n18918 DVSS.n18917 0.107643
R25334 DVSS.n18913 DVSS.n18912 0.107643
R25335 DVSS.n18912 DVSS.n18911 0.107643
R25336 DVSS.n18909 DVSS.n18908 0.107643
R25337 DVSS.n18910 DVSS.n18909 0.107643
R25338 DVSS.n18907 DVSS.n18906 0.107643
R25339 DVSS.n18906 DVSS.n18905 0.107643
R25340 DVSS.n18893 DVSS.n18892 0.107643
R25341 DVSS.n7288 DVSS.n7287 0.107643
R25342 DVSS.n7283 DVSS.n7282 0.107643
R25343 DVSS.n7284 DVSS.n7283 0.107643
R25344 DVSS.n7281 DVSS.n7280 0.107643
R25345 DVSS.n7280 DVSS.n7279 0.107643
R25346 DVSS.n7277 DVSS.n7276 0.107643
R25347 DVSS.n7278 DVSS.n7277 0.107643
R25348 DVSS.n7275 DVSS.n7274 0.107643
R25349 DVSS.n7274 DVSS.n7273 0.107643
R25350 DVSS.n7271 DVSS.n7270 0.107643
R25351 DVSS.n7272 DVSS.n7271 0.107643
R25352 DVSS.n7269 DVSS.n7268 0.107643
R25353 DVSS.n7268 DVSS.n7267 0.107643
R25354 DVSS.n7265 DVSS.n7264 0.107643
R25355 DVSS.n7266 DVSS.n7265 0.107643
R25356 DVSS.n7263 DVSS.n7262 0.107643
R25357 DVSS.n7262 DVSS.n7261 0.107643
R25358 DVSS.n7259 DVSS.n7258 0.107643
R25359 DVSS.n7260 DVSS.n7259 0.107643
R25360 DVSS.n7257 DVSS.n7256 0.107643
R25361 DVSS.n7256 DVSS.n7255 0.107643
R25362 DVSS.n7253 DVSS.n7252 0.107643
R25363 DVSS.n7254 DVSS.n7253 0.107643
R25364 DVSS.n7251 DVSS.n7250 0.107643
R25365 DVSS.n7250 DVSS.n7249 0.107643
R25366 DVSS.n7247 DVSS.n7246 0.107643
R25367 DVSS.n7248 DVSS.n7247 0.107643
R25368 DVSS.n7234 DVSS.n7233 0.107643
R25369 DVSS.n7231 DVSS.n7229 0.107643
R25370 DVSS.n7232 DVSS.n7231 0.107643
R25371 DVSS.n3723 DVSS.n3722 0.107643
R25372 DVSS.n3722 DVSS.n3721 0.107643
R25373 DVSS.n3716 DVSS.n3715 0.107643
R25374 DVSS.n3717 DVSS.n3716 0.107643
R25375 DVSS.n3711 DVSS.n3710 0.107643
R25376 DVSS.n3710 DVSS.n3709 0.107643
R25377 DVSS.n3707 DVSS.n3706 0.107643
R25378 DVSS.n3708 DVSS.n3707 0.107643
R25379 DVSS.n3705 DVSS.n3704 0.107643
R25380 DVSS.n3704 DVSS.n3703 0.107643
R25381 DVSS.n3700 DVSS.n3699 0.107643
R25382 DVSS.n3701 DVSS.n3700 0.107643
R25383 DVSS.n1306 DVSS.n1305 0.107643
R25384 DVSS.n3527 DVSS.n3525 0.107643
R25385 DVSS.n3528 DVSS.n3527 0.107643
R25386 DVSS.n3666 DVSS.n3665 0.107643
R25387 DVSS.n3665 DVSS.n3664 0.107643
R25388 DVSS.n3669 DVSS.n3668 0.107643
R25389 DVSS.n3670 DVSS.n3669 0.107643
R25390 DVSS.n3674 DVSS.n3673 0.107643
R25391 DVSS.n3673 DVSS.n3672 0.107643
R25392 DVSS.n3676 DVSS.n3675 0.107643
R25393 DVSS.n3677 DVSS.n3676 0.107643
R25394 DVSS.n3680 DVSS.n3679 0.107643
R25395 DVSS.n3679 DVSS.n3678 0.107643
R25396 DVSS.n3682 DVSS.n3681 0.107643
R25397 DVSS.n3683 DVSS.n3682 0.107643
R25398 DVSS.n3686 DVSS.n3685 0.107643
R25399 DVSS.n3685 DVSS.n3684 0.107643
R25400 DVSS.n3695 DVSS.n3693 0.107643
R25401 DVSS.n3696 DVSS.n3695 0.107643
R25402 DVSS.n3725 DVSS.n3724 0.107643
R25403 DVSS.n3726 DVSS.n3725 0.107643
R25404 DVSS.n19849 DVSS.n19847 0.107643
R25405 DVSS.n19850 DVSS.n19849 0.107643
R25406 DVSS.n20049 DVSS.n20048 0.107643
R25407 DVSS.n20048 DVSS.n20047 0.107643
R25408 DVSS.n20051 DVSS.n20050 0.107643
R25409 DVSS.n20052 DVSS.n20051 0.107643
R25410 DVSS.n20055 DVSS.n20054 0.107643
R25411 DVSS.n20054 DVSS.n20053 0.107643
R25412 DVSS.n20057 DVSS.n20056 0.107643
R25413 DVSS.n20058 DVSS.n20057 0.107643
R25414 DVSS.n20061 DVSS.n20060 0.107643
R25415 DVSS.n20060 DVSS.n20059 0.107643
R25416 DVSS.n20063 DVSS.n20062 0.107643
R25417 DVSS.n20064 DVSS.n20063 0.107643
R25418 DVSS.n20067 DVSS.n20066 0.107643
R25419 DVSS.n20066 DVSS.n20065 0.107643
R25420 DVSS.n20069 DVSS.n20068 0.107643
R25421 DVSS.n20070 DVSS.n20069 0.107643
R25422 DVSS.n20073 DVSS.n20072 0.107643
R25423 DVSS.n20072 DVSS.n20071 0.107643
R25424 DVSS.n20077 DVSS.n20075 0.107643
R25425 DVSS.n20078 DVSS.n20077 0.107643
R25426 DVSS.n20082 DVSS.n20081 0.107643
R25427 DVSS.n20081 DVSS.n20080 0.107643
R25428 DVSS.n20084 DVSS.n20083 0.107643
R25429 DVSS.n20085 DVSS.n20084 0.107643
R25430 DVSS.n20088 DVSS.n20087 0.107643
R25431 DVSS.n20087 DVSS.n20086 0.107643
R25432 DVSS.n20090 DVSS.n20089 0.107643
R25433 DVSS.n20091 DVSS.n20090 0.107643
R25434 DVSS.n20102 DVSS.n20101 0.107643
R25435 DVSS.n20101 DVSS.n20100 0.107643
R25436 DVSS.n20111 DVSS.n20109 0.107643
R25437 DVSS.n20112 DVSS.n20111 0.107643
R25438 DVSS.n20329 DVSS.n20328 0.107643
R25439 DVSS.n20328 DVSS.n20327 0.107643
R25440 DVSS.n20331 DVSS.n20330 0.107643
R25441 DVSS.n20332 DVSS.n20331 0.107643
R25442 DVSS.n20335 DVSS.n20334 0.107643
R25443 DVSS.n20334 DVSS.n20333 0.107643
R25444 DVSS.n20337 DVSS.n20336 0.107643
R25445 DVSS.n20338 DVSS.n20337 0.107643
R25446 DVSS.n20341 DVSS.n20340 0.107643
R25447 DVSS.n20340 DVSS.n20339 0.107643
R25448 DVSS.n20343 DVSS.n20342 0.107643
R25449 DVSS.n20344 DVSS.n20343 0.107643
R25450 DVSS.n20347 DVSS.n20346 0.107643
R25451 DVSS.n20346 DVSS.n20345 0.107643
R25452 DVSS.n20349 DVSS.n20348 0.107643
R25453 DVSS.n20350 DVSS.n20349 0.107643
R25454 DVSS.n20353 DVSS.n20352 0.107643
R25455 DVSS.n20352 DVSS.n20351 0.107643
R25456 DVSS.n20355 DVSS.n20354 0.107643
R25457 DVSS.n20356 DVSS.n20355 0.107643
R25458 DVSS.n20359 DVSS.n20358 0.107643
R25459 DVSS.n20358 DVSS.n20357 0.107643
R25460 DVSS.n20361 DVSS.n20360 0.107643
R25461 DVSS.n20362 DVSS.n20361 0.107643
R25462 DVSS.n20365 DVSS.n20364 0.107643
R25463 DVSS.n20364 DVSS.n20363 0.107643
R25464 DVSS.n20367 DVSS.n20366 0.107643
R25465 DVSS.n20379 DVSS.n20378 0.107643
R25466 DVSS.n20378 DVSS.n20377 0.107643
R25467 DVSS.n20597 DVSS.n20595 0.107643
R25468 DVSS.n20598 DVSS.n20597 0.107643
R25469 DVSS.n20614 DVSS.n20613 0.107643
R25470 DVSS.n20613 DVSS.n20612 0.107643
R25471 DVSS.n20618 DVSS.n20616 0.107643
R25472 DVSS.n20619 DVSS.n20618 0.107643
R25473 DVSS.n20672 DVSS.n20671 0.107643
R25474 DVSS.n20671 DVSS.n20670 0.107643
R25475 DVSS.n20668 DVSS.n20667 0.107643
R25476 DVSS.n20669 DVSS.n20668 0.107643
R25477 DVSS.n20666 DVSS.n20665 0.107643
R25478 DVSS.n20665 DVSS.n20664 0.107643
R25479 DVSS.n20662 DVSS.n20661 0.107643
R25480 DVSS.n20663 DVSS.n20662 0.107643
R25481 DVSS.n20660 DVSS.n20659 0.107643
R25482 DVSS.n20659 DVSS.n20658 0.107643
R25483 DVSS.n20648 DVSS.n20646 0.107643
R25484 DVSS.n20649 DVSS.n20648 0.107643
R25485 DVSS.n20636 DVSS.n20635 0.107643
R25486 DVSS.n20635 DVSS.n20634 0.107643
R25487 DVSS.n20624 DVSS.n20623 0.107643
R25488 DVSS.n20625 DVSS.n20624 0.107643
R25489 DVSS.n20622 DVSS.n20621 0.107643
R25490 DVSS.n20621 DVSS.n20620 0.107643
R25491 DVSS.n1 DVSS.n0 0.107643
R25492 DVSS.n2 DVSS.n1 0.107643
R25493 DVSS.n21578 DVSS.n21577 0.107643
R25494 DVSS.n21577 DVSS.n21576 0.107643
R25495 DVSS.n21574 DVSS.n21564 0.107643
R25496 DVSS.n21575 DVSS.n21574 0.107643
R25497 DVSS.n21572 DVSS.n21563 0.107643
R25498 DVSS.n21572 DVSS.n21571 0.107643
R25499 DVSS.n21561 DVSS.n21559 0.107643
R25500 DVSS.n21562 DVSS.n21561 0.107643
R25501 DVSS.n13 DVSS.n12 0.107643
R25502 DVSS.n12 DVSS.n11 0.107643
R25503 DVSS.n19838 DVSS.n19836 0.107643
R25504 DVSS.n19839 DVSS.n19838 0.107643
R25505 DVSS.n19581 DVSS.n19580 0.107643
R25506 DVSS.n19582 DVSS.n19581 0.107643
R25507 DVSS.n19585 DVSS.n19584 0.107643
R25508 DVSS.n19584 DVSS.n19583 0.107643
R25509 DVSS.n19587 DVSS.n19586 0.107643
R25510 DVSS.n19588 DVSS.n19587 0.107643
R25511 DVSS.n19593 DVSS.n19592 0.107643
R25512 DVSS.n19592 DVSS.n19591 0.107643
R25513 DVSS.n19596 DVSS.n19595 0.107643
R25514 DVSS.n19597 DVSS.n19596 0.107643
R25515 DVSS.n19600 DVSS.n19599 0.107643
R25516 DVSS.n19599 DVSS.n19598 0.107643
R25517 DVSS.n19602 DVSS.n19601 0.107643
R25518 DVSS.n19603 DVSS.n19602 0.107643
R25519 DVSS.n19606 DVSS.n19605 0.107643
R25520 DVSS.n19605 DVSS.n19604 0.107643
R25521 DVSS.n19608 DVSS.n19607 0.107643
R25522 DVSS.n19609 DVSS.n19608 0.107643
R25523 DVSS.n19612 DVSS.n19611 0.107643
R25524 DVSS.n19611 DVSS.n19610 0.107643
R25525 DVSS.n19614 DVSS.n19613 0.107643
R25526 DVSS.n19615 DVSS.n19614 0.107643
R25527 DVSS.n19618 DVSS.n19617 0.107643
R25528 DVSS.n19617 DVSS.n19616 0.107643
R25529 DVSS.n19620 DVSS.n19619 0.107643
R25530 DVSS.n19621 DVSS.n19620 0.107643
R25531 DVSS.n19631 DVSS.n19630 0.107643
R25532 DVSS.n19630 DVSS.n19629 0.107643
R25533 DVSS.n19817 DVSS.n19815 0.107643
R25534 DVSS.n19818 DVSS.n19817 0.107643
R25535 DVSS.n19831 DVSS.n19830 0.107643
R25536 DVSS.n19830 DVSS.n19829 0.107643
R25537 DVSS.n18929 DVSS.n18928 0.107643
R25538 DVSS.n18928 DVSS.n18927 0.107643
R25539 DVSS.n18937 DVSS.n18935 0.107643
R25540 DVSS.n18938 DVSS.n18937 0.107643
R25541 DVSS.n19023 DVSS.n19022 0.107643
R25542 DVSS.n19022 DVSS.n19021 0.107643
R25543 DVSS.n19026 DVSS.n19025 0.107643
R25544 DVSS.n19027 DVSS.n19026 0.107643
R25545 DVSS.n19030 DVSS.n19029 0.107643
R25546 DVSS.n19029 DVSS.n19028 0.107643
R25547 DVSS.n19032 DVSS.n19031 0.107643
R25548 DVSS.n19033 DVSS.n19032 0.107643
R25549 DVSS.n19036 DVSS.n19035 0.107643
R25550 DVSS.n19035 DVSS.n19034 0.107643
R25551 DVSS.n19038 DVSS.n19037 0.107643
R25552 DVSS.n19039 DVSS.n19038 0.107643
R25553 DVSS.n19049 DVSS.n19048 0.107643
R25554 DVSS.n19048 DVSS.n19047 0.107643
R25555 DVSS.n19059 DVSS.n19057 0.107643
R25556 DVSS.n19060 DVSS.n19059 0.107643
R25557 DVSS.n19066 DVSS.n19065 0.107643
R25558 DVSS.n19065 DVSS.n19064 0.107643
R25559 DVSS.n19071 DVSS.n19070 0.107643
R25560 DVSS.n19072 DVSS.n19071 0.107643
R25561 DVSS.n19075 DVSS.n19074 0.107643
R25562 DVSS.n19074 DVSS.n19073 0.107643
R25563 DVSS.n19077 DVSS.n19076 0.107643
R25564 DVSS.n19078 DVSS.n19077 0.107643
R25565 DVSS.n19081 DVSS.n19080 0.107643
R25566 DVSS.n19080 DVSS.n19079 0.107643
R25567 DVSS.n19086 DVSS.n19085 0.107643
R25568 DVSS.n19087 DVSS.n19086 0.107643
R25569 DVSS.n19091 DVSS.n19090 0.107643
R25570 DVSS.n19306 DVSS.n19304 0.107643
R25571 DVSS.n19307 DVSS.n19306 0.107643
R25572 DVSS.n19314 DVSS.n19313 0.107643
R25573 DVSS.n19313 DVSS.n19312 0.107643
R25574 DVSS.n19316 DVSS.n19315 0.107643
R25575 DVSS.n19317 DVSS.n19316 0.107643
R25576 DVSS.n19320 DVSS.n19319 0.107643
R25577 DVSS.n19319 DVSS.n19318 0.107643
R25578 DVSS.n19322 DVSS.n19321 0.107643
R25579 DVSS.n19323 DVSS.n19322 0.107643
R25580 DVSS.n19326 DVSS.n19325 0.107643
R25581 DVSS.n19325 DVSS.n19324 0.107643
R25582 DVSS.n19328 DVSS.n19327 0.107643
R25583 DVSS.n19329 DVSS.n19328 0.107643
R25584 DVSS.n19332 DVSS.n19331 0.107643
R25585 DVSS.n19331 DVSS.n19330 0.107643
R25586 DVSS.n19334 DVSS.n19333 0.107643
R25587 DVSS.n19335 DVSS.n19334 0.107643
R25588 DVSS.n19338 DVSS.n19337 0.107643
R25589 DVSS.n19337 DVSS.n19336 0.107643
R25590 DVSS.n19340 DVSS.n19339 0.107643
R25591 DVSS.n19341 DVSS.n19340 0.107643
R25592 DVSS.n19344 DVSS.n19343 0.107643
R25593 DVSS.n19343 DVSS.n19342 0.107643
R25594 DVSS.n19346 DVSS.n19345 0.107643
R25595 DVSS.n19347 DVSS.n19346 0.107643
R25596 DVSS.n19350 DVSS.n19349 0.107643
R25597 DVSS.n19349 DVSS.n19348 0.107643
R25598 DVSS.n19352 DVSS.n19351 0.107643
R25599 DVSS.n19353 DVSS.n19352 0.107643
R25600 DVSS.n19357 DVSS.n19356 0.107643
R25601 DVSS.n19375 DVSS.n19373 0.107643
R25602 DVSS.n19376 DVSS.n19375 0.107643
R25603 DVSS.n19576 DVSS.n19575 0.107643
R25604 DVSS.n19575 DVSS.n19574 0.107643
R25605 DVSS.n21380 DVSS.n21379 0.107643
R25606 DVSS.n627 DVSS.n625 0.107643
R25607 DVSS.n628 DVSS.n627 0.107643
R25608 DVSS.n632 DVSS.n631 0.107643
R25609 DVSS.n631 DVSS.n630 0.107643
R25610 DVSS.n635 DVSS.n634 0.107643
R25611 DVSS.n636 DVSS.n635 0.107643
R25612 DVSS.n639 DVSS.n638 0.107643
R25613 DVSS.n638 DVSS.n637 0.107643
R25614 DVSS.n641 DVSS.n640 0.107643
R25615 DVSS.n642 DVSS.n641 0.107643
R25616 DVSS.n645 DVSS.n644 0.107643
R25617 DVSS.n644 DVSS.n643 0.107643
R25618 DVSS.n647 DVSS.n646 0.107643
R25619 DVSS.n648 DVSS.n647 0.107643
R25620 DVSS.n684 DVSS.n683 0.107643
R25621 DVSS.n683 DVSS.n682 0.107643
R25622 DVSS.n724 DVSS.n722 0.107643
R25623 DVSS.n725 DVSS.n724 0.107643
R25624 DVSS.n795 DVSS.n794 0.107643
R25625 DVSS.n794 DVSS.n793 0.107643
R25626 DVSS.n808 DVSS.n807 0.107643
R25627 DVSS.n809 DVSS.n808 0.107643
R25628 DVSS.n812 DVSS.n811 0.107643
R25629 DVSS.n811 DVSS.n810 0.107643
R25630 DVSS.n814 DVSS.n813 0.107643
R25631 DVSS.n815 DVSS.n814 0.107643
R25632 DVSS.n818 DVSS.n817 0.107643
R25633 DVSS.n817 DVSS.n816 0.107643
R25634 DVSS.n823 DVSS.n822 0.107643
R25635 DVSS.n824 DVSS.n823 0.107643
R25636 DVSS.n828 DVSS.n827 0.107643
R25637 DVSS.n1062 DVSS.n1060 0.107643
R25638 DVSS.n1063 DVSS.n1062 0.107643
R25639 DVSS.n1069 DVSS.n1068 0.107643
R25640 DVSS.n1068 DVSS.n1067 0.107643
R25641 DVSS.n1074 DVSS.n1073 0.107643
R25642 DVSS.n1075 DVSS.n1074 0.107643
R25643 DVSS.n1078 DVSS.n1077 0.107643
R25644 DVSS.n1077 DVSS.n1076 0.107643
R25645 DVSS.n1080 DVSS.n1079 0.107643
R25646 DVSS.n1081 DVSS.n1080 0.107643
R25647 DVSS.n1084 DVSS.n1083 0.107643
R25648 DVSS.n1083 DVSS.n1082 0.107643
R25649 DVSS.n1086 DVSS.n1085 0.107643
R25650 DVSS.n1087 DVSS.n1086 0.107643
R25651 DVSS.n1090 DVSS.n1089 0.107643
R25652 DVSS.n1089 DVSS.n1088 0.107643
R25653 DVSS.n1092 DVSS.n1091 0.107643
R25654 DVSS.n1093 DVSS.n1092 0.107643
R25655 DVSS.n1096 DVSS.n1095 0.107643
R25656 DVSS.n1095 DVSS.n1094 0.107643
R25657 DVSS.n1098 DVSS.n1097 0.107643
R25658 DVSS.n1099 DVSS.n1098 0.107643
R25659 DVSS.n1102 DVSS.n1101 0.107643
R25660 DVSS.n1101 DVSS.n1100 0.107643
R25661 DVSS.n1104 DVSS.n1103 0.107643
R25662 DVSS.n1105 DVSS.n1104 0.107643
R25663 DVSS.n1108 DVSS.n1107 0.107643
R25664 DVSS.n1107 DVSS.n1106 0.107643
R25665 DVSS.n1110 DVSS.n1109 0.107643
R25666 DVSS.n1111 DVSS.n1110 0.107643
R25667 DVSS.n1115 DVSS.n1114 0.107643
R25668 DVSS.n1277 DVSS.n1275 0.107643
R25669 DVSS.n1278 DVSS.n1277 0.107643
R25670 DVSS.n1284 DVSS.n1283 0.107643
R25671 DVSS.n1283 DVSS.n1282 0.107643
R25672 DVSS.n1289 DVSS.n1288 0.107643
R25673 DVSS.n1290 DVSS.n1289 0.107643
R25674 DVSS.n1293 DVSS.n1292 0.107643
R25675 DVSS.n1292 DVSS.n1291 0.107643
R25676 DVSS.n1295 DVSS.n1294 0.107643
R25677 DVSS.n1296 DVSS.n1295 0.107643
R25678 DVSS.n1301 DVSS.n1300 0.107643
R25679 DVSS.n1300 DVSS.n1299 0.107643
R25680 DVSS.n83 DVSS.n82 0.107643
R25681 DVSS.n84 DVSS.n83 0.107643
R25682 DVSS.n87 DVSS.n86 0.107643
R25683 DVSS.n86 DVSS.n85 0.107643
R25684 DVSS.n89 DVSS.n88 0.107643
R25685 DVSS.n90 DVSS.n89 0.107643
R25686 DVSS.n93 DVSS.n92 0.107643
R25687 DVSS.n92 DVSS.n91 0.107643
R25688 DVSS.n95 DVSS.n94 0.107643
R25689 DVSS.n96 DVSS.n95 0.107643
R25690 DVSS.n99 DVSS.n98 0.107643
R25691 DVSS.n98 DVSS.n97 0.107643
R25692 DVSS.n101 DVSS.n100 0.107643
R25693 DVSS.n102 DVSS.n101 0.107643
R25694 DVSS.n105 DVSS.n104 0.107643
R25695 DVSS.n104 DVSS.n103 0.107643
R25696 DVSS.n107 DVSS.n106 0.107643
R25697 DVSS.n108 DVSS.n107 0.107643
R25698 DVSS.n118 DVSS.n117 0.107643
R25699 DVSS.n117 DVSS.n116 0.107643
R25700 DVSS.n122 DVSS.n121 0.107643
R25701 DVSS.n267 DVSS.n266 0.107643
R25702 DVSS.n266 DVSS.n265 0.107643
R25703 DVSS.n274 DVSS.n272 0.107643
R25704 DVSS.n275 DVSS.n274 0.107643
R25705 DVSS.n286 DVSS.n285 0.107643
R25706 DVSS.n285 DVSS.n284 0.107643
R25707 DVSS.n473 DVSS.n471 0.107643
R25708 DVSS.n474 DVSS.n473 0.107643
R25709 DVSS.n477 DVSS.n476 0.107643
R25710 DVSS.n476 DVSS.n475 0.107643
R25711 DVSS.n479 DVSS.n478 0.107643
R25712 DVSS.n480 DVSS.n479 0.107643
R25713 DVSS.n483 DVSS.n482 0.107643
R25714 DVSS.n482 DVSS.n481 0.107643
R25715 DVSS.n485 DVSS.n484 0.107643
R25716 DVSS.n486 DVSS.n485 0.107643
R25717 DVSS.n489 DVSS.n488 0.107643
R25718 DVSS.n488 DVSS.n487 0.107643
R25719 DVSS.n491 DVSS.n490 0.107643
R25720 DVSS.n492 DVSS.n491 0.107643
R25721 DVSS.n495 DVSS.n494 0.107643
R25722 DVSS.n494 DVSS.n493 0.107643
R25723 DVSS.n497 DVSS.n496 0.107643
R25724 DVSS.n498 DVSS.n497 0.107643
R25725 DVSS.n503 DVSS.n502 0.107643
R25726 DVSS.n502 DVSS.n501 0.107643
R25727 DVSS.n20675 DVSS.n20674 0.107643
R25728 DVSS.n20676 DVSS.n20675 0.107643
R25729 DVSS.n20679 DVSS.n20678 0.107643
R25730 DVSS.n20678 DVSS.n20677 0.107643
R25731 DVSS.n20681 DVSS.n20680 0.107643
R25732 DVSS.n20682 DVSS.n20681 0.107643
R25733 DVSS.n20684 DVSS.n20683 0.107643
R25734 DVSS.n20695 DVSS.n20693 0.107643
R25735 DVSS.n20696 DVSS.n20695 0.107643
R25736 DVSS.n20707 DVSS.n20706 0.107643
R25737 DVSS.n20706 DVSS.n20705 0.107643
R25738 DVSS.n20874 DVSS.n20872 0.107643
R25739 DVSS.n20875 DVSS.n20874 0.107643
R25740 DVSS.n20878 DVSS.n20877 0.107643
R25741 DVSS.n20877 DVSS.n20876 0.107643
R25742 DVSS.n20880 DVSS.n20879 0.107643
R25743 DVSS.n20881 DVSS.n20880 0.107643
R25744 DVSS.n20884 DVSS.n20883 0.107643
R25745 DVSS.n20883 DVSS.n20882 0.107643
R25746 DVSS.n20886 DVSS.n20885 0.107643
R25747 DVSS.n20887 DVSS.n20886 0.107643
R25748 DVSS.n20890 DVSS.n20889 0.107643
R25749 DVSS.n20889 DVSS.n20888 0.107643
R25750 DVSS.n20892 DVSS.n20891 0.107643
R25751 DVSS.n20893 DVSS.n20892 0.107643
R25752 DVSS.n20896 DVSS.n20895 0.107643
R25753 DVSS.n20895 DVSS.n20894 0.107643
R25754 DVSS.n20898 DVSS.n20897 0.107643
R25755 DVSS.n20899 DVSS.n20898 0.107643
R25756 DVSS.n20902 DVSS.n20901 0.107643
R25757 DVSS.n20901 DVSS.n20900 0.107643
R25758 DVSS.n20904 DVSS.n20903 0.107643
R25759 DVSS.n20905 DVSS.n20904 0.107643
R25760 DVSS.n20908 DVSS.n20907 0.107643
R25761 DVSS.n20907 DVSS.n20906 0.107643
R25762 DVSS.n20910 DVSS.n20909 0.107643
R25763 DVSS.n20911 DVSS.n20910 0.107643
R25764 DVSS.n20914 DVSS.n20913 0.107643
R25765 DVSS.n20913 DVSS.n20912 0.107643
R25766 DVSS.n20924 DVSS.n20922 0.107643
R25767 DVSS.n20925 DVSS.n20924 0.107643
R25768 DVSS.n20936 DVSS.n20935 0.107643
R25769 DVSS.n20935 DVSS.n20934 0.107643
R25770 DVSS.n21100 DVSS.n21098 0.107643
R25771 DVSS.n21101 DVSS.n21100 0.107643
R25772 DVSS.n21106 DVSS.n21105 0.107643
R25773 DVSS.n21105 DVSS.n21104 0.107643
R25774 DVSS.n21109 DVSS.n21108 0.107643
R25775 DVSS.n21110 DVSS.n21109 0.107643
R25776 DVSS.n21113 DVSS.n21112 0.107643
R25777 DVSS.n21112 DVSS.n21111 0.107643
R25778 DVSS.n21115 DVSS.n21114 0.107643
R25779 DVSS.n21116 DVSS.n21115 0.107643
R25780 DVSS.n21121 DVSS.n21120 0.107643
R25781 DVSS.n21120 DVSS.n21119 0.107643
R25782 DVSS.n21258 DVSS.n21256 0.107643
R25783 DVSS.n21259 DVSS.n21258 0.107643
R25784 DVSS.n21274 DVSS.n21273 0.107643
R25785 DVSS.n21273 DVSS.n21272 0.107643
R25786 DVSS.n21349 DVSS.n21347 0.107643
R25787 DVSS.n21350 DVSS.n21349 0.107643
R25788 DVSS.n21353 DVSS.n21352 0.107643
R25789 DVSS.n21352 DVSS.n21351 0.107643
R25790 DVSS.n21355 DVSS.n21354 0.107643
R25791 DVSS.n21356 DVSS.n21355 0.107643
R25792 DVSS.n21359 DVSS.n21358 0.107643
R25793 DVSS.n21358 DVSS.n21357 0.107643
R25794 DVSS.n21365 DVSS.n21360 0.107643
R25795 DVSS.n21366 DVSS.n21365 0.107643
R25796 DVSS.n21364 DVSS.n21363 0.107643
R25797 DVSS.n21370 DVSS.n21369 0.107643
R25798 DVSS.n21369 DVSS.n21368 0.107643
R25799 DVSS.n21389 DVSS.n21388 0.107643
R25800 DVSS.n21390 DVSS.n21389 0.107643
R25801 DVSS.n514 DVSS.n513 0.107643
R25802 DVSS.n513 DVSS.n512 0.107643
R25803 DVSS.n13914 DVSS.t9 0.1076
R25804 DVSS.n16798 DVSS.t13 0.1076
R25805 DVSS.n15113 DVSS.t16 0.1076
R25806 DVSS.n7636 DVSS.t15 0.1076
R25807 DVSS.n16006 DVSS.t10 0.1076
R25808 DVSS.n15303 DVSS.t34 0.1076
R25809 DVSS.n18296 DVSS.t12 0.1076
R25810 DVSS.n18005 DVSS.t6 0.1076
R25811 DVSS.n17864 DVSS.t14 0.1076
R25812 DVSS.n13829 DVSS.n13828 0.107508
R25813 DVSS.n18603 DVSS.n18602 0.107508
R25814 DVSS.n13706 DVSS.n13705 0.107331
R25815 DVSS.n18689 DVSS.n18688 0.107331
R25816 DVSS.n13810 DVSS.n13809 0.101041
R25817 DVSS.n7408 DVSS.n7407 0.101041
R25818 DVSS.n7387 DVSS.n7384 0.101041
R25819 DVSS.n13770 DVSS.n13767 0.101041
R25820 DVSS.n13730 DVSS.n13723 0.101041
R25821 DVSS.n7360 DVSS.n7352 0.101041
R25822 DVSS.n7360 DVSS.n7359 0.101041
R25823 DVSS.n13730 DVSS.n13729 0.101041
R25824 DVSS DVSS.n18563 0.0977905
R25825 DVSS DVSS.n14927 0.0975391
R25826 DVSS.n8046 DVSS.n8043 0.0945223
R25827 DVSS.n6907 DVSS.n6904 0.0945223
R25828 DVSS.n5387 DVSS.n5386 0.093014
R25829 DVSS.n10266 DVSS.n10264 0.093014
R25830 DVSS.n11527 DVSS.n11526 0.0929803
R25831 DVSS.n6574 DVSS.n6573 0.0929803
R25832 DVSS.n5386 DVSS.n5384 0.0915056
R25833 DVSS.n10267 DVSS.n10266 0.0915056
R25834 DVSS.n1799 DVSS.n1798 0.0913803
R25835 DVSS.n1885 DVSS.n1884 0.0913803
R25836 DVSS.n1538 DVSS.n1537 0.0913803
R25837 DVSS.n13171 DVSS.n13169 0.0889916
R25838 DVSS.n6928 DVSS.n6926 0.0889916
R25839 DVSS.n4470 DVSS.n4469 0.087311
R25840 DVSS.n9489 DVSS.n8953 0.087311
R25841 DVSS.n15708 DVSS.n15707 0.087311
R25842 DVSS.n9705 DVSS.n9704 0.087311
R25843 DVSS.n16220 DVSS.n16219 0.087311
R25844 DVSS.n5364 DVSS.n5363 0.0859749
R25845 DVSS.n10245 DVSS.n10243 0.0859749
R25846 DVSS.n10246 DVSS.n10245 0.0859749
R25847 DVSS.n1769 DVSS.n1768 0.081839
R25848 DVSS.n1776 DVSS.n1775 0.081839
R25849 DVSS.n1783 DVSS.n1782 0.081839
R25850 DVSS.n1791 DVSS.n1790 0.081839
R25851 DVSS.n1806 DVSS.n1805 0.081839
R25852 DVSS.n1812 DVSS.n1811 0.081839
R25853 DVSS.n1819 DVSS.n1818 0.081839
R25854 DVSS.n1826 DVSS.n1825 0.081839
R25855 DVSS.n1862 DVSS.n1861 0.081839
R25856 DVSS.n1868 DVSS.n1867 0.081839
R25857 DVSS.n1875 DVSS.n1874 0.081839
R25858 DVSS.n1881 DVSS.n1880 0.081839
R25859 DVSS.n1889 DVSS.n1888 0.081839
R25860 DVSS.n1893 DVSS.n1892 0.081839
R25861 DVSS.n2468 DVSS.n2466 0.081839
R25862 DVSS.n1508 DVSS.n1507 0.081839
R25863 DVSS.n1514 DVSS.n1513 0.081839
R25864 DVSS.n1522 DVSS.n1521 0.081839
R25865 DVSS.n1529 DVSS.n1528 0.081839
R25866 DVSS.n1534 DVSS.n1533 0.081839
R25867 DVSS.n1542 DVSS.n1541 0.081839
R25868 DVSS.n1546 DVSS.n1545 0.081839
R25869 DVSS.n1551 DVSS.n1549 0.081839
R25870 DVSS.n952 DVSS.n949 0.0797308
R25871 DVSS DVSS.n17449 0.0796667
R25872 DVSS.n17552 DVSS 0.0796667
R25873 DVSS DVSS.n18401 0.0796667
R25874 DVSS.n14962 DVSS 0.0796667
R25875 DVSS.n18369 DVSS 0.0796667
R25876 DVSS.n15591 DVSS 0.0796667
R25877 DVSS.n16240 DVSS 0.0796667
R25878 DVSS DVSS.n15727 0.0796667
R25879 DVSS.n16340 DVSS 0.0796667
R25880 DVSS DVSS.n17659 0.0796667
R25881 DVSS.n16279 DVSS 0.0796667
R25882 DVSS.n15837 DVSS 0.0796667
R25883 DVSS.n7491 DVSS 0.0796667
R25884 DVSS DVSS.n15051 0.0796667
R25885 DVSS.n17248 DVSS 0.0796667
R25886 DVSS DVSS.n17105 0.0796667
R25887 DVSS.n8043 DVSS.n8041 0.075919
R25888 DVSS.n6904 DVSS.n6902 0.075919
R25889 DVSS.n5825 DVSS.n5823 0.0728611
R25890 DVSS.n6554 DVSS.n6553 0.0728611
R25891 DVSS.n6485 DVSS.n6483 0.0728611
R25892 DVSS.n6418 DVSS.n6417 0.0728611
R25893 DVSS.n154 DVSS.n153 0.0693732
R25894 DVSS.n314 DVSS.n313 0.0693732
R25895 DVSS.n1728 DVSS.n1727 0.0687349
R25896 DVSS.n1755 DVSS.n1754 0.0682096
R25897 DVSS.n1846 DVSS.n1845 0.0682096
R25898 DVSS.n7405 DVSS.n7403 0.0673919
R25899 DVSS.n13807 DVSS.n13805 0.0669865
R25900 DVSS.n20503 DVSS.n20500 0.0599231
R25901 DVSS.n20946 DVSS.n20945 0.0599231
R25902 DVSS.n19217 DVSS.n19214 0.0597308
R25903 DVSS.n955 DVSS.n952 0.0597308
R25904 DVSS.n863 DVSS.n862 0.0582559
R25905 DVSS.n20848 DVSS.n20847 0.0582559
R25906 DVSS.n64 DVSS.n63 0.0582559
R25907 DVSS.n21481 DVSS.n21480 0.0582559
R25908 DVSS.n21074 DVSS.n21073 0.0582559
R25909 DVSS.n1150 DVSS.n1149 0.0582559
R25910 DVSS.n18963 DVSS.n18962 0.0582559
R25911 DVSS.n541 DVSS.n540 0.0582559
R25912 DVSS.n19157 DVSS.n19156 0.0576622
R25913 DVSS.n20389 DVSS.n20388 0.0576622
R25914 DVSS.n7020 DVSS.n7018 0.0576622
R25915 DVSS.n13290 DVSS.n13288 0.0576622
R25916 DVSS.n13974 DVSS.n13973 0.056075
R25917 DVSS.n2461 DVSS.n2460 0.0550258
R25918 DVSS.n17451 DVSS 0.0548056
R25919 DVSS.n18403 DVSS 0.0548056
R25920 DVSS DVSS.n18368 0.0548056
R25921 DVSS DVSS.n16239 0.0548056
R25922 DVSS DVSS.n16338 0.0548056
R25923 DVSS DVSS.n16278 0.0548056
R25924 DVSS DVSS.n7490 0.0548056
R25925 DVSS DVSS.n17246 0.0548056
R25926 DVSS.n1832 DVSS.n1831 0.0546818
R25927 DVSS DVSS.n17547 0.0546667
R25928 DVSS DVSS.n14959 0.0546667
R25929 DVSS DVSS.n15588 0.0546667
R25930 DVSS.n15729 DVSS 0.0546667
R25931 DVSS.n17661 DVSS 0.0546667
R25932 DVSS DVSS.n15834 0.0546667
R25933 DVSS.n15053 DVSS 0.0546667
R25934 DVSS.n17107 DVSS 0.0546667
R25935 DVSS.n11034 DVSS.n11032 0.0545278
R25936 DVSS.n9135 DVSS.n9134 0.0545278
R25937 DVSS.n8983 DVSS.n8982 0.0545278
R25938 DVSS.n9747 DVSS.n9746 0.0545278
R25939 DVSS.n11206 DVSS.n11205 0.0545278
R25940 DVSS.n8950 DVSS.n8949 0.0545278
R25941 DVSS.n8056 DVSS.n8055 0.0545278
R25942 DVSS.n5520 DVSS.n5517 0.0545278
R25943 DVSS.n10045 DVSS.n10044 0.0545278
R25944 DVSS.n1762 DVSS.n1761 0.0545
R25945 DVSS.n1490 DVSS.n1489 0.0545
R25946 DVSS.n1854 DVSS.n1853 0.0545
R25947 DVSS.n1502 DVSS.n1501 0.0545
R25948 DVSS.n17946 DVSS.n17945 0.0539507
R25949 DVSS.n18087 DVSS.n18086 0.0539507
R25950 DVSS.n7607 DVSS.n7606 0.0539507
R25951 DVSS.n18418 DVSS.n18417 0.0539507
R25952 DVSS.n18526 DVSS.n18525 0.0539507
R25953 DVSS.n15778 DVSS.n15777 0.0539507
R25954 DVSS.n15371 DVSS.n7673 0.0539507
R25955 DVSS.n15370 DVSS.n15369 0.0539507
R25956 DVSS.n15220 DVSS.n15219 0.0539507
R25957 DVSS.n13855 DVSS.n13854 0.0539507
R25958 DVSS.n17476 DVSS.n17475 0.0537394
R25959 DVSS.n17883 DVSS.n17882 0.0537394
R25960 DVSS.n18024 DVSS.n18023 0.0537394
R25961 DVSS.n7575 DVSS.n7574 0.0537394
R25962 DVSS.n18513 DVSS.n18512 0.0537394
R25963 DVSS.n16817 DVSS.n16816 0.0537394
R25964 DVSS.n15816 DVSS.n15815 0.0537394
R25965 DVSS.n15746 DVSS.n15745 0.0537394
R25966 DVSS.n15234 DVSS.n15233 0.0537394
R25967 DVSS.n7754 DVSS.n7753 0.0537394
R25968 DVSS.n11054 DVSS.n11052 0.0535556
R25969 DVSS.n4113 DVSS.n4112 0.0535556
R25970 DVSS.n9122 DVSS.n9119 0.0535556
R25971 DVSS.n4359 DVSS.n4357 0.0535556
R25972 DVSS.n9597 DVSS.n9595 0.0535556
R25973 DVSS.n9734 DVSS.n9731 0.0535556
R25974 DVSS.n11170 DVSS.n11167 0.0535556
R25975 DVSS.n9789 DVSS.n9787 0.0535556
R25976 DVSS.n4015 DVSS.n4013 0.0535556
R25977 DVSS.n9032 DVSS.n9030 0.0535556
R25978 DVSS.n5536 DVSS.n5534 0.0535556
R25979 DVSS.n10004 DVSS.n10002 0.0535556
R25980 DVSS.n16503 DVSS.n16502 0.0535282
R25981 DVSS.n16849 DVSS.n16848 0.0535282
R25982 DVSS.n18558 DVSS.n18557 0.0526831
R25983 DVSS.n13975 DVSS.n13851 0.0526831
R25984 DVSS.n5832 DVSS.n5830 0.0524444
R25985 DVSS.n6568 DVSS.n6566 0.0524444
R25986 DVSS.n6479 DVSS.n6476 0.0524444
R25987 DVSS.n6432 DVSS.n6430 0.0524444
R25988 DVSS.n1326 DVSS.n1325 0.0510053
R25989 DVSS.n13339 DVSS.n13338 0.0510053
R25990 DVSS.n7024 DVSS.n7023 0.0510053
R25991 DVSS.n13327 DVSS.n13326 0.0510053
R25992 DVSS.n13174 DVSS 0.0487682
R25993 DVSS.n6931 DVSS 0.0487682
R25994 DVSS.n2344 DVSS.n2343 0.04775
R25995 DVSS.n2348 DVSS.n2347 0.04775
R25996 DVSS.n2359 DVSS.n2358 0.04775
R25997 DVSS.n2363 DVSS.n2362 0.04775
R25998 DVSS.n2382 DVSS.n2381 0.04775
R25999 DVSS.n2386 DVSS.n2385 0.04775
R26000 DVSS.n2407 DVSS.n2406 0.04775
R26001 DVSS.n2403 DVSS.n2402 0.04775
R26002 DVSS.n13915 DVSS.n13913 0.0467
R26003 DVSS.n16799 DVSS.n16797 0.0467
R26004 DVSS.n15114 DVSS.n15112 0.0467
R26005 DVSS.n7637 DVSS.n7635 0.0467
R26006 DVSS.n16007 DVSS.n16005 0.0467
R26007 DVSS.n15304 DVSS.n15302 0.0467
R26008 DVSS.n18297 DVSS.n18295 0.0467
R26009 DVSS.n18006 DVSS.n18004 0.0467
R26010 DVSS.n17865 DVSS.n17863 0.0467
R26011 DVSS.n2355 DVSS.n2354 0.0455
R26012 DVSS.n2412 DVSS.n2390 0.0451759
R26013 DVSS.n2353 DVSS.n2352 0.0449197
R26014 DVSS.n6561 DVSS.n6560 0.0449145
R26015 DVSS.n6425 DVSS.n6424 0.0449145
R26016 DVSS.n6565 DVSS.n6564 0.0445103
R26017 DVSS.n6429 DVSS.n6428 0.0445103
R26018 DVSS.n2412 DVSS.n2411 0.0443278
R26019 DVSS.n11032 DVSS.n11030 0.04425
R26020 DVSS.n6767 DVSS.n6766 0.04425
R26021 DVSS.n6712 DVSS.n6711 0.04425
R26022 DVSS.n11205 DVSS.n11203 0.04425
R26023 DVSS.n6894 DVSS.n6893 0.04425
R26024 DVSS.n5517 DVSS.n5515 0.04425
R26025 DVSS.n10044 DVSS.n10042 0.04425
R26026 DVSS.n5833 DVSS.n5832 0.0421667
R26027 DVSS.n6569 DVSS.n6568 0.0421667
R26028 DVSS.n6476 DVSS.n6474 0.0421667
R26029 DVSS.n6433 DVSS.n6432 0.0421667
R26030 DVSS.n5823 DVSS 0.0420278
R26031 DVSS.n6553 DVSS 0.0420278
R26032 DVSS DVSS.n6485 0.0420278
R26033 DVSS.n6417 DVSS 0.0420278
R26034 DVSS DVSS.n13171 0.0407235
R26035 DVSS DVSS.n6928 0.0407235
R26036 DVSS.n1411 DVSS.n1409 0.0403361
R26037 DVSS.n1415 DVSS.n1411 0.0403361
R26038 DVSS.n1418 DVSS.n1415 0.0403361
R26039 DVSS.n1423 DVSS.n1418 0.0403361
R26040 DVSS.n1425 DVSS.n1423 0.0403361
R26041 DVSS.n1429 DVSS.n1425 0.0403361
R26042 DVSS.n1432 DVSS.n1429 0.0403361
R26043 DVSS.n1436 DVSS.n1432 0.0403361
R26044 DVSS.n1439 DVSS.n1436 0.0403361
R26045 DVSS.n1443 DVSS.n1439 0.0403361
R26046 DVSS.n1445 DVSS.n1443 0.0403361
R26047 DVSS.n1449 DVSS.n1445 0.0403361
R26048 DVSS.n1451 DVSS.n1449 0.0403361
R26049 DVSS.n1456 DVSS.n1451 0.0403361
R26050 DVSS.n1458 DVSS.n1456 0.0403361
R26051 DVSS.n1463 DVSS.n1458 0.0403361
R26052 DVSS.n1466 DVSS.n1463 0.0403361
R26053 DVSS.n1470 DVSS.n1466 0.0403361
R26054 DVSS.n1473 DVSS.n1470 0.0403361
R26055 DVSS.n1478 DVSS.n1473 0.0403361
R26056 DVSS.n1480 DVSS.n1478 0.0403361
R26057 DVSS.n1485 DVSS.n1480 0.0403361
R26058 DVSS.n1488 DVSS.n1485 0.0403361
R26059 DVSS.n1492 DVSS.n1488 0.0403361
R26060 DVSS.n1500 DVSS.n1498 0.0403361
R26061 DVSS.n1504 DVSS.n1500 0.0403361
R26062 DVSS.n1506 DVSS.n1504 0.0403361
R26063 DVSS.n1510 DVSS.n1506 0.0403361
R26064 DVSS.n1512 DVSS.n1510 0.0403361
R26065 DVSS.n1517 DVSS.n1512 0.0403361
R26066 DVSS.n1520 DVSS.n1517 0.0403361
R26067 DVSS.n1525 DVSS.n1520 0.0403361
R26068 DVSS.n1527 DVSS.n1525 0.0403361
R26069 DVSS.n1531 DVSS.n1527 0.0403361
R26070 DVSS.n1532 DVSS.n1531 0.0403361
R26071 DVSS.n1535 DVSS.n1532 0.0403361
R26072 DVSS.n1536 DVSS.n1535 0.0403361
R26073 DVSS.n1539 DVSS.n1536 0.0403361
R26074 DVSS.n1540 DVSS.n1539 0.0403361
R26075 DVSS.n1543 DVSS.n1540 0.0403361
R26076 DVSS.n1544 DVSS.n1543 0.0403361
R26077 DVSS.n1547 DVSS.n1544 0.0403361
R26078 DVSS.n1548 DVSS.n1547 0.0403361
R26079 DVSS.n1740 DVSS.n1548 0.0403361
R26080 DVSS.n1740 DVSS.n1739 0.0403361
R26081 DVSS.n1739 DVSS.n1738 0.0403361
R26082 DVSS.n1738 DVSS.n1736 0.0403361
R26083 DVSS.n1736 DVSS.n1733 0.0403361
R26084 DVSS.n1753 DVSS.n1750 0.0403361
R26085 DVSS.n1758 DVSS.n1753 0.0403361
R26086 DVSS.n1760 DVSS.n1758 0.0403361
R26087 DVSS.n1764 DVSS.n1760 0.0403361
R26088 DVSS.n1767 DVSS.n1764 0.0403361
R26089 DVSS.n1772 DVSS.n1767 0.0403361
R26090 DVSS.n1774 DVSS.n1772 0.0403361
R26091 DVSS.n1779 DVSS.n1774 0.0403361
R26092 DVSS.n1781 DVSS.n1779 0.0403361
R26093 DVSS.n1786 DVSS.n1781 0.0403361
R26094 DVSS.n1789 DVSS.n1786 0.0403361
R26095 DVSS.n1794 DVSS.n1789 0.0403361
R26096 DVSS.n1797 DVSS.n1794 0.0403361
R26097 DVSS.n1801 DVSS.n1797 0.0403361
R26098 DVSS.n1804 DVSS.n1801 0.0403361
R26099 DVSS.n1808 DVSS.n1804 0.0403361
R26100 DVSS.n1810 DVSS.n1808 0.0403361
R26101 DVSS.n1815 DVSS.n1810 0.0403361
R26102 DVSS.n1817 DVSS.n1815 0.0403361
R26103 DVSS.n1821 DVSS.n1817 0.0403361
R26104 DVSS.n1824 DVSS.n1821 0.0403361
R26105 DVSS.n1828 DVSS.n1824 0.0403361
R26106 DVSS.n1830 DVSS.n1828 0.0403361
R26107 DVSS.n1835 DVSS.n1830 0.0403361
R26108 DVSS.n1844 DVSS.n1841 0.0403361
R26109 DVSS.n1849 DVSS.n1844 0.0403361
R26110 DVSS.n1852 DVSS.n1849 0.0403361
R26111 DVSS.n1857 DVSS.n1852 0.0403361
R26112 DVSS.n1860 DVSS.n1857 0.0403361
R26113 DVSS.n1864 DVSS.n1860 0.0403361
R26114 DVSS.n1866 DVSS.n1864 0.0403361
R26115 DVSS.n1870 DVSS.n1866 0.0403361
R26116 DVSS.n1873 DVSS.n1870 0.0403361
R26117 DVSS.n1878 DVSS.n1873 0.0403361
R26118 DVSS.n1879 DVSS.n1878 0.0403361
R26119 DVSS.n1882 DVSS.n1879 0.0403361
R26120 DVSS.n1883 DVSS.n1882 0.0403361
R26121 DVSS.n1886 DVSS.n1883 0.0403361
R26122 DVSS.n1887 DVSS.n1886 0.0403361
R26123 DVSS.n1890 DVSS.n1887 0.0403361
R26124 DVSS.n1891 DVSS.n1890 0.0403361
R26125 DVSS.n1894 DVSS.n1891 0.0403361
R26126 DVSS.n1895 DVSS.n1894 0.0403361
R26127 DVSS.n2469 DVSS.n1895 0.0403361
R26128 DVSS.n2469 DVSS.n2465 0.0403361
R26129 DVSS.n2465 DVSS.n2464 0.0403361
R26130 DVSS.n2464 DVSS.n1901 0.0403361
R26131 DVSS.n1901 DVSS.n1899 0.0403361
R26132 DVSS.n17805 DVSS.n17804 0.0402183
R26133 DVSS.n15784 DVSS.n15783 0.0402183
R26134 DVSS.n17235 DVSS.n17231 0.0401
R26135 DVSS.n15065 DVSS.n15064 0.0401
R26136 DVSS.n17679 DVSS.n17678 0.0401
R26137 DVSS.n17532 DVSS.n17529 0.0401
R26138 DVSS.n15262 DVSS.n15261 0.0401
R26139 DVSS.n18359 DVSS.n18356 0.0401
R26140 DVSS.n18080 DVSS.n18077 0.0401
R26141 DVSS.n17939 DVSS.n17936 0.0401
R26142 DVSS DVSS.n17432 0.039875
R26143 DVSS DVSS.n16889 0.039875
R26144 DVSS DVSS.n7460 0.039875
R26145 DVSS DVSS.n14973 0.039875
R26146 DVSS DVSS.n7549 0.039875
R26147 DVSS DVSS.n15602 0.039875
R26148 DVSS DVSS.n16221 0.039875
R26149 DVSS DVSS.n7689 0.039875
R26150 DVSS DVSS.n16305 0.039875
R26151 DVSS DVSS.n17642 0.039875
R26152 DVSS DVSS.n16260 0.039875
R26153 DVSS DVSS.n15848 0.039875
R26154 DVSS DVSS.n14942 0.039875
R26155 DVSS DVSS.n7470 0.039875
R26156 DVSS DVSS.n7777 0.039875
R26157 DVSS DVSS.n16425 0.039875
R26158 DVSS DVSS.n16879 0.039875
R26159 DVSS DVSS.n7432 0.039875
R26160 DVSS.n6424 DVSS.n6423 0.037361
R26161 DVSS.n6560 DVSS.n6559 0.037361
R26162 DVSS.n6428 DVSS.n6427 0.0372894
R26163 DVSS.n6564 DVSS.n6563 0.0372894
R26164 DVSS.n2378 DVSS.n2377 0.03515
R26165 DVSS.n2399 DVSS.n2398 0.03515
R26166 DVSS.n13288 DVSS.n13287 0.0337432
R26167 DVSS.n13980 DVSS.n13978 0.0333378
R26168 DVSS.n14049 DVSS.n14047 0.0333378
R26169 DVSS.n7018 DVSS.n7017 0.0333378
R26170 DVSS.n14790 DVSS.n14786 0.0333378
R26171 DVSS.n6141 DVSS.n6140 0.03245
R26172 DVSS.n6135 DVSS.n6134 0.032
R26173 DVSS.n6121 DVSS.n6120 0.032
R26174 DVSS.n6115 DVSS.n6114 0.032
R26175 DVSS.n2352 DVSS.n2351 0.0319852
R26176 DVSS.n2390 DVSS.n2389 0.0319852
R26177 DVSS DVSS.n5821 0.0313333
R26178 DVSS.n11056 DVSS 0.0313333
R26179 DVSS DVSS.n4110 0.0313333
R26180 DVSS DVSS.n9117 0.0313333
R26181 DVSS.n4362 DVSS 0.0313333
R26182 DVSS.n9598 DVSS 0.0313333
R26183 DVSS DVSS.n6551 0.0313333
R26184 DVSS DVSS.n9729 0.0313333
R26185 DVSS.n6502 DVSS 0.0313333
R26186 DVSS DVSS.n11165 0.0313333
R26187 DVSS DVSS.n6415 0.0313333
R26188 DVSS.n9790 DVSS 0.0313333
R26189 DVSS.n4018 DVSS 0.0313333
R26190 DVSS.n9033 DVSS 0.0313333
R26191 DVSS.n5553 DVSS 0.0313333
R26192 DVSS DVSS.n10000 0.0313333
R26193 DVSS.n2411 DVSS.n2410 0.0308013
R26194 DVSS.n6010 DVSS.n6009 0.03065
R26195 DVSS.n6017 DVSS.n6016 0.03065
R26196 DVSS.n6019 DVSS.n6018 0.03065
R26197 DVSS.n19893 DVSS.n19892 0.0300946
R26198 DVSS.n2354 DVSS.n2353 0.0291833
R26199 DVSS.n6429 DVSS.n6426 0.0291833
R26200 DVSS.n6565 DVSS.n6562 0.0291833
R26201 DVSS.n6021 DVSS.n6020 0.0291833
R26202 DVSS.n16803 DVSS.n16802 0.0290496
R26203 DVSS.n15071 DVSS.n15070 0.0290496
R26204 DVSS.n7641 DVSS.n7640 0.0290496
R26205 DVSS.n16010 DVSS.n16009 0.0290496
R26206 DVSS.n15307 DVSS.n15306 0.0290496
R26207 DVSS.n18352 DVSS.n18351 0.0290496
R26208 DVSS.n18009 DVSS.n18008 0.0290496
R26209 DVSS.n17868 DVSS.n17867 0.0290496
R26210 DVSS.n13968 DVSS.n13967 0.0290496
R26211 DVSS.n6425 DVSS.n6421 0.0289271
R26212 DVSS.n6561 DVSS.n6557 0.0289271
R26213 DVSS.n6142 DVSS.n6141 0.0289271
R26214 DVSS.n5912 DVSS.n5911 0.0289271
R26215 DVSS.n6144 DVSS.n6143 0.0289271
R26216 DVSS.n20390 DVSS.n20389 0.0288784
R26217 DVSS.n2371 DVSS.n2370 0.0285987
R26218 DVSS.n2394 DVSS.n2393 0.0285987
R26219 DVSS.n19158 DVSS.n19157 0.028473
R26220 DVSS.n1413 DVSS.n1412 0.027839
R26221 DVSS.n1420 DVSS.n1419 0.027839
R26222 DVSS.n1427 DVSS.n1426 0.027839
R26223 DVSS.n1434 DVSS.n1433 0.027839
R26224 DVSS.n1441 DVSS.n1440 0.027839
R26225 DVSS.n1453 DVSS.n1452 0.027839
R26226 DVSS.n1460 DVSS.n1459 0.027839
R26227 DVSS.n1468 DVSS.n1467 0.027839
R26228 DVSS.n1475 DVSS.n1474 0.027839
R26229 DVSS.n1482 DVSS.n1481 0.027839
R26230 DVSS.n2468 DVSS.n2467 0.027839
R26231 DVSS.n1551 DVSS.n1550 0.027839
R26232 DVSS.n6009 DVSS.n6008 0.02615
R26233 DVSS.n6011 DVSS.n6010 0.02615
R26234 DVSS.n6018 DVSS.n6017 0.02615
R26235 DVSS.n6020 DVSS.n6019 0.02615
R26236 DVSS.n8034 DVSS.n8033 0.0248803
R26237 DVSS.n17435 DVSS.n17434 0.0246667
R26238 DVSS.n7463 DVSS.n7462 0.0246667
R26239 DVSS.n7552 DVSS.n7551 0.0246667
R26240 DVSS.n16224 DVSS.n16223 0.0246667
R26241 DVSS.n16308 DVSS.n16307 0.0246667
R26242 DVSS.n16263 DVSS.n16262 0.0246667
R26243 DVSS.n7473 DVSS.n7472 0.0246667
R26244 DVSS.n7780 DVSS.n7779 0.0246667
R26245 DVSS.n16428 DVSS.n16427 0.0246667
R26246 DVSS.n2341 DVSS.n2340 0.024601
R26247 DVSS.n2370 DVSS.n2369 0.0245016
R26248 DVSS.n2395 DVSS.n2394 0.0245016
R26249 DVSS.n2367 DVSS.n2366 0.0243765
R26250 DVSS.n2366 DVSS.n2365 0.0237031
R26251 DVSS.n2340 DVSS.n2339 0.0234786
R26252 DVSS.n14915 DVSS.n14912 0.02345
R26253 DVSS.n19951 DVSS.n19948 0.0233846
R26254 DVSS.n19966 DVSS.n19951 0.0233846
R26255 DVSS.n359 DVSS.n341 0.0233846
R26256 DVSS.n362 DVSS.n359 0.0233846
R26257 DVSS.n16616 DVSS.n16612 0.0233169
R26258 DVSS.n16620 DVSS.n16616 0.0233169
R26259 DVSS.n16624 DVSS.n16620 0.0233169
R26260 DVSS.n16625 DVSS.n16624 0.0233169
R26261 DVSS.n16626 DVSS.n16625 0.0233169
R26262 DVSS.n16630 DVSS.n16626 0.0233169
R26263 DVSS.n16631 DVSS.n16630 0.0233169
R26264 DVSS.n16632 DVSS.n16631 0.0233169
R26265 DVSS.n16633 DVSS.n16632 0.0233169
R26266 DVSS.n16634 DVSS.n16633 0.0233169
R26267 DVSS.n16635 DVSS.n16634 0.0233169
R26268 DVSS.n16636 DVSS.n16635 0.0233169
R26269 DVSS.n16637 DVSS.n16636 0.0233169
R26270 DVSS.n16638 DVSS.n16637 0.0233169
R26271 DVSS.n16639 DVSS.n16638 0.0233169
R26272 DVSS.n16640 DVSS.n16639 0.0233169
R26273 DVSS.n16499 DVSS.n16492 0.0233169
R26274 DVSS.n16492 DVSS.n16488 0.0233169
R26275 DVSS.n16488 DVSS.n16484 0.0233169
R26276 DVSS.n16484 DVSS.n16480 0.0233169
R26277 DVSS.n16480 DVSS.n16476 0.0233169
R26278 DVSS.n16476 DVSS.n16472 0.0233169
R26279 DVSS.n16472 DVSS.n16468 0.0233169
R26280 DVSS.n16468 DVSS.n16464 0.0233169
R26281 DVSS.n16464 DVSS.n16460 0.0233169
R26282 DVSS.n16460 DVSS.n16456 0.0233169
R26283 DVSS.n16456 DVSS.n16452 0.0233169
R26284 DVSS.n16452 DVSS.n16448 0.0233169
R26285 DVSS.n16448 DVSS.n16014 0.0233169
R26286 DVSS.n17490 DVSS.n16014 0.0233169
R26287 DVSS.n17490 DVSS.n17489 0.0233169
R26288 DVSS.n17489 DVSS.n17488 0.0233169
R26289 DVSS.n17488 DVSS.n17487 0.0233169
R26290 DVSS.n17487 DVSS.n17486 0.0233169
R26291 DVSS.n17486 DVSS.n17485 0.0233169
R26292 DVSS.n17485 DVSS.n17484 0.0233169
R26293 DVSS.n17484 DVSS.n17483 0.0233169
R26294 DVSS.n17483 DVSS.n17482 0.0233169
R26295 DVSS.n17482 DVSS.n17481 0.0233169
R26296 DVSS.n17481 DVSS.n17480 0.0233169
R26297 DVSS.n17480 DVSS.n17479 0.0233169
R26298 DVSS.n16058 DVSS.n16042 0.0233169
R26299 DVSS.n16042 DVSS.n16038 0.0233169
R26300 DVSS.n16038 DVSS.n16034 0.0233169
R26301 DVSS.n16034 DVSS.n16030 0.0233169
R26302 DVSS.n16030 DVSS.n16026 0.0233169
R26303 DVSS.n16026 DVSS.n16022 0.0233169
R26304 DVSS.n16022 DVSS.n16018 0.0233169
R26305 DVSS.n16018 DVSS.n7644 0.0233169
R26306 DVSS.n17721 DVSS.n7644 0.0233169
R26307 DVSS.n17722 DVSS.n17721 0.0233169
R26308 DVSS.n17723 DVSS.n17722 0.0233169
R26309 DVSS.n17724 DVSS.n17723 0.0233169
R26310 DVSS.n17725 DVSS.n17724 0.0233169
R26311 DVSS.n17726 DVSS.n17725 0.0233169
R26312 DVSS.n17727 DVSS.n17726 0.0233169
R26313 DVSS.n17728 DVSS.n17727 0.0233169
R26314 DVSS.n17818 DVSS.n17814 0.0233169
R26315 DVSS.n17822 DVSS.n17818 0.0233169
R26316 DVSS.n17826 DVSS.n17822 0.0233169
R26317 DVSS.n17830 DVSS.n17826 0.0233169
R26318 DVSS.n17834 DVSS.n17830 0.0233169
R26319 DVSS.n17838 DVSS.n17834 0.0233169
R26320 DVSS.n17842 DVSS.n17838 0.0233169
R26321 DVSS.n17846 DVSS.n17842 0.0233169
R26322 DVSS.n17850 DVSS.n17846 0.0233169
R26323 DVSS.n17854 DVSS.n17850 0.0233169
R26324 DVSS.n17858 DVSS.n17854 0.0233169
R26325 DVSS.n17862 DVSS.n17858 0.0233169
R26326 DVSS.n17872 DVSS.n17862 0.0233169
R26327 DVSS.n17897 DVSS.n17872 0.0233169
R26328 DVSS.n17897 DVSS.n17896 0.0233169
R26329 DVSS.n17896 DVSS.n17895 0.0233169
R26330 DVSS.n17895 DVSS.n17894 0.0233169
R26331 DVSS.n17894 DVSS.n17893 0.0233169
R26332 DVSS.n17893 DVSS.n17892 0.0233169
R26333 DVSS.n17892 DVSS.n17891 0.0233169
R26334 DVSS.n17891 DVSS.n17890 0.0233169
R26335 DVSS.n17890 DVSS.n17889 0.0233169
R26336 DVSS.n17889 DVSS.n17888 0.0233169
R26337 DVSS.n17888 DVSS.n17887 0.0233169
R26338 DVSS.n17887 DVSS.n17886 0.0233169
R26339 DVSS.n17959 DVSS.n17955 0.0233169
R26340 DVSS.n17963 DVSS.n17959 0.0233169
R26341 DVSS.n17967 DVSS.n17963 0.0233169
R26342 DVSS.n17971 DVSS.n17967 0.0233169
R26343 DVSS.n17975 DVSS.n17971 0.0233169
R26344 DVSS.n17979 DVSS.n17975 0.0233169
R26345 DVSS.n17983 DVSS.n17979 0.0233169
R26346 DVSS.n17987 DVSS.n17983 0.0233169
R26347 DVSS.n17991 DVSS.n17987 0.0233169
R26348 DVSS.n17995 DVSS.n17991 0.0233169
R26349 DVSS.n17999 DVSS.n17995 0.0233169
R26350 DVSS.n18003 DVSS.n17999 0.0233169
R26351 DVSS.n18013 DVSS.n18003 0.0233169
R26352 DVSS.n18038 DVSS.n18013 0.0233169
R26353 DVSS.n18038 DVSS.n18037 0.0233169
R26354 DVSS.n18037 DVSS.n18036 0.0233169
R26355 DVSS.n18036 DVSS.n18035 0.0233169
R26356 DVSS.n18035 DVSS.n18034 0.0233169
R26357 DVSS.n18034 DVSS.n18033 0.0233169
R26358 DVSS.n18033 DVSS.n18032 0.0233169
R26359 DVSS.n18032 DVSS.n18031 0.0233169
R26360 DVSS.n18031 DVSS.n18030 0.0233169
R26361 DVSS.n18030 DVSS.n18029 0.0233169
R26362 DVSS.n18029 DVSS.n18028 0.0233169
R26363 DVSS.n18028 DVSS.n18027 0.0233169
R26364 DVSS.n7603 DVSS.n7602 0.0233169
R26365 DVSS.n7602 DVSS.n7601 0.0233169
R26366 DVSS.n7601 DVSS.n7600 0.0233169
R26367 DVSS.n7600 DVSS.n7599 0.0233169
R26368 DVSS.n7599 DVSS.n7598 0.0233169
R26369 DVSS.n7598 DVSS.n7597 0.0233169
R26370 DVSS.n7597 DVSS.n7596 0.0233169
R26371 DVSS.n7596 DVSS.n7595 0.0233169
R26372 DVSS.n7595 DVSS.n7594 0.0233169
R26373 DVSS.n7594 DVSS.n7593 0.0233169
R26374 DVSS.n7593 DVSS.n7592 0.0233169
R26375 DVSS.n7592 DVSS.n7591 0.0233169
R26376 DVSS.n7591 DVSS.n7590 0.0233169
R26377 DVSS.n7590 DVSS.n7589 0.0233169
R26378 DVSS.n7589 DVSS.n7588 0.0233169
R26379 DVSS.n7588 DVSS.n7587 0.0233169
R26380 DVSS.n7587 DVSS.n7586 0.0233169
R26381 DVSS.n7586 DVSS.n7585 0.0233169
R26382 DVSS.n7585 DVSS.n7584 0.0233169
R26383 DVSS.n7584 DVSS.n7583 0.0233169
R26384 DVSS.n7583 DVSS.n7582 0.0233169
R26385 DVSS.n7582 DVSS.n7581 0.0233169
R26386 DVSS.n7581 DVSS.n7580 0.0233169
R26387 DVSS.n7580 DVSS.n7579 0.0233169
R26388 DVSS.n7579 DVSS.n7578 0.0233169
R26389 DVSS.n18422 DVSS.n18421 0.0233169
R26390 DVSS.n18500 DVSS.n18499 0.0233169
R26391 DVSS.n18501 DVSS.n18500 0.0233169
R26392 DVSS.n18502 DVSS.n18501 0.0233169
R26393 DVSS.n18503 DVSS.n18502 0.0233169
R26394 DVSS.n18504 DVSS.n18503 0.0233169
R26395 DVSS.n18505 DVSS.n18504 0.0233169
R26396 DVSS.n18506 DVSS.n18505 0.0233169
R26397 DVSS.n18507 DVSS.n18506 0.0233169
R26398 DVSS.n18508 DVSS.n18507 0.0233169
R26399 DVSS.n18509 DVSS.n18508 0.0233169
R26400 DVSS.n18530 DVSS.n18529 0.0233169
R26401 DVSS.n18531 DVSS.n18530 0.0233169
R26402 DVSS.n18532 DVSS.n18531 0.0233169
R26403 DVSS.n18533 DVSS.n18532 0.0233169
R26404 DVSS.n18534 DVSS.n18533 0.0233169
R26405 DVSS.n18535 DVSS.n18534 0.0233169
R26406 DVSS.n18536 DVSS.n18535 0.0233169
R26407 DVSS.n18537 DVSS.n18536 0.0233169
R26408 DVSS.n18538 DVSS.n18537 0.0233169
R26409 DVSS.n18539 DVSS.n18538 0.0233169
R26410 DVSS.n18540 DVSS.n18539 0.0233169
R26411 DVSS.n18541 DVSS.n18540 0.0233169
R26412 DVSS.n18542 DVSS.n18541 0.0233169
R26413 DVSS.n18543 DVSS.n18542 0.0233169
R26414 DVSS.n18544 DVSS.n18543 0.0233169
R26415 DVSS.n18545 DVSS.n18544 0.0233169
R26416 DVSS.n18546 DVSS.n18545 0.0233169
R26417 DVSS.n18547 DVSS.n18546 0.0233169
R26418 DVSS.n18548 DVSS.n18547 0.0233169
R26419 DVSS.n18549 DVSS.n18548 0.0233169
R26420 DVSS.n18550 DVSS.n18549 0.0233169
R26421 DVSS.n18551 DVSS.n18550 0.0233169
R26422 DVSS.n18552 DVSS.n18551 0.0233169
R26423 DVSS.n18553 DVSS.n18552 0.0233169
R26424 DVSS.n18554 DVSS.n18553 0.0233169
R26425 DVSS.n16777 DVSS.n16776 0.0233169
R26426 DVSS.n16778 DVSS.n16777 0.0233169
R26427 DVSS.n16779 DVSS.n16778 0.0233169
R26428 DVSS.n16783 DVSS.n16779 0.0233169
R26429 DVSS.n16787 DVSS.n16783 0.0233169
R26430 DVSS.n16788 DVSS.n16787 0.0233169
R26431 DVSS.n16792 DVSS.n16788 0.0233169
R26432 DVSS.n16796 DVSS.n16792 0.0233169
R26433 DVSS.n16806 DVSS.n16796 0.0233169
R26434 DVSS.n17188 DVSS.n16806 0.0233169
R26435 DVSS.n17188 DVSS.n17187 0.0233169
R26436 DVSS.n17187 DVSS.n17186 0.0233169
R26437 DVSS.n17186 DVSS.n17185 0.0233169
R26438 DVSS.n17185 DVSS.n17184 0.0233169
R26439 DVSS.n17184 DVSS.n17183 0.0233169
R26440 DVSS.n17183 DVSS.n17182 0.0233169
R26441 DVSS.n16845 DVSS.n16844 0.0233169
R26442 DVSS.n16844 DVSS.n16843 0.0233169
R26443 DVSS.n16843 DVSS.n16842 0.0233169
R26444 DVSS.n16842 DVSS.n16841 0.0233169
R26445 DVSS.n16841 DVSS.n16840 0.0233169
R26446 DVSS.n16840 DVSS.n16839 0.0233169
R26447 DVSS.n16839 DVSS.n16838 0.0233169
R26448 DVSS.n16838 DVSS.n16837 0.0233169
R26449 DVSS.n16837 DVSS.n16836 0.0233169
R26450 DVSS.n16836 DVSS.n16835 0.0233169
R26451 DVSS.n16835 DVSS.n16834 0.0233169
R26452 DVSS.n16834 DVSS.n16833 0.0233169
R26453 DVSS.n16833 DVSS.n16832 0.0233169
R26454 DVSS.n16832 DVSS.n16831 0.0233169
R26455 DVSS.n16831 DVSS.n16830 0.0233169
R26456 DVSS.n16830 DVSS.n16829 0.0233169
R26457 DVSS.n16829 DVSS.n16828 0.0233169
R26458 DVSS.n16828 DVSS.n16827 0.0233169
R26459 DVSS.n16827 DVSS.n16826 0.0233169
R26460 DVSS.n16826 DVSS.n16825 0.0233169
R26461 DVSS.n16825 DVSS.n16824 0.0233169
R26462 DVSS.n16824 DVSS.n16823 0.0233169
R26463 DVSS.n16823 DVSS.n16822 0.0233169
R26464 DVSS.n16822 DVSS.n16821 0.0233169
R26465 DVSS.n16821 DVSS.n16820 0.0233169
R26466 DVSS.n15950 DVSS.n15949 0.0233169
R26467 DVSS.n15949 DVSS.n15948 0.0233169
R26468 DVSS.n15948 DVSS.n15947 0.0233169
R26469 DVSS.n15947 DVSS.n15946 0.0233169
R26470 DVSS.n15946 DVSS.n15945 0.0233169
R26471 DVSS.n15945 DVSS.n15944 0.0233169
R26472 DVSS.n15944 DVSS.n15943 0.0233169
R26473 DVSS.n15943 DVSS.n15942 0.0233169
R26474 DVSS.n15942 DVSS.n15941 0.0233169
R26475 DVSS.n15941 DVSS.n15940 0.0233169
R26476 DVSS.n15940 DVSS.n15939 0.0233169
R26477 DVSS.n15939 DVSS.n15938 0.0233169
R26478 DVSS.n15938 DVSS.n15937 0.0233169
R26479 DVSS.n15937 DVSS.n15936 0.0233169
R26480 DVSS.n15936 DVSS.n15935 0.0233169
R26481 DVSS.n15935 DVSS.n15934 0.0233169
R26482 DVSS.n15788 DVSS.n15787 0.0233169
R26483 DVSS.n15789 DVSS.n15788 0.0233169
R26484 DVSS.n15790 DVSS.n15789 0.0233169
R26485 DVSS.n15791 DVSS.n15790 0.0233169
R26486 DVSS.n15792 DVSS.n15791 0.0233169
R26487 DVSS.n15793 DVSS.n15792 0.0233169
R26488 DVSS.n15794 DVSS.n15793 0.0233169
R26489 DVSS.n15795 DVSS.n15794 0.0233169
R26490 DVSS.n15796 DVSS.n15795 0.0233169
R26491 DVSS.n15797 DVSS.n15796 0.0233169
R26492 DVSS.n15798 DVSS.n15797 0.0233169
R26493 DVSS.n15799 DVSS.n15798 0.0233169
R26494 DVSS.n15800 DVSS.n15799 0.0233169
R26495 DVSS.n15801 DVSS.n15800 0.0233169
R26496 DVSS.n15802 DVSS.n15801 0.0233169
R26497 DVSS.n15803 DVSS.n15802 0.0233169
R26498 DVSS.n15804 DVSS.n15803 0.0233169
R26499 DVSS.n15805 DVSS.n15804 0.0233169
R26500 DVSS.n15806 DVSS.n15805 0.0233169
R26501 DVSS.n15807 DVSS.n15806 0.0233169
R26502 DVSS.n15808 DVSS.n15807 0.0233169
R26503 DVSS.n15809 DVSS.n15808 0.0233169
R26504 DVSS.n15810 DVSS.n15809 0.0233169
R26505 DVSS.n15811 DVSS.n15810 0.0233169
R26506 DVSS.n15812 DVSS.n15811 0.0233169
R26507 DVSS.n15774 DVSS.n15773 0.0233169
R26508 DVSS.n15773 DVSS.n15772 0.0233169
R26509 DVSS.n15772 DVSS.n15771 0.0233169
R26510 DVSS.n15771 DVSS.n15770 0.0233169
R26511 DVSS.n15770 DVSS.n15769 0.0233169
R26512 DVSS.n15769 DVSS.n15768 0.0233169
R26513 DVSS.n15768 DVSS.n15767 0.0233169
R26514 DVSS.n15767 DVSS.n15766 0.0233169
R26515 DVSS.n15766 DVSS.n15765 0.0233169
R26516 DVSS.n15765 DVSS.n15764 0.0233169
R26517 DVSS.n15764 DVSS.n15763 0.0233169
R26518 DVSS.n15763 DVSS.n15762 0.0233169
R26519 DVSS.n15762 DVSS.n15761 0.0233169
R26520 DVSS.n15761 DVSS.n15760 0.0233169
R26521 DVSS.n15760 DVSS.n15759 0.0233169
R26522 DVSS.n15759 DVSS.n15758 0.0233169
R26523 DVSS.n15758 DVSS.n15757 0.0233169
R26524 DVSS.n15757 DVSS.n15756 0.0233169
R26525 DVSS.n15756 DVSS.n15755 0.0233169
R26526 DVSS.n15755 DVSS.n15754 0.0233169
R26527 DVSS.n15754 DVSS.n15753 0.0233169
R26528 DVSS.n15753 DVSS.n15752 0.0233169
R26529 DVSS.n15752 DVSS.n15751 0.0233169
R26530 DVSS.n15751 DVSS.n15750 0.0233169
R26531 DVSS.n15750 DVSS.n15749 0.0233169
R26532 DVSS.n15366 DVSS.n15359 0.0233169
R26533 DVSS.n15359 DVSS.n15355 0.0233169
R26534 DVSS.n15355 DVSS.n15351 0.0233169
R26535 DVSS.n15351 DVSS.n15347 0.0233169
R26536 DVSS.n15347 DVSS.n15343 0.0233169
R26537 DVSS.n15343 DVSS.n15339 0.0233169
R26538 DVSS.n15339 DVSS.n15335 0.0233169
R26539 DVSS.n15335 DVSS.n15331 0.0233169
R26540 DVSS.n15331 DVSS.n15327 0.0233169
R26541 DVSS.n15327 DVSS.n15323 0.0233169
R26542 DVSS.n15323 DVSS.n15319 0.0233169
R26543 DVSS.n15319 DVSS.n15315 0.0233169
R26544 DVSS.n15315 DVSS.n15311 0.0233169
R26545 DVSS.n15311 DVSS.n15301 0.0233169
R26546 DVSS.n15301 DVSS.n7702 0.0233169
R26547 DVSS.n15221 DVSS.n7702 0.0233169
R26548 DVSS.n15222 DVSS.n15221 0.0233169
R26549 DVSS.n15223 DVSS.n15222 0.0233169
R26550 DVSS.n15224 DVSS.n15223 0.0233169
R26551 DVSS.n15225 DVSS.n15224 0.0233169
R26552 DVSS.n15226 DVSS.n15225 0.0233169
R26553 DVSS.n15227 DVSS.n15226 0.0233169
R26554 DVSS.n15228 DVSS.n15227 0.0233169
R26555 DVSS.n15229 DVSS.n15228 0.0233169
R26556 DVSS.n15230 DVSS.n15229 0.0233169
R26557 DVSS.n15216 DVSS.n15209 0.0233169
R26558 DVSS.n7741 DVSS.n7740 0.0233169
R26559 DVSS.n7742 DVSS.n7741 0.0233169
R26560 DVSS.n7743 DVSS.n7742 0.0233169
R26561 DVSS.n7744 DVSS.n7743 0.0233169
R26562 DVSS.n7745 DVSS.n7744 0.0233169
R26563 DVSS.n7746 DVSS.n7745 0.0233169
R26564 DVSS.n7747 DVSS.n7746 0.0233169
R26565 DVSS.n7748 DVSS.n7747 0.0233169
R26566 DVSS.n7749 DVSS.n7748 0.0233169
R26567 DVSS.n7750 DVSS.n7749 0.0233169
R26568 DVSS.n13868 DVSS.n13864 0.0233169
R26569 DVSS.n13872 DVSS.n13868 0.0233169
R26570 DVSS.n13876 DVSS.n13872 0.0233169
R26571 DVSS.n13880 DVSS.n13876 0.0233169
R26572 DVSS.n13884 DVSS.n13880 0.0233169
R26573 DVSS.n13888 DVSS.n13884 0.0233169
R26574 DVSS.n13892 DVSS.n13888 0.0233169
R26575 DVSS.n13896 DVSS.n13892 0.0233169
R26576 DVSS.n13900 DVSS.n13896 0.0233169
R26577 DVSS.n13904 DVSS.n13900 0.0233169
R26578 DVSS.n13908 DVSS.n13904 0.0233169
R26579 DVSS.n13912 DVSS.n13908 0.0233169
R26580 DVSS.n13918 DVSS.n13912 0.0233169
R26581 DVSS.n13932 DVSS.n13918 0.0233169
R26582 DVSS.n13932 DVSS.n13931 0.0233169
R26583 DVSS.n13931 DVSS.n13930 0.0233169
R26584 DVSS.n13930 DVSS.n13929 0.0233169
R26585 DVSS.n13929 DVSS.n13928 0.0233169
R26586 DVSS.n13928 DVSS.n13927 0.0233169
R26587 DVSS.n13927 DVSS.n13926 0.0233169
R26588 DVSS.n13926 DVSS.n13925 0.0233169
R26589 DVSS.n13925 DVSS.n13924 0.0233169
R26590 DVSS.n13924 DVSS.n13923 0.0233169
R26591 DVSS.n13923 DVSS.n13922 0.0233169
R26592 DVSS.n13922 DVSS.n13921 0.0233169
R26593 DVSS DVSS.n11054 0.0227222
R26594 DVSS.n4112 DVSS 0.0227222
R26595 DVSS.n9119 DVSS 0.0227222
R26596 DVSS DVSS.n4359 0.0227222
R26597 DVSS DVSS.n9597 0.0227222
R26598 DVSS.n9731 DVSS 0.0227222
R26599 DVSS.n11167 DVSS 0.0227222
R26600 DVSS DVSS.n9789 0.0227222
R26601 DVSS DVSS.n4015 0.0227222
R26602 DVSS DVSS.n9032 0.0227222
R26603 DVSS DVSS.n5536 0.0227222
R26604 DVSS.n10002 DVSS 0.0227222
R26605 DVSS.n14376 DVSS.n14375 0.0226831
R26606 DVSS.n14380 DVSS.n14379 0.0226831
R26607 DVSS.n14414 DVSS.n14413 0.0226831
R26608 DVSS.n14423 DVSS.n14422 0.0226831
R26609 DVSS.n14520 DVSS.n14519 0.0226831
R26610 DVSS.n14516 DVSS.n14515 0.0226831
R26611 DVSS.n14512 DVSS.n14511 0.0226831
R26612 DVSS.n19648 DVSS.n19647 0.0226831
R26613 DVSS.n19697 DVSS.n19696 0.0226831
R26614 DVSS.n19701 DVSS.n19700 0.0226831
R26615 DVSS.n19710 DVSS.n19709 0.0226831
R26616 DVSS.n19714 DVSS.n19713 0.0226831
R26617 DVSS.n19758 DVSS.n19757 0.0226831
R26618 DVSS.n19810 DVSS.n19809 0.0226831
R26619 DVSS.n19806 DVSS.n19805 0.0226831
R26620 DVSS.n19802 DVSS.n19801 0.0226831
R26621 DVSS.n19793 DVSS.n19792 0.0226831
R26622 DVSS.n19789 DVSS.n19788 0.0226831
R26623 DVSS.n19780 DVSS.n19779 0.0226831
R26624 DVSS.n19776 DVSS.n19775 0.0226831
R26625 DVSS.n132 DVSS.n131 0.0226831
R26626 DVSS.n141 DVSS.n140 0.0226831
R26627 DVSS.n145 DVSS.n144 0.0226831
R26628 DVSS.n158 DVSS.n157 0.0226831
R26629 DVSS.n162 DVSS.n161 0.0226831
R26630 DVSS.n251 DVSS.n250 0.0226831
R26631 DVSS.n247 DVSS.n246 0.0226831
R26632 DVSS.n243 DVSS.n242 0.0226831
R26633 DVSS.n234 DVSS.n233 0.0226831
R26634 DVSS.n230 DVSS.n229 0.0226831
R26635 DVSS.n221 DVSS.n220 0.0226831
R26636 DVSS.n217 DVSS.n216 0.0226831
R26637 DVSS.n204 DVSS.n203 0.0226831
R26638 DVSS.n200 DVSS.n199 0.0226831
R26639 DVSS.n191 DVSS.n190 0.0226831
R26640 DVSS.n187 DVSS.n186 0.0226831
R26641 DVSS.n14774 DVSS.n14773 0.0226831
R26642 DVSS.n14770 DVSS.n14769 0.0226831
R26643 DVSS.n14714 DVSS.n14713 0.0226831
R26644 DVSS.n14705 DVSS.n14704 0.0226831
R26645 DVSS.n14617 DVSS.n14616 0.0226831
R26646 DVSS.n14613 DVSS.n14612 0.0226831
R26647 DVSS.n14609 DVSS.n14608 0.0226831
R26648 DVSS.n19857 DVSS.n19856 0.0226831
R26649 DVSS.n19916 DVSS.n19915 0.0226831
R26650 DVSS.n19920 DVSS.n19919 0.0226831
R26651 DVSS.n19929 DVSS.n19928 0.0226831
R26652 DVSS.n19933 DVSS.n19932 0.0226831
R26653 DVSS.n19983 DVSS.n19982 0.0226831
R26654 DVSS.n20035 DVSS.n20034 0.0226831
R26655 DVSS.n20031 DVSS.n20030 0.0226831
R26656 DVSS.n20027 DVSS.n20026 0.0226831
R26657 DVSS.n20018 DVSS.n20017 0.0226831
R26658 DVSS.n20014 DVSS.n20013 0.0226831
R26659 DVSS.n20005 DVSS.n20004 0.0226831
R26660 DVSS.n20001 DVSS.n20000 0.0226831
R26661 DVSS.n292 DVSS.n291 0.0226831
R26662 DVSS.n301 DVSS.n300 0.0226831
R26663 DVSS.n305 DVSS.n304 0.0226831
R26664 DVSS.n318 DVSS.n317 0.0226831
R26665 DVSS.n322 DVSS.n321 0.0226831
R26666 DVSS.n459 DVSS.n458 0.0226831
R26667 DVSS.n455 DVSS.n454 0.0226831
R26668 DVSS.n451 DVSS.n450 0.0226831
R26669 DVSS.n442 DVSS.n441 0.0226831
R26670 DVSS.n438 DVSS.n437 0.0226831
R26671 DVSS.n429 DVSS.n428 0.0226831
R26672 DVSS.n425 DVSS.n424 0.0226831
R26673 DVSS.n412 DVSS.n411 0.0226831
R26674 DVSS.n408 DVSS.n407 0.0226831
R26675 DVSS.n399 DVSS.n398 0.0226831
R26676 DVSS.n395 DVSS.n394 0.0226831
R26677 DVSS.n18594 DVSS.n18592 0.0223919
R26678 DVSS.n18598 DVSS.n18594 0.0223919
R26679 DVSS.n18598 DVSS.n18597 0.0223919
R26680 DVSS.n7426 DVSS.n7424 0.0223919
R26681 DVSS.n7430 DVSS.n7426 0.0223919
R26682 DVSS.n7430 DVSS.n7429 0.0223919
R26683 DVSS.n14212 DVSS.n14211 0.0223919
R26684 DVSS.n14235 DVSS.n14229 0.0223919
R26685 DVSS.n14235 DVSS.n14234 0.0223919
R26686 DVSS.n14234 DVSS.n14232 0.0223919
R26687 DVSS.n13982 DVSS.n13980 0.0223919
R26688 DVSS.n13986 DVSS.n13982 0.0223919
R26689 DVSS.n13986 DVSS.n13985 0.0223919
R26690 DVSS.n13990 DVSS.n13988 0.0223919
R26691 DVSS.n7799 DVSS.n7793 0.0223919
R26692 DVSS.n7799 DVSS.n7798 0.0223919
R26693 DVSS.n7798 DVSS.n7796 0.0223919
R26694 DVSS.n7791 DVSS.n7785 0.0223919
R26695 DVSS.n7791 DVSS.n7790 0.0223919
R26696 DVSS.n7790 DVSS.n7788 0.0223919
R26697 DVSS.n18701 DVSS.n18697 0.0223919
R26698 DVSS.n18701 DVSS.n18699 0.0223919
R26699 DVSS.n7338 DVSS.n7336 0.0223919
R26700 DVSS.n7346 DVSS.n7338 0.0223919
R26701 DVSS.n7346 DVSS.n7344 0.0223919
R26702 DVSS.n7344 DVSS.n7342 0.0223919
R26703 DVSS.n14341 DVSS.n14340 0.0223919
R26704 DVSS.n14340 DVSS.n14338 0.0223919
R26705 DVSS.n14333 DVSS.n14327 0.0223919
R26706 DVSS.n14333 DVSS.n14331 0.0223919
R26707 DVSS.n14331 DVSS.n14329 0.0223919
R26708 DVSS.n14805 DVSS.n14801 0.0223919
R26709 DVSS.n14805 DVSS.n14803 0.0223919
R26710 DVSS.n14045 DVSS.n14043 0.0223919
R26711 DVSS.n13695 DVSS.n13693 0.0223919
R26712 DVSS.n7838 DVSS.n7837 0.0223919
R26713 DVSS.n7842 DVSS.n7840 0.0223919
R26714 DVSS.n7850 DVSS.n7842 0.0223919
R26715 DVSS.n7850 DVSS.n7849 0.0223919
R26716 DVSS.n7849 DVSS.n7847 0.0223919
R26717 DVSS.n19141 DVSS.n19139 0.0223919
R26718 DVSS.n19415 DVSS.n19413 0.0223919
R26719 DVSS.n19640 DVSS.n19638 0.0223919
R26720 DVSS.n19663 DVSS.n19661 0.0223919
R26721 DVSS.n19898 DVSS.n19896 0.0223919
R26722 DVSS.n19878 DVSS.n19870 0.0223919
R26723 DVSS.n19878 DVSS.n19877 0.0223919
R26724 DVSS.n20152 DVSS.n20138 0.0223919
R26725 DVSS.n20152 DVSS.n20151 0.0223919
R26726 DVSS.n20423 DVSS.n20421 0.0223919
R26727 DVSS.n7017 DVSS.n7016 0.0223919
R26728 DVSS.n7016 DVSS.n7014 0.0223919
R26729 DVSS.n7014 DVSS.n7013 0.0223919
R26730 DVSS.n7013 DVSS.n7011 0.0223919
R26731 DVSS.n7011 DVSS.n7010 0.0223919
R26732 DVSS.n7010 DVSS.n7008 0.0223919
R26733 DVSS.n7008 DVSS.n7007 0.0223919
R26734 DVSS.n7007 DVSS.n7005 0.0223919
R26735 DVSS.n18720 DVSS.n18718 0.0223919
R26736 DVSS.n18724 DVSS.n18720 0.0223919
R26737 DVSS.n18724 DVSS.n18723 0.0223919
R26738 DVSS.n18730 DVSS.n18728 0.0223919
R26739 DVSS.n18734 DVSS.n18730 0.0223919
R26740 DVSS.n18734 DVSS.n18733 0.0223919
R26741 DVSS.n14354 DVSS.n14352 0.0223919
R26742 DVSS.n14364 DVSS.n14360 0.0223919
R26743 DVSS.n14364 DVSS.n14362 0.0223919
R26744 DVSS.n14790 DVSS.n14788 0.0223919
R26745 DVSS.n14059 DVSS.n14053 0.0223919
R26746 DVSS.n14059 DVSS.n14057 0.0223919
R26747 DVSS.n14057 DVSS.n14055 0.0223919
R26748 DVSS.n7856 DVSS.n7852 0.0223919
R26749 DVSS.n7856 DVSS.n7854 0.0223919
R26750 DVSS.n7860 DVSS.n7858 0.0223919
R26751 DVSS.n7864 DVSS.n7860 0.0223919
R26752 DVSS.n7864 DVSS.n7862 0.0223919
R26753 DVSS.n13196 DVSS.n13194 0.0223919
R26754 DVSS.n13198 DVSS.n13196 0.0223919
R26755 DVSS.n13278 DVSS.n13276 0.0223919
R26756 DVSS.n13280 DVSS.n13278 0.0223919
R26757 DVSS.n13282 DVSS.n13280 0.0223919
R26758 DVSS.n13284 DVSS.n13282 0.0223919
R26759 DVSS.n13287 DVSS.n13284 0.0223919
R26760 DVSS.n11615 DVSS.n11614 0.0217598
R26761 DVSS.n6656 DVSS.n6655 0.0217598
R26762 DVSS.n19762 DVSS.n19761 0.0214155
R26763 DVSS.n166 DVSS.n165 0.0214155
R26764 DVSS.n19987 DVSS.n19986 0.0214155
R26765 DVSS.n326 DVSS.n325 0.0214155
R26766 DVSS.n17479 DVSS.n17478 0.0212042
R26767 DVSS.n17886 DVSS.n17885 0.0212042
R26768 DVSS.n18027 DVSS.n18026 0.0212042
R26769 DVSS.n7578 DVSS.n7577 0.0212042
R26770 DVSS.n18510 DVSS.n18509 0.0212042
R26771 DVSS.n18555 DVSS.n18554 0.0212042
R26772 DVSS.n19652 DVSS.n19651 0.0212042
R26773 DVSS.n19706 DVSS.n19705 0.0212042
R26774 DVSS.n19785 DVSS.n19784 0.0212042
R26775 DVSS.n137 DVSS.n136 0.0212042
R26776 DVSS.n226 DVSS.n225 0.0212042
R26777 DVSS.n195 DVSS.n194 0.0212042
R26778 DVSS.n16820 DVSS.n16819 0.0212042
R26779 DVSS.n15813 DVSS.n15812 0.0212042
R26780 DVSS.n15749 DVSS.n15748 0.0212042
R26781 DVSS.n15231 DVSS.n15230 0.0212042
R26782 DVSS.n7751 DVSS.n7750 0.0212042
R26783 DVSS.n13921 DVSS.n13920 0.0212042
R26784 DVSS.n19861 DVSS.n19860 0.0212042
R26785 DVSS.n19925 DVSS.n19924 0.0212042
R26786 DVSS.n20010 DVSS.n20009 0.0212042
R26787 DVSS.n297 DVSS.n296 0.0212042
R26788 DVSS.n434 DVSS.n433 0.0212042
R26789 DVSS.n403 DVSS.n402 0.0212042
R26790 DVSS.n6129 DVSS.n6128 0.0212
R26791 DVSS.n1371 DVSS.n1370 0.0211145
R26792 DVSS.n13967 DVSS.n13966 0.0210354
R26793 DVSS.n16802 DVSS.n16801 0.0210354
R26794 DVSS.n15070 DVSS.n15069 0.0210354
R26795 DVSS.n7640 DVSS.n7639 0.0210354
R26796 DVSS.n16009 DVSS.n16008 0.0210354
R26797 DVSS.n15306 DVSS.n15305 0.0210354
R26798 DVSS.n18351 DVSS.n18350 0.0210354
R26799 DVSS.n18008 DVSS.n18007 0.0210354
R26800 DVSS.n17867 DVSS.n17866 0.0210354
R26801 DVSS.n16500 DVSS.n16499 0.020993
R26802 DVSS.n17814 DVSS.n17807 0.020993
R26803 DVSS.n17955 DVSS.n17948 0.020993
R26804 DVSS.n18096 DVSS.n18089 0.020993
R26805 DVSS.n7604 DVSS.n7603 0.020993
R26806 DVSS.n18421 DVSS.n18420 0.020993
R26807 DVSS.n18529 DVSS.n18528 0.020993
R26808 DVSS.n19653 DVSS.n19652 0.020993
R26809 DVSS.n19705 DVSS.n19704 0.020993
R26810 DVSS.n19784 DVSS.n19783 0.020993
R26811 DVSS.n136 DVSS.n135 0.020993
R26812 DVSS.n225 DVSS.n224 0.020993
R26813 DVSS.n196 DVSS.n195 0.020993
R26814 DVSS.n16846 DVSS.n16845 0.020993
R26815 DVSS.n15787 DVSS.n15786 0.020993
R26816 DVSS.n15775 DVSS.n15774 0.020993
R26817 DVSS.n15374 DVSS.n15373 0.020993
R26818 DVSS.n15367 DVSS.n15366 0.020993
R26819 DVSS.n15217 DVSS.n15216 0.020993
R26820 DVSS.n13864 DVSS.n13857 0.020993
R26821 DVSS.n19862 DVSS.n19861 0.020993
R26822 DVSS.n19924 DVSS.n19923 0.020993
R26823 DVSS.n20009 DVSS.n20008 0.020993
R26824 DVSS.n296 DVSS.n295 0.020993
R26825 DVSS.n433 DVSS.n432 0.020993
R26826 DVSS.n404 DVSS.n403 0.020993
R26827 DVSS.n18423 DVSS.n18422 0.0207817
R26828 DVSS.n15209 DVSS.n15205 0.0207817
R26829 DVSS.n19165 DVSS.n19163 0.0207703
R26830 DVSS.n19114 DVSS.n19113 0.0207703
R26831 DVSS.n19435 DVSS.n19433 0.0207703
R26832 DVSS.n19389 DVSS.n19388 0.0207703
R26833 DVSS.n20173 DVSS.n20171 0.0207703
R26834 DVSS.n20146 DVSS.n20145 0.0207703
R26835 DVSS.n20443 DVSS.n20441 0.0207703
R26836 DVSS.n20397 DVSS.n20396 0.0207703
R26837 DVSS.n18097 DVSS.n18096 0.0205704
R26838 DVSS.n15375 DVSS.n15374 0.0205704
R26839 DVSS.n18499 DVSS.n18498 0.0203592
R26840 DVSS.n7740 DVSS.n7739 0.0203592
R26841 DVSS.n10638 DVSS.n10637 0.0203552
R26842 DVSS.n13347 DVSS.n13344 0.0201277
R26843 DVSS.n14457 DVSS.n14456 0.0199366
R26844 DVSS.n14665 DVSS.n14664 0.0199366
R26845 DVSS.n14208 DVSS.n14207 0.0198883
R26846 DVSS.n14200 DVSS.n14198 0.0198883
R26847 DVSS.n14192 DVSS.n14191 0.0198883
R26848 DVSS.n1334 DVSS.n1331 0.0198883
R26849 DVSS.n14690 DVSS.n14678 0.0198883
R26850 DVSS.n6012 DVSS.n6011 0.01985
R26851 DVSS.n12393 DVSS.n12392 0.0196339
R26852 DVSS.n3019 DVSS.n3018 0.0196339
R26853 DVSS.n14410 DVSS.n14409 0.0193028
R26854 DVSS.n14718 DVSS.n14717 0.0193028
R26855 DVSS.n14521 DVSS.n14502 0.0191189
R26856 DVSS.n8041 DVSS.n8040 0.0191034
R26857 DVSS.n6902 DVSS.n6901 0.0191034
R26858 DVSS.n5618 DVSS.n5617 0.0191024
R26859 DVSS.n5622 DVSS.n5621 0.0191024
R26860 DVSS.n5633 DVSS.n5632 0.0191024
R26861 DVSS.n5640 DVSS.n5639 0.0191024
R26862 DVSS.n5644 DVSS.n5643 0.0191024
R26863 DVSS.n5786 DVSS.n5785 0.0191024
R26864 DVSS.n5782 DVSS.n5781 0.0191024
R26865 DVSS.n5775 DVSS.n5774 0.0191024
R26866 DVSS.n5764 DVSS.n5763 0.0191024
R26867 DVSS.n5760 DVSS.n5759 0.0191024
R26868 DVSS.n4466 DVSS.n4465 0.0191024
R26869 DVSS.n4462 DVSS.n4461 0.0191024
R26870 DVSS.n4455 DVSS.n4454 0.0191024
R26871 DVSS.n4451 DVSS.n4450 0.0191024
R26872 DVSS.n4447 DVSS.n4446 0.0191024
R26873 DVSS.n4440 DVSS.n4439 0.0191024
R26874 DVSS.n4436 DVSS.n4435 0.0191024
R26875 DVSS.n4427 DVSS.n4426 0.0191024
R26876 DVSS.n4423 DVSS.n4422 0.0191024
R26877 DVSS.n4419 DVSS.n4418 0.0191024
R26878 DVSS.n4413 DVSS.n4412 0.0191024
R26879 DVSS.n4409 DVSS.n4408 0.0191024
R26880 DVSS.n4400 DVSS.n4399 0.0191024
R26881 DVSS.n4396 DVSS.n4395 0.0191024
R26882 DVSS.n4075 DVSS.n4074 0.0191024
R26883 DVSS.n4071 DVSS.n4070 0.0191024
R26884 DVSS.n4060 DVSS.n4059 0.0191024
R26885 DVSS.n4056 DVSS.n4055 0.0191024
R26886 DVSS.n4049 DVSS.n4048 0.0191024
R26887 DVSS.n6977 DVSS.n6976 0.0191024
R26888 DVSS.n6981 DVSS.n6980 0.0191024
R26889 DVSS.n7101 DVSS.n7100 0.0191024
R26890 DVSS.n7108 DVSS.n7107 0.0191024
R26891 DVSS.n7213 DVSS.n7212 0.0191024
R26892 DVSS.n7209 DVSS.n7208 0.0191024
R26893 DVSS.n7205 DVSS.n7204 0.0191024
R26894 DVSS.n19121 DVSS.n19120 0.0191024
R26895 DVSS.n19125 DVSS.n19124 0.0191024
R26896 DVSS.n19180 DVSS.n19179 0.0191024
R26897 DVSS.n19184 DVSS.n19183 0.0191024
R26898 DVSS.n19193 DVSS.n19192 0.0191024
R26899 DVSS.n19197 DVSS.n19196 0.0191024
R26900 DVSS.n19252 DVSS.n19251 0.0191024
R26901 DVSS.n19299 DVSS.n19298 0.0191024
R26902 DVSS.n19295 DVSS.n19294 0.0191024
R26903 DVSS.n19291 DVSS.n19290 0.0191024
R26904 DVSS.n19284 DVSS.n19283 0.0191024
R26905 DVSS.n19280 DVSS.n19279 0.0191024
R26906 DVSS.n19271 DVSS.n19270 0.0191024
R26907 DVSS.n19267 DVSS.n19266 0.0191024
R26908 DVSS.n843 DVSS.n842 0.0191024
R26909 DVSS.n852 DVSS.n851 0.0191024
R26910 DVSS.n856 DVSS.n855 0.0191024
R26911 DVSS.n867 DVSS.n866 0.0191024
R26912 DVSS.n871 DVSS.n870 0.0191024
R26913 DVSS.n1054 DVSS.n1053 0.0191024
R26914 DVSS.n1050 DVSS.n1049 0.0191024
R26915 DVSS.n1046 DVSS.n1045 0.0191024
R26916 DVSS.n1039 DVSS.n1038 0.0191024
R26917 DVSS.n1035 DVSS.n1034 0.0191024
R26918 DVSS.n1026 DVSS.n1025 0.0191024
R26919 DVSS.n1022 DVSS.n1021 0.0191024
R26920 DVSS.n1012 DVSS.n1011 0.0191024
R26921 DVSS.n1008 DVSS.n1007 0.0191024
R26922 DVSS.n999 DVSS.n998 0.0191024
R26923 DVSS.n995 DVSS.n994 0.0191024
R26924 DVSS.n10907 DVSS.n10906 0.0191024
R26925 DVSS.n10911 DVSS.n10910 0.0191024
R26926 DVSS.n10924 DVSS.n10923 0.0191024
R26927 DVSS.n10933 DVSS.n10932 0.0191024
R26928 DVSS.n10937 DVSS.n10936 0.0191024
R26929 DVSS.n11293 DVSS.n11292 0.0191024
R26930 DVSS.n11289 DVSS.n11288 0.0191024
R26931 DVSS.n11280 DVSS.n11279 0.0191024
R26932 DVSS.n11267 DVSS.n11266 0.0191024
R26933 DVSS.n11263 DVSS.n11262 0.0191024
R26934 DVSS.n9493 DVSS.n9492 0.0191024
R26935 DVSS.n9497 DVSS.n9496 0.0191024
R26936 DVSS.n9504 DVSS.n9503 0.0191024
R26937 DVSS.n9508 DVSS.n9507 0.0191024
R26938 DVSS.n9512 DVSS.n9511 0.0191024
R26939 DVSS.n9521 DVSS.n9520 0.0191024
R26940 DVSS.n9525 DVSS.n9524 0.0191024
R26941 DVSS.n9534 DVSS.n9533 0.0191024
R26942 DVSS.n9538 DVSS.n9537 0.0191024
R26943 DVSS.n9551 DVSS.n9550 0.0191024
R26944 DVSS.n9555 DVSS.n9554 0.0191024
R26945 DVSS.n9564 DVSS.n9563 0.0191024
R26946 DVSS.n9568 DVSS.n9567 0.0191024
R26947 DVSS.n8994 DVSS.n8993 0.0191024
R26948 DVSS.n8990 DVSS.n8989 0.0191024
R26949 DVSS.n13121 DVSS.n13120 0.0191024
R26950 DVSS.n13125 DVSS.n13124 0.0191024
R26951 DVSS.n13134 DVSS.n13133 0.0191024
R26952 DVSS.n12957 DVSS.n12956 0.0191024
R26953 DVSS.n12961 DVSS.n12960 0.0191024
R26954 DVSS.n12937 DVSS.n12936 0.0191024
R26955 DVSS.n12933 DVSS.n12932 0.0191024
R26956 DVSS.n12924 DVSS.n12923 0.0191024
R26957 DVSS.n12916 DVSS.n12915 0.0191024
R26958 DVSS.n12912 DVSS.n12911 0.0191024
R26959 DVSS.n12905 DVSS.n12904 0.0191024
R26960 DVSS.n12901 DVSS.n12900 0.0191024
R26961 DVSS.n12897 DVSS.n12896 0.0191024
R26962 DVSS.n12888 DVSS.n12887 0.0191024
R26963 DVSS.n12884 DVSS.n12883 0.0191024
R26964 DVSS.n12875 DVSS.n12874 0.0191024
R26965 DVSS.n12871 DVSS.n12870 0.0191024
R26966 DVSS.n12858 DVSS.n12857 0.0191024
R26967 DVSS.n12854 DVSS.n12853 0.0191024
R26968 DVSS.n12845 DVSS.n12844 0.0191024
R26969 DVSS.n12841 DVSS.n12840 0.0191024
R26970 DVSS.n17040 DVSS.n17039 0.0191024
R26971 DVSS.n17044 DVSS.n17043 0.0191024
R26972 DVSS.n17057 DVSS.n17056 0.0191024
R26973 DVSS.n17066 DVSS.n17065 0.0191024
R26974 DVSS.n17070 DVSS.n17069 0.0191024
R26975 DVSS.n17572 DVSS.n17571 0.0191024
R26976 DVSS.n17576 DVSS.n17575 0.0191024
R26977 DVSS.n17585 DVSS.n17584 0.0191024
R26978 DVSS.n17598 DVSS.n17597 0.0191024
R26979 DVSS.n17602 DVSS.n17601 0.0191024
R26980 DVSS.n15704 DVSS.n15703 0.0191024
R26981 DVSS.n15700 DVSS.n15699 0.0191024
R26982 DVSS.n15693 DVSS.n15692 0.0191024
R26983 DVSS.n15689 DVSS.n15688 0.0191024
R26984 DVSS.n15685 DVSS.n15684 0.0191024
R26985 DVSS.n15676 DVSS.n15675 0.0191024
R26986 DVSS.n15672 DVSS.n15671 0.0191024
R26987 DVSS.n15663 DVSS.n15662 0.0191024
R26988 DVSS.n15659 DVSS.n15658 0.0191024
R26989 DVSS.n15646 DVSS.n15645 0.0191024
R26990 DVSS.n15642 DVSS.n15641 0.0191024
R26991 DVSS.n15633 DVSS.n15632 0.0191024
R26992 DVSS.n15629 DVSS.n15628 0.0191024
R26993 DVSS.n15001 DVSS.n15000 0.0191024
R26994 DVSS.n15005 DVSS.n15004 0.0191024
R26995 DVSS.n15016 DVSS.n15015 0.0191024
R26996 DVSS.n15020 DVSS.n15019 0.0191024
R26997 DVSS.n15029 DVSS.n15028 0.0191024
R26998 DVSS.n13661 DVSS.n13660 0.0191024
R26999 DVSS.n13657 DVSS.n13656 0.0191024
R27000 DVSS.n13582 DVSS.n13581 0.0191024
R27001 DVSS.n13573 DVSS.n13572 0.0191024
R27002 DVSS.n13516 DVSS.n13515 0.0191024
R27003 DVSS.n13512 DVSS.n13511 0.0191024
R27004 DVSS.n13508 DVSS.n13507 0.0191024
R27005 DVSS.n20121 DVSS.n20120 0.0191024
R27006 DVSS.n20125 DVSS.n20124 0.0191024
R27007 DVSS.n20191 DVSS.n20190 0.0191024
R27008 DVSS.n20195 DVSS.n20194 0.0191024
R27009 DVSS.n20204 DVSS.n20203 0.0191024
R27010 DVSS.n20208 DVSS.n20207 0.0191024
R27011 DVSS.n20263 DVSS.n20262 0.0191024
R27012 DVSS.n20315 DVSS.n20314 0.0191024
R27013 DVSS.n20311 DVSS.n20310 0.0191024
R27014 DVSS.n20307 DVSS.n20306 0.0191024
R27015 DVSS.n20298 DVSS.n20297 0.0191024
R27016 DVSS.n20294 DVSS.n20293 0.0191024
R27017 DVSS.n20285 DVSS.n20284 0.0191024
R27018 DVSS.n20281 DVSS.n20280 0.0191024
R27019 DVSS.n20826 DVSS.n20825 0.0191024
R27020 DVSS.n20835 DVSS.n20834 0.0191024
R27021 DVSS.n20839 DVSS.n20838 0.0191024
R27022 DVSS.n20852 DVSS.n20851 0.0191024
R27023 DVSS.n20856 DVSS.n20855 0.0191024
R27024 DVSS.n20821 DVSS.n20820 0.0191024
R27025 DVSS.n20817 DVSS.n20816 0.0191024
R27026 DVSS.n20813 DVSS.n20812 0.0191024
R27027 DVSS.n20804 DVSS.n20803 0.0191024
R27028 DVSS.n20800 DVSS.n20799 0.0191024
R27029 DVSS.n20791 DVSS.n20790 0.0191024
R27030 DVSS.n20787 DVSS.n20786 0.0191024
R27031 DVSS.n20774 DVSS.n20773 0.0191024
R27032 DVSS.n20770 DVSS.n20769 0.0191024
R27033 DVSS.n20761 DVSS.n20760 0.0191024
R27034 DVSS.n20757 DVSS.n20756 0.0191024
R27035 DVSS.n10855 DVSS.n10854 0.0191024
R27036 DVSS.n10851 DVSS.n10850 0.0191024
R27037 DVSS.n10838 DVSS.n10837 0.0191024
R27038 DVSS.n10829 DVSS.n10828 0.0191024
R27039 DVSS.n10825 DVSS.n10824 0.0191024
R27040 DVSS.n11369 DVSS.n11368 0.0191024
R27041 DVSS.n11373 DVSS.n11372 0.0191024
R27042 DVSS.n11382 DVSS.n11381 0.0191024
R27043 DVSS.n11395 DVSS.n11394 0.0191024
R27044 DVSS.n11399 DVSS.n11398 0.0191024
R27045 DVSS.n11531 DVSS.n11530 0.0191024
R27046 DVSS.n11535 DVSS.n11534 0.0191024
R27047 DVSS.n11542 DVSS.n11541 0.0191024
R27048 DVSS.n11546 DVSS.n11545 0.0191024
R27049 DVSS.n11550 DVSS.n11549 0.0191024
R27050 DVSS.n11559 DVSS.n11558 0.0191024
R27051 DVSS.n11563 DVSS.n11562 0.0191024
R27052 DVSS.n11572 DVSS.n11571 0.0191024
R27053 DVSS.n11576 DVSS.n11575 0.0191024
R27054 DVSS.n11589 DVSS.n11588 0.0191024
R27055 DVSS.n11593 DVSS.n11592 0.0191024
R27056 DVSS.n11602 DVSS.n11601 0.0191024
R27057 DVSS.n11606 DVSS.n11605 0.0191024
R27058 DVSS.n11698 DVSS.n11697 0.0191024
R27059 DVSS.n11702 DVSS.n11701 0.0191024
R27060 DVSS.n13080 DVSS.n13079 0.0191024
R27061 DVSS.n13076 DVSS.n13075 0.0191024
R27062 DVSS.n13067 DVSS.n13066 0.0191024
R27063 DVSS.n13035 DVSS.n13034 0.0191024
R27064 DVSS.n13031 DVSS.n13030 0.0191024
R27065 DVSS.n12035 DVSS.n12034 0.0191024
R27066 DVSS.n12039 DVSS.n12038 0.0191024
R27067 DVSS.n12048 DVSS.n12047 0.0191024
R27068 DVSS.n12056 DVSS.n12055 0.0191024
R27069 DVSS.n12060 DVSS.n12059 0.0191024
R27070 DVSS.n12090 DVSS.n12089 0.0191024
R27071 DVSS.n12086 DVSS.n12085 0.0191024
R27072 DVSS.n12082 DVSS.n12081 0.0191024
R27073 DVSS.n12073 DVSS.n12072 0.0191024
R27074 DVSS.n12069 DVSS.n12068 0.0191024
R27075 DVSS.n21 DVSS.n20 0.0191024
R27076 DVSS.n25 DVSS.n24 0.0191024
R27077 DVSS.n38 DVSS.n37 0.0191024
R27078 DVSS.n42 DVSS.n41 0.0191024
R27079 DVSS.n51 DVSS.n50 0.0191024
R27080 DVSS.n55 DVSS.n54 0.0191024
R27081 DVSS.n68 DVSS.n67 0.0191024
R27082 DVSS.n72 DVSS.n71 0.0191024
R27083 DVSS.n21554 DVSS.n21553 0.0191024
R27084 DVSS.n21550 DVSS.n21549 0.0191024
R27085 DVSS.n21546 DVSS.n21545 0.0191024
R27086 DVSS.n21537 DVSS.n21536 0.0191024
R27087 DVSS.n21533 DVSS.n21532 0.0191024
R27088 DVSS.n21524 DVSS.n21523 0.0191024
R27089 DVSS.n21520 DVSS.n21519 0.0191024
R27090 DVSS.n21507 DVSS.n21506 0.0191024
R27091 DVSS.n21503 DVSS.n21502 0.0191024
R27092 DVSS.n21494 DVSS.n21493 0.0191024
R27093 DVSS.n21490 DVSS.n21489 0.0191024
R27094 DVSS.n21477 DVSS.n21476 0.0191024
R27095 DVSS.n21473 DVSS.n21472 0.0191024
R27096 DVSS.n21466 DVSS.n21465 0.0191024
R27097 DVSS.n21462 DVSS.n21461 0.0191024
R27098 DVSS.n21458 DVSS.n21457 0.0191024
R27099 DVSS.n21449 DVSS.n21448 0.0191024
R27100 DVSS.n21445 DVSS.n21444 0.0191024
R27101 DVSS.n21436 DVSS.n21435 0.0191024
R27102 DVSS.n21432 DVSS.n21431 0.0191024
R27103 DVSS.n21419 DVSS.n21418 0.0191024
R27104 DVSS.n21415 DVSS.n21414 0.0191024
R27105 DVSS.n21406 DVSS.n21405 0.0191024
R27106 DVSS.n21402 DVSS.n21401 0.0191024
R27107 DVSS.n5202 DVSS.n5201 0.0191024
R27108 DVSS.n5198 DVSS.n5197 0.0191024
R27109 DVSS.n4703 DVSS.n4702 0.0191024
R27110 DVSS.n4710 DVSS.n4709 0.0191024
R27111 DVSS.n4714 DVSS.n4713 0.0191024
R27112 DVSS.n4264 DVSS.n4263 0.0191024
R27113 DVSS.n4268 DVSS.n4267 0.0191024
R27114 DVSS.n4275 DVSS.n4274 0.0191024
R27115 DVSS.n4279 DVSS.n4278 0.0191024
R27116 DVSS.n4283 DVSS.n4282 0.0191024
R27117 DVSS.n4290 DVSS.n4289 0.0191024
R27118 DVSS.n4294 DVSS.n4293 0.0191024
R27119 DVSS.n4303 DVSS.n4302 0.0191024
R27120 DVSS.n4307 DVSS.n4306 0.0191024
R27121 DVSS.n4317 DVSS.n4316 0.0191024
R27122 DVSS.n4321 DVSS.n4320 0.0191024
R27123 DVSS.n4330 DVSS.n4329 0.0191024
R27124 DVSS.n4334 DVSS.n4333 0.0191024
R27125 DVSS.n3798 DVSS.n3797 0.0191024
R27126 DVSS.n3802 DVSS.n3801 0.0191024
R27127 DVSS.n3975 DVSS.n3974 0.0191024
R27128 DVSS.n3979 DVSS.n3978 0.0191024
R27129 DVSS.n3986 DVSS.n3985 0.0191024
R27130 DVSS.n3774 DVSS.n3773 0.0191024
R27131 DVSS.n3770 DVSS.n3769 0.0191024
R27132 DVSS.n3759 DVSS.n3758 0.0191024
R27133 DVSS.n3755 DVSS.n3754 0.0191024
R27134 DVSS.n3748 DVSS.n3747 0.0191024
R27135 DVSS.n3740 DVSS.n3739 0.0191024
R27136 DVSS.n3736 DVSS.n3735 0.0191024
R27137 DVSS.n3512 DVSS.n3511 0.0191024
R27138 DVSS.n3508 DVSS.n3507 0.0191024
R27139 DVSS.n3504 DVSS.n3503 0.0191024
R27140 DVSS.n3497 DVSS.n3496 0.0191024
R27141 DVSS.n3493 DVSS.n3492 0.0191024
R27142 DVSS.n3484 DVSS.n3483 0.0191024
R27143 DVSS.n3480 DVSS.n3479 0.0191024
R27144 DVSS.n3476 DVSS.n3475 0.0191024
R27145 DVSS.n3470 DVSS.n3469 0.0191024
R27146 DVSS.n3466 DVSS.n3465 0.0191024
R27147 DVSS.n3457 DVSS.n3456 0.0191024
R27148 DVSS.n3453 DVSS.n3452 0.0191024
R27149 DVSS.n9929 DVSS.n9928 0.0191024
R27150 DVSS.n9933 DVSS.n9932 0.0191024
R27151 DVSS.n9946 DVSS.n9945 0.0191024
R27152 DVSS.n9955 DVSS.n9954 0.0191024
R27153 DVSS.n9959 DVSS.n9958 0.0191024
R27154 DVSS.n11095 DVSS.n11094 0.0191024
R27155 DVSS.n11099 DVSS.n11098 0.0191024
R27156 DVSS.n11108 DVSS.n11107 0.0191024
R27157 DVSS.n11121 DVSS.n11120 0.0191024
R27158 DVSS.n11125 DVSS.n11124 0.0191024
R27159 DVSS.n9701 DVSS.n9700 0.0191024
R27160 DVSS.n9697 DVSS.n9696 0.0191024
R27161 DVSS.n9690 DVSS.n9689 0.0191024
R27162 DVSS.n9686 DVSS.n9685 0.0191024
R27163 DVSS.n9682 DVSS.n9681 0.0191024
R27164 DVSS.n9673 DVSS.n9672 0.0191024
R27165 DVSS.n9669 DVSS.n9668 0.0191024
R27166 DVSS.n9660 DVSS.n9659 0.0191024
R27167 DVSS.n9656 DVSS.n9655 0.0191024
R27168 DVSS.n9643 DVSS.n9642 0.0191024
R27169 DVSS.n9639 DVSS.n9638 0.0191024
R27170 DVSS.n9630 DVSS.n9629 0.0191024
R27171 DVSS.n9626 DVSS.n9625 0.0191024
R27172 DVSS.n9084 DVSS.n9083 0.0191024
R27173 DVSS.n9080 DVSS.n9079 0.0191024
R27174 DVSS.n9069 DVSS.n9068 0.0191024
R27175 DVSS.n9065 DVSS.n9064 0.0191024
R27176 DVSS.n9056 DVSS.n9055 0.0191024
R27177 DVSS.n13214 DVSS.n13213 0.0191024
R27178 DVSS.n13218 DVSS.n13217 0.0191024
R27179 DVSS.n13250 DVSS.n13249 0.0191024
R27180 DVSS.n13259 DVSS.n13258 0.0191024
R27181 DVSS.n13418 DVSS.n13417 0.0191024
R27182 DVSS.n13414 DVSS.n13413 0.0191024
R27183 DVSS.n13410 DVSS.n13409 0.0191024
R27184 DVSS.n20404 DVSS.n20403 0.0191024
R27185 DVSS.n20408 DVSS.n20407 0.0191024
R27186 DVSS.n20462 DVSS.n20461 0.0191024
R27187 DVSS.n20466 DVSS.n20465 0.0191024
R27188 DVSS.n20475 DVSS.n20474 0.0191024
R27189 DVSS.n20479 DVSS.n20478 0.0191024
R27190 DVSS.n20537 DVSS.n20536 0.0191024
R27191 DVSS.n20589 DVSS.n20588 0.0191024
R27192 DVSS.n20585 DVSS.n20584 0.0191024
R27193 DVSS.n20581 DVSS.n20580 0.0191024
R27194 DVSS.n20572 DVSS.n20571 0.0191024
R27195 DVSS.n20568 DVSS.n20567 0.0191024
R27196 DVSS.n20559 DVSS.n20558 0.0191024
R27197 DVSS.n20555 DVSS.n20554 0.0191024
R27198 DVSS.n21052 DVSS.n21051 0.0191024
R27199 DVSS.n21061 DVSS.n21060 0.0191024
R27200 DVSS.n21065 DVSS.n21064 0.0191024
R27201 DVSS.n21078 DVSS.n21077 0.0191024
R27202 DVSS.n21082 DVSS.n21081 0.0191024
R27203 DVSS.n21047 DVSS.n21046 0.0191024
R27204 DVSS.n21043 DVSS.n21042 0.0191024
R27205 DVSS.n21039 DVSS.n21038 0.0191024
R27206 DVSS.n21030 DVSS.n21029 0.0191024
R27207 DVSS.n21026 DVSS.n21025 0.0191024
R27208 DVSS.n21017 DVSS.n21016 0.0191024
R27209 DVSS.n21013 DVSS.n21012 0.0191024
R27210 DVSS.n21000 DVSS.n20999 0.0191024
R27211 DVSS.n20996 DVSS.n20995 0.0191024
R27212 DVSS.n20987 DVSS.n20986 0.0191024
R27213 DVSS.n20983 DVSS.n20982 0.0191024
R27214 DVSS.n17337 DVSS.n17336 0.0191024
R27215 DVSS.n17341 DVSS.n17340 0.0191024
R27216 DVSS.n17352 DVSS.n17351 0.0191024
R27217 DVSS.n17359 DVSS.n17358 0.0191024
R27218 DVSS.n17363 DVSS.n17362 0.0191024
R27219 DVSS.n16407 DVSS.n16406 0.0191024
R27220 DVSS.n16403 DVSS.n16402 0.0191024
R27221 DVSS.n16396 DVSS.n16395 0.0191024
R27222 DVSS.n16385 DVSS.n16384 0.0191024
R27223 DVSS.n16381 DVSS.n16380 0.0191024
R27224 DVSS.n16216 DVSS.n16215 0.0191024
R27225 DVSS.n16212 DVSS.n16211 0.0191024
R27226 DVSS.n16205 DVSS.n16204 0.0191024
R27227 DVSS.n16201 DVSS.n16200 0.0191024
R27228 DVSS.n16197 DVSS.n16196 0.0191024
R27229 DVSS.n16190 DVSS.n16189 0.0191024
R27230 DVSS.n16186 DVSS.n16185 0.0191024
R27231 DVSS.n16177 DVSS.n16176 0.0191024
R27232 DVSS.n16173 DVSS.n16172 0.0191024
R27233 DVSS.n16162 DVSS.n16161 0.0191024
R27234 DVSS.n16158 DVSS.n16157 0.0191024
R27235 DVSS.n16149 DVSS.n16148 0.0191024
R27236 DVSS.n16145 DVSS.n16144 0.0191024
R27237 DVSS.n7540 DVSS.n7539 0.0191024
R27238 DVSS.n7536 DVSS.n7535 0.0191024
R27239 DVSS.n7525 DVSS.n7524 0.0191024
R27240 DVSS.n7521 DVSS.n7520 0.0191024
R27241 DVSS.n7514 DVSS.n7513 0.0191024
R27242 DVSS.n18744 DVSS.n18743 0.0191024
R27243 DVSS.n18748 DVSS.n18747 0.0191024
R27244 DVSS.n18780 DVSS.n18779 0.0191024
R27245 DVSS.n18787 DVSS.n18786 0.0191024
R27246 DVSS.n18873 DVSS.n18872 0.0191024
R27247 DVSS.n18869 DVSS.n18868 0.0191024
R27248 DVSS.n18865 DVSS.n18864 0.0191024
R27249 DVSS.n19395 DVSS.n19394 0.0191024
R27250 DVSS.n19399 DVSS.n19398 0.0191024
R27251 DVSS.n19451 DVSS.n19450 0.0191024
R27252 DVSS.n19455 DVSS.n19454 0.0191024
R27253 DVSS.n19464 DVSS.n19463 0.0191024
R27254 DVSS.n19468 DVSS.n19467 0.0191024
R27255 DVSS.n19523 DVSS.n19522 0.0191024
R27256 DVSS.n19570 DVSS.n19569 0.0191024
R27257 DVSS.n19566 DVSS.n19565 0.0191024
R27258 DVSS.n19562 DVSS.n19561 0.0191024
R27259 DVSS.n19555 DVSS.n19554 0.0191024
R27260 DVSS.n19551 DVSS.n19550 0.0191024
R27261 DVSS.n19542 DVSS.n19541 0.0191024
R27262 DVSS.n19538 DVSS.n19537 0.0191024
R27263 DVSS.n1130 DVSS.n1129 0.0191024
R27264 DVSS.n1139 DVSS.n1138 0.0191024
R27265 DVSS.n1143 DVSS.n1142 0.0191024
R27266 DVSS.n1154 DVSS.n1153 0.0191024
R27267 DVSS.n1158 DVSS.n1157 0.0191024
R27268 DVSS.n1269 DVSS.n1268 0.0191024
R27269 DVSS.n1265 DVSS.n1264 0.0191024
R27270 DVSS.n1261 DVSS.n1260 0.0191024
R27271 DVSS.n1254 DVSS.n1253 0.0191024
R27272 DVSS.n1250 DVSS.n1249 0.0191024
R27273 DVSS.n1241 DVSS.n1240 0.0191024
R27274 DVSS.n1237 DVSS.n1236 0.0191024
R27275 DVSS.n1227 DVSS.n1226 0.0191024
R27276 DVSS.n1223 DVSS.n1222 0.0191024
R27277 DVSS.n1214 DVSS.n1213 0.0191024
R27278 DVSS.n1210 DVSS.n1209 0.0191024
R27279 DVSS.n5413 DVSS.n5412 0.0191024
R27280 DVSS.n5417 DVSS.n5416 0.0191024
R27281 DVSS.n5428 DVSS.n5427 0.0191024
R27282 DVSS.n5435 DVSS.n5434 0.0191024
R27283 DVSS.n5439 DVSS.n5438 0.0191024
R27284 DVSS.n6056 DVSS.n6055 0.0191024
R27285 DVSS.n6060 DVSS.n6059 0.0191024
R27286 DVSS.n6067 DVSS.n6066 0.0191024
R27287 DVSS.n6078 DVSS.n6077 0.0191024
R27288 DVSS.n6082 DVSS.n6081 0.0191024
R27289 DVSS.n6578 DVSS.n6577 0.0191024
R27290 DVSS.n6582 DVSS.n6581 0.0191024
R27291 DVSS.n6589 DVSS.n6588 0.0191024
R27292 DVSS.n6593 DVSS.n6592 0.0191024
R27293 DVSS.n6597 DVSS.n6596 0.0191024
R27294 DVSS.n6604 DVSS.n6603 0.0191024
R27295 DVSS.n6608 DVSS.n6607 0.0191024
R27296 DVSS.n6617 DVSS.n6616 0.0191024
R27297 DVSS.n6621 DVSS.n6620 0.0191024
R27298 DVSS.n6632 DVSS.n6631 0.0191024
R27299 DVSS.n6636 DVSS.n6635 0.0191024
R27300 DVSS.n6645 DVSS.n6644 0.0191024
R27301 DVSS.n6649 DVSS.n6648 0.0191024
R27302 DVSS.n6779 DVSS.n6778 0.0191024
R27303 DVSS.n6783 DVSS.n6782 0.0191024
R27304 DVSS.n6823 DVSS.n6822 0.0191024
R27305 DVSS.n6827 DVSS.n6826 0.0191024
R27306 DVSS.n6834 DVSS.n6833 0.0191024
R27307 DVSS.n3587 DVSS.n3586 0.0191024
R27308 DVSS.n3591 DVSS.n3590 0.0191024
R27309 DVSS.n3632 DVSS.n3631 0.0191024
R27310 DVSS.n3636 DVSS.n3635 0.0191024
R27311 DVSS.n3643 DVSS.n3642 0.0191024
R27312 DVSS.n3651 DVSS.n3650 0.0191024
R27313 DVSS.n3655 DVSS.n3654 0.0191024
R27314 DVSS.n3574 DVSS.n3573 0.0191024
R27315 DVSS.n3570 DVSS.n3569 0.0191024
R27316 DVSS.n3566 DVSS.n3565 0.0191024
R27317 DVSS.n3559 DVSS.n3558 0.0191024
R27318 DVSS.n3555 DVSS.n3554 0.0191024
R27319 DVSS.n3546 DVSS.n3545 0.0191024
R27320 DVSS.n3542 DVSS.n3541 0.0191024
R27321 DVSS.n3538 DVSS.n3537 0.0191024
R27322 DVSS.n18943 DVSS.n18942 0.0191024
R27323 DVSS.n18952 DVSS.n18951 0.0191024
R27324 DVSS.n18956 DVSS.n18955 0.0191024
R27325 DVSS.n18967 DVSS.n18966 0.0191024
R27326 DVSS.n18971 DVSS.n18970 0.0191024
R27327 DVSS.n19018 DVSS.n19017 0.0191024
R27328 DVSS.n19014 DVSS.n19013 0.0191024
R27329 DVSS.n19010 DVSS.n19009 0.0191024
R27330 DVSS.n19003 DVSS.n19002 0.0191024
R27331 DVSS.n18999 DVSS.n18998 0.0191024
R27332 DVSS.n18990 DVSS.n18989 0.0191024
R27333 DVSS.n18986 DVSS.n18985 0.0191024
R27334 DVSS.n521 DVSS.n520 0.0191024
R27335 DVSS.n530 DVSS.n529 0.0191024
R27336 DVSS.n534 DVSS.n533 0.0191024
R27337 DVSS.n545 DVSS.n544 0.0191024
R27338 DVSS.n549 DVSS.n548 0.0191024
R27339 DVSS.n620 DVSS.n619 0.0191024
R27340 DVSS.n616 DVSS.n615 0.0191024
R27341 DVSS.n612 DVSS.n611 0.0191024
R27342 DVSS.n605 DVSS.n604 0.0191024
R27343 DVSS.n601 DVSS.n600 0.0191024
R27344 DVSS.n592 DVSS.n591 0.0191024
R27345 DVSS.n588 DVSS.n587 0.0191024
R27346 DVSS.n578 DVSS.n577 0.0191024
R27347 DVSS.n574 DVSS.n573 0.0191024
R27348 DVSS.n565 DVSS.n564 0.0191024
R27349 DVSS.n561 DVSS.n560 0.0191024
R27350 DVSS.n16641 DVSS.n16640 0.0190915
R27351 DVSS.n18170 DVSS.n18169 0.0190915
R27352 DVSS.n17182 DVSS.n17181 0.0190915
R27353 DVSS.n15570 DVSS.n15569 0.0190915
R27354 DVSS.n15818 DVSS.n15817 0.0190636
R27355 DVSS.n15744 DVSS.n15743 0.0190636
R27356 DVSS.n15572 DVSS.n15571 0.0190636
R27357 DVSS.n15236 DVSS.n15235 0.0190636
R27358 DVSS.n18515 DVSS.n18514 0.0190636
R27359 DVSS.n5756 DVSS.n5755 0.0189252
R27360 DVSS.n4067 DVSS.n4066 0.0189252
R27361 DVSS.n11259 DVSS.n11258 0.0189252
R27362 DVSS.n8986 DVSS.n8060 0.0189252
R27363 DVSS.n12965 DVSS.n12964 0.0189252
R27364 DVSS.n17606 DVSS.n17605 0.0189252
R27365 DVSS.n15009 DVSS.n15008 0.0189252
R27366 DVSS.n11403 DVSS.n11402 0.0189252
R27367 DVSS.n11706 DVSS.n11705 0.0189252
R27368 DVSS.n13027 DVSS.n13026 0.0189252
R27369 DVSS.n3806 DVSS.n3805 0.0189252
R27370 DVSS.n3766 DVSS.n3765 0.0189252
R27371 DVSS.n11129 DVSS.n11128 0.0189252
R27372 DVSS.n9076 DVSS.n9075 0.0189252
R27373 DVSS.n16377 DVSS.n16376 0.0189252
R27374 DVSS.n7532 DVSS.n7531 0.0189252
R27375 DVSS.n6086 DVSS.n6085 0.0189252
R27376 DVSS.n6787 DVSS.n6786 0.0189252
R27377 DVSS.n3595 DVSS.n3594 0.0189252
R27378 DVSS.n1447 DVSS.n1446 0.0188571
R27379 DVSS.n16971 DVSS.n16970 0.018852
R27380 DVSS.n381 DVSS.n380 0.0187841
R27381 DVSS.n17729 DVSS.n17728 0.018669
R27382 DVSS.n14384 DVSS.n14383 0.018669
R27383 DVSS.n15934 DVSS.n15933 0.018669
R27384 DVSS.n14766 DVSS.n14765 0.018669
R27385 DVSS.n13049 DVSS.n13048 0.0185709
R27386 DVSS.n3575 DVSS.n1378 0.0185709
R27387 DVSS.n19684 DVSS.n19683 0.0184577
R27388 DVSS.n19903 DVSS.n19902 0.0184577
R27389 DVSS.n14619 DVSS.n14618 0.0184525
R27390 DVSS.n17881 DVSS.n17880 0.0183973
R27391 DVSS.n18022 DVSS.n18021 0.0183973
R27392 DVSS.n18168 DVSS.n18167 0.0183973
R27393 DVSS.n7573 DVSS.n7572 0.0183973
R27394 DVSS.n7756 DVSS.n7755 0.0183973
R27395 DVSS.n170 DVSS.n169 0.0183973
R27396 DVSS.n169 DVSS.n168 0.0183973
R27397 DVSS.n5614 DVSS.n5613 0.0183937
R27398 DVSS.n10903 DVSS.n10902 0.0183937
R27399 DVSS.n17036 DVSS.n17035 0.0183937
R27400 DVSS.n10859 DVSS.n10858 0.0183937
R27401 DVSS.n5206 DVSS.n5205 0.0183937
R27402 DVSS.n9925 DVSS.n9924 0.0183937
R27403 DVSS.n17333 DVSS.n17332 0.0183937
R27404 DVSS.n5409 DVSS.n5408 0.0183937
R27405 DVSS.n16683 DVSS.n16682 0.0182575
R27406 DVSS.n17140 DVSS.n17139 0.0182575
R27407 DVSS.n16059 DVSS.n16058 0.0182465
R27408 DVSS.n15951 DVSS.n15950 0.0182465
R27409 DVSS.n5790 DVSS.n5789 0.0182165
R27410 DVSS.n4064 DVSS.n4063 0.0182165
R27411 DVSS.n11297 DVSS.n11296 0.0182165
R27412 DVSS.n13117 DVSS.n13116 0.0182165
R27413 DVSS.n12941 DVSS.n12940 0.0182165
R27414 DVSS.n17568 DVSS.n17567 0.0182165
R27415 DVSS.n15012 DVSS.n15011 0.0182165
R27416 DVSS.n11365 DVSS.n11364 0.0182165
R27417 DVSS.n13084 DVSS.n13083 0.0182165
R27418 DVSS.n12031 DVSS.n11732 0.0182165
R27419 DVSS.n3971 DVSS.n3970 0.0182165
R27420 DVSS.n3763 DVSS.n3762 0.0182165
R27421 DVSS.n11091 DVSS.n11090 0.0182165
R27422 DVSS.n9073 DVSS.n9072 0.0182165
R27423 DVSS.n16411 DVSS.n16410 0.0182165
R27424 DVSS.n7529 DVSS.n7528 0.0182165
R27425 DVSS.n6052 DVSS.n6051 0.0182165
R27426 DVSS.n6819 DVSS.n6818 0.0182165
R27427 DVSS.n3628 DVSS.n3627 0.0182165
R27428 DVSS.n173 DVSS.n172 0.0181177
R27429 DVSS.n5648 DVSS.n5647 0.0180394
R27430 DVSS.n4458 DVSS.n4457 0.0180394
R27431 DVSS.n19256 DVSS.n19255 0.0180394
R27432 DVSS.n875 DVSS.n874 0.0180394
R27433 DVSS.n10941 DVSS.n10940 0.0180394
R27434 DVSS.n9501 DVSS.n9500 0.0180394
R27435 DVSS.n12908 DVSS.n12907 0.0180394
R27436 DVSS.n17074 DVSS.n17073 0.0180394
R27437 DVSS.n15696 DVSS.n15695 0.0180394
R27438 DVSS.n20267 DVSS.n20266 0.0180394
R27439 DVSS.n20860 DVSS.n20859 0.0180394
R27440 DVSS.n10821 DVSS.n10820 0.0180394
R27441 DVSS.n11539 DVSS.n11538 0.0180394
R27442 DVSS.n12064 DVSS.n12063 0.0180394
R27443 DVSS.n76 DVSS.n75 0.0180394
R27444 DVSS.n21469 DVSS.n21468 0.0180394
R27445 DVSS.n4718 DVSS.n4717 0.0180394
R27446 DVSS.n4272 DVSS.n4271 0.0180394
R27447 DVSS.n3732 DVSS.n3731 0.0180394
R27448 DVSS.n9963 DVSS.n9962 0.0180394
R27449 DVSS.n9693 DVSS.n9692 0.0180394
R27450 DVSS.n20541 DVSS.n20540 0.0180394
R27451 DVSS.n21086 DVSS.n21085 0.0180394
R27452 DVSS.n17367 DVSS.n17366 0.0180394
R27453 DVSS.n16208 DVSS.n16207 0.0180394
R27454 DVSS.n19527 DVSS.n19526 0.0180394
R27455 DVSS.n1162 DVSS.n1161 0.0180394
R27456 DVSS.n5443 DVSS.n5442 0.0180394
R27457 DVSS.n6586 DVSS.n6585 0.0180394
R27458 DVSS.n3659 DVSS.n3658 0.0180394
R27459 DVSS.n18975 DVSS.n18974 0.0180394
R27460 DVSS.n553 DVSS.n552 0.0180394
R27461 DVSS.n16612 DVSS.n16588 0.0180352
R27462 DVSS.n16776 DVSS.n16775 0.0180352
R27463 DVSS.n14078 DVSS.n14077 0.0179734
R27464 DVSS.n14732 DVSS.n14731 0.0179734
R27465 DVSS.n4432 DVSS.n4431 0.0178622
R27466 DVSS.n4404 DVSS.n4403 0.0178622
R27467 DVSS.n19129 DVSS.n19128 0.0178622
R27468 DVSS.n19189 DVSS.n19188 0.0178622
R27469 DVSS.n19276 DVSS.n19275 0.0178622
R27470 DVSS.n848 DVSS.n847 0.0178622
R27471 DVSS.n1031 DVSS.n1030 0.0178622
R27472 DVSS.n1003 DVSS.n1002 0.0178622
R27473 DVSS.n9529 DVSS.n9528 0.0178622
R27474 DVSS.n9560 DVSS.n9559 0.0178622
R27475 DVSS.n12880 DVSS.n12879 0.0178622
R27476 DVSS.n12849 DVSS.n12848 0.0178622
R27477 DVSS.n15668 DVSS.n15667 0.0178622
R27478 DVSS.n15637 DVSS.n15636 0.0178622
R27479 DVSS.n20129 DVSS.n20128 0.0178622
R27480 DVSS.n20200 DVSS.n20199 0.0178622
R27481 DVSS.n20290 DVSS.n20289 0.0178622
R27482 DVSS.n20831 DVSS.n20830 0.0178622
R27483 DVSS.n20796 DVSS.n20795 0.0178622
R27484 DVSS.n20765 DVSS.n20764 0.0178622
R27485 DVSS.n11567 DVSS.n11566 0.0178622
R27486 DVSS.n11598 DVSS.n11597 0.0178622
R27487 DVSS.n47 DVSS.n46 0.0178622
R27488 DVSS.n21529 DVSS.n21528 0.0178622
R27489 DVSS.n21498 DVSS.n21497 0.0178622
R27490 DVSS.n21441 DVSS.n21440 0.0178622
R27491 DVSS.n21410 DVSS.n21409 0.0178622
R27492 DVSS.n4298 DVSS.n4297 0.0178622
R27493 DVSS.n4326 DVSS.n4325 0.0178622
R27494 DVSS.n3489 DVSS.n3488 0.0178622
R27495 DVSS.n3461 DVSS.n3460 0.0178622
R27496 DVSS.n9665 DVSS.n9664 0.0178622
R27497 DVSS.n9634 DVSS.n9633 0.0178622
R27498 DVSS.n20412 DVSS.n20411 0.0178622
R27499 DVSS.n20471 DVSS.n20470 0.0178622
R27500 DVSS.n20564 DVSS.n20563 0.0178622
R27501 DVSS.n21057 DVSS.n21056 0.0178622
R27502 DVSS.n21022 DVSS.n21021 0.0178622
R27503 DVSS.n20991 DVSS.n20990 0.0178622
R27504 DVSS.n16182 DVSS.n16181 0.0178622
R27505 DVSS.n16153 DVSS.n16152 0.0178622
R27506 DVSS.n19403 DVSS.n19402 0.0178622
R27507 DVSS.n19460 DVSS.n19459 0.0178622
R27508 DVSS.n19547 DVSS.n19546 0.0178622
R27509 DVSS.n1135 DVSS.n1134 0.0178622
R27510 DVSS.n1246 DVSS.n1245 0.0178622
R27511 DVSS.n1218 DVSS.n1217 0.0178622
R27512 DVSS.n6612 DVSS.n6611 0.0178622
R27513 DVSS.n6641 DVSS.n6640 0.0178622
R27514 DVSS.n3551 DVSS.n3550 0.0178622
R27515 DVSS.n18948 DVSS.n18947 0.0178622
R27516 DVSS.n18995 DVSS.n18994 0.0178622
R27517 DVSS.n526 DVSS.n525 0.0178622
R27518 DVSS.n597 DVSS.n596 0.0178622
R27519 DVSS.n569 DVSS.n568 0.0178622
R27520 DVSS.n4431 DVSS.n4430 0.017685
R27521 DVSS.n4405 DVSS.n4404 0.017685
R27522 DVSS.n19130 DVSS.n19129 0.017685
R27523 DVSS.n19188 DVSS.n19187 0.017685
R27524 DVSS.n19275 DVSS.n19274 0.017685
R27525 DVSS.n847 DVSS.n846 0.017685
R27526 DVSS.n1030 DVSS.n1029 0.017685
R27527 DVSS.n1004 DVSS.n1003 0.017685
R27528 DVSS.n9530 DVSS.n9529 0.017685
R27529 DVSS.n9559 DVSS.n9558 0.017685
R27530 DVSS.n12879 DVSS.n12878 0.017685
R27531 DVSS.n12850 DVSS.n12849 0.017685
R27532 DVSS.n15667 DVSS.n15666 0.017685
R27533 DVSS.n15638 DVSS.n15637 0.017685
R27534 DVSS.n20130 DVSS.n20129 0.017685
R27535 DVSS.n20199 DVSS.n20198 0.017685
R27536 DVSS.n20289 DVSS.n20288 0.017685
R27537 DVSS.n20830 DVSS.n20829 0.017685
R27538 DVSS.n20795 DVSS.n20794 0.017685
R27539 DVSS.n20766 DVSS.n20765 0.017685
R27540 DVSS.n11568 DVSS.n11567 0.017685
R27541 DVSS.n11597 DVSS.n11596 0.017685
R27542 DVSS.n17 DVSS.n16 0.017685
R27543 DVSS.n46 DVSS.n45 0.017685
R27544 DVSS.n21528 DVSS.n21527 0.017685
R27545 DVSS.n21499 DVSS.n21498 0.017685
R27546 DVSS.n21440 DVSS.n21439 0.017685
R27547 DVSS.n21411 DVSS.n21410 0.017685
R27548 DVSS.n4299 DVSS.n4298 0.017685
R27549 DVSS.n4325 DVSS.n4324 0.017685
R27550 DVSS.n3488 DVSS.n3487 0.017685
R27551 DVSS.n3462 DVSS.n3461 0.017685
R27552 DVSS.n9664 DVSS.n9663 0.017685
R27553 DVSS.n9635 DVSS.n9634 0.017685
R27554 DVSS.n20413 DVSS.n20412 0.017685
R27555 DVSS.n20470 DVSS.n20469 0.017685
R27556 DVSS.n20563 DVSS.n20562 0.017685
R27557 DVSS.n21056 DVSS.n21055 0.017685
R27558 DVSS.n21021 DVSS.n21020 0.017685
R27559 DVSS.n20992 DVSS.n20991 0.017685
R27560 DVSS.n16181 DVSS.n16180 0.017685
R27561 DVSS.n16154 DVSS.n16153 0.017685
R27562 DVSS.n19404 DVSS.n19403 0.017685
R27563 DVSS.n19459 DVSS.n19458 0.017685
R27564 DVSS.n19546 DVSS.n19545 0.017685
R27565 DVSS.n1134 DVSS.n1133 0.017685
R27566 DVSS.n1245 DVSS.n1244 0.017685
R27567 DVSS.n1219 DVSS.n1218 0.017685
R27568 DVSS.n6613 DVSS.n6612 0.017685
R27569 DVSS.n6640 DVSS.n6639 0.017685
R27570 DVSS.n3550 DVSS.n3549 0.017685
R27571 DVSS.n18947 DVSS.n18946 0.017685
R27572 DVSS.n18994 DVSS.n18993 0.017685
R27573 DVSS.n525 DVSS.n524 0.017685
R27574 DVSS.n596 DVSS.n595 0.017685
R27575 DVSS.n570 DVSS.n569 0.017685
R27576 DVSS.n7412 DVSS.n7409 0.0174947
R27577 DVSS.n7391 DVSS.n7388 0.0174947
R27578 DVSS.n7366 DVSS.n7361 0.0174947
R27579 DVSS.n1331 DVSS.n1326 0.0174947
R27580 DVSS.n7160 DVSS.n7156 0.0174947
R27581 DVSS.n7028 DVSS.n7024 0.0174947
R27582 DVSS.n13814 DVSS.n13811 0.0172553
R27583 DVSS.n13774 DVSS.n13771 0.0172553
R27584 DVSS.n13736 DVSS.n13731 0.0172553
R27585 DVSS.n13344 DVSS.n13339 0.0172553
R27586 DVSS.n7971 DVSS.n7970 0.0172553
R27587 DVSS.n7970 DVSS.n7966 0.0172553
R27588 DVSS.n13325 DVSS.n13321 0.0172553
R27589 DVSS.n13326 DVSS.n13325 0.0172553
R27590 DVSS.n19970 DVSS.n19969 0.0171062
R27591 DVSS.n19745 DVSS.n19744 0.0171062
R27592 DVSS.n17536 DVSS.n17532 0.0170278
R27593 DVSS.n15261 DVSS.n15249 0.0170278
R27594 DVSS.n18360 DVSS.n18359 0.0170278
R27595 DVSS.n18081 DVSS.n18080 0.0170278
R27596 DVSS.n17678 DVSS.n17675 0.0170278
R27597 DVSS.n17940 DVSS.n17939 0.0170278
R27598 DVSS.n15064 DVSS.n15060 0.0170278
R27599 DVSS.n17236 DVSS.n17235 0.0170278
R27600 DVSS.n7161 DVSS.n7160 0.017016
R27601 DVSS.n7029 DVSS.n7028 0.017016
R27602 DVSS.n12394 DVSS.n12393 0.0169764
R27603 DVSS.n3020 DVSS.n3019 0.0169764
R27604 DVSS.n18462 DVSS.n18461 0.0169489
R27605 DVSS.n15140 DVSS.n15139 0.0169489
R27606 DVSS.n5397 DVSS.n5396 0.0168408
R27607 DVSS.n7145 DVSS.n7144 0.0167992
R27608 DVSS.n13548 DVSS.n13547 0.0167992
R27609 DVSS.n13366 DVSS.n13365 0.0167992
R27610 DVSS.n18827 DVSS.n18826 0.0167992
R27611 DVSS.n16681 DVSS.n16680 0.0167676
R27612 DVSS.n17142 DVSS.n17141 0.0167676
R27613 DVSS.n18247 DVSS.n18246 0.0167379
R27614 DVSS.n15493 DVSS.n15492 0.0167379
R27615 DVSS.n19166 DVSS.n19165 0.0167162
R27616 DVSS.n19113 DVSS.n19111 0.0167162
R27617 DVSS.n19436 DVSS.n19435 0.0167162
R27618 DVSS.n19388 DVSS.n19386 0.0167162
R27619 DVSS.n20174 DVSS.n20173 0.0167162
R27620 DVSS.n20145 DVSS.n20143 0.0167162
R27621 DVSS.n20444 DVSS.n20443 0.0167162
R27622 DVSS.n20396 DVSS.n20394 0.0167162
R27623 DVSS.n18197 DVSS.n18196 0.0166324
R27624 DVSS.n15543 DVSS.n15542 0.0166324
R27625 DVSS.n18210 DVSS.n18209 0.0163158
R27626 DVSS.n15530 DVSS.n15529 0.0163158
R27627 DVSS.n7097 DVSS.n7096 0.0162677
R27628 DVSS.n13586 DVSS.n13585 0.0162677
R27629 DVSS.n13246 DVSS.n13245 0.0162677
R27630 DVSS.n18776 DVSS.n18775 0.0162677
R27631 DVSS.n18260 DVSS.n18259 0.0162103
R27632 DVSS.n15480 DVSS.n15479 0.0162103
R27633 DVSS.n9965 DVSS.n9964 0.0161472
R27634 DVSS.n17369 DVSS.n17368 0.0161472
R27635 DVSS.n18136 DVSS.n18135 0.0161047
R27636 DVSS.n18453 DVSS.n18452 0.0161047
R27637 DVSS.n15441 DVSS.n15440 0.0161047
R27638 DVSS.n15164 DVSS.n15163 0.0161047
R27639 DVSS.n4389 DVSS.n4388 0.0160906
R27640 DVSS.n9577 DVSS.n9576 0.0160906
R27641 DVSS.n15620 DVSS.n15619 0.0160906
R27642 DVSS.n4341 DVSS.n4340 0.0160906
R27643 DVSS.n9617 DVSS.n9616 0.0160906
R27644 DVSS.n16138 DVSS.n16137 0.0160906
R27645 DVSS.n12796 DVSS.n12795 0.0160769
R27646 DVSS.n20968 DVSS.n20967 0.0160299
R27647 DVSS.n980 DVSS.n979 0.0160299
R27648 DVSS.n18125 DVSS.n18124 0.0159992
R27649 DVSS.n15415 DVSS.n15414 0.0159992
R27650 DVSS.n14883 DVSS.n14882 0.0159869
R27651 DVSS.n11406 DVSS.n11405 0.0159134
R27652 DVSS.n6329 DVSS.n6328 0.0159134
R27653 DVSS.n3391 DVSS.n3390 0.0158846
R27654 DVSS.n6985 DVSS.n6984 0.0157362
R27655 DVSS.n13653 DVSS.n13652 0.0157362
R27656 DVSS.n13222 DVSS.n13221 0.0157362
R27657 DVSS.n18752 DVSS.n18751 0.0157362
R27658 DVSS.n16108 DVSS.n16107 0.0157113
R27659 DVSS.n19726 DVSS.n19725 0.0157113
R27660 DVSS.n15989 DVSS.n15988 0.0157113
R27661 DVSS.n19945 DVSS.n19944 0.0157113
R27662 DVSS.n18470 DVSS.n18469 0.0156825
R27663 DVSS.n15132 DVSS.n15131 0.0156825
R27664 DVSS.n3992 DVSS.n3991 0.0155982
R27665 DVSS.n9807 DVSS.n9806 0.0155982
R27666 DVSS.n9708 DVSS.n9707 0.0155982
R27667 DVSS.n9615 DVSS.n9614 0.0155982
R27668 DVSS.n9096 DVSS.n9095 0.0155982
R27669 DVSS.n9050 DVSS.n9049 0.0155982
R27670 DVSS.n20955 DVSS.n20954 0.0155982
R27671 DVSS.n20965 DVSS.n20955 0.0155982
R27672 DVSS.n16296 DVSS.n16295 0.0155982
R27673 DVSS.n16257 DVSS.n16256 0.0155982
R27674 DVSS.n16136 DVSS.n16135 0.0155982
R27675 DVSS.n18380 DVSS.n18379 0.0155982
R27676 DVSS.n7508 DVSS.n7507 0.0155982
R27677 DVSS.n18189 DVSS.n18188 0.015577
R27678 DVSS.n15551 DVSS.n15550 0.015577
R27679 DVSS.n17874 DVSS.n17873 0.015567
R27680 DVSS.n18015 DVSS.n18014 0.015567
R27681 DVSS.n18161 DVSS.n18160 0.015567
R27682 DVSS.n7566 DVSS.n7565 0.015567
R27683 DVSS.n15825 DVSS.n15824 0.015567
R27684 DVSS.n15737 DVSS.n15736 0.015567
R27685 DVSS.n15579 DVSS.n15578 0.015567
R27686 DVSS.n15243 DVSS.n15242 0.015567
R27687 DVSS.n18522 DVSS.n18521 0.015567
R27688 DVSS.n7763 DVSS.n7762 0.015567
R27689 DVSS.n6439 DVSS.n6438 0.0155658
R27690 DVSS.n6350 DVSS.n6349 0.0155658
R27691 DVSS.n6663 DVSS.n6662 0.0155658
R27692 DVSS.n6724 DVSS.n6723 0.0155658
R27693 DVSS.n6845 DVSS.n6844 0.0155658
R27694 DVSS.n19170 DVSS.n19169 0.0155591
R27695 DVSS.n20178 DVSS.n20177 0.0155591
R27696 DVSS.n20449 DVSS.n20448 0.0155591
R27697 DVSS.n19441 DVSS.n19440 0.0155591
R27698 DVSS.n17764 DVSS.n17763 0.0155
R27699 DVSS.n15899 DVSS.n15898 0.0155
R27700 DVSS.n10943 DVSS.n10942 0.0154808
R27701 DVSS.n17076 DVSS.n17075 0.0154808
R27702 DVSS.n4719 DVSS.n4698 0.0154808
R27703 DVSS.n5650 DVSS.n5649 0.0154808
R27704 DVSS.n20742 DVSS.n20741 0.0153635
R27705 DVSS.n1196 DVSS.n1195 0.0153635
R27706 DVSS.n14214 DVSS.n14213 0.0153205
R27707 DVSS.n16553 DVSS.n16552 0.0152887
R27708 DVSS.n16740 DVSS.n16739 0.0152887
R27709 DVSS.n18120 DVSS.n18119 0.0151547
R27710 DVSS.n18268 DVSS.n18267 0.0151547
R27711 DVSS.n15410 DVSS.n15409 0.0151547
R27712 DVSS.n15472 DVSS.n15471 0.0151547
R27713 DVSS.n19641 DVSS.n19640 0.0150946
R27714 DVSS.n19678 DVSS.n19677 0.0150946
R27715 DVSS.n19899 DVSS.n19898 0.0150946
R27716 DVSS.n19877 DVSS.n19875 0.0150946
R27717 DVSS.n16672 DVSS.n16671 0.0149435
R27718 DVSS.n18239 DVSS.n18238 0.0149435
R27719 DVSS.n17151 DVSS.n17150 0.0149435
R27720 DVSS.n15501 DVSS.n15500 0.0149435
R27721 DVSS.n6016 DVSS.n6015 0.0149
R27722 DVSS.n17797 DVSS.n17796 0.0148662
R27723 DVSS.n17671 DVSS.n17670 0.0148662
R27724 DVSS.n12392 DVSS.n12391 0.0148504
R27725 DVSS.n3018 DVSS.n3017 0.0148504
R27726 DVSS.n16067 DVSS.n16066 0.0148379
R27727 DVSS.n15959 DVSS.n15958 0.0148379
R27728 DVSS.n18874 DVSS.n18861 0.0147386
R27729 DVSS.n7214 DVSS.n7201 0.0147386
R27730 DVSS.n13419 DVSS.n13405 0.0147386
R27731 DVSS.n13518 DVSS.n13517 0.0147386
R27732 DVSS.n17771 DVSS.n17770 0.0146549
R27733 DVSS.n15892 DVSS.n15891 0.0146549
R27734 DVSS.n17944 DVSS.n7620 0.0146478
R27735 DVSS.n18085 DVSS.n7612 0.0146478
R27736 DVSS.n18159 DVSS.n7608 0.0146478
R27737 DVSS.n18416 DVSS.n7459 0.0146478
R27738 DVSS.n16110 DVSS.n16109 0.0146478
R27739 DVSS.n17762 DVSS.n17761 0.0146478
R27740 DVSS.n16555 DVSS.n16554 0.0146478
R27741 DVSS.n15827 DVSS.n15778 0.0146478
R27742 DVSS.n15734 DVSS.n7673 0.0146478
R27743 DVSS.n15581 DVSS.n15370 0.0146478
R27744 DVSS.n15245 DVSS.n15220 0.0146478
R27745 DVSS.n15991 DVSS.n15990 0.0146478
R27746 DVSS.n15901 DVSS.n15900 0.0146478
R27747 DVSS.n16741 DVSS.n16740 0.0146478
R27748 DVSS.n7765 DVSS.n7764 0.0146478
R27749 DVSS.n18525 DVSS.n18524 0.0146478
R27750 DVSS.n19742 DVSS.n19726 0.0146478
R27751 DVSS.n19967 DVSS.n19945 0.0146478
R27752 DVSS.n376 DVSS.n375 0.0146478
R27753 DVSS.n379 DVSS.n378 0.0146478
R27754 DVSS.n19811 DVSS.n19762 0.0146478
R27755 DVSS.n20036 DVSS.n19987 0.0146478
R27756 DVSS.n252 DVSS.n166 0.0146478
R27757 DVSS.n460 DVSS.n326 0.0146478
R27758 DVSS.n16099 DVSS.n16098 0.0146267
R27759 DVSS.n15980 DVSS.n15979 0.0146267
R27760 DVSS.n20249 DVSS.n20248 0.0146212
R27761 DVSS.n20523 DVSS.n20522 0.0146212
R27762 DVSS.n19510 DVSS.n19509 0.0146212
R27763 DVSS.n16649 DVSS.n16648 0.0145211
R27764 DVSS.n18218 DVSS.n18217 0.0145211
R27765 DVSS.n17174 DVSS.n17173 0.0145211
R27766 DVSS.n15522 DVSS.n15521 0.0145211
R27767 DVSS.n10734 DVSS.n8337 0.0144961
R27768 DVSS.n5859 DVSS.n5858 0.0144961
R27769 DVSS.n18445 DVSS.n18444 0.0144155
R27770 DVSS.n15172 DVSS.n15171 0.0144155
R27771 DVSS.n17945 DVSS.n17944 0.0143948
R27772 DVSS.n18086 DVSS.n18085 0.0143948
R27773 DVSS.n7608 DVSS.n7607 0.0143948
R27774 DVSS.n18417 DVSS.n18416 0.0143948
R27775 DVSS.n16554 DVSS.n16553 0.0143948
R27776 DVSS.n16109 DVSS.n16108 0.0143948
R27777 DVSS.n17763 DVSS.n17762 0.0143948
R27778 DVSS.n15735 DVSS.n15734 0.0143948
R27779 DVSS.n15827 DVSS.n15826 0.0143948
R27780 DVSS.n15245 DVSS.n15244 0.0143948
R27781 DVSS.n15581 DVSS.n15580 0.0143948
R27782 DVSS.n16742 DVSS.n16741 0.0143948
R27783 DVSS.n15990 DVSS.n15989 0.0143948
R27784 DVSS.n15900 DVSS.n15899 0.0143948
R27785 DVSS.n18524 DVSS.n18523 0.0143948
R27786 DVSS.n13854 DVSS.n7765 0.0143948
R27787 DVSS.n19743 DVSS.n19742 0.0143948
R27788 DVSS.n19968 DVSS.n19967 0.0143948
R27789 DVSS.n377 DVSS.n376 0.0143948
R27790 DVSS.n378 DVSS.n377 0.0143948
R27791 DVSS.n19811 DVSS.n19810 0.0143948
R27792 DVSS.n20036 DVSS.n20035 0.0143948
R27793 DVSS.n460 DVSS.n459 0.0143948
R27794 DVSS.n252 DVSS.n251 0.0143948
R27795 DVSS.n17737 DVSS.n17736 0.0143098
R27796 DVSS.n18144 DVSS.n18143 0.0143098
R27797 DVSS.n15926 DVSS.n15925 0.0143098
R27798 DVSS.n15449 DVSS.n15448 0.0143098
R27799 DVSS.n16582 DVSS.n16581 0.0142042
R27800 DVSS.n16769 DVSS.n16768 0.0142042
R27801 DVSS.n6442 DVSS.n6441 0.0141909
R27802 DVSS.n6353 DVSS.n6352 0.0141909
R27803 DVSS.n6660 DVSS.n6659 0.0141909
R27804 DVSS.n6721 DVSS.n6720 0.0141909
R27805 DVSS.n6842 DVSS.n6841 0.0141909
R27806 DVSS.n11486 DVSS.n11485 0.0141618
R27807 DVSS.n11523 DVSS.n11522 0.0141618
R27808 DVSS.n11648 DVSS.n11647 0.0141618
R27809 DVSS.n11685 DVSS.n11684 0.0141618
R27810 DVSS.n13056 DVSS.n13055 0.0141618
R27811 DVSS.n991 DVSS.n990 0.0141417
R27812 DVSS.n10818 DVSS.n10817 0.0141417
R27813 DVSS.n16166 DVSS.n16165 0.0141417
R27814 DVSS.n5446 DVSS.n5445 0.0141417
R27815 DVSS.n6628 DVSS.n6627 0.0141417
R27816 DVSS.n7438 DVSS.n7436 0.0140754
R27817 DVSS.n7441 DVSS.n7438 0.0140754
R27818 DVSS.n7443 DVSS.n7441 0.0140754
R27819 DVSS.n7446 DVSS.n7443 0.0140754
R27820 DVSS.n7448 DVSS.n7446 0.0140754
R27821 DVSS.n18571 DVSS.n7448 0.0140754
R27822 DVSS.n18571 DVSS.n18568 0.0140754
R27823 DVSS.n18568 DVSS.n18566 0.0140754
R27824 DVSS.n18561 DVSS.n7450 0.0140754
R27825 DVSS.n14888 DVSS.n14886 0.0140754
R27826 DVSS.n5376 DVSS.n5374 0.0140754
R27827 DVSS.n5374 DVSS.n5373 0.0140754
R27828 DVSS.n5600 DVSS.n5594 0.0140754
R27829 DVSS.n5600 DVSS.n5597 0.0140754
R27830 DVSS.n17318 DVSS.n17312 0.0140754
R27831 DVSS.n17318 DVSS.n17315 0.0140754
R27832 DVSS.n17296 DVSS.n17294 0.0140754
R27833 DVSS.n17294 DVSS.n17293 0.0140754
R27834 DVSS.n17293 DVSS.n17291 0.0140754
R27835 DVSS.n17291 DVSS.n17290 0.0140754
R27836 DVSS.n16980 DVSS.n16977 0.0140754
R27837 DVSS.n16982 DVSS.n16980 0.0140754
R27838 DVSS.n16985 DVSS.n16982 0.0140754
R27839 DVSS.n16987 DVSS.n16985 0.0140754
R27840 DVSS.n17022 DVSS.n17017 0.0140754
R27841 DVSS.n17022 DVSS.n17021 0.0140754
R27842 DVSS.n10230 DVSS.n10227 0.0140754
R27843 DVSS.n10232 DVSS.n10230 0.0140754
R27844 DVSS.n10283 DVSS.n10278 0.0140754
R27845 DVSS.n10283 DVSS.n10282 0.0140754
R27846 DVSS.n14922 DVSS.n14920 0.0140754
R27847 DVSS.n14925 DVSS.n14922 0.0140754
R27848 DVSS.n14931 DVSS.n14929 0.0140754
R27849 DVSS.n14934 DVSS.n14931 0.0140754
R27850 DVSS.n14936 DVSS.n14934 0.0140754
R27851 DVSS.n14939 DVSS.n14936 0.0140754
R27852 DVSS.n14941 DVSS.n14939 0.0140754
R27853 DVSS.n14952 DVSS.n14941 0.0140754
R27854 DVSS.n14952 DVSS.n14949 0.0140754
R27855 DVSS.n14949 DVSS.n14947 0.0140754
R27856 DVSS.n8010 DVSS.n8008 0.0140754
R27857 DVSS.n8013 DVSS.n8010 0.0140754
R27858 DVSS.n8015 DVSS.n8013 0.0140754
R27859 DVSS.n8018 DVSS.n8015 0.0140754
R27860 DVSS.n8020 DVSS.n8018 0.0140754
R27861 DVSS.n13179 DVSS.n8020 0.0140754
R27862 DVSS.n13179 DVSS.n13176 0.0140754
R27863 DVSS.n13176 DVSS.n13174 0.0140754
R27864 DVSS.n13169 DVSS.n13167 0.0140754
R27865 DVSS.n13167 DVSS.n13165 0.0140754
R27866 DVSS.n13165 DVSS.n13162 0.0140754
R27867 DVSS.n13162 DVSS.n13160 0.0140754
R27868 DVSS.n13160 DVSS.n13157 0.0140754
R27869 DVSS.n13157 DVSS.n13155 0.0140754
R27870 DVSS.n13155 DVSS.n8048 0.0140754
R27871 DVSS.n8048 DVSS.n8046 0.0140754
R27872 DVSS.n8040 DVSS.n8038 0.0140754
R27873 DVSS.n8038 DVSS.n8036 0.0140754
R27874 DVSS.n6901 DVSS.n1376 0.0140754
R27875 DVSS.n6909 DVSS.n6907 0.0140754
R27876 DVSS.n6912 DVSS.n6909 0.0140754
R27877 DVSS.n6914 DVSS.n6912 0.0140754
R27878 DVSS.n6917 DVSS.n6914 0.0140754
R27879 DVSS.n6919 DVSS.n6917 0.0140754
R27880 DVSS.n6922 DVSS.n6919 0.0140754
R27881 DVSS.n6924 DVSS.n6922 0.0140754
R27882 DVSS.n6926 DVSS.n6924 0.0140754
R27883 DVSS.n6933 DVSS.n6931 0.0140754
R27884 DVSS.n6936 DVSS.n6933 0.0140754
R27885 DVSS.n6938 DVSS.n6936 0.0140754
R27886 DVSS.n6941 DVSS.n6938 0.0140754
R27887 DVSS.n6943 DVSS.n6941 0.0140754
R27888 DVSS.n6950 DVSS.n6943 0.0140754
R27889 DVSS.n6950 DVSS.n6947 0.0140754
R27890 DVSS.n6947 DVSS.n6945 0.0140754
R27891 DVSS.n19239 DVSS.n19238 0.0139547
R27892 DVSS.n5402 DVSS.n5400 0.013824
R27893 DVSS.n1376 DVSS.n1374 0.013824
R27894 DVSS.n12828 DVSS.n12827 0.0137198
R27895 DVSS.n21138 DVSS.n21137 0.0137198
R27896 DVSS.n21137 DVSS.n21136 0.0137198
R27897 DVSS.n3788 DVSS.n3787 0.0137198
R27898 DVSS.n13849 DVSS.n13848 0.0136815
R27899 DVSS.n12943 DVSS.n12942 0.0136815
R27900 DVSS.n13183 DVSS.n13182 0.0136815
R27901 DVSS.n18575 DVSS.n18574 0.0136815
R27902 DVSS.n6954 DVSS.n6953 0.0136815
R27903 DVSS.n16533 DVSS.n16532 0.0135986
R27904 DVSS.n16575 DVSS.n16574 0.0135986
R27905 DVSS.n16085 DVSS.n16080 0.0135986
R27906 DVSS.n17744 DVSS.n17743 0.0135986
R27907 DVSS.n18104 DVSS.n18103 0.0135986
R27908 DVSS.n18130 DVSS.n18129 0.0135986
R27909 DVSS.n18255 DVSS.n18254 0.0135986
R27910 DVSS.n18202 DVSS.n18201 0.0135986
R27911 DVSS.n18458 DVSS.n18457 0.0135986
R27912 DVSS.n14393 DVSS.n14392 0.0135986
R27913 DVSS.n19668 DVSS.n19667 0.0135986
R27914 DVSS.n16720 DVSS.n16719 0.0135986
R27915 DVSS.n16762 DVSS.n16761 0.0135986
R27916 DVSS.n15973 DVSS.n15972 0.0135986
R27917 DVSS.n15919 DVSS.n15918 0.0135986
R27918 DVSS.n15382 DVSS.n15381 0.0135986
R27919 DVSS.n15420 DVSS.n15419 0.0135986
R27920 DVSS.n15485 DVSS.n15484 0.0135986
R27921 DVSS.n15538 DVSS.n15537 0.0135986
R27922 DVSS.n15159 DVSS.n15158 0.0135986
R27923 DVSS.n14757 DVSS.n14756 0.0135986
R27924 DVSS.n19883 DVSS.n19882 0.0135986
R27925 DVSS.n11457 DVSS.n11456 0.0135244
R27926 DVSS.n11494 DVSS.n11493 0.0135244
R27927 DVSS.n11619 DVSS.n11618 0.0135244
R27928 DVSS.n11656 DVSS.n11655 0.0135244
R27929 DVSS.n13059 DVSS.n13058 0.0135244
R27930 DVSS.n19139 DVSS.n19137 0.013473
R27931 DVSS.n19107 DVSS.n19106 0.013473
R27932 DVSS.n19413 DVSS.n19411 0.013473
R27933 DVSS.n19379 DVSS.n19378 0.013473
R27934 DVSS.n20138 DVSS.n20136 0.013473
R27935 DVSS.n20151 DVSS.n20149 0.013473
R27936 DVSS.n20421 DVSS.n20419 0.013473
R27937 DVSS.n20384 DVSS.n20383 0.013473
R27938 DVSS.n6515 DVSS.n6514 0.0134466
R27939 DVSS.n9773 DVSS.n9772 0.0134466
R27940 DVSS.n9759 DVSS.n9758 0.0134466
R27941 DVSS.n9581 DVSS.n9580 0.0134466
R27942 DVSS.n9147 DVSS.n9146 0.0134466
R27943 DVSS.n15862 DVSS.n15861 0.0134466
R27944 DVSS.n15713 DVSS.n15712 0.0134466
R27945 DVSS.n15616 DVSS.n15615 0.0134466
R27946 DVSS.n14983 DVSS.n14982 0.0134466
R27947 DVSS.n13142 DVSS.n13141 0.0134466
R27948 DVSS.n15037 DVSS.n15036 0.0134466
R27949 DVSS.n4041 DVSS.n4040 0.0134466
R27950 DVSS.n4345 DVSS.n4344 0.0134466
R27951 DVSS.n4125 DVSS.n4124 0.0134466
R27952 DVSS.n12830 DVSS.n12829 0.0134331
R27953 DVSS.n3442 DVSS.n3441 0.0134331
R27954 DVSS.n7416 DVSS.n7414 0.0134255
R27955 DVSS.n7422 DVSS.n7416 0.0134255
R27956 DVSS.n7422 DVSS.n7421 0.0134255
R27957 DVSS.n7421 DVSS.n7419 0.0134255
R27958 DVSS.n18619 DVSS.n18611 0.0134255
R27959 DVSS.n18619 DVSS.n18618 0.0134255
R27960 DVSS.n18618 DVSS.n18616 0.0134255
R27961 DVSS.n14250 DVSS.n14248 0.0134255
R27962 DVSS.n14254 DVSS.n14250 0.0134255
R27963 DVSS.n14254 DVSS.n14253 0.0134255
R27964 DVSS.n14204 DVSS.n14202 0.0134255
R27965 DVSS.n14208 DVSS.n14204 0.0134255
R27966 DVSS.n13994 DVSS.n13992 0.0134255
R27967 DVSS.n13998 DVSS.n13994 0.0134255
R27968 DVSS.n13998 DVSS.n13997 0.0134255
R27969 DVSS.n14002 DVSS.n14000 0.0134255
R27970 DVSS.n14004 DVSS.n14002 0.0134255
R27971 DVSS.n7805 DVSS.n7803 0.0134255
R27972 DVSS.n7809 DVSS.n7805 0.0134255
R27973 DVSS.n7809 DVSS.n7808 0.0134255
R27974 DVSS.n13801 DVSS.n13799 0.0134255
R27975 DVSS.n13818 DVSS.n13801 0.0134255
R27976 DVSS.n13818 DVSS.n13817 0.0134255
R27977 DVSS.n13817 DVSS.n13815 0.0134255
R27978 DVSS.n7395 DVSS.n7393 0.0134255
R27979 DVSS.n7401 DVSS.n7395 0.0134255
R27980 DVSS.n7401 DVSS.n7399 0.0134255
R27981 DVSS.n7399 DVSS.n7397 0.0134255
R27982 DVSS.n18646 DVSS.n18638 0.0134255
R27983 DVSS.n18646 DVSS.n18644 0.0134255
R27984 DVSS.n18644 DVSS.n18642 0.0134255
R27985 DVSS.n14275 DVSS.n14273 0.0134255
R27986 DVSS.n14279 DVSS.n14275 0.0134255
R27987 DVSS.n14279 DVSS.n14277 0.0134255
R27988 DVSS.n14196 DVSS.n14194 0.0134255
R27989 DVSS.n14200 DVSS.n14196 0.0134255
R27990 DVSS.n14008 DVSS.n14006 0.0134255
R27991 DVSS.n14012 DVSS.n14008 0.0134255
R27992 DVSS.n14012 DVSS.n14010 0.0134255
R27993 DVSS.n14016 DVSS.n14014 0.0134255
R27994 DVSS.n14018 DVSS.n14016 0.0134255
R27995 DVSS.n7815 DVSS.n7813 0.0134255
R27996 DVSS.n7819 DVSS.n7815 0.0134255
R27997 DVSS.n7819 DVSS.n7817 0.0134255
R27998 DVSS.n13764 DVSS.n13762 0.0134255
R27999 DVSS.n13780 DVSS.n13764 0.0134255
R28000 DVSS.n13780 DVSS.n13778 0.0134255
R28001 DVSS.n13778 DVSS.n13776 0.0134255
R28002 DVSS.n7372 DVSS.n7369 0.0134255
R28003 DVSS.n7381 DVSS.n7372 0.0134255
R28004 DVSS.n7381 DVSS.n7380 0.0134255
R28005 DVSS.n7380 DVSS.n7377 0.0134255
R28006 DVSS.n18678 DVSS.n18666 0.0134255
R28007 DVSS.n18678 DVSS.n18677 0.0134255
R28008 DVSS.n18677 DVSS.n18674 0.0134255
R28009 DVSS.n14302 DVSS.n14299 0.0134255
R28010 DVSS.n14308 DVSS.n14302 0.0134255
R28011 DVSS.n14308 DVSS.n14307 0.0134255
R28012 DVSS.n14186 DVSS.n14183 0.0134255
R28013 DVSS.n14192 DVSS.n14186 0.0134255
R28014 DVSS.n14024 DVSS.n14021 0.0134255
R28015 DVSS.n14030 DVSS.n14024 0.0134255
R28016 DVSS.n14030 DVSS.n14029 0.0134255
R28017 DVSS.n14036 DVSS.n14033 0.0134255
R28018 DVSS.n14039 DVSS.n14036 0.0134255
R28019 DVSS.n7828 DVSS.n7825 0.0134255
R28020 DVSS.n7834 DVSS.n7828 0.0134255
R28021 DVSS.n7834 DVSS.n7833 0.0134255
R28022 DVSS.n13718 DVSS.n13715 0.0134255
R28023 DVSS.n13743 DVSS.n13718 0.0134255
R28024 DVSS.n13743 DVSS.n13742 0.0134255
R28025 DVSS.n13742 DVSS.n13739 0.0134255
R28026 DVSS.n1337 DVSS.n1334 0.0134255
R28027 DVSS.n1346 DVSS.n1337 0.0134255
R28028 DVSS.n1346 DVSS.n1343 0.0134255
R28029 DVSS.n1343 DVSS.n1340 0.0134255
R28030 DVSS.n7130 DVSS.n7121 0.0134255
R28031 DVSS.n7130 DVSS.n7127 0.0134255
R28032 DVSS.n7127 DVSS.n7124 0.0134255
R28033 DVSS.n7325 DVSS.n7322 0.0134255
R28034 DVSS.n7334 DVSS.n7325 0.0134255
R28035 DVSS.n7334 DVSS.n7333 0.0134255
R28036 DVSS.n7333 DVSS.n7330 0.0134255
R28037 DVSS.n18812 DVSS.n18800 0.0134255
R28038 DVSS.n18812 DVSS.n18811 0.0134255
R28039 DVSS.n18811 DVSS.n18808 0.0134255
R28040 DVSS.n14151 DVSS.n14148 0.0134255
R28041 DVSS.n14148 DVSS.n14145 0.0134255
R28042 DVSS.n14145 DVSS.n14142 0.0134255
R28043 DVSS.n14439 DVSS.n14436 0.0134255
R28044 DVSS.n14442 DVSS.n14439 0.0134255
R28045 DVSS.n14690 DVSS.n14689 0.0134255
R28046 DVSS.n14689 DVSS.n14686 0.0134255
R28047 DVSS.n14686 DVSS.n14685 0.0134255
R28048 DVSS.n14065 DVSS.n14062 0.0134255
R28049 DVSS.n14075 DVSS.n14065 0.0134255
R28050 DVSS.n14069 DVSS.n14067 0.0134255
R28051 DVSS.n7977 DVSS.n7975 0.0134255
R28052 DVSS.n7979 DVSS.n7977 0.0134255
R28053 DVSS.n7981 DVSS.n7979 0.0134255
R28054 DVSS.n7983 DVSS.n7981 0.0134255
R28055 DVSS.n7985 DVSS.n7983 0.0134255
R28056 DVSS.n7987 DVSS.n7985 0.0134255
R28057 DVSS.n7996 DVSS.n7993 0.0134255
R28058 DVSS.n8005 DVSS.n7996 0.0134255
R28059 DVSS.n8005 DVSS.n8004 0.0134255
R28060 DVSS.n8004 DVSS.n8001 0.0134255
R28061 DVSS.n13351 DVSS.n13272 0.0134255
R28062 DVSS.n13351 DVSS.n13350 0.0134255
R28063 DVSS.n13350 DVSS.n13347 0.0134255
R28064 DVSS.n7195 DVSS.n7191 0.0134255
R28065 DVSS.n7195 DVSS.n7193 0.0134255
R28066 DVSS.n18855 DVSS.n18853 0.0134255
R28067 DVSS.n14496 DVSS.n14494 0.0134255
R28068 DVSS.n14139 DVSS.n14137 0.0134255
R28069 DVSS.n14629 DVSS.n14625 0.0134255
R28070 DVSS.n14629 DVSS.n14628 0.0134255
R28071 DVSS.n14643 DVSS.n14641 0.0134255
R28072 DVSS.n7890 DVSS.n7886 0.0134255
R28073 DVSS.n7890 DVSS.n7888 0.0134255
R28074 DVSS.n13399 DVSS.n13394 0.0134255
R28075 DVSS.n13399 DVSS.n13397 0.0134255
R28076 DVSS.n7084 DVSS.n7042 0.0134255
R28077 DVSS.n7084 DVSS.n7082 0.0134255
R28078 DVSS.n7057 DVSS.n7055 0.0134255
R28079 DVSS.n7055 DVSS.n7054 0.0134255
R28080 DVSS.n14167 DVSS.n14165 0.0134255
R28081 DVSS.n14169 DVSS.n14167 0.0134255
R28082 DVSS.n14178 DVSS.n14169 0.0134255
R28083 DVSS.n14178 DVSS.n14176 0.0134255
R28084 DVSS.n14751 DVSS.n14738 0.0134255
R28085 DVSS.n14751 DVSS.n14749 0.0134255
R28086 DVSS.n14749 DVSS.n14747 0.0134255
R28087 DVSS.n14747 DVSS.n14745 0.0134255
R28088 DVSS.n13639 DVSS.n13616 0.0134255
R28089 DVSS.n13639 DVSS.n13636 0.0134255
R28090 DVSS.n13307 DVSS.n13305 0.0134255
R28091 DVSS.n13309 DVSS.n13307 0.0134255
R28092 DVSS.n16702 DVSS.n16701 0.0133873
R28093 DVSS.n17121 DVSS.n17120 0.0133873
R28094 DVSS.n6533 DVSS.n6532 0.0133291
R28095 DVSS.n4380 DVSS.n4379 0.0133291
R28096 DVSS.n4092 DVSS.n4091 0.0133291
R28097 DVSS.n6520 DVSS.n6519 0.0133291
R28098 DVSS.n9142 DVSS.n9141 0.0133291
R28099 DVSS.n9586 DVSS.n9585 0.0133291
R28100 DVSS.n9754 DVSS.n9753 0.0133291
R28101 DVSS.n9778 DVSS.n9777 0.0133291
R28102 DVSS.n15718 DVSS.n15717 0.0133291
R28103 DVSS.n15857 DVSS.n15856 0.0133291
R28104 DVSS.n14988 DVSS.n14987 0.0133291
R28105 DVSS.n15611 DVSS.n15610 0.0133291
R28106 DVSS.n13147 DVSS.n13146 0.0133291
R28107 DVSS.n4036 DVSS.n4035 0.0133291
R28108 DVSS.n15042 DVSS.n15041 0.0133291
R28109 DVSS.n4120 DVSS.n4119 0.0133291
R28110 DVSS.n4350 DVSS.n4349 0.0133291
R28111 DVSS.n3999 DVSS.n3998 0.0133291
R28112 DVSS.n9800 DVSS.n9799 0.0133291
R28113 DVSS.n9715 DVSS.n9714 0.0133291
R28114 DVSS.n9608 DVSS.n9607 0.0133291
R28115 DVSS.n9103 DVSS.n9102 0.0133291
R28116 DVSS.n9043 DVSS.n9042 0.0133291
R28117 DVSS.n16289 DVSS.n16288 0.0133291
R28118 DVSS.n16250 DVSS.n16249 0.0133291
R28119 DVSS.n16129 DVSS.n16128 0.0133291
R28120 DVSS.n18387 DVSS.n18386 0.0133291
R28121 DVSS.n7501 DVSS.n7500 0.0133291
R28122 DVSS.n19211 DVSS.n19210 0.0132559
R28123 DVSS.n20221 DVSS.n20220 0.0132559
R28124 DVSS.n20492 DVSS.n20491 0.0132559
R28125 DVSS.n19482 DVSS.n19481 0.0132559
R28126 DVSS.n18477 DVSS.n18476 0.0131761
R28127 DVSS.n15125 DVSS.n15124 0.0131761
R28128 DVSS.n5753 DVSS.n5752 0.0130787
R28129 DVSS.n11256 DVSS.n11255 0.0130787
R28130 DVSS.n17609 DVSS.n17608 0.0130787
R28131 DVSS.n11132 DVSS.n11131 0.0130787
R28132 DVSS.n16374 DVSS.n16373 0.0130787
R28133 DVSS.n5381 DVSS.n5379 0.0130698
R28134 DVSS.n5369 DVSS.n5368 0.0130698
R28135 DVSS.n5579 DVSS.n5578 0.0130698
R28136 DVSS.n17001 DVSS.n17000 0.0130698
R28137 DVSS.n17029 DVSS.n17028 0.0130698
R28138 DVSS.n10221 DVSS.n10220 0.0130698
R28139 DVSS.n10239 DVSS.n10237 0.0130698
R28140 DVSS.n10253 DVSS.n10252 0.0130698
R28141 DVSS.n10290 DVSS.n10289 0.0130698
R28142 DVSS.n18559 DVSS.n7451 0.0129759
R28143 DVSS.n14917 DVSS.n13975 0.0129759
R28144 DVSS.n18492 DVSS.n18491 0.0129648
R28145 DVSS.n7733 DVSS.n7732 0.0129648
R28146 DVSS.n5611 DVSS.n5610 0.0129016
R28147 DVSS.n10294 DVSS.n10293 0.0129016
R28148 DVSS.n12837 DVSS.n12836 0.0129016
R28149 DVSS.n17033 DVSS.n17032 0.0129016
R28150 DVSS.n10643 DVSS.n10642 0.0129016
R28151 DVSS.n5234 DVSS.n5233 0.0129016
R28152 DVSS.n3449 DVSS.n3448 0.0129016
R28153 DVSS.n9922 DVSS.n9921 0.0129016
R28154 DVSS.n17330 DVSS.n17329 0.0129016
R28155 DVSS.n5406 DVSS.n5405 0.0129016
R28156 DVSS.n3438 DVSS.n3437 0.0128976
R28157 DVSS.n6528 DVSS.n6527 0.0127801
R28158 DVSS.n4385 DVSS.n4384 0.0127801
R28159 DVSS.n4087 DVSS.n4086 0.0127801
R28160 DVSS.n18437 DVSS.n18436 0.0127535
R28161 DVSS.n14482 DVSS.n14481 0.0127535
R28162 DVSS.n15192 DVSS.n15191 0.0127535
R28163 DVSS.n14634 DVSS.n14633 0.0127535
R28164 DVSS.n18559 DVSS.n18558 0.0127233
R28165 DVSS.n14917 DVSS.n14916 0.0127233
R28166 DVSS.n17193 DVSS.n17192 0.01265
R28167 DVSS.n17196 DVSS.n17195 0.01265
R28168 DVSS.n17199 DVSS.n17198 0.01265
R28169 DVSS.n17202 DVSS.n17201 0.01265
R28170 DVSS.n17205 DVSS.n17204 0.01265
R28171 DVSS.n17208 DVSS.n17207 0.01265
R28172 DVSS.n17221 DVSS.n17220 0.01265
R28173 DVSS.n15215 DVSS.n15214 0.01265
R28174 DVSS.n15208 DVSS.n15207 0.01265
R28175 DVSS.n15116 DVSS.n15115 0.01265
R28176 DVSS.n15104 DVSS.n15103 0.01265
R28177 DVSS.n15101 DVSS.n15100 0.01265
R28178 DVSS.n15098 DVSS.n15097 0.01265
R28179 DVSS.n15095 DVSS.n15094 0.01265
R28180 DVSS.n15092 DVSS.n15091 0.01265
R28181 DVSS.n15089 DVSS.n15088 0.01265
R28182 DVSS.n15086 DVSS.n15085 0.01265
R28183 DVSS.n15083 DVSS.n15082 0.01265
R28184 DVSS.n15080 DVSS.n15079 0.01265
R28185 DVSS.n15077 DVSS.n15076 0.01265
R28186 DVSS.n15074 DVSS.n15073 0.01265
R28187 DVSS.n17717 DVSS.n17716 0.01265
R28188 DVSS.n17714 DVSS.n17713 0.01265
R28189 DVSS.n17711 DVSS.n17710 0.01265
R28190 DVSS.n17708 DVSS.n17707 0.01265
R28191 DVSS.n17705 DVSS.n17704 0.01265
R28192 DVSS.n17702 DVSS.n17701 0.01265
R28193 DVSS.n17699 DVSS.n17698 0.01265
R28194 DVSS.n17684 DVSS.n17683 0.01265
R28195 DVSS.n16498 DVSS.n16497 0.01265
R28196 DVSS.n16491 DVSS.n16490 0.01265
R28197 DVSS.n16487 DVSS.n16486 0.01265
R28198 DVSS.n16483 DVSS.n16482 0.01265
R28199 DVSS.n16479 DVSS.n16478 0.01265
R28200 DVSS.n16475 DVSS.n16474 0.01265
R28201 DVSS.n16471 DVSS.n16470 0.01265
R28202 DVSS.n16467 DVSS.n16466 0.01265
R28203 DVSS.n16463 DVSS.n16462 0.01265
R28204 DVSS.n16459 DVSS.n16458 0.01265
R28205 DVSS.n16455 DVSS.n16454 0.01265
R28206 DVSS.n16451 DVSS.n16450 0.01265
R28207 DVSS.n16447 DVSS.n16446 0.01265
R28208 DVSS.n16013 DVSS.n16012 0.01265
R28209 DVSS.n17491 DVSS.n16004 0.01265
R28210 DVSS.n17495 DVSS.n17494 0.01265
R28211 DVSS.n17498 DVSS.n17497 0.01265
R28212 DVSS.n17501 DVSS.n17500 0.01265
R28213 DVSS.n17504 DVSS.n17503 0.01265
R28214 DVSS.n17507 DVSS.n17506 0.01265
R28215 DVSS.n17510 DVSS.n17509 0.01265
R28216 DVSS.n17513 DVSS.n17512 0.01265
R28217 DVSS.n17516 DVSS.n17515 0.01265
R28218 DVSS.n17519 DVSS.n17518 0.01265
R28219 DVSS.n17522 DVSS.n17521 0.01265
R28220 DVSS.n17525 DVSS.n17524 0.01265
R28221 DVSS.n15365 DVSS.n15364 0.01265
R28222 DVSS.n15358 DVSS.n15357 0.01265
R28223 DVSS.n15354 DVSS.n15353 0.01265
R28224 DVSS.n15350 DVSS.n15349 0.01265
R28225 DVSS.n15346 DVSS.n15345 0.01265
R28226 DVSS.n15342 DVSS.n15341 0.01265
R28227 DVSS.n15338 DVSS.n15337 0.01265
R28228 DVSS.n15334 DVSS.n15333 0.01265
R28229 DVSS.n15330 DVSS.n15329 0.01265
R28230 DVSS.n15326 DVSS.n15325 0.01265
R28231 DVSS.n15322 DVSS.n15321 0.01265
R28232 DVSS.n15318 DVSS.n15317 0.01265
R28233 DVSS.n15314 DVSS.n15313 0.01265
R28234 DVSS.n15310 DVSS.n15309 0.01265
R28235 DVSS.n15300 DVSS.n7704 0.01265
R28236 DVSS.n15297 DVSS.n15296 0.01265
R28237 DVSS.n15294 DVSS.n15293 0.01265
R28238 DVSS.n15291 DVSS.n15290 0.01265
R28239 DVSS.n15288 DVSS.n15287 0.01265
R28240 DVSS.n15285 DVSS.n15284 0.01265
R28241 DVSS.n15282 DVSS.n15281 0.01265
R28242 DVSS.n15279 DVSS.n15278 0.01265
R28243 DVSS.n15276 DVSS.n15275 0.01265
R28244 DVSS.n15273 DVSS.n15272 0.01265
R28245 DVSS.n15270 DVSS.n15269 0.01265
R28246 DVSS.n15267 DVSS.n15266 0.01265
R28247 DVSS.n18095 DVSS.n18094 0.01265
R28248 DVSS.n18291 DVSS.n18290 0.01265
R28249 DVSS.n18325 DVSS.n18324 0.01265
R28250 DVSS.n17954 DVSS.n17953 0.01265
R28251 DVSS.n17958 DVSS.n17957 0.01265
R28252 DVSS.n17962 DVSS.n17961 0.01265
R28253 DVSS.n17966 DVSS.n17965 0.01265
R28254 DVSS.n17970 DVSS.n17969 0.01265
R28255 DVSS.n17974 DVSS.n17973 0.01265
R28256 DVSS.n17978 DVSS.n17977 0.01265
R28257 DVSS.n17982 DVSS.n17981 0.01265
R28258 DVSS.n17986 DVSS.n17985 0.01265
R28259 DVSS.n17990 DVSS.n17989 0.01265
R28260 DVSS.n17994 DVSS.n17993 0.01265
R28261 DVSS.n17998 DVSS.n17997 0.01265
R28262 DVSS.n18002 DVSS.n18001 0.01265
R28263 DVSS.n18012 DVSS.n18011 0.01265
R28264 DVSS.n18039 DVSS.n7619 0.01265
R28265 DVSS.n18043 DVSS.n18042 0.01265
R28266 DVSS.n18046 DVSS.n18045 0.01265
R28267 DVSS.n18049 DVSS.n18048 0.01265
R28268 DVSS.n18052 DVSS.n18051 0.01265
R28269 DVSS.n18055 DVSS.n18054 0.01265
R28270 DVSS.n18058 DVSS.n18057 0.01265
R28271 DVSS.n18061 DVSS.n18060 0.01265
R28272 DVSS.n18064 DVSS.n18063 0.01265
R28273 DVSS.n18067 DVSS.n18066 0.01265
R28274 DVSS.n18070 DVSS.n18069 0.01265
R28275 DVSS.n18073 DVSS.n18072 0.01265
R28276 DVSS.n17813 DVSS.n17812 0.01265
R28277 DVSS.n17817 DVSS.n17816 0.01265
R28278 DVSS.n17821 DVSS.n17820 0.01265
R28279 DVSS.n17825 DVSS.n17824 0.01265
R28280 DVSS.n17829 DVSS.n17828 0.01265
R28281 DVSS.n17833 DVSS.n17832 0.01265
R28282 DVSS.n17837 DVSS.n17836 0.01265
R28283 DVSS.n17841 DVSS.n17840 0.01265
R28284 DVSS.n17845 DVSS.n17844 0.01265
R28285 DVSS.n17849 DVSS.n17848 0.01265
R28286 DVSS.n17853 DVSS.n17852 0.01265
R28287 DVSS.n17857 DVSS.n17856 0.01265
R28288 DVSS.n17861 DVSS.n17860 0.01265
R28289 DVSS.n17871 DVSS.n17870 0.01265
R28290 DVSS.n17898 DVSS.n7627 0.01265
R28291 DVSS.n17902 DVSS.n17901 0.01265
R28292 DVSS.n17905 DVSS.n17904 0.01265
R28293 DVSS.n17908 DVSS.n17907 0.01265
R28294 DVSS.n17911 DVSS.n17910 0.01265
R28295 DVSS.n17914 DVSS.n17913 0.01265
R28296 DVSS.n17917 DVSS.n17916 0.01265
R28297 DVSS.n17920 DVSS.n17919 0.01265
R28298 DVSS.n17923 DVSS.n17922 0.01265
R28299 DVSS.n17926 DVSS.n17925 0.01265
R28300 DVSS.n17929 DVSS.n17928 0.01265
R28301 DVSS.n17932 DVSS.n17931 0.01265
R28302 DVSS.n13917 DVSS.n13916 0.01265
R28303 DVSS.n13933 DVSS.n13853 0.01265
R28304 DVSS.n13935 DVSS.n13934 0.01265
R28305 DVSS.n13938 DVSS.n13937 0.01265
R28306 DVSS.n13941 DVSS.n13940 0.01265
R28307 DVSS.n13944 DVSS.n13943 0.01265
R28308 DVSS.n13947 DVSS.n13946 0.01265
R28309 DVSS.n13950 DVSS.n13949 0.01265
R28310 DVSS.n13953 DVSS.n13952 0.01265
R28311 DVSS.n13956 DVSS.n13955 0.01265
R28312 DVSS.n13959 DVSS.n13958 0.01265
R28313 DVSS.n13962 DVSS.n13961 0.01265
R28314 DVSS.n13965 DVSS.n13964 0.01265
R28315 DVSS.n6526 DVSS.n6525 0.0125559
R28316 DVSS.n4387 DVSS.n4386 0.0125559
R28317 DVSS.n4085 DVSS.n4084 0.0125559
R28318 DVSS.n6512 DVSS.n6511 0.0125559
R28319 DVSS.n6523 DVSS.n6522 0.0125559
R28320 DVSS.n9771 DVSS.n9770 0.0125559
R28321 DVSS.n9780 DVSS.n9763 0.0125559
R28322 DVSS.n9761 DVSS.n9760 0.0125559
R28323 DVSS.n9751 DVSS.n8953 0.0125559
R28324 DVSS.n9579 DVSS.n9578 0.0125559
R28325 DVSS.n9588 DVSS.n9151 0.0125559
R28326 DVSS.n9149 DVSS.n9148 0.0125559
R28327 DVSS.n9139 DVSS.n9003 0.0125559
R28328 DVSS.n12966 DVSS.n12941 0.0125559
R28329 DVSS.n13115 DVSS.n8060 0.0125559
R28330 DVSS.n9503 DVSS.n9502 0.0125559
R28331 DVSS.n10901 DVSS.n10294 0.0125559
R28332 DVSS.n11298 DVSS.n8586 0.0125559
R28333 DVSS.n11258 DVSS.n11257 0.0125559
R28334 DVSS.n5755 DVSS.n5754 0.0125559
R28335 DVSS.n15864 DVSS.n15863 0.0125559
R28336 DVSS.n15854 DVSS.n7665 0.0125559
R28337 DVSS.n15711 DVSS.n15710 0.0125559
R28338 DVSS.n15720 DVSS.n15708 0.0125559
R28339 DVSS.n15618 DVSS.n15617 0.0125559
R28340 DVSS.n15608 DVSS.n7694 0.0125559
R28341 DVSS.n14981 DVSS.n14980 0.0125559
R28342 DVSS.n14991 DVSS.n14990 0.0125559
R28343 DVSS.n15694 DVSS.n15693 0.0125559
R28344 DVSS.n15011 DVSS.n15010 0.0125559
R28345 DVSS.n17607 DVSS.n17606 0.0125559
R28346 DVSS.n17034 DVSS.n17033 0.0125559
R28347 DVSS.n17566 DVSS.n17565 0.0125559
R28348 DVSS.n13025 DVSS.n11732 0.0125559
R28349 DVSS.n13085 DVSS.n11706 0.0125559
R28350 DVSS.n11541 DVSS.n11540 0.0125559
R28351 DVSS.n11405 DVSS.n11404 0.0125559
R28352 DVSS.n11363 DVSS.n8337 0.0125559
R28353 DVSS.n10860 DVSS.n10643 0.0125559
R28354 DVSS.n10820 DVSS.n10819 0.0125559
R28355 DVSS.n13140 DVSS.n13139 0.0125559
R28356 DVSS.n15035 DVSS.n15034 0.0125559
R28357 DVSS.n4043 DVSS.n4042 0.0125559
R28358 DVSS.n4033 DVSS.n2574 0.0125559
R28359 DVSS.n15044 DVSS.n14955 0.0125559
R28360 DVSS.n13150 DVSS.n13149 0.0125559
R28361 DVSS.n5235 DVSS.n5206 0.0125559
R28362 DVSS.n4343 DVSS.n4342 0.0125559
R28363 DVSS.n4352 DVSS.n4129 0.0125559
R28364 DVSS.n4127 DVSS.n4126 0.0125559
R28365 DVSS.n4117 DVSS.n2559 0.0125559
R28366 DVSS.n4001 DVSS.n4000 0.0125559
R28367 DVSS.n3765 DVSS.n3764 0.0125559
R28368 DVSS.n3969 DVSS.n3806 0.0125559
R28369 DVSS.n4274 DVSS.n4273 0.0125559
R28370 DVSS.n20246 DVSS.n20221 0.0125559
R28371 DVSS.n19236 DVSS.n19211 0.0125559
R28372 DVSS.n9798 DVSS.n9797 0.0125559
R28373 DVSS.n9717 DVSS.n9716 0.0125559
R28374 DVSS.n9606 DVSS.n9605 0.0125559
R28375 DVSS.n9105 DVSS.n9104 0.0125559
R28376 DVSS.n9041 DVSS.n9040 0.0125559
R28377 DVSS.n9691 DVSS.n9690 0.0125559
R28378 DVSS.n9075 DVSS.n9074 0.0125559
R28379 DVSS.n11130 DVSS.n11129 0.0125559
R28380 DVSS.n9923 DVSS.n9922 0.0125559
R28381 DVSS.n11089 DVSS.n11088 0.0125559
R28382 DVSS.n20737 DVSS.n20724 0.0125559
R28383 DVSS.n978 DVSS.n977 0.0125559
R28384 DVSS.n20740 DVSS.n20739 0.0125559
R28385 DVSS.n976 DVSS.n975 0.0125559
R28386 DVSS.n1182 DVSS.n1163 0.0125559
R28387 DVSS.n16287 DVSS.n16286 0.0125559
R28388 DVSS.n16248 DVSS.n16247 0.0125559
R28389 DVSS.n18376 DVSS.n7548 0.0125559
R28390 DVSS.n18389 DVSS.n18388 0.0125559
R28391 DVSS.n7499 DVSS.n7498 0.0125559
R28392 DVSS.n16412 DVSS.n16411 0.0125559
R28393 DVSS.n16206 DVSS.n16205 0.0125559
R28394 DVSS.n7531 DVSS.n7530 0.0125559
R28395 DVSS.n16376 DVSS.n16375 0.0125559
R28396 DVSS.n17332 DVSS.n17331 0.0125559
R28397 DVSS.n19507 DVSS.n19482 0.0125559
R28398 DVSS.n5408 DVSS.n5407 0.0125559
R28399 DVSS.n5445 DVSS.n5444 0.0125559
R28400 DVSS.n6327 DVSS.n6086 0.0125559
R28401 DVSS.n6588 DVSS.n6587 0.0125559
R28402 DVSS.n6817 DVSS.n6787 0.0125559
R28403 DVSS.n3626 DVSS.n3595 0.0125559
R28404 DVSS.n6050 DVSS.n5859 0.0125559
R28405 DVSS.n3660 DVSS.n3574 0.0125559
R28406 DVSS.n3730 DVSS.n3512 0.0125559
R28407 DVSS.n12091 DVSS.n12064 0.0125559
R28408 DVSS.n12907 DVSS.n12906 0.0125559
R28409 DVSS.n19019 DVSS.n18975 0.0125559
R28410 DVSS.n20316 DVSS.n20267 0.0125559
R28411 DVSS.n20590 DVSS.n20541 0.0125559
R28412 DVSS.n21555 DVSS.n76 0.0125559
R28413 DVSS.n19300 DVSS.n19256 0.0125559
R28414 DVSS.n19571 DVSS.n19527 0.0125559
R28415 DVSS.n1270 DVSS.n1162 0.0125559
R28416 DVSS.n21468 DVSS.n21467 0.0125559
R28417 DVSS.n1055 DVSS.n875 0.0125559
R28418 DVSS.n21087 DVSS.n21047 0.0125559
R28419 DVSS.n20861 DVSS.n20821 0.0125559
R28420 DVSS.n621 DVSS.n553 0.0125559
R28421 DVSS.n5713 DVSS.n4478 0.0125472
R28422 DVSS.n11217 DVSS.n11216 0.0125472
R28423 DVSS.n17652 DVSS.n17651 0.0125472
R28424 DVSS.n9834 DVSS.n9833 0.0125472
R28425 DVSS.n16325 DVSS.n16324 0.0125472
R28426 DVSS.n16544 DVSS.n16543 0.0125423
R28427 DVSS.n16567 DVSS.n16566 0.0125423
R28428 DVSS.n16111 DVSS.n16110 0.0125423
R28429 DVSS.n17761 DVSS.n17760 0.0125423
R28430 DVSS.n16731 DVSS.n16730 0.0125423
R28431 DVSS.n16754 DVSS.n16753 0.0125423
R28432 DVSS.n15992 DVSS.n15991 0.0125423
R28433 DVSS.n15902 DVSS.n15901 0.0125423
R28434 DVSS.n7167 DVSS.n7166 0.0124681
R28435 DVSS.n7184 DVSS.n7183 0.0124681
R28436 DVSS.n7302 DVSS.n7301 0.0124681
R28437 DVSS.n7871 DVSS.n7870 0.0124681
R28438 DVSS.n7881 DVSS.n7880 0.0124681
R28439 DVSS.n7959 DVSS.n7958 0.0124681
R28440 DVSS.n7036 DVSS.n7035 0.0124681
R28441 DVSS.n7077 DVSS.n7076 0.0124681
R28442 DVSS.n7063 DVSS.n7061 0.0124681
R28443 DVSS.n7050 DVSS.n7049 0.0124681
R28444 DVSS.n13608 DVSS.n13607 0.0124681
R28445 DVSS.n13628 DVSS.n13627 0.0124681
R28446 DVSS.n13300 DVSS.n13299 0.0124681
R28447 DVSS.n13316 DVSS.n13314 0.0124681
R28448 DVSS.n19173 DVSS.n19172 0.0124644
R28449 DVSS.n19264 DVSS.n19263 0.0124644
R28450 DVSS.n1019 DVSS.n1018 0.0124644
R28451 DVSS.n4310 DVSS.n4309 0.0124644
R28452 DVSS.n16170 DVSS.n16169 0.0124644
R28453 DVSS.n19444 DVSS.n19443 0.0124644
R28454 DVSS.n19535 DVSS.n19534 0.0124644
R28455 DVSS.n1234 DVSS.n1233 0.0124644
R28456 DVSS.n6624 DVSS.n6623 0.0124644
R28457 DVSS.n18983 DVSS.n18982 0.0124644
R28458 DVSS.n585 DVSS.n584 0.0124644
R28459 DVSS.n16597 DVSS.n16596 0.012425
R28460 DVSS.n16606 DVSS.n16605 0.012425
R28461 DVSS.n18310 DVSS.n18309 0.012425
R28462 DVSS.n18319 DVSS.n18318 0.012425
R28463 DVSS.n19220 DVSS.n19217 0.0124231
R28464 DVSS.n19223 DVSS.n19220 0.0124231
R28465 DVSS.n19226 DVSS.n19223 0.0124231
R28466 DVSS.n19235 DVSS.n19226 0.0124231
R28467 DVSS.n19235 DVSS.n19234 0.0124231
R28468 DVSS.n19234 DVSS.n19231 0.0124231
R28469 DVSS.n19506 DVSS.n19505 0.0124231
R28470 DVSS.n19505 DVSS.n19502 0.0124231
R28471 DVSS.n19502 DVSS.n19499 0.0124231
R28472 DVSS.n19499 DVSS.n19496 0.0124231
R28473 DVSS.n19496 DVSS.n19495 0.0124231
R28474 DVSS.n19495 DVSS.n19492 0.0124231
R28475 DVSS.n19741 DVSS.n19738 0.0124231
R28476 DVSS.n19738 DVSS.n19735 0.0124231
R28477 DVSS.n19735 DVSS.n19734 0.0124231
R28478 DVSS.n19966 DVSS.n19963 0.0124231
R28479 DVSS.n19963 DVSS.n19960 0.0124231
R28480 DVSS.n19960 DVSS.n19959 0.0124231
R28481 DVSS.n19959 DVSS.n19956 0.0124231
R28482 DVSS.n20230 DVSS.n20227 0.0124231
R28483 DVSS.n20233 DVSS.n20230 0.0124231
R28484 DVSS.n20236 DVSS.n20233 0.0124231
R28485 DVSS.n20245 DVSS.n20236 0.0124231
R28486 DVSS.n20245 DVSS.n20244 0.0124231
R28487 DVSS.n20244 DVSS.n20241 0.0124231
R28488 DVSS.n20519 DVSS.n20516 0.0124231
R28489 DVSS.n20516 DVSS.n20513 0.0124231
R28490 DVSS.n20513 DVSS.n20510 0.0124231
R28491 DVSS.n20510 DVSS.n20507 0.0124231
R28492 DVSS.n20507 DVSS.n20506 0.0124231
R28493 DVSS.n20506 DVSS.n20503 0.0124231
R28494 DVSS.n958 DVSS.n955 0.0124231
R28495 DVSS.n961 DVSS.n958 0.0124231
R28496 DVSS.n964 DVSS.n961 0.0124231
R28497 DVSS.n973 DVSS.n964 0.0124231
R28498 DVSS.n973 DVSS.n970 0.0124231
R28499 DVSS.n970 DVSS.n967 0.0124231
R28500 DVSS.n1192 DVSS.n1189 0.0124231
R28501 DVSS.n1181 DVSS.n1178 0.0124231
R28502 DVSS.n1178 DVSS.n1175 0.0124231
R28503 DVSS.n1175 DVSS.n1172 0.0124231
R28504 DVSS.n1172 DVSS.n1169 0.0124231
R28505 DVSS.n332 DVSS.n329 0.0124231
R28506 DVSS.n335 DVSS.n332 0.0124231
R28507 DVSS.n338 DVSS.n335 0.0124231
R28508 DVSS.n341 DVSS.n338 0.0124231
R28509 DVSS.n365 DVSS.n362 0.0124231
R28510 DVSS.n368 DVSS.n365 0.0124231
R28511 DVSS.n371 DVSS.n368 0.0124231
R28512 DVSS.n374 DVSS.n371 0.0124231
R28513 DVSS.n20733 DVSS.n20730 0.0124231
R28514 DVSS.n20736 DVSS.n20733 0.0124231
R28515 DVSS.n20723 DVSS.n20711 0.0124231
R28516 DVSS.n20723 DVSS.n20720 0.0124231
R28517 DVSS.n20720 DVSS.n20717 0.0124231
R28518 DVSS.n20961 DVSS.n20958 0.0124231
R28519 DVSS.n20964 DVSS.n20961 0.0124231
R28520 DVSS.n20952 DVSS.n20940 0.0124231
R28521 DVSS.n20952 DVSS.n20949 0.0124231
R28522 DVSS.n20949 DVSS.n20946 0.0124231
R28523 DVSS.n5744 DVSS.n5743 0.0123701
R28524 DVSS.n11247 DVSS.n11246 0.0123701
R28525 DVSS.n17618 DVSS.n17617 0.0123701
R28526 DVSS.n11141 DVSS.n11140 0.0123701
R28527 DVSS.n16365 DVSS.n16364 0.0123701
R28528 DVSS.n16664 DVSS.n16663 0.012331
R28529 DVSS.n16117 DVSS.n16116 0.012331
R28530 DVSS.n17752 DVSS.n17751 0.012331
R28531 DVSS.n18113 DVSS.n18112 0.012331
R28532 DVSS.n17159 DVSS.n17158 0.012331
R28533 DVSS.n15998 DVSS.n15997 0.012331
R28534 DVSS.n15911 DVSS.n15910 0.012331
R28535 DVSS.n15403 DVSS.n15402 0.012331
R28536 DVSS.n6513 DVSS.n6512 0.0123034
R28537 DVSS.n19237 DVSS.n19236 0.0123034
R28538 DVSS.n19300 DVSS.n19299 0.0123034
R28539 DVSS.n4084 DVSS.n4083 0.0123034
R28540 DVSS.n4388 DVSS.n4387 0.0123034
R28541 DVSS.n6525 DVSS.n6524 0.0123034
R28542 DVSS.n6522 DVSS.n6521 0.0123034
R28543 DVSS.n11298 DVSS.n11297 0.0123034
R28544 DVSS.n12906 DVSS.n12905 0.0123034
R28545 DVSS.n12966 DVSS.n12965 0.0123034
R28546 DVSS.n9140 DVSS.n9139 0.0123034
R28547 DVSS.n9150 DVSS.n9149 0.0123034
R28548 DVSS.n9588 DVSS.n9587 0.0123034
R28549 DVSS.n9578 DVSS.n9577 0.0123034
R28550 DVSS.n9752 DVSS.n9751 0.0123034
R28551 DVSS.n9762 DVSS.n9761 0.0123034
R28552 DVSS.n9780 DVSS.n9779 0.0123034
R28553 DVSS.n9770 DVSS.n9769 0.0123034
R28554 DVSS.n9502 DVSS.n9501 0.0123034
R28555 DVSS.n13116 DVSS.n13115 0.0123034
R28556 DVSS.n10902 DVSS.n10901 0.0123034
R28557 DVSS.n5754 DVSS.n5753 0.0123034
R28558 DVSS.n11257 DVSS.n11256 0.0123034
R28559 DVSS.n17567 DVSS.n17566 0.0123034
R28560 DVSS.n15695 DVSS.n15694 0.0123034
R28561 DVSS.n15720 DVSS.n15719 0.0123034
R28562 DVSS.n15710 DVSS.n15709 0.0123034
R28563 DVSS.n15855 DVSS.n15854 0.0123034
R28564 DVSS.n15865 DVSS.n15864 0.0123034
R28565 DVSS.n15010 DVSS.n15009 0.0123034
R28566 DVSS.n14990 DVSS.n14989 0.0123034
R28567 DVSS.n14980 DVSS.n14979 0.0123034
R28568 DVSS.n15609 DVSS.n15608 0.0123034
R28569 DVSS.n15619 DVSS.n15618 0.0123034
R28570 DVSS.n17035 DVSS.n17034 0.0123034
R28571 DVSS.n17608 DVSS.n17607 0.0123034
R28572 DVSS.n11364 DVSS.n11363 0.0123034
R28573 DVSS.n12091 DVSS.n12090 0.0123034
R28574 DVSS.n21555 DVSS.n21554 0.0123034
R28575 DVSS.n13026 DVSS.n13025 0.0123034
R28576 DVSS.n11540 DVSS.n11539 0.0123034
R28577 DVSS.n13085 DVSS.n13084 0.0123034
R28578 DVSS.n11404 DVSS.n11403 0.0123034
R28579 DVSS.n10819 DVSS.n10818 0.0123034
R28580 DVSS.n10860 DVSS.n10859 0.0123034
R28581 DVSS.n13149 DVSS.n13148 0.0123034
R28582 DVSS.n13139 DVSS.n13138 0.0123034
R28583 DVSS.n4034 DVSS.n4033 0.0123034
R28584 DVSS.n4044 DVSS.n4043 0.0123034
R28585 DVSS.n15044 DVSS.n15043 0.0123034
R28586 DVSS.n15034 DVSS.n15033 0.0123034
R28587 DVSS.n5235 DVSS.n5234 0.0123034
R28588 DVSS.n4118 DVSS.n4117 0.0123034
R28589 DVSS.n4128 DVSS.n4127 0.0123034
R28590 DVSS.n4352 DVSS.n4351 0.0123034
R28591 DVSS.n4342 DVSS.n4341 0.0123034
R28592 DVSS.n4273 DVSS.n4272 0.0123034
R28593 DVSS.n3970 DVSS.n3969 0.0123034
R28594 DVSS.n4001 DVSS.n3790 0.0123034
R28595 DVSS.n3764 DVSS.n3763 0.0123034
R28596 DVSS.n20247 DVSS.n20246 0.0123034
R28597 DVSS.n11090 DVSS.n11089 0.0123034
R28598 DVSS.n9074 DVSS.n9073 0.0123034
R28599 DVSS.n9797 DVSS.n8928 0.0123034
R28600 DVSS.n9717 DVSS.n9705 0.0123034
R28601 DVSS.n9605 DVSS.n8961 0.0123034
R28602 DVSS.n9105 DVSS.n9093 0.0123034
R28603 DVSS.n9040 DVSS.n9011 0.0123034
R28604 DVSS.n9692 DVSS.n9691 0.0123034
R28605 DVSS.n9924 DVSS.n9923 0.0123034
R28606 DVSS.n11131 DVSS.n11130 0.0123034
R28607 DVSS.n20739 DVSS.n20738 0.0123034
R28608 DVSS.n20738 DVSS.n20737 0.0123034
R28609 DVSS.n977 DVSS.n976 0.0123034
R28610 DVSS.n975 DVSS.n974 0.0123034
R28611 DVSS.n7530 DVSS.n7529 0.0123034
R28612 DVSS.n19571 DVSS.n19570 0.0123034
R28613 DVSS.n16286 DVSS.n16259 0.0123034
R28614 DVSS.n16247 DVSS.n16220 0.0123034
R28615 DVSS.n16207 DVSS.n16206 0.0123034
R28616 DVSS.n18377 DVSS.n18376 0.0123034
R28617 DVSS.n18389 DVSS.n7547 0.0123034
R28618 DVSS.n7498 DVSS.n7469 0.0123034
R28619 DVSS.n16413 DVSS.n16412 0.0123034
R28620 DVSS.n17331 DVSS.n17330 0.0123034
R28621 DVSS.n16375 DVSS.n16374 0.0123034
R28622 DVSS.n19508 DVSS.n19507 0.0123034
R28623 DVSS.n1183 DVSS.n1182 0.0123034
R28624 DVSS.n6051 DVSS.n6050 0.0123034
R28625 DVSS.n6818 DVSS.n6817 0.0123034
R28626 DVSS.n621 DVSS.n620 0.0123034
R28627 DVSS.n5407 DVSS.n5406 0.0123034
R28628 DVSS.n6587 DVSS.n6586 0.0123034
R28629 DVSS.n5444 DVSS.n5443 0.0123034
R28630 DVSS.n3627 DVSS.n3626 0.0123034
R28631 DVSS.n6328 DVSS.n6327 0.0123034
R28632 DVSS.n3660 DVSS.n3659 0.0123034
R28633 DVSS.n3731 DVSS.n3730 0.0123034
R28634 DVSS.n20590 DVSS.n20589 0.0123034
R28635 DVSS.n20316 DVSS.n20315 0.0123034
R28636 DVSS.n19019 DVSS.n19018 0.0123034
R28637 DVSS.n21467 DVSS.n21466 0.0123034
R28638 DVSS.n1270 DVSS.n1269 0.0123034
R28639 DVSS.n1055 DVSS.n1054 0.0123034
R28640 DVSS.n21087 DVSS.n21086 0.0123034
R28641 DVSS.n20861 DVSS.n20860 0.0123034
R28642 DVSS.n2020 DVSS.n2019 0.0122524
R28643 DVSS.n7721 DVSS.n7720 0.0122
R28644 DVSS.n16052 DVSS.n16051 0.0122
R28645 DVSS.n19688 DVSS.n19687 0.0120643
R28646 DVSS.n19772 DVSS.n19771 0.0120643
R28647 DVSS.n213 DVSS.n212 0.0120643
R28648 DVSS.n19907 DVSS.n19906 0.0120643
R28649 DVSS.n19997 DVSS.n19996 0.0120643
R28650 DVSS.n421 DVSS.n420 0.0120643
R28651 DVSS.n19689 DVSS.n19688 0.0120643
R28652 DVSS.n19908 DVSS.n19907 0.0120643
R28653 DVSS.n19771 DVSS.n19770 0.0120643
R28654 DVSS.n19996 DVSS.n19995 0.0120643
R28655 DVSS.n212 DVSS.n211 0.0120643
R28656 DVSS.n420 DVSS.n419 0.0120643
R28657 DVSS.n15427 DVSS.n15426 0.011975
R28658 DVSS.n18285 DVSS.n18284 0.011975
R28659 DVSS.n18334 DVSS.n18333 0.011975
R28660 DVSS.n18341 DVSS.n18340 0.011975
R28661 DVSS.n5612 DVSS.n5611 0.0119309
R28662 DVSS.n5791 DVSS.n5790 0.0119309
R28663 DVSS.n6535 DVSS.n4470 0.0119309
R28664 DVSS.n4457 DVSS.n4456 0.0119309
R28665 DVSS.n4377 DVSS.n2546 0.0119309
R28666 DVSS.n4094 DVSS.n4082 0.0119309
R28667 DVSS.n4066 DVSS.n4065 0.0119309
R28668 DVSS.n6535 DVSS.n6534 0.0119309
R28669 DVSS.n4378 DVSS.n4377 0.0119309
R28670 DVSS.n4094 DVSS.n4093 0.0119309
R28671 DVSS.n5792 DVSS.n5791 0.0119309
R28672 DVSS.n4065 DVSS.n4064 0.0119309
R28673 DVSS.n4456 DVSS.n4455 0.0119309
R28674 DVSS.n5613 DVSS.n5612 0.0119309
R28675 DVSS.n20521 DVSS.n20520 0.0119309
R28676 DVSS.n20520 DVSS.n20492 0.0119309
R28677 DVSS.n1193 DVSS.n1183 0.0119309
R28678 DVSS.n1194 DVSS.n1193 0.0119309
R28679 DVSS.n18430 DVSS.n18429 0.0119085
R28680 DVSS.n15199 DVSS.n15198 0.0119085
R28681 DVSS.n4520 DVSS.n4519 0.0117632
R28682 DVSS.n17217 DVSS.n17216 0.01175
R28683 DVSS.n17227 DVSS.n17226 0.01175
R28684 DVSS.n15185 DVSS.n15184 0.01175
R28685 DVSS.n15146 DVSS.n15145 0.01175
R28686 DVSS.n17695 DVSS.n17694 0.01175
R28687 DVSS.n16556 DVSS.n16555 0.0116972
R28688 DVSS.n18275 DVSS.n18158 0.0116972
R28689 DVSS.n18232 DVSS.n18231 0.0116972
R28690 DVSS.n19718 DVSS.n19717 0.0116972
R28691 DVSS.n16743 DVSS.n16742 0.0116972
R28692 DVSS.n15464 DVSS.n15463 0.0116972
R28693 DVSS.n15508 DVSS.n15507 0.0116972
R28694 DVSS.n19937 DVSS.n19936 0.0116972
R28695 DVSS.n11023 DVSS.n11022 0.0116937
R28696 DVSS.n11193 DVSS.n11192 0.0116937
R28697 DVSS.n10033 DVSS.n10032 0.0116937
R28698 DVSS.n17879 DVSS.n17878 0.0115386
R28699 DVSS.n18020 DVSS.n18019 0.0115386
R28700 DVSS.n18166 DVSS.n18165 0.0115386
R28701 DVSS.n7571 DVSS.n7570 0.0115386
R28702 DVSS.n18517 DVSS.n18516 0.0115386
R28703 DVSS.n17880 DVSS.n17879 0.0115386
R28704 DVSS.n18021 DVSS.n18020 0.0115386
R28705 DVSS.n18167 DVSS.n18166 0.0115386
R28706 DVSS.n7572 DVSS.n7571 0.0115386
R28707 DVSS.n15820 DVSS.n15819 0.0115386
R28708 DVSS.n15742 DVSS.n15741 0.0115386
R28709 DVSS.n15574 DVSS.n15573 0.0115386
R28710 DVSS.n15238 DVSS.n15237 0.0115386
R28711 DVSS.n7758 DVSS.n7757 0.0115386
R28712 DVSS.n15743 DVSS.n15742 0.0115386
R28713 DVSS.n15819 DVSS.n15818 0.0115386
R28714 DVSS.n15237 DVSS.n15236 0.0115386
R28715 DVSS.n15573 DVSS.n15572 0.0115386
R28716 DVSS.n18516 DVSS.n18515 0.0115386
R28717 DVSS.n7757 DVSS.n7756 0.0115386
R28718 DVSS.n15396 DVSS.n15395 0.011525
R28719 DVSS.n18298 DVSS.n18294 0.011525
R28720 DVSS.n18303 DVSS.n18302 0.011525
R28721 DVSS.n16692 DVSS.n16691 0.0114859
R28722 DVSS.n16074 DVSS.n16073 0.0114859
R28723 DVSS.n18275 DVSS.n18274 0.0114859
R28724 DVSS.n17131 DVSS.n17130 0.0114859
R28725 DVSS.n15966 DVSS.n15965 0.0114859
R28726 DVSS.n15465 DVSS.n15464 0.0114859
R28727 DVSS.n5561 DVSS.n5560 0.0114843
R28728 DVSS.n6993 DVSS.n6992 0.0114843
R28729 DVSS.n19146 DVSS.n19145 0.0114843
R28730 DVSS.n10202 DVSS.n10201 0.0114843
R28731 DVSS.n12763 DVSS.n12762 0.0114843
R28732 DVSS.n12754 DVSS.n12753 0.0114843
R28733 DVSS.n12748 DVSS.n12747 0.0114843
R28734 DVSS.n12733 DVSS.n12732 0.0114843
R28735 DVSS.n12724 DVSS.n12723 0.0114843
R28736 DVSS.n12687 DVSS.n12686 0.0114843
R28737 DVSS.n12678 DVSS.n12677 0.0114843
R28738 DVSS.n12497 DVSS.n12496 0.0114843
R28739 DVSS.n12488 DVSS.n12487 0.0114843
R28740 DVSS.n12479 DVSS.n12478 0.0114843
R28741 DVSS.n12453 DVSS.n12452 0.0114843
R28742 DVSS.n12444 DVSS.n12443 0.0114843
R28743 DVSS.n12430 DVSS.n12429 0.0114843
R28744 DVSS.n12421 DVSS.n12420 0.0114843
R28745 DVSS.n12213 DVSS.n12212 0.0114843
R28746 DVSS.n12206 DVSS.n12205 0.0114843
R28747 DVSS.n12177 DVSS.n12176 0.0114843
R28748 DVSS.n12170 DVSS.n12169 0.0114843
R28749 DVSS.n12154 DVSS.n12153 0.0114843
R28750 DVSS.n21289 DVSS.n21288 0.0114843
R28751 DVSS.n21280 DVSS.n21279 0.0114843
R28752 DVSS.n16947 DVSS.n16946 0.0114843
R28753 DVSS.n13645 DVSS.n13644 0.0114843
R28754 DVSS.n20157 DVSS.n20156 0.0114843
R28755 DVSS.n10606 DVSS.n10605 0.0114843
R28756 DVSS.n10744 DVSS.n10743 0.0114843
R28757 DVSS.n11416 DVSS.n11415 0.0114843
R28758 DVSS.n5214 DVSS.n5213 0.0114843
R28759 DVSS.n3375 DVSS.n3374 0.0114843
R28760 DVSS.n3367 DVSS.n3366 0.0114843
R28761 DVSS.n3361 DVSS.n3360 0.0114843
R28762 DVSS.n3355 DVSS.n3354 0.0114843
R28763 DVSS.n3347 DVSS.n3346 0.0114843
R28764 DVSS.n3310 DVSS.n3309 0.0114843
R28765 DVSS.n3302 DVSS.n3301 0.0114843
R28766 DVSS.n3121 DVSS.n3120 0.0114843
R28767 DVSS.n3113 DVSS.n3112 0.0114843
R28768 DVSS.n3105 DVSS.n3104 0.0114843
R28769 DVSS.n3079 DVSS.n3078 0.0114843
R28770 DVSS.n3071 DVSS.n3070 0.0114843
R28771 DVSS.n3056 DVSS.n3055 0.0114843
R28772 DVSS.n3048 DVSS.n3047 0.0114843
R28773 DVSS.n2843 DVSS.n2842 0.0114843
R28774 DVSS.n2836 DVSS.n2835 0.0114843
R28775 DVSS.n2805 DVSS.n2804 0.0114843
R28776 DVSS.n2798 DVSS.n2797 0.0114843
R28777 DVSS.n739 DVSS.n738 0.0114843
R28778 DVSS.n657 DVSS.n656 0.0114843
R28779 DVSS.n9903 DVSS.n9902 0.0114843
R28780 DVSS.n13230 DVSS.n13229 0.0114843
R28781 DVSS.n20428 DVSS.n20427 0.0114843
R28782 DVSS.n17256 DVSS.n17255 0.0114843
R28783 DVSS.n18760 DVSS.n18759 0.0114843
R28784 DVSS.n19420 DVSS.n19419 0.0114843
R28785 DVSS.n5319 DVSS.n5318 0.0114843
R28786 DVSS.n5850 DVSS.n5849 0.0114843
R28787 DVSS.n6338 DVSS.n6337 0.0114843
R28788 DVSS.n14915 DVSS.n14888 0.0113101
R28789 DVSS.n14915 DVSS.n14914 0.0113101
R28790 DVSS.n5670 DVSS.n5669 0.0113071
R28791 DVSS.n10962 DVSS.n10961 0.0113071
R28792 DVSS.n12818 DVSS.n12817 0.0113071
R28793 DVSS.n12696 DVSS.n12695 0.0113071
R28794 DVSS.n12436 DVSS.n12435 0.0113071
R28795 DVSS.n12161 DVSS.n12160 0.0113071
R28796 DVSS.n17095 DVSS.n17094 0.0113071
R28797 DVSS.n11449 DVSS.n11448 0.0113071
R28798 DVSS.n4679 DVSS.n4678 0.0113071
R28799 DVSS.n3430 DVSS.n3429 0.0113071
R28800 DVSS.n3319 DVSS.n3318 0.0113071
R28801 DVSS.n3062 DVSS.n3061 0.0113071
R28802 DVSS.n2789 DVSS.n2788 0.0113071
R28803 DVSS.n9984 DVSS.n9983 0.0113071
R28804 DVSS.n17389 DVSS.n17388 0.0113071
R28805 DVSS.n6450 DVSS.n6449 0.0113071
R28806 DVSS.n17212 DVSS.n17211 0.0113
R28807 DVSS.n15151 DVSS.n15150 0.0113
R28808 DVSS.n15109 DVSS.n15108 0.0113
R28809 DVSS.n2410 DVSS.n2409 0.0113
R28810 DVSS.n17690 DVSS.n17689 0.0113
R28811 DVSS.n16512 DVSS.n16511 0.0112746
R28812 DVSS.n16858 DVSS.n16857 0.0112746
R28813 DVSS.n19753 DVSS.n19752 0.0112232
R28814 DVSS.n19979 DVSS.n19978 0.0112232
R28815 DVSS.n19978 DVSS.n19977 0.0112232
R28816 DVSS.n19754 DVSS.n19753 0.0112232
R28817 DVSS.n14953 DVSS.n13850 0.0111514
R28818 DVSS.n13152 DVSS.n8049 0.0111514
R28819 DVSS.n13051 DVSS.n13050 0.0111514
R28820 DVSS.n11687 DVSS.n11686 0.0111514
R28821 DVSS.n11653 DVSS.n11652 0.0111514
R28822 DVSS.n11650 DVSS.n11649 0.0111514
R28823 DVSS.n11616 DVSS.n11615 0.0111514
R28824 DVSS.n11525 DVSS.n11524 0.0111514
R28825 DVSS.n11491 DVSS.n11490 0.0111514
R28826 DVSS.n11488 DVSS.n11487 0.0111514
R28827 DVSS.n11454 DVSS.n11453 0.0111514
R28828 DVSS.n13062 DVSS.n13061 0.0111514
R28829 DVSS.n690 DVSS.n689 0.0111514
R28830 DVSS.n3441 DVSS.n3440 0.0111514
R28831 DVSS.n13180 DVSS.n8006 0.0111514
R28832 DVSS.n21140 DVSS.n21139 0.0111514
R28833 DVSS.n694 DVSS.n693 0.0111514
R28834 DVSS.n692 DVSS.n691 0.0111514
R28835 DVSS.n18572 DVSS.n7431 0.0111514
R28836 DVSS.n6952 DVSS.n6951 0.0111514
R28837 DVSS.n19249 DVSS.n19248 0.0111389
R28838 DVSS.n19520 DVSS.n19519 0.0111389
R28839 DVSS.n15432 DVSS.n15431 0.011075
R28840 DVSS.n18280 DVSS.n18279 0.011075
R28841 DVSS.n18329 DVSS.n18328 0.011075
R28842 DVSS.n18346 DVSS.n18345 0.011075
R28843 DVSS.n17475 DVSS.n17474 0.0110634
R28844 DVSS.n16816 DVSS.n16815 0.0110634
R28845 DVSS.n12469 DVSS.n12468 0.0109528
R28846 DVSS.n12411 DVSS.n12410 0.0109528
R28847 DVSS.n12191 DVSS.n12190 0.0109528
R28848 DVSS.n21142 DVSS.n21141 0.0109528
R28849 DVSS.n10787 DVSS.n10786 0.0109528
R28850 DVSS.n3095 DVSS.n3094 0.0109528
R28851 DVSS.n3038 DVSS.n3037 0.0109528
R28852 DVSS.n2820 DVSS.n2819 0.0109528
R28853 DVSS.n695 DVSS.n694 0.0109528
R28854 DVSS.n5477 DVSS.n5476 0.0109528
R28855 DVSS.n14954 DVSS.n14953 0.0108992
R28856 DVSS.n13152 DVSS.n13151 0.0108992
R28857 DVSS.n11455 DVSS.n11454 0.0108992
R28858 DVSS.n11489 DVSS.n11488 0.0108992
R28859 DVSS.n11492 DVSS.n11491 0.0108992
R28860 DVSS.n11526 DVSS.n11525 0.0108992
R28861 DVSS.n11617 DVSS.n11616 0.0108992
R28862 DVSS.n11651 DVSS.n11650 0.0108992
R28863 DVSS.n11654 DVSS.n11653 0.0108992
R28864 DVSS.n11688 DVSS.n11687 0.0108992
R28865 DVSS.n13050 DVSS.n13049 0.0108992
R28866 DVSS.n13061 DVSS.n13060 0.0108992
R28867 DVSS.n3440 DVSS.n3439 0.0108992
R28868 DVSS.n693 DVSS.n692 0.0108992
R28869 DVSS.n13181 DVSS.n13180 0.0108992
R28870 DVSS.n21141 DVSS.n21140 0.0108992
R28871 DVSS.n691 DVSS.n690 0.0108992
R28872 DVSS.n689 DVSS.n688 0.0108992
R28873 DVSS.n18573 DVSS.n18572 0.0108992
R28874 DVSS.n6951 DVSS.n1347 0.0108992
R28875 DVSS.n12816 DVSS.n12801 0.0108846
R28876 DVSS.n12523 DVSS.n12518 0.0108846
R28877 DVSS.n12524 DVSS.n12523 0.0108846
R28878 DVSS.n12673 DVSS.n12548 0.0108846
R28879 DVSS.n12673 DVSS.n12672 0.0108846
R28880 DVSS.n12648 DVSS.n12647 0.0108846
R28881 DVSS.n12647 DVSS.n12642 0.0108846
R28882 DVSS.n12586 DVSS.n12585 0.0108846
R28883 DVSS.n12585 DVSS.n12580 0.0108846
R28884 DVSS.n12564 DVSS.n12563 0.0108846
R28885 DVSS.n12563 DVSS.n12558 0.0108846
R28886 DVSS.n12558 DVSS.n12557 0.0108846
R28887 DVSS.n12385 DVSS.n12215 0.0108846
R28888 DVSS.n12385 DVSS.n12384 0.0108846
R28889 DVSS.n12360 DVSS.n12359 0.0108846
R28890 DVSS.n12359 DVSS.n12354 0.0108846
R28891 DVSS.n12298 DVSS.n12297 0.0108846
R28892 DVSS.n12297 DVSS.n12292 0.0108846
R28893 DVSS.n12244 DVSS.n12243 0.0108846
R28894 DVSS.n12243 DVSS.n12238 0.0108846
R28895 DVSS.n3428 DVSS.n3413 0.0108846
R28896 DVSS.n3147 DVSS.n3142 0.0108846
R28897 DVSS.n3148 DVSS.n3147 0.0108846
R28898 DVSS.n3297 DVSS.n3172 0.0108846
R28899 DVSS.n3297 DVSS.n3296 0.0108846
R28900 DVSS.n3272 DVSS.n3271 0.0108846
R28901 DVSS.n3271 DVSS.n3266 0.0108846
R28902 DVSS.n3210 DVSS.n3209 0.0108846
R28903 DVSS.n3209 DVSS.n3204 0.0108846
R28904 DVSS.n3188 DVSS.n3187 0.0108846
R28905 DVSS.n3187 DVSS.n3182 0.0108846
R28906 DVSS.n3182 DVSS.n3181 0.0108846
R28907 DVSS.n3012 DVSS.n2845 0.0108846
R28908 DVSS.n3012 DVSS.n3011 0.0108846
R28909 DVSS.n2987 DVSS.n2986 0.0108846
R28910 DVSS.n2986 DVSS.n2981 0.0108846
R28911 DVSS.n2925 DVSS.n2924 0.0108846
R28912 DVSS.n2924 DVSS.n2919 0.0108846
R28913 DVSS.n2871 DVSS.n2870 0.0108846
R28914 DVSS.n2870 DVSS.n2865 0.0108846
R28915 DVSS.n16656 DVSS.n16655 0.0108521
R28916 DVSS.n16665 DVSS.n16664 0.0108521
R28917 DVSS.n16116 DVSS.n16115 0.0108521
R28918 DVSS.n17753 DVSS.n17752 0.0108521
R28919 DVSS.n17789 DVSS.n17788 0.0108521
R28920 DVSS.n18112 DVSS.n18111 0.0108521
R28921 DVSS.n17167 DVSS.n17166 0.0108521
R28922 DVSS.n17158 DVSS.n17157 0.0108521
R28923 DVSS.n15997 DVSS.n15996 0.0108521
R28924 DVSS.n15910 DVSS.n15909 0.0108521
R28925 DVSS.n15874 DVSS.n7655 0.0108521
R28926 DVSS.n15402 DVSS.n15389 0.0108521
R28927 DVSS.n7716 DVSS.n7715 0.01085
R28928 DVSS.n16047 DVSS.n16046 0.01085
R28929 DVSS.n4417 DVSS.n4416 0.0107895
R28930 DVSS.n19176 DVSS.n19175 0.0107895
R28931 DVSS.n19261 DVSS.n19260 0.0107895
R28932 DVSS.n1016 DVSS.n1015 0.0107895
R28933 DVSS.n4313 DVSS.n4312 0.0107895
R28934 DVSS.n3474 DVSS.n3473 0.0107895
R28935 DVSS.n19447 DVSS.n19446 0.0107895
R28936 DVSS.n19532 DVSS.n19531 0.0107895
R28937 DVSS.n1231 DVSS.n1230 0.0107895
R28938 DVSS.n3536 DVSS.n3535 0.0107895
R28939 DVSS.n18980 DVSS.n18979 0.0107895
R28940 DVSS.n582 DVSS.n581 0.0107895
R28941 DVSS.n6769 DVSS.n6767 0.0107778
R28942 DVSS.n11660 DVSS.n11657 0.0107778
R28943 DVSS.n6714 DVSS.n6712 0.0107778
R28944 DVSS.n11623 DVSS.n11620 0.0107778
R28945 DVSS.n6571 DVSS.n6569 0.0107778
R28946 DVSS.n11498 DVSS.n11495 0.0107778
R28947 DVSS.n6435 DVSS.n6433 0.0107778
R28948 DVSS.n11461 DVSS.n11458 0.0107778
R28949 DVSS.n6896 DVSS.n6894 0.0107778
R28950 DVSS.n11709 DVSS.n11707 0.0107778
R28951 DVSS.n7180 DVSS.n7179 0.0107756
R28952 DVSS.n12715 DVSS.n12714 0.0107756
R28953 DVSS.n13527 DVSS.n13526 0.0107756
R28954 DVSS.n10807 DVSS.n10806 0.0107756
R28955 DVSS.n3338 DVSS.n3337 0.0107756
R28956 DVSS.n13390 DVSS.n13389 0.0107756
R28957 DVSS.n18848 DVSS.n18847 0.0107756
R28958 DVSS.n5456 DVSS.n5455 0.0107756
R28959 DVSS.n4444 DVSS.n4443 0.010701
R28960 DVSS.n4392 DVSS.n4391 0.010701
R28961 DVSS.n19288 DVSS.n19287 0.010701
R28962 DVSS.n1043 DVSS.n1042 0.010701
R28963 DVSS.n4286 DVSS.n4285 0.010701
R28964 DVSS.n4338 DVSS.n4337 0.010701
R28965 DVSS.n3501 DVSS.n3500 0.010701
R28966 DVSS.n16194 DVSS.n16193 0.010701
R28967 DVSS.n19559 DVSS.n19558 0.010701
R28968 DVSS.n1258 DVSS.n1257 0.010701
R28969 DVSS.n16141 DVSS.n16140 0.010701
R28970 DVSS.n6600 DVSS.n6599 0.010701
R28971 DVSS.n3563 DVSS.n3562 0.010701
R28972 DVSS.n19007 DVSS.n19006 0.010701
R28973 DVSS.n609 DVSS.n608 0.010701
R28974 DVSS.n6653 DVSS.n6652 0.010701
R28975 DVSS.n18960 DVSS.n18959 0.010701
R28976 DVSS.n1147 DVSS.n1146 0.010701
R28977 DVSS.n860 DVSS.n859 0.010701
R28978 DVSS.n538 DVSS.n537 0.010701
R28979 DVSS.n557 DVSS.n556 0.010701
R28980 DVSS.n12766 DVSS.n12765 0.0106923
R28981 DVSS.n12611 DVSS.n12610 0.0106923
R28982 DVSS.n12594 DVSS.n12593 0.0106923
R28983 DVSS.n12323 DVSS.n12322 0.0106923
R28984 DVSS.n12306 DVSS.n12305 0.0106923
R28985 DVSS.n12231 DVSS.n12230 0.0106923
R28986 DVSS.n21341 DVSS.n21331 0.0106923
R28987 DVSS.n3378 DVSS.n3377 0.0106923
R28988 DVSS.n3235 DVSS.n3234 0.0106923
R28989 DVSS.n3218 DVSS.n3217 0.0106923
R28990 DVSS.n2950 DVSS.n2949 0.0106923
R28991 DVSS.n2933 DVSS.n2932 0.0106923
R28992 DVSS.n2858 DVSS.n2857 0.0106923
R28993 DVSS.n885 DVSS.n884 0.0106923
R28994 DVSS.n21172 DVSS.n21171 0.0106727
R28995 DVSS.n16545 DVSS.n16544 0.0106408
R28996 DVSS.n18225 DVSS.n18224 0.0106408
R28997 DVSS.n18182 DVSS.n18181 0.0106408
R28998 DVSS.n16732 DVSS.n16731 0.0106408
R28999 DVSS.n15515 DVSS.n15514 0.0106408
R29000 DVSS.n15558 DVSS.n15557 0.0106408
R29001 DVSS.n16601 DVSS.n16600 0.010625
R29002 DVSS.n16602 DVSS.n16601 0.010625
R29003 DVSS.n18314 DVSS.n18313 0.010625
R29004 DVSS.n18315 DVSS.n18314 0.010625
R29005 DVSS.n5636 DVSS.n5635 0.0106125
R29006 DVSS.n5767 DVSS.n5766 0.0106125
R29007 DVSS.n6974 DVSS.n6973 0.0106125
R29008 DVSS.n4078 DVSS.n4077 0.0106125
R29009 DVSS.n4706 DVSS.n4705 0.0106125
R29010 DVSS.n3795 DVSS.n3794 0.0106125
R29011 DVSS.n3777 DVSS.n3776 0.0106125
R29012 DVSS.n17355 DVSS.n17354 0.0106125
R29013 DVSS.n16388 DVSS.n16387 0.0106125
R29014 DVSS.n7543 DVSS.n7542 0.0106125
R29015 DVSS.n18741 DVSS.n18740 0.0106125
R29016 DVSS.n5431 DVSS.n5430 0.0106125
R29017 DVSS.n6075 DVSS.n6074 0.0106125
R29018 DVSS.n6776 DVSS.n6775 0.0106125
R29019 DVSS.n3584 DVSS.n3583 0.0106125
R29020 DVSS.n1206 DVSS.n1205 0.0106125
R29021 DVSS.n5586 DVSS.n5571 0.0105984
R29022 DVSS.n5793 DVSS.n5792 0.0105984
R29023 DVSS.n10270 DVSS.n10211 0.0105984
R29024 DVSS.n9841 DVSS.n8586 0.0105984
R29025 DVSS.n12192 DVSS.n12191 0.0105984
R29026 DVSS.n17009 DVSS.n16956 0.0105984
R29027 DVSS.n17565 DVSS.n17564 0.0105984
R29028 DVSS.n10630 DVSS.n10618 0.0105984
R29029 DVSS.n5225 DVSS.n5224 0.0105984
R29030 DVSS.n2821 DVSS.n2820 0.0105984
R29031 DVSS.n9913 DVSS.n9912 0.0105984
R29032 DVSS.n11088 DVSS.n11087 0.0105984
R29033 DVSS.n17304 DVSS.n17266 0.0105984
R29034 DVSS.n16414 DVSS.n16413 0.0105984
R29035 DVSS.n5389 DVSS.n5331 0.0105984
R29036 DVSS.n930 DVSS.n929 0.01057
R29037 DVSS.n5382 DVSS.n5381 0.0105559
R29038 DVSS.n5368 DVSS.n5366 0.0105559
R29039 DVSS.n5607 DVSS.n5606 0.0105559
R29040 DVSS.n17325 DVSS.n17324 0.0105559
R29041 DVSS.n17277 DVSS.n17276 0.0105559
R29042 DVSS.n10220 DVSS.n10218 0.0105559
R29043 DVSS.n10240 DVSS.n10239 0.0105559
R29044 DVSS.n13053 DVSS.n13052 0.0105466
R29045 DVSS.n13054 DVSS.n13053 0.0105466
R29046 DVSS.n6445 DVSS.n6444 0.0105264
R29047 DVSS.n6437 DVSS.n6436 0.0105264
R29048 DVSS.n6356 DVSS.n6355 0.0105264
R29049 DVSS.n6572 DVSS.n1402 0.0105264
R29050 DVSS.n6657 DVSS.n6656 0.0105264
R29051 DVSS.n6715 DVSS.n6664 0.0105264
R29052 DVSS.n6718 DVSS.n6717 0.0105264
R29053 DVSS.n6770 DVSS.n6725 0.0105264
R29054 DVSS.n6839 DVSS.n6838 0.0105264
R29055 DVSS.n6897 DVSS.n6846 0.0105264
R29056 DVSS.n6900 DVSS.n1378 0.0105264
R29057 DVSS.n6444 DVSS.n6443 0.0105264
R29058 DVSS.n6436 DVSS.n6357 0.0105264
R29059 DVSS.n6355 DVSS.n6354 0.0105264
R29060 DVSS.n6573 DVSS.n6572 0.0105264
R29061 DVSS.n6658 DVSS.n6657 0.0105264
R29062 DVSS.n6716 DVSS.n6715 0.0105264
R29063 DVSS.n6719 DVSS.n6718 0.0105264
R29064 DVSS.n6771 DVSS.n6770 0.0105264
R29065 DVSS.n6840 DVSS.n6839 0.0105264
R29066 DVSS.n6898 DVSS.n6897 0.0105264
R29067 DVSS.n6900 DVSS.n6899 0.0105264
R29068 DVSS.n5558 DVSS.n5557 0.010524
R29069 DVSS.n4052 DVSS.n4051 0.010524
R29070 DVSS.n7105 DVSS.n7104 0.010524
R29071 DVSS.n5778 DVSS.n5777 0.010524
R29072 DVSS.n5211 DVSS.n5210 0.010524
R29073 DVSS.n3751 DVSS.n3750 0.010524
R29074 DVSS.n3983 DVSS.n3982 0.010524
R29075 DVSS.n17253 DVSS.n17252 0.010524
R29076 DVSS.n16399 DVSS.n16398 0.010524
R29077 DVSS.n18784 DVSS.n18783 0.010524
R29078 DVSS.n7517 DVSS.n7516 0.010524
R29079 DVSS.n5316 DVSS.n5315 0.010524
R29080 DVSS.n6064 DVSS.n6063 0.010524
R29081 DVSS.n3640 DVSS.n3639 0.010524
R29082 DVSS.n6831 DVSS.n6830 0.010524
R29083 DVSS.n5258 DVSS.n5257 0.0105
R29084 DVSS.n5257 DVSS.n5256 0.0105
R29085 DVSS.n5256 DVSS.n5255 0.0105
R29086 DVSS.n5255 DVSS.n5254 0.0105
R29087 DVSS.n5169 DVSS.n5168 0.0105
R29088 DVSS.n5137 DVSS.n5136 0.0105
R29089 DVSS.n5131 DVSS.n5130 0.0105
R29090 DVSS.n5130 DVSS.n5129 0.0105
R29091 DVSS.n5125 DVSS.n5124 0.0105
R29092 DVSS.n5124 DVSS.n5123 0.0105
R29093 DVSS.n5119 DVSS.n5118 0.0105
R29094 DVSS.n5118 DVSS.n5117 0.0105
R29095 DVSS.n5083 DVSS.n5082 0.0105
R29096 DVSS.n5082 DVSS.n5081 0.0105
R29097 DVSS.n5081 DVSS.n5080 0.0105
R29098 DVSS.n5080 DVSS.n5079 0.0105
R29099 DVSS.n5079 DVSS.n5078 0.0105
R29100 DVSS.n5078 DVSS.n5077 0.0105
R29101 DVSS.n10299 DVSS.n10298 0.0105
R29102 DVSS.n10300 DVSS.n10299 0.0105
R29103 DVSS.n10301 DVSS.n10300 0.0105
R29104 DVSS.n10305 DVSS.n10304 0.0105
R29105 DVSS.n10371 DVSS.n10370 0.0105
R29106 DVSS.n10376 DVSS.n10375 0.0105
R29107 DVSS.n10377 DVSS.n10376 0.0105
R29108 DVSS.n10383 DVSS.n10382 0.0105
R29109 DVSS.n10392 DVSS.n10391 0.0105
R29110 DVSS.n10393 DVSS.n10392 0.0105
R29111 DVSS.n10430 DVSS.n10429 0.0105
R29112 DVSS.n10439 DVSS.n10438 0.0105
R29113 DVSS.n10440 DVSS.n10439 0.0105
R29114 DVSS.n10448 DVSS.n10447 0.0105
R29115 DVSS.n10449 DVSS.n10448 0.0105
R29116 DVSS.n10450 DVSS.n10449 0.0105
R29117 DVSS.n10451 DVSS.n10450 0.0105
R29118 DVSS.n10452 DVSS.n10451 0.0105
R29119 DVSS.n10492 DVSS.n10491 0.0105
R29120 DVSS.n10493 DVSS.n10492 0.0105
R29121 DVSS.n10494 DVSS.n10493 0.0105
R29122 DVSS.n10495 DVSS.n10494 0.0105
R29123 DVSS.n10588 DVSS.n10587 0.0105
R29124 DVSS.n10589 DVSS.n10588 0.0105
R29125 DVSS.n5259 DVSS.n5252 0.0105
R29126 DVSS.n5252 DVSS.n5251 0.0105
R29127 DVSS.n5251 DVSS.n5250 0.0105
R29128 DVSS.n5250 DVSS.n5249 0.0105
R29129 DVSS.n5176 DVSS.n5174 0.0105
R29130 DVSS.n5174 DVSS.n5172 0.0105
R29131 DVSS.n5172 DVSS.n5170 0.0105
R29132 DVSS.n5170 DVSS.n5166 0.0105
R29133 DVSS.n5138 DVSS.n5135 0.0105
R29134 DVSS.n5135 DVSS.n5134 0.0105
R29135 DVSS.n5134 DVSS.n5132 0.0105
R29136 DVSS.n5132 DVSS.n5128 0.0105
R29137 DVSS.n5128 DVSS.n5127 0.0105
R29138 DVSS.n5127 DVSS.n5126 0.0105
R29139 DVSS.n5126 DVSS.n5122 0.0105
R29140 DVSS.n5122 DVSS.n5121 0.0105
R29141 DVSS.n5121 DVSS.n5120 0.0105
R29142 DVSS.n5120 DVSS.n5116 0.0105
R29143 DVSS.n5116 DVSS.n5115 0.0105
R29144 DVSS.n5115 DVSS.n5114 0.0105
R29145 DVSS.n5084 DVSS.n5076 0.0105
R29146 DVSS.n5076 DVSS.n5075 0.0105
R29147 DVSS.n5075 DVSS.n5074 0.0105
R29148 DVSS.n5074 DVSS.n5073 0.0105
R29149 DVSS.n5073 DVSS.n5072 0.0105
R29150 DVSS.n5072 DVSS.n5071 0.0105
R29151 DVSS.n10296 DVSS.n10295 0.0105
R29152 DVSS.n10297 DVSS.n10296 0.0105
R29153 DVSS.n10302 DVSS.n10297 0.0105
R29154 DVSS.n10303 DVSS.n10302 0.0105
R29155 DVSS.n10306 DVSS.n10303 0.0105
R29156 DVSS.n10372 DVSS.n10369 0.0105
R29157 DVSS.n10373 DVSS.n10372 0.0105
R29158 DVSS.n10374 DVSS.n10373 0.0105
R29159 DVSS.n10378 DVSS.n10374 0.0105
R29160 DVSS.n10380 DVSS.n10378 0.0105
R29161 DVSS.n10381 DVSS.n10380 0.0105
R29162 DVSS.n10384 DVSS.n10381 0.0105
R29163 DVSS.n10386 DVSS.n10384 0.0105
R29164 DVSS.n10388 DVSS.n10386 0.0105
R29165 DVSS.n10389 DVSS.n10388 0.0105
R29166 DVSS.n10390 DVSS.n10389 0.0105
R29167 DVSS.n10394 DVSS.n10390 0.0105
R29168 DVSS.n10431 DVSS.n10427 0.0105
R29169 DVSS.n10433 DVSS.n10431 0.0105
R29170 DVSS.n10435 DVSS.n10433 0.0105
R29171 DVSS.n10436 DVSS.n10435 0.0105
R29172 DVSS.n10437 DVSS.n10436 0.0105
R29173 DVSS.n10441 DVSS.n10437 0.0105
R29174 DVSS.n10442 DVSS.n10441 0.0105
R29175 DVSS.n10443 DVSS.n10442 0.0105
R29176 DVSS.n10444 DVSS.n10443 0.0105
R29177 DVSS.n10445 DVSS.n10444 0.0105
R29178 DVSS.n10446 DVSS.n10445 0.0105
R29179 DVSS.n10453 DVSS.n10446 0.0105
R29180 DVSS.n10487 DVSS.n10486 0.0105
R29181 DVSS.n10488 DVSS.n10487 0.0105
R29182 DVSS.n10489 DVSS.n10488 0.0105
R29183 DVSS.n10496 DVSS.n10489 0.0105
R29184 DVSS.n10586 DVSS.n10583 0.0105
R29185 DVSS.n10586 DVSS.n10585 0.0105
R29186 DVSS.n10585 DVSS.n10584 0.0105
R29187 DVSS.n5626 DVSS.n5625 0.0104355
R29188 DVSS.n5194 DVSS.n5193 0.0104355
R29189 DVSS.n17345 DVSS.n17344 0.0104355
R29190 DVSS.n5421 DVSS.n5420 0.0104355
R29191 DVSS.n16519 DVSS.n16518 0.0104296
R29192 DVSS.n16112 DVSS.n16111 0.0104296
R29193 DVSS.n18151 DVSS.n18150 0.0104296
R29194 DVSS.n16864 DVSS.n16863 0.0104296
R29195 DVSS.n15993 DVSS.n15992 0.0104296
R29196 DVSS.n15456 DVSS.n15455 0.0104296
R29197 DVSS.n5799 DVSS.n5798 0.0104213
R29198 DVSS.n9847 DVSS.n9846 0.0104213
R29199 DVSS.n21188 DVSS.n21187 0.0104213
R29200 DVSS.n17559 DVSS.n17558 0.0104213
R29201 DVSS.n10767 DVSS.n10766 0.0104213
R29202 DVSS.n702 DVSS.n701 0.0104213
R29203 DVSS.n11082 DVSS.n11081 0.0104213
R29204 DVSS.n16420 DVSS.n16419 0.0104213
R29205 DVSS.n5493 DVSS.n5492 0.0104213
R29206 DVSS.n7717 DVSS.n7716 0.0104
R29207 DVSS.n15068 DVSS.n15067 0.0104
R29208 DVSS.n16048 DVSS.n16047 0.0104
R29209 DVSS.n13971 DVSS.n13970 0.0104
R29210 DVSS.n5625 DVSS.n5624 0.010347
R29211 DVSS.n5195 DVSS.n5194 0.010347
R29212 DVSS.n17344 DVSS.n17343 0.010347
R29213 DVSS.n5420 DVSS.n5419 0.010347
R29214 DVSS.n11483 DVSS.n11482 0.0103395
R29215 DVSS.n11520 DVSS.n11519 0.0103395
R29216 DVSS.n11645 DVSS.n11644 0.0103395
R29217 DVSS.n11682 DVSS.n11681 0.0103395
R29218 DVSS.n11731 DVSS.n11730 0.0103395
R29219 DVSS.n12532 DVSS.n12531 0.0103077
R29220 DVSS.n12656 DVSS.n12655 0.0103077
R29221 DVSS.n12368 DVSS.n12367 0.0103077
R29222 DVSS.n12276 DVSS.n12275 0.0103077
R29223 DVSS.n12261 DVSS.n12260 0.0103077
R29224 DVSS.n3156 DVSS.n3155 0.0103077
R29225 DVSS.n3280 DVSS.n3279 0.0103077
R29226 DVSS.n2995 DVSS.n2994 0.0103077
R29227 DVSS.n2903 DVSS.n2902 0.0103077
R29228 DVSS.n2888 DVSS.n2887 0.0103077
R29229 DVSS.n9542 DVSS.n9541 0.010282
R29230 DVSS.n12867 DVSS.n12866 0.010282
R29231 DVSS.n9543 DVSS.n9542 0.010282
R29232 DVSS.n15655 DVSS.n15654 0.010282
R29233 DVSS.n20182 DVSS.n20181 0.010282
R29234 DVSS.n20277 DVSS.n20276 0.010282
R29235 DVSS.n20783 DVSS.n20782 0.010282
R29236 DVSS.n15654 DVSS.n15653 0.010282
R29237 DVSS.n11580 DVSS.n11579 0.010282
R29238 DVSS.n29 DVSS.n28 0.010282
R29239 DVSS.n21515 DVSS.n21514 0.010282
R29240 DVSS.n21427 DVSS.n21426 0.010282
R29241 DVSS.n11581 DVSS.n11580 0.010282
R29242 DVSS.n4311 DVSS.n4310 0.010282
R29243 DVSS.n9652 DVSS.n9651 0.010282
R29244 DVSS.n20453 DVSS.n20452 0.010282
R29245 DVSS.n20551 DVSS.n20550 0.010282
R29246 DVSS.n21009 DVSS.n21008 0.010282
R29247 DVSS.n9651 DVSS.n9650 0.010282
R29248 DVSS.n16169 DVSS.n16168 0.010282
R29249 DVSS.n6625 DVSS.n6624 0.010282
R29250 DVSS.n19174 DVSS.n19173 0.010282
R29251 DVSS.n20454 DVSS.n20453 0.010282
R29252 DVSS.n12866 DVSS.n12865 0.010282
R29253 DVSS.n19445 DVSS.n19444 0.010282
R29254 DVSS.n20183 DVSS.n20182 0.010282
R29255 DVSS.n30 DVSS.n29 0.010282
R29256 DVSS.n18982 DVSS.n18981 0.010282
R29257 DVSS.n19534 DVSS.n19533 0.010282
R29258 DVSS.n19263 DVSS.n19262 0.010282
R29259 DVSS.n21516 DVSS.n21515 0.010282
R29260 DVSS.n20550 DVSS.n20549 0.010282
R29261 DVSS.n20276 DVSS.n20275 0.010282
R29262 DVSS.n584 DVSS.n583 0.010282
R29263 DVSS.n1233 DVSS.n1232 0.010282
R29264 DVSS.n1018 DVSS.n1017 0.010282
R29265 DVSS.n21428 DVSS.n21427 0.010282
R29266 DVSS.n21008 DVSS.n21007 0.010282
R29267 DVSS.n20782 DVSS.n20781 0.010282
R29268 DVSS.n4053 DVSS.n4052 0.0102585
R29269 DVSS.n7104 DVSS.n7103 0.0102585
R29270 DVSS.n5779 DVSS.n5778 0.0102585
R29271 DVSS.n5557 DVSS.n5556 0.0102585
R29272 DVSS.n5210 DVSS.n5209 0.0102585
R29273 DVSS.n3982 DVSS.n3981 0.0102585
R29274 DVSS.n3752 DVSS.n3751 0.0102585
R29275 DVSS.n17252 DVSS.n17251 0.0102585
R29276 DVSS.n16400 DVSS.n16399 0.0102585
R29277 DVSS.n7518 DVSS.n7517 0.0102585
R29278 DVSS.n18783 DVSS.n18782 0.0102585
R29279 DVSS.n5315 DVSS.n5314 0.0102585
R29280 DVSS.n6063 DVSS.n6062 0.0102585
R29281 DVSS.n6830 DVSS.n6829 0.0102585
R29282 DVSS.n3639 DVSS.n3638 0.0102585
R29283 DVSS.n12462 DVSS.n12461 0.0102441
R29284 DVSS.n12185 DVSS.n12184 0.0102441
R29285 DVSS.n3088 DVSS.n3087 0.0102441
R29286 DVSS.n2814 DVSS.n2813 0.0102441
R29287 DVSS.n17471 DVSS.n17470 0.0102183
R29288 DVSS.n16812 DVSS.n16811 0.0102183
R29289 DVSS.n15431 DVSS.n15430 0.010175
R29290 DVSS.n18281 DVSS.n18280 0.010175
R29291 DVSS.n18330 DVSS.n18329 0.010175
R29292 DVSS.n18345 DVSS.n18344 0.010175
R29293 DVSS.n13861 DVSS.n13860 0.010175
R29294 DVSS.n5637 DVSS.n5636 0.01017
R29295 DVSS.n5768 DVSS.n5767 0.01017
R29296 DVSS.n4079 DVSS.n4078 0.01017
R29297 DVSS.n6973 DVSS.n6972 0.01017
R29298 DVSS.n4707 DVSS.n4706 0.01017
R29299 DVSS.n3794 DVSS.n3793 0.01017
R29300 DVSS.n3778 DVSS.n3777 0.01017
R29301 DVSS.n17356 DVSS.n17355 0.01017
R29302 DVSS.n16389 DVSS.n16388 0.01017
R29303 DVSS.n18740 DVSS.n18739 0.01017
R29304 DVSS.n7544 DVSS.n7543 0.01017
R29305 DVSS.n5432 DVSS.n5431 0.01017
R29306 DVSS.n6074 DVSS.n6073 0.01017
R29307 DVSS.n6775 DVSS.n6774 0.01017
R29308 DVSS.n3583 DVSS.n3582 0.01017
R29309 DVSS.n6760 DVSS.n6759 0.0101595
R29310 DVSS.n6705 DVSS.n6704 0.0101595
R29311 DVSS.n2537 DVSS.n2536 0.0101595
R29312 DVSS.n6398 DVSS.n6397 0.0101595
R29313 DVSS.n6887 DVSS.n6886 0.0101595
R29314 DVSS.n4443 DVSS.n4442 0.0100815
R29315 DVSS.n19287 DVSS.n19286 0.0100815
R29316 DVSS.n859 DVSS.n858 0.0100815
R29317 DVSS.n4393 DVSS.n4392 0.0100815
R29318 DVSS.n4337 DVSS.n4336 0.0100815
R29319 DVSS.n4287 DVSS.n4286 0.0100815
R29320 DVSS.n16142 DVSS.n16141 0.0100815
R29321 DVSS.n1146 DVSS.n1145 0.0100815
R29322 DVSS.n16193 DVSS.n16192 0.0100815
R29323 DVSS.n6652 DVSS.n6651 0.0100815
R29324 DVSS.n18959 DVSS.n18958 0.0100815
R29325 DVSS.n19006 DVSS.n19005 0.0100815
R29326 DVSS.n537 DVSS.n536 0.0100815
R29327 DVSS.n558 DVSS.n557 0.0100815
R29328 DVSS.n6601 DVSS.n6600 0.0100815
R29329 DVSS.n19392 DVSS.n19391 0.0100815
R29330 DVSS.n19118 DVSS.n19117 0.0100815
R29331 DVSS.n3500 DVSS.n3499 0.0100815
R29332 DVSS.n3562 DVSS.n3561 0.0100815
R29333 DVSS.n19558 DVSS.n19557 0.0100815
R29334 DVSS.n1257 DVSS.n1256 0.0100815
R29335 DVSS.n1042 DVSS.n1041 0.0100815
R29336 DVSS.n608 DVSS.n607 0.0100815
R29337 DVSS.n1207 DVSS.n1206 0.0100815
R29338 DVSS.n7166 DVSS.n7164 0.0100745
R29339 DVSS.n7301 DVSS.n7299 0.0100745
R29340 DVSS.n7310 DVSS.n7309 0.0100745
R29341 DVSS.n7870 DVSS.n7868 0.0100745
R29342 DVSS.n7880 DVSS.n7878 0.0100745
R29343 DVSS.n7958 DVSS.n7956 0.0100745
R29344 DVSS.n7965 DVSS.n7964 0.0100745
R29345 DVSS.n7035 DVSS.n7033 0.0100745
R29346 DVSS.n7076 DVSS.n7074 0.0100745
R29347 DVSS.n7064 DVSS.n7063 0.0100745
R29348 DVSS.n13607 DVSS.n13604 0.0100745
R29349 DVSS.n13627 DVSS.n13624 0.0100745
R29350 DVSS.n13299 DVSS.n13297 0.0100745
R29351 DVSS.n13317 DVSS.n13316 0.0100745
R29352 DVSS.n15745 DVSS.n15744 0.0100303
R29353 DVSS.n15817 DVSS.n15816 0.0100303
R29354 DVSS.n15235 DVSS.n15234 0.0100303
R29355 DVSS.n15571 DVSS.n15570 0.0100303
R29356 DVSS.n18514 DVSS.n18513 0.0100303
R29357 DVSS.n3786 DVSS.n3785 0.0100173
R29358 DVSS.n3787 DVSS.n3786 0.0100173
R29359 DVSS.n4416 DVSS.n4415 0.00999298
R29360 DVSS.n19177 DVSS.n19176 0.00999298
R29361 DVSS.n3473 DVSS.n3472 0.00999298
R29362 DVSS.n4314 DVSS.n4313 0.00999298
R29363 DVSS.n19448 DVSS.n19447 0.00999298
R29364 DVSS.n3535 DVSS.n3534 0.00999298
R29365 DVSS.n19531 DVSS.n19530 0.00999298
R29366 DVSS.n19260 DVSS.n19259 0.00999298
R29367 DVSS.n18979 DVSS.n18978 0.00999298
R29368 DVSS.n1230 DVSS.n1229 0.00999298
R29369 DVSS.n1015 DVSS.n1014 0.00999298
R29370 DVSS.n581 DVSS.n580 0.00999298
R29371 DVSS.n17213 DVSS.n17212 0.00995
R29372 DVSS.n15181 DVSS.n15180 0.00995
R29373 DVSS.n15150 DVSS.n15149 0.00995
R29374 DVSS.n15108 DVSS.n15107 0.00995
R29375 DVSS.n17691 DVSS.n17690 0.00995
R29376 DVSS.n5834 DVSS.n5833 0.00994444
R29377 DVSS.n11030 DVSS.n11029 0.00994444
R29378 DVSS.n6474 DVSS.n6473 0.00994444
R29379 DVSS.n11203 DVSS.n11202 0.00994444
R29380 DVSS.n5515 DVSS.n5514 0.00994444
R29381 DVSS.n10042 DVSS.n10041 0.00994444
R29382 DVSS.n10339 DVSS.n10338 0.00993662
R29383 DVSS.n10337 DVSS.n10336 0.00993662
R29384 DVSS.n12826 DVSS.n12825 0.0099291
R29385 DVSS.n12827 DVSS.n12826 0.0099291
R29386 DVSS.n12502 DVSS.n12501 0.00992308
R29387 DVSS.n12511 DVSS.n12510 0.00992308
R29388 DVSS.n12635 DVSS.n12634 0.00992308
R29389 DVSS.n12626 DVSS.n12625 0.00992308
R29390 DVSS.n12347 DVSS.n12346 0.00992308
R29391 DVSS.n12338 DVSS.n12337 0.00992308
R29392 DVSS.n21325 DVSS.n21324 0.00992308
R29393 DVSS.n3126 DVSS.n3125 0.00992308
R29394 DVSS.n3135 DVSS.n3134 0.00992308
R29395 DVSS.n3259 DVSS.n3258 0.00992308
R29396 DVSS.n3250 DVSS.n3249 0.00992308
R29397 DVSS.n2974 DVSS.n2973 0.00992308
R29398 DVSS.n2965 DVSS.n2964 0.00992308
R29399 DVSS.n900 DVSS.n899 0.00992308
R29400 DVSS.n909 DVSS.n908 0.00992308
R29401 DVSS.n380 DVSS.n379 0.00989057
R29402 DVSS.n19201 DVSS.n19200 0.00988976
R29403 DVSS.n20212 DVSS.n20211 0.00988976
R29404 DVSS.n20483 DVSS.n20482 0.00988976
R29405 DVSS.n19472 DVSS.n19471 0.00988976
R29406 DVSS.n3994 DVSS.n3993 0.00984086
R29407 DVSS.n3993 DVSS.n3992 0.00984086
R29408 DVSS.n9805 DVSS.n9804 0.00984086
R29409 DVSS.n9710 DVSS.n9709 0.00984086
R29410 DVSS.n9613 DVSS.n9612 0.00984086
R29411 DVSS.n9098 DVSS.n9097 0.00984086
R29412 DVSS.n9048 DVSS.n9047 0.00984086
R29413 DVSS.n9806 DVSS.n9805 0.00984086
R29414 DVSS.n9709 DVSS.n9708 0.00984086
R29415 DVSS.n9614 DVSS.n9613 0.00984086
R29416 DVSS.n9097 DVSS.n9096 0.00984086
R29417 DVSS.n9049 DVSS.n9048 0.00984086
R29418 DVSS.n16294 DVSS.n16293 0.00984086
R29419 DVSS.n16255 DVSS.n16254 0.00984086
R29420 DVSS.n16134 DVSS.n16133 0.00984086
R29421 DVSS.n18382 DVSS.n18381 0.00984086
R29422 DVSS.n7506 DVSS.n7505 0.00984086
R29423 DVSS.n16295 DVSS.n16294 0.00984086
R29424 DVSS.n16256 DVSS.n16255 0.00984086
R29425 DVSS.n16135 DVSS.n16134 0.00984086
R29426 DVSS.n18381 DVSS.n18380 0.00984086
R29427 DVSS.n7507 DVSS.n7506 0.00984086
R29428 DVSS.n18438 DVSS.n18437 0.00979577
R29429 DVSS.n15191 DVSS.n15178 0.00979577
R29430 DVSS.n17190 DVSS 0.009725
R29431 DVSS DVSS.n17719 0.009725
R29432 DVSS.n17492 DVSS 0.009725
R29433 DVSS DVSS.n15299 0.009725
R29434 DVSS.n15392 DVSS.n15391 0.009725
R29435 DVSS.n15395 DVSS.n15394 0.009725
R29436 DVSS.n18299 DVSS.n18298 0.009725
R29437 DVSS.n18302 DVSS.n18301 0.009725
R29438 DVSS.n18040 DVSS 0.009725
R29439 DVSS.n17899 DVSS 0.009725
R29440 DVSS.n13934 DVSS 0.009725
R29441 DVSS.n5659 DVSS.n5658 0.0097126
R29442 DVSS.n10952 DVSS.n10951 0.0097126
R29443 DVSS.n17085 DVSS.n17084 0.0097126
R29444 DVSS.n4690 DVSS.n4689 0.0097126
R29445 DVSS.n9974 DVSS.n9973 0.0097126
R29446 DVSS.n17378 DVSS.n17377 0.0097126
R29447 DVSS.n17882 DVSS.n17881 0.00969863
R29448 DVSS.n18023 DVSS.n18022 0.00969863
R29449 DVSS.n18169 DVSS.n18168 0.00969863
R29450 DVSS.n7574 DVSS.n7573 0.00969863
R29451 DVSS.n171 DVSS.n170 0.00969863
R29452 DVSS.n168 DVSS.n167 0.00969863
R29453 DVSS.n7755 DVSS.n7754 0.00969863
R29454 DVSS.n14227 DVSS.n14226 0.00964533
R29455 DVSS.n14246 DVSS.n14245 0.00964533
R29456 DVSS.n14260 DVSS.n14259 0.00964533
R29457 DVSS.n14271 DVSS.n14270 0.00964533
R29458 DVSS.n14285 DVSS.n14284 0.00964533
R29459 DVSS.n14296 DVSS.n14295 0.00964533
R29460 DVSS.n14314 DVSS.n14313 0.00964533
R29461 DVSS.n14325 DVSS.n14324 0.00964533
R29462 DVSS.n14356 DVSS.n14355 0.00964533
R29463 DVSS.n14433 DVSS.n14432 0.00964533
R29464 DVSS.n14448 DVSS.n14447 0.00964533
R29465 DVSS.n14324 DVSS.n14323 0.00964533
R29466 DVSS.n14259 DVSS.n14258 0.00964533
R29467 DVSS.n14270 DVSS.n14269 0.00964533
R29468 DVSS.n14284 DVSS.n14283 0.00964533
R29469 DVSS.n14295 DVSS.n14294 0.00964533
R29470 DVSS.n14313 DVSS.n14312 0.00964533
R29471 DVSS.n14245 DVSS.n14244 0.00964533
R29472 DVSS.n14226 DVSS.n14223 0.00964533
R29473 DVSS.n14447 DVSS.n14446 0.00964533
R29474 DVSS.n14432 DVSS.n14431 0.00964533
R29475 DVSS.n14355 DVSS.n14350 0.00964533
R29476 DVSS.n14872 DVSS.n14871 0.00964533
R29477 DVSS.n14861 DVSS.n14860 0.00964533
R29478 DVSS.n14855 DVSS.n14854 0.00964533
R29479 DVSS.n14844 DVSS.n14843 0.00964533
R29480 DVSS.n14838 DVSS.n14837 0.00964533
R29481 DVSS.n14827 DVSS.n14826 0.00964533
R29482 DVSS.n14821 DVSS.n14820 0.00964533
R29483 DVSS.n14810 DVSS.n14809 0.00964533
R29484 DVSS.n14793 DVSS.n14792 0.00964533
R29485 DVSS.n14695 DVSS.n14694 0.00964533
R29486 DVSS.n14674 DVSS.n14673 0.00964533
R29487 DVSS.n14811 DVSS.n14810 0.00964533
R29488 DVSS.n14856 DVSS.n14855 0.00964533
R29489 DVSS.n14845 DVSS.n14844 0.00964533
R29490 DVSS.n14839 DVSS.n14838 0.00964533
R29491 DVSS.n14828 DVSS.n14827 0.00964533
R29492 DVSS.n14822 DVSS.n14821 0.00964533
R29493 DVSS.n14862 DVSS.n14861 0.00964533
R29494 DVSS.n14873 DVSS.n14872 0.00964533
R29495 DVSS.n14794 DVSS.n14793 0.00964533
R29496 DVSS.n14675 DVSS.n14674 0.00964533
R29497 DVSS.n14696 DVSS.n14695 0.00964533
R29498 DVSS.n16682 DVSS.n16681 0.00962875
R29499 DVSS.n17141 DVSS.n17140 0.00962875
R29500 DVSS.n2434 DVSS.n2433 0.00962857
R29501 DVSS.n2433 DVSS.n2432 0.00962857
R29502 DVSS.n2432 DVSS.n2431 0.00962857
R29503 DVSS.n2431 DVSS.n2430 0.00962857
R29504 DVSS.n2430 DVSS.n2429 0.00962857
R29505 DVSS.n2429 DVSS.n2428 0.00962857
R29506 DVSS.n2428 DVSS.n2427 0.00962857
R29507 DVSS.n2427 DVSS.n2426 0.00962857
R29508 DVSS.n2426 DVSS.n2425 0.00962857
R29509 DVSS.n1971 DVSS.n1970 0.00962857
R29510 DVSS.n1970 DVSS.n1969 0.00962857
R29511 DVSS.n1961 DVSS.n1960 0.00962857
R29512 DVSS.n1947 DVSS.n1946 0.00962857
R29513 DVSS.n1946 DVSS.n1945 0.00962857
R29514 DVSS.n2143 DVSS.n2142 0.00962857
R29515 DVSS.n2147 DVSS.n2146 0.00962857
R29516 DVSS.n2217 DVSS.n2216 0.00962857
R29517 DVSS.n2231 DVSS.n2230 0.00962857
R29518 DVSS.n2235 DVSS.n2234 0.00962857
R29519 DVSS.n2056 DVSS.n2054 0.00962857
R29520 DVSS.n2021 DVSS.n2012 0.00962857
R29521 DVSS.n2023 DVSS.n2021 0.00962857
R29522 DVSS.n2025 DVSS.n2023 0.00962857
R29523 DVSS.n2027 DVSS.n2025 0.00962857
R29524 DVSS.n2029 DVSS.n2027 0.00962857
R29525 DVSS.n2031 DVSS.n2029 0.00962857
R29526 DVSS.n2033 DVSS.n2031 0.00962857
R29527 DVSS.n2035 DVSS.n2033 0.00962857
R29528 DVSS.n2037 DVSS.n2035 0.00962857
R29529 DVSS.n2042 DVSS.n2037 0.00962857
R29530 DVSS.n2071 DVSS.n2069 0.00962857
R29531 DVSS.n2073 DVSS.n2071 0.00962857
R29532 DVSS.n2075 DVSS.n2073 0.00962857
R29533 DVSS.n2077 DVSS.n2075 0.00962857
R29534 DVSS.n2079 DVSS.n2077 0.00962857
R29535 DVSS.n2081 DVSS.n2079 0.00962857
R29536 DVSS.n2083 DVSS.n2081 0.00962857
R29537 DVSS.n2085 DVSS.n2083 0.00962857
R29538 DVSS.n2087 DVSS.n2085 0.00962857
R29539 DVSS.n2089 DVSS.n2087 0.00962857
R29540 DVSS.n2091 DVSS.n2089 0.00962857
R29541 DVSS.n2093 DVSS.n2091 0.00962857
R29542 DVSS.n2095 DVSS.n2093 0.00962857
R29543 DVSS.n2097 DVSS.n2095 0.00962857
R29544 DVSS.n2099 DVSS.n2097 0.00962857
R29545 DVSS.n2101 DVSS.n2099 0.00962857
R29546 DVSS.n2103 DVSS.n2101 0.00962857
R29547 DVSS.n2105 DVSS.n2103 0.00962857
R29548 DVSS.n2107 DVSS.n2105 0.00962857
R29549 DVSS.n2109 DVSS.n2107 0.00962857
R29550 DVSS.n2111 DVSS.n2109 0.00962857
R29551 DVSS.n2113 DVSS.n2111 0.00962857
R29552 DVSS.n2115 DVSS.n2113 0.00962857
R29553 DVSS.n2117 DVSS.n2115 0.00962857
R29554 DVSS.n2119 DVSS.n2117 0.00962857
R29555 DVSS.n2121 DVSS.n2119 0.00962857
R29556 DVSS.n2123 DVSS.n2121 0.00962857
R29557 DVSS.n2125 DVSS.n2123 0.00962857
R29558 DVSS.n2127 DVSS.n2125 0.00962857
R29559 DVSS.n2129 DVSS.n2127 0.00962857
R29560 DVSS.n2131 DVSS.n2129 0.00962857
R29561 DVSS.n2133 DVSS.n2131 0.00962857
R29562 DVSS.n2135 DVSS.n2133 0.00962857
R29563 DVSS.n2137 DVSS.n2135 0.00962857
R29564 DVSS.n2139 DVSS.n2137 0.00962857
R29565 DVSS.n2141 DVSS.n2139 0.00962857
R29566 DVSS.n2144 DVSS.n2141 0.00962857
R29567 DVSS.n2145 DVSS.n2144 0.00962857
R29568 DVSS.n2148 DVSS.n2145 0.00962857
R29569 DVSS.n2149 DVSS.n2148 0.00962857
R29570 DVSS.n2151 DVSS.n2149 0.00962857
R29571 DVSS.n2153 DVSS.n2151 0.00962857
R29572 DVSS.n2155 DVSS.n2153 0.00962857
R29573 DVSS.n2157 DVSS.n2155 0.00962857
R29574 DVSS.n2159 DVSS.n2157 0.00962857
R29575 DVSS.n2161 DVSS.n2159 0.00962857
R29576 DVSS.n2163 DVSS.n2161 0.00962857
R29577 DVSS.n2165 DVSS.n2163 0.00962857
R29578 DVSS.n2167 DVSS.n2165 0.00962857
R29579 DVSS.n2169 DVSS.n2167 0.00962857
R29580 DVSS.n2171 DVSS.n2169 0.00962857
R29581 DVSS.n2173 DVSS.n2171 0.00962857
R29582 DVSS.n2175 DVSS.n2173 0.00962857
R29583 DVSS.n2177 DVSS.n2175 0.00962857
R29584 DVSS.n2179 DVSS.n2177 0.00962857
R29585 DVSS.n2181 DVSS.n2179 0.00962857
R29586 DVSS.n2183 DVSS.n2181 0.00962857
R29587 DVSS.n2185 DVSS.n2183 0.00962857
R29588 DVSS.n2187 DVSS.n2185 0.00962857
R29589 DVSS.n2189 DVSS.n2187 0.00962857
R29590 DVSS.n2191 DVSS.n2189 0.00962857
R29591 DVSS.n2193 DVSS.n2191 0.00962857
R29592 DVSS.n2195 DVSS.n2193 0.00962857
R29593 DVSS.n2197 DVSS.n2195 0.00962857
R29594 DVSS.n2199 DVSS.n2197 0.00962857
R29595 DVSS.n2201 DVSS.n2199 0.00962857
R29596 DVSS.n2203 DVSS.n2201 0.00962857
R29597 DVSS.n2205 DVSS.n2203 0.00962857
R29598 DVSS.n2207 DVSS.n2205 0.00962857
R29599 DVSS.n2209 DVSS.n2207 0.00962857
R29600 DVSS.n2211 DVSS.n2209 0.00962857
R29601 DVSS.n2213 DVSS.n2211 0.00962857
R29602 DVSS.n2215 DVSS.n2213 0.00962857
R29603 DVSS.n2218 DVSS.n2215 0.00962857
R29604 DVSS.n2219 DVSS.n2218 0.00962857
R29605 DVSS.n2221 DVSS.n2219 0.00962857
R29606 DVSS.n2223 DVSS.n2221 0.00962857
R29607 DVSS.n2225 DVSS.n2223 0.00962857
R29608 DVSS.n2227 DVSS.n2225 0.00962857
R29609 DVSS.n2229 DVSS.n2227 0.00962857
R29610 DVSS.n2232 DVSS.n2229 0.00962857
R29611 DVSS.n2233 DVSS.n2232 0.00962857
R29612 DVSS.n2236 DVSS.n2233 0.00962857
R29613 DVSS.n2237 DVSS.n2236 0.00962857
R29614 DVSS.n2239 DVSS.n2237 0.00962857
R29615 DVSS.n2457 DVSS.n2435 0.00962857
R29616 DVSS.n2435 DVSS.n2423 0.00962857
R29617 DVSS.n2423 DVSS.n2422 0.00962857
R29618 DVSS.n2422 DVSS.n2421 0.00962857
R29619 DVSS.n2421 DVSS.n2420 0.00962857
R29620 DVSS.n2420 DVSS.n2419 0.00962857
R29621 DVSS.n2419 DVSS.n2418 0.00962857
R29622 DVSS.n2418 DVSS.n2417 0.00962857
R29623 DVSS.n2417 DVSS.n2416 0.00962857
R29624 DVSS.n2416 DVSS.n2415 0.00962857
R29625 DVSS.n1994 DVSS.n1992 0.00962857
R29626 DVSS.n1992 DVSS.n1990 0.00962857
R29627 DVSS.n1990 DVSS.n1988 0.00962857
R29628 DVSS.n1988 DVSS.n1986 0.00962857
R29629 DVSS.n1986 DVSS.n1984 0.00962857
R29630 DVSS.n1984 DVSS.n1982 0.00962857
R29631 DVSS.n1982 DVSS.n1980 0.00962857
R29632 DVSS.n1980 DVSS.n1978 0.00962857
R29633 DVSS.n1978 DVSS.n1976 0.00962857
R29634 DVSS.n1976 DVSS.n1974 0.00962857
R29635 DVSS.n1974 DVSS.n1972 0.00962857
R29636 DVSS.n1972 DVSS.n1968 0.00962857
R29637 DVSS.n1968 DVSS.n1967 0.00962857
R29638 DVSS.n1967 DVSS.n1966 0.00962857
R29639 DVSS.n1966 DVSS.n1964 0.00962857
R29640 DVSS.n1964 DVSS.n1962 0.00962857
R29641 DVSS.n1962 DVSS.n1959 0.00962857
R29642 DVSS.n1959 DVSS.n1958 0.00962857
R29643 DVSS.n1958 DVSS.n1956 0.00962857
R29644 DVSS.n1956 DVSS.n1954 0.00962857
R29645 DVSS.n1954 DVSS.n1952 0.00962857
R29646 DVSS.n1952 DVSS.n1950 0.00962857
R29647 DVSS.n1950 DVSS.n1948 0.00962857
R29648 DVSS.n1948 DVSS.n1944 0.00962857
R29649 DVSS.n1944 DVSS.n1943 0.00962857
R29650 DVSS.n1943 DVSS.n1942 0.00962857
R29651 DVSS.n1942 DVSS.n1940 0.00962857
R29652 DVSS.n1940 DVSS.n1938 0.00962857
R29653 DVSS.n1938 DVSS.n1937 0.00962857
R29654 DVSS.n1937 DVSS.n1936 0.00962857
R29655 DVSS.n1936 DVSS.n1935 0.00962857
R29656 DVSS.n1935 DVSS.n1934 0.00962857
R29657 DVSS.n1934 DVSS.n1933 0.00962857
R29658 DVSS.n1933 DVSS.n1932 0.00962857
R29659 DVSS.n1932 DVSS.n1931 0.00962857
R29660 DVSS.n1931 DVSS.n1930 0.00962857
R29661 DVSS.n1930 DVSS.n1929 0.00962857
R29662 DVSS.n1929 DVSS.n1928 0.00962857
R29663 DVSS.n1928 DVSS.n1927 0.00962857
R29664 DVSS.n1927 DVSS.n1926 0.00962857
R29665 DVSS.n1926 DVSS.n1925 0.00962857
R29666 DVSS.n1925 DVSS.n1924 0.00962857
R29667 DVSS.n1924 DVSS.n1923 0.00962857
R29668 DVSS.n1923 DVSS.n1922 0.00962857
R29669 DVSS.n1922 DVSS.n1921 0.00962857
R29670 DVSS.n1921 DVSS.n1920 0.00962857
R29671 DVSS.n1920 DVSS.n1919 0.00962857
R29672 DVSS.n1919 DVSS.n1918 0.00962857
R29673 DVSS.n1918 DVSS.n1917 0.00962857
R29674 DVSS.n1917 DVSS.n1916 0.00962857
R29675 DVSS.n1916 DVSS.n1915 0.00962857
R29676 DVSS.n1915 DVSS.n1914 0.00962857
R29677 DVSS.n1914 DVSS.n1913 0.00962857
R29678 DVSS.n1913 DVSS.n1912 0.00962857
R29679 DVSS.n1912 DVSS.n1911 0.00962857
R29680 DVSS.n1911 DVSS.n1910 0.00962857
R29681 DVSS.n1910 DVSS.n1909 0.00962857
R29682 DVSS.n1909 DVSS.n1908 0.00962857
R29683 DVSS.n1908 DVSS.n1907 0.00962857
R29684 DVSS.n1907 DVSS.n1906 0.00962857
R29685 DVSS.n1906 DVSS.n1905 0.00962857
R29686 DVSS.n1905 DVSS.n1904 0.00962857
R29687 DVSS.n1716 DVSS.n1715 0.00962857
R29688 DVSS.n1715 DVSS.n1713 0.00962857
R29689 DVSS.n1713 DVSS.n1553 0.00962857
R29690 DVSS.n1722 DVSS.n1553 0.00962857
R29691 DVSS.n4985 DVSS.n4984 0.00962857
R29692 DVSS.n4984 DVSS.n4983 0.00962857
R29693 DVSS.n4983 DVSS.n4982 0.00962857
R29694 DVSS.n4982 DVSS.n4981 0.00962857
R29695 DVSS.n4941 DVSS.n4940 0.00962857
R29696 DVSS.n4940 DVSS.n4939 0.00962857
R29697 DVSS.n4939 DVSS.n4938 0.00962857
R29698 DVSS.n4938 DVSS.n4937 0.00962857
R29699 DVSS.n4897 DVSS.n4896 0.00962857
R29700 DVSS.n4896 DVSS.n4895 0.00962857
R29701 DVSS.n4895 DVSS.n4894 0.00962857
R29702 DVSS.n4894 DVSS.n4893 0.00962857
R29703 DVSS.n4893 DVSS.n4892 0.00962857
R29704 DVSS.n4892 DVSS.n4891 0.00962857
R29705 DVSS.n4891 DVSS.n4890 0.00962857
R29706 DVSS.n4881 DVSS.n4880 0.00962857
R29707 DVSS.n4880 DVSS.n4879 0.00962857
R29708 DVSS.n4875 DVSS.n4874 0.00962857
R29709 DVSS.n4833 DVSS.n4832 0.00962857
R29710 DVSS.n4823 DVSS.n4822 0.00962857
R29711 DVSS.n4822 DVSS.n4821 0.00962857
R29712 DVSS.n4821 DVSS.n4820 0.00962857
R29713 DVSS.n4820 DVSS.n4819 0.00962857
R29714 DVSS.n4819 DVSS.n4818 0.00962857
R29715 DVSS.n4742 DVSS.n4741 0.00962857
R29716 DVSS.n4741 DVSS.n4740 0.00962857
R29717 DVSS.n4740 DVSS.n4739 0.00962857
R29718 DVSS.n4739 DVSS.n4738 0.00962857
R29719 DVSS.n4738 DVSS.n4737 0.00962857
R29720 DVSS.n4730 DVSS.n4729 0.00962857
R29721 DVSS.n4729 DVSS.n4728 0.00962857
R29722 DVSS.n4728 DVSS.n4727 0.00962857
R29723 DVSS.n4727 DVSS.n4726 0.00962857
R29724 DVSS.n4726 DVSS.n4725 0.00962857
R29725 DVSS.n10107 DVSS.n10106 0.00962857
R29726 DVSS.n10108 DVSS.n10107 0.00962857
R29727 DVSS.n10109 DVSS.n10108 0.00962857
R29728 DVSS.n10110 DVSS.n10109 0.00962857
R29729 DVSS.n10111 DVSS.n10110 0.00962857
R29730 DVSS.n10112 DVSS.n10111 0.00962857
R29731 DVSS.n10113 DVSS.n10112 0.00962857
R29732 DVSS.n10114 DVSS.n10113 0.00962857
R29733 DVSS.n10115 DVSS.n10114 0.00962857
R29734 DVSS.n10116 DVSS.n10115 0.00962857
R29735 DVSS.n10117 DVSS.n10116 0.00962857
R29736 DVSS.n10118 DVSS.n10117 0.00962857
R29737 DVSS.n10161 DVSS.n10160 0.00962857
R29738 DVSS.n10162 DVSS.n10161 0.00962857
R29739 DVSS.n10709 DVSS.n10708 0.00962857
R29740 DVSS.n4986 DVSS.n4980 0.00962857
R29741 DVSS.n4980 DVSS.n4979 0.00962857
R29742 DVSS.n4979 DVSS.n4978 0.00962857
R29743 DVSS.n4978 DVSS.n4977 0.00962857
R29744 DVSS.n4942 DVSS.n4936 0.00962857
R29745 DVSS.n4936 DVSS.n4935 0.00962857
R29746 DVSS.n4935 DVSS.n4934 0.00962857
R29747 DVSS.n4934 DVSS.n4933 0.00962857
R29748 DVSS.n4898 DVSS.n4889 0.00962857
R29749 DVSS.n4889 DVSS.n4888 0.00962857
R29750 DVSS.n4888 DVSS.n4887 0.00962857
R29751 DVSS.n4887 DVSS.n4886 0.00962857
R29752 DVSS.n4886 DVSS.n4885 0.00962857
R29753 DVSS.n4885 DVSS.n4884 0.00962857
R29754 DVSS.n4884 DVSS.n4883 0.00962857
R29755 DVSS.n4883 DVSS.n4882 0.00962857
R29756 DVSS.n4882 DVSS.n4878 0.00962857
R29757 DVSS.n4878 DVSS.n4877 0.00962857
R29758 DVSS.n4877 DVSS.n4876 0.00962857
R29759 DVSS.n4876 DVSS.n4873 0.00962857
R29760 DVSS.n4838 DVSS.n4836 0.00962857
R29761 DVSS.n4836 DVSS.n4834 0.00962857
R29762 DVSS.n4834 DVSS.n4831 0.00962857
R29763 DVSS.n4831 DVSS.n4830 0.00962857
R29764 DVSS.n4830 DVSS.n4828 0.00962857
R29765 DVSS.n4828 DVSS.n4826 0.00962857
R29766 DVSS.n4826 DVSS.n4824 0.00962857
R29767 DVSS.n4824 DVSS.n4817 0.00962857
R29768 DVSS.n4817 DVSS.n4816 0.00962857
R29769 DVSS.n4816 DVSS.n4815 0.00962857
R29770 DVSS.n4815 DVSS.n4814 0.00962857
R29771 DVSS.n4814 DVSS.n4813 0.00962857
R29772 DVSS.n4743 DVSS.n4736 0.00962857
R29773 DVSS.n4736 DVSS.n4735 0.00962857
R29774 DVSS.n4735 DVSS.n4734 0.00962857
R29775 DVSS.n4734 DVSS.n4733 0.00962857
R29776 DVSS.n4733 DVSS.n4732 0.00962857
R29777 DVSS.n4732 DVSS.n4731 0.00962857
R29778 DVSS.n4731 DVSS.n4724 0.00962857
R29779 DVSS.n4724 DVSS.n4723 0.00962857
R29780 DVSS.n4723 DVSS.n4722 0.00962857
R29781 DVSS.n4722 DVSS.n4721 0.00962857
R29782 DVSS.n4721 DVSS.n4720 0.00962857
R29783 DVSS.n10091 DVSS.n10090 0.00962857
R29784 DVSS.n10092 DVSS.n10091 0.00962857
R29785 DVSS.n10093 DVSS.n10092 0.00962857
R29786 DVSS.n10094 DVSS.n10093 0.00962857
R29787 DVSS.n10095 DVSS.n10094 0.00962857
R29788 DVSS.n10096 DVSS.n10095 0.00962857
R29789 DVSS.n10097 DVSS.n10096 0.00962857
R29790 DVSS.n10098 DVSS.n10097 0.00962857
R29791 DVSS.n10099 DVSS.n10098 0.00962857
R29792 DVSS.n10100 DVSS.n10099 0.00962857
R29793 DVSS.n10101 DVSS.n10100 0.00962857
R29794 DVSS.n10119 DVSS.n10101 0.00962857
R29795 DVSS.n10158 DVSS.n10157 0.00962857
R29796 DVSS.n10163 DVSS.n10158 0.00962857
R29797 DVSS.n10165 DVSS.n10163 0.00962857
R29798 DVSS.n10167 DVSS.n10165 0.00962857
R29799 DVSS.n10711 DVSS.n10710 0.00962857
R29800 DVSS.n10713 DVSS.n10711 0.00962857
R29801 DVSS.n10714 DVSS.n10713 0.00962857
R29802 DVSS.n3833 DVSS.n3832 0.00962857
R29803 DVSS.n3832 DVSS.n3831 0.00962857
R29804 DVSS.n6802 DVSS.n6800 0.00962857
R29805 DVSS.n3810 DVSS.n3808 0.00962857
R29806 DVSS.n3812 DVSS.n3810 0.00962857
R29807 DVSS.n3924 DVSS.n3922 0.00962857
R29808 DVSS.n3922 DVSS.n3920 0.00962857
R29809 DVSS.n3920 DVSS.n3918 0.00962857
R29810 DVSS.n3918 DVSS.n3916 0.00962857
R29811 DVSS.n3894 DVSS.n3892 0.00962857
R29812 DVSS.n3892 DVSS.n3890 0.00962857
R29813 DVSS.n3890 DVSS.n3888 0.00962857
R29814 DVSS.n3888 DVSS.n3886 0.00962857
R29815 DVSS.n3886 DVSS.n3884 0.00962857
R29816 DVSS.n3884 DVSS.n3882 0.00962857
R29817 DVSS.n3882 DVSS.n3880 0.00962857
R29818 DVSS.n3880 DVSS.n3878 0.00962857
R29819 DVSS.n3878 DVSS.n3876 0.00962857
R29820 DVSS.n3876 DVSS.n3874 0.00962857
R29821 DVSS.n3874 DVSS.n3872 0.00962857
R29822 DVSS.n3872 DVSS.n3870 0.00962857
R29823 DVSS.n3848 DVSS.n3846 0.00962857
R29824 DVSS.n3846 DVSS.n3844 0.00962857
R29825 DVSS.n3844 DVSS.n3842 0.00962857
R29826 DVSS.n3842 DVSS.n3840 0.00962857
R29827 DVSS.n3840 DVSS.n3838 0.00962857
R29828 DVSS.n3838 DVSS.n3836 0.00962857
R29829 DVSS.n3836 DVSS.n3834 0.00962857
R29830 DVSS.n3834 DVSS.n3830 0.00962857
R29831 DVSS.n3830 DVSS.n3829 0.00962857
R29832 DVSS.n3829 DVSS.n3828 0.00962857
R29833 DVSS.n8064 DVSS.n8062 0.00962857
R29834 DVSS.n8122 DVSS.n8120 0.00962857
R29835 DVSS.n8124 DVSS.n8122 0.00962857
R29836 DVSS.n8126 DVSS.n8124 0.00962857
R29837 DVSS.n8128 DVSS.n8126 0.00962857
R29838 DVSS.n8130 DVSS.n8128 0.00962857
R29839 DVSS.n8132 DVSS.n8130 0.00962857
R29840 DVSS.n8134 DVSS.n8132 0.00962857
R29841 DVSS.n8136 DVSS.n8134 0.00962857
R29842 DVSS.n8138 DVSS.n8136 0.00962857
R29843 DVSS.n8140 DVSS.n8138 0.00962857
R29844 DVSS.n8142 DVSS.n8140 0.00962857
R29845 DVSS.n8144 DVSS.n8142 0.00962857
R29846 DVSS.n8173 DVSS.n8171 0.00962857
R29847 DVSS.n8175 DVSS.n8173 0.00962857
R29848 DVSS.n8177 DVSS.n8175 0.00962857
R29849 DVSS.n8179 DVSS.n8177 0.00962857
R29850 DVSS.n8181 DVSS.n8179 0.00962857
R29851 DVSS.n8183 DVSS.n8181 0.00962857
R29852 DVSS.n8185 DVSS.n8183 0.00962857
R29853 DVSS.n8187 DVSS.n8185 0.00962857
R29854 DVSS.n8189 DVSS.n8187 0.00962857
R29855 DVSS.n8191 DVSS.n8189 0.00962857
R29856 DVSS.n8193 DVSS.n8191 0.00962857
R29857 DVSS.n8195 DVSS.n8193 0.00962857
R29858 DVSS.n8224 DVSS.n8222 0.00962857
R29859 DVSS.n8226 DVSS.n8224 0.00962857
R29860 DVSS.n8228 DVSS.n8226 0.00962857
R29861 DVSS.n8230 DVSS.n8228 0.00962857
R29862 DVSS.n8308 DVSS.n8306 0.00962857
R29863 DVSS.n8310 DVSS.n8308 0.00962857
R29864 DVSS.n8311 DVSS.n8310 0.00962857
R29865 DVSS.n3618 DVSS.n3616 0.00962857
R29866 DVSS.n2583 DVSS.n2581 0.00962857
R29867 DVSS.n2585 DVSS.n2583 0.00962857
R29868 DVSS.n2720 DVSS.n2718 0.00962857
R29869 DVSS.n2718 DVSS.n2716 0.00962857
R29870 DVSS.n2716 DVSS.n2714 0.00962857
R29871 DVSS.n2714 DVSS.n2712 0.00962857
R29872 DVSS.n2682 DVSS.n2680 0.00962857
R29873 DVSS.n2680 DVSS.n2678 0.00962857
R29874 DVSS.n2678 DVSS.n2676 0.00962857
R29875 DVSS.n2676 DVSS.n2674 0.00962857
R29876 DVSS.n2674 DVSS.n2672 0.00962857
R29877 DVSS.n2672 DVSS.n2670 0.00962857
R29878 DVSS.n2670 DVSS.n2668 0.00962857
R29879 DVSS.n2668 DVSS.n2666 0.00962857
R29880 DVSS.n2666 DVSS.n2664 0.00962857
R29881 DVSS.n2664 DVSS.n2662 0.00962857
R29882 DVSS.n2662 DVSS.n2660 0.00962857
R29883 DVSS.n2660 DVSS.n2658 0.00962857
R29884 DVSS.n2628 DVSS.n2626 0.00962857
R29885 DVSS.n2626 DVSS.n2624 0.00962857
R29886 DVSS.n2624 DVSS.n2622 0.00962857
R29887 DVSS.n2622 DVSS.n2620 0.00962857
R29888 DVSS.n2620 DVSS.n2618 0.00962857
R29889 DVSS.n2618 DVSS.n2616 0.00962857
R29890 DVSS.n2616 DVSS.n2614 0.00962857
R29891 DVSS.n2614 DVSS.n2612 0.00962857
R29892 DVSS.n2612 DVSS.n2610 0.00962857
R29893 DVSS.n2610 DVSS.n2608 0.00962857
R29894 DVSS.n11741 DVSS.n11739 0.00962857
R29895 DVSS.n11801 DVSS.n11799 0.00962857
R29896 DVSS.n11803 DVSS.n11801 0.00962857
R29897 DVSS.n11805 DVSS.n11803 0.00962857
R29898 DVSS.n11807 DVSS.n11805 0.00962857
R29899 DVSS.n11809 DVSS.n11807 0.00962857
R29900 DVSS.n11811 DVSS.n11809 0.00962857
R29901 DVSS.n11813 DVSS.n11811 0.00962857
R29902 DVSS.n11815 DVSS.n11813 0.00962857
R29903 DVSS.n11817 DVSS.n11815 0.00962857
R29904 DVSS.n11819 DVSS.n11817 0.00962857
R29905 DVSS.n11821 DVSS.n11819 0.00962857
R29906 DVSS.n11823 DVSS.n11821 0.00962857
R29907 DVSS.n11860 DVSS.n11858 0.00962857
R29908 DVSS.n11862 DVSS.n11860 0.00962857
R29909 DVSS.n11864 DVSS.n11862 0.00962857
R29910 DVSS.n11866 DVSS.n11864 0.00962857
R29911 DVSS.n11868 DVSS.n11866 0.00962857
R29912 DVSS.n11870 DVSS.n11868 0.00962857
R29913 DVSS.n11872 DVSS.n11870 0.00962857
R29914 DVSS.n11874 DVSS.n11872 0.00962857
R29915 DVSS.n11876 DVSS.n11874 0.00962857
R29916 DVSS.n11878 DVSS.n11876 0.00962857
R29917 DVSS.n11880 DVSS.n11878 0.00962857
R29918 DVSS.n11882 DVSS.n11880 0.00962857
R29919 DVSS.n11919 DVSS.n11917 0.00962857
R29920 DVSS.n11921 DVSS.n11919 0.00962857
R29921 DVSS.n11923 DVSS.n11921 0.00962857
R29922 DVSS.n11925 DVSS.n11923 0.00962857
R29923 DVSS.n12980 DVSS.n12978 0.00962857
R29924 DVSS.n12978 DVSS.n12976 0.00962857
R29925 DVSS.n12976 DVSS.n12974 0.00962857
R29926 DVSS.n6033 DVSS.n6032 0.00962857
R29927 DVSS.n5969 DVSS.n5968 0.00962857
R29928 DVSS.n5925 DVSS.n5924 0.00962857
R29929 DVSS.n8429 DVSS.n8428 0.00962857
R29930 DVSS.n8478 DVSS.n8477 0.00962857
R29931 DVSS.n8486 DVSS.n8485 0.00962857
R29932 DVSS.n11311 DVSS.n11310 0.00962857
R29933 DVSS.n6036 DVSS.n6034 0.00962857
R29934 DVSS.n6034 DVSS.n6031 0.00962857
R29935 DVSS.n6031 DVSS.n6030 0.00962857
R29936 DVSS.n6030 DVSS.n6028 0.00962857
R29937 DVSS.n6006 DVSS.n6004 0.00962857
R29938 DVSS.n6004 DVSS.n6002 0.00962857
R29939 DVSS.n6002 DVSS.n6000 0.00962857
R29940 DVSS.n6000 DVSS.n5998 0.00962857
R29941 DVSS.n5998 DVSS.n5996 0.00962857
R29942 DVSS.n5996 DVSS.n5994 0.00962857
R29943 DVSS.n5972 DVSS.n5970 0.00962857
R29944 DVSS.n5970 DVSS.n5967 0.00962857
R29945 DVSS.n5967 DVSS.n5966 0.00962857
R29946 DVSS.n5966 DVSS.n5964 0.00962857
R29947 DVSS.n5964 DVSS.n5962 0.00962857
R29948 DVSS.n5962 DVSS.n5960 0.00962857
R29949 DVSS.n5960 DVSS.n5958 0.00962857
R29950 DVSS.n5958 DVSS.n5956 0.00962857
R29951 DVSS.n5956 DVSS.n5954 0.00962857
R29952 DVSS.n5954 DVSS.n5952 0.00962857
R29953 DVSS.n5952 DVSS.n5950 0.00962857
R29954 DVSS.n5950 DVSS.n5948 0.00962857
R29955 DVSS.n5926 DVSS.n5923 0.00962857
R29956 DVSS.n5923 DVSS.n5922 0.00962857
R29957 DVSS.n5922 DVSS.n5920 0.00962857
R29958 DVSS.n5920 DVSS.n5918 0.00962857
R29959 DVSS.n5918 DVSS.n5916 0.00962857
R29960 DVSS.n8346 DVSS.n8344 0.00962857
R29961 DVSS.n8348 DVSS.n8346 0.00962857
R29962 DVSS.n8350 DVSS.n8348 0.00962857
R29963 DVSS.n8352 DVSS.n8350 0.00962857
R29964 DVSS.n8354 DVSS.n8352 0.00962857
R29965 DVSS.n8356 DVSS.n8354 0.00962857
R29966 DVSS.n8414 DVSS.n8412 0.00962857
R29967 DVSS.n8416 DVSS.n8414 0.00962857
R29968 DVSS.n8418 DVSS.n8416 0.00962857
R29969 DVSS.n8420 DVSS.n8418 0.00962857
R29970 DVSS.n8422 DVSS.n8420 0.00962857
R29971 DVSS.n8424 DVSS.n8422 0.00962857
R29972 DVSS.n8426 DVSS.n8424 0.00962857
R29973 DVSS.n8427 DVSS.n8426 0.00962857
R29974 DVSS.n8430 DVSS.n8427 0.00962857
R29975 DVSS.n8432 DVSS.n8430 0.00962857
R29976 DVSS.n8434 DVSS.n8432 0.00962857
R29977 DVSS.n8436 DVSS.n8434 0.00962857
R29978 DVSS.n8465 DVSS.n8463 0.00962857
R29979 DVSS.n8467 DVSS.n8465 0.00962857
R29980 DVSS.n8469 DVSS.n8467 0.00962857
R29981 DVSS.n8471 DVSS.n8469 0.00962857
R29982 DVSS.n8473 DVSS.n8471 0.00962857
R29983 DVSS.n8475 DVSS.n8473 0.00962857
R29984 DVSS.n8476 DVSS.n8475 0.00962857
R29985 DVSS.n8479 DVSS.n8476 0.00962857
R29986 DVSS.n8481 DVSS.n8479 0.00962857
R29987 DVSS.n8483 DVSS.n8481 0.00962857
R29988 DVSS.n8484 DVSS.n8483 0.00962857
R29989 DVSS.n8487 DVSS.n8484 0.00962857
R29990 DVSS.n8516 DVSS.n8514 0.00962857
R29991 DVSS.n8518 DVSS.n8516 0.00962857
R29992 DVSS.n8520 DVSS.n8518 0.00962857
R29993 DVSS.n8522 DVSS.n8520 0.00962857
R29994 DVSS.n11314 DVSS.n11312 0.00962857
R29995 DVSS.n11312 DVSS.n11309 0.00962857
R29996 DVSS.n11309 DVSS.n11308 0.00962857
R29997 DVSS.n6284 DVSS.n6277 0.00962857
R29998 DVSS.n6277 DVSS.n6276 0.00962857
R29999 DVSS.n6276 DVSS.n6275 0.00962857
R30000 DVSS.n6275 DVSS.n6274 0.00962857
R30001 DVSS.n6261 DVSS.n6253 0.00962857
R30002 DVSS.n6253 DVSS.n6252 0.00962857
R30003 DVSS.n6252 DVSS.n6251 0.00962857
R30004 DVSS.n6251 DVSS.n6250 0.00962857
R30005 DVSS.n6250 DVSS.n6249 0.00962857
R30006 DVSS.n6249 DVSS.n6248 0.00962857
R30007 DVSS.n6215 DVSS.n6210 0.00962857
R30008 DVSS.n6210 DVSS.n6209 0.00962857
R30009 DVSS.n6209 DVSS.n6208 0.00962857
R30010 DVSS.n6208 DVSS.n6207 0.00962857
R30011 DVSS.n6207 DVSS.n6204 0.00962857
R30012 DVSS.n6204 DVSS.n6203 0.00962857
R30013 DVSS.n6203 DVSS.n6201 0.00962857
R30014 DVSS.n6201 DVSS.n6199 0.00962857
R30015 DVSS.n6199 DVSS.n6197 0.00962857
R30016 DVSS.n6197 DVSS.n6195 0.00962857
R30017 DVSS.n6195 DVSS.n6192 0.00962857
R30018 DVSS.n6192 DVSS.n6191 0.00962857
R30019 DVSS.n6157 DVSS.n6153 0.00962857
R30020 DVSS.n6153 DVSS.n6152 0.00962857
R30021 DVSS.n6152 DVSS.n6151 0.00962857
R30022 DVSS.n6151 DVSS.n6148 0.00962857
R30023 DVSS.n6148 DVSS.n6147 0.00962857
R30024 DVSS.n8590 DVSS.n8587 0.00962857
R30025 DVSS.n8591 DVSS.n8590 0.00962857
R30026 DVSS.n8594 DVSS.n8591 0.00962857
R30027 DVSS.n8596 DVSS.n8594 0.00962857
R30028 DVSS.n8598 DVSS.n8596 0.00962857
R30029 DVSS.n8600 DVSS.n8598 0.00962857
R30030 DVSS.n8668 DVSS.n8666 0.00962857
R30031 DVSS.n8669 DVSS.n8668 0.00962857
R30032 DVSS.n8672 DVSS.n8669 0.00962857
R30033 DVSS.n8674 DVSS.n8672 0.00962857
R30034 DVSS.n8676 DVSS.n8674 0.00962857
R30035 DVSS.n8678 DVSS.n8676 0.00962857
R30036 DVSS.n8679 DVSS.n8678 0.00962857
R30037 DVSS.n8680 DVSS.n8679 0.00962857
R30038 DVSS.n8681 DVSS.n8680 0.00962857
R30039 DVSS.n8686 DVSS.n8681 0.00962857
R30040 DVSS.n8687 DVSS.n8686 0.00962857
R30041 DVSS.n8690 DVSS.n8687 0.00962857
R30042 DVSS.n8726 DVSS.n8725 0.00962857
R30043 DVSS.n8727 DVSS.n8726 0.00962857
R30044 DVSS.n8728 DVSS.n8727 0.00962857
R30045 DVSS.n8729 DVSS.n8728 0.00962857
R30046 DVSS.n8730 DVSS.n8729 0.00962857
R30047 DVSS.n8731 DVSS.n8730 0.00962857
R30048 DVSS.n8732 DVSS.n8731 0.00962857
R30049 DVSS.n8733 DVSS.n8732 0.00962857
R30050 DVSS.n8734 DVSS.n8733 0.00962857
R30051 DVSS.n8735 DVSS.n8734 0.00962857
R30052 DVSS.n8749 DVSS.n8735 0.00962857
R30053 DVSS.n8751 DVSS.n8749 0.00962857
R30054 DVSS.n8790 DVSS.n8786 0.00962857
R30055 DVSS.n8792 DVSS.n8790 0.00962857
R30056 DVSS.n8794 DVSS.n8792 0.00962857
R30057 DVSS.n8796 DVSS.n8794 0.00962857
R30058 DVSS.n8884 DVSS.n8882 0.00962857
R30059 DVSS.n8886 DVSS.n8884 0.00962857
R30060 DVSS.n8887 DVSS.n8886 0.00962857
R30061 DVSS.n6283 DVSS.n6282 0.00962857
R30062 DVSS.n6282 DVSS.n6281 0.00962857
R30063 DVSS.n6281 DVSS.n6280 0.00962857
R30064 DVSS.n6280 DVSS.n6279 0.00962857
R30065 DVSS.n6279 DVSS.n6278 0.00962857
R30066 DVSS.n6260 DVSS.n6259 0.00962857
R30067 DVSS.n6259 DVSS.n6258 0.00962857
R30068 DVSS.n6258 DVSS.n6257 0.00962857
R30069 DVSS.n6257 DVSS.n6256 0.00962857
R30070 DVSS.n6256 DVSS.n6255 0.00962857
R30071 DVSS.n6255 DVSS.n6254 0.00962857
R30072 DVSS.n6214 DVSS.n6213 0.00962857
R30073 DVSS.n6213 DVSS.n6212 0.00962857
R30074 DVSS.n6212 DVSS.n6211 0.00962857
R30075 DVSS.n6206 DVSS.n6205 0.00962857
R30076 DVSS.n6194 DVSS.n6193 0.00962857
R30077 DVSS.n6156 DVSS.n6155 0.00962857
R30078 DVSS.n6155 DVSS.n6154 0.00962857
R30079 DVSS.n6150 DVSS.n6149 0.00962857
R30080 DVSS.n8589 DVSS.n8588 0.00962857
R30081 DVSS.n8593 DVSS.n8592 0.00962857
R30082 DVSS.n8671 DVSS.n8670 0.00962857
R30083 DVSS.n8683 DVSS.n8682 0.00962857
R30084 DVSS.n8684 DVSS.n8683 0.00962857
R30085 DVSS.n8685 DVSS.n8684 0.00962857
R30086 DVSS.n8689 DVSS.n8688 0.00962857
R30087 DVSS.n8738 DVSS.n8737 0.00962857
R30088 DVSS.n8739 DVSS.n8738 0.00962857
R30089 DVSS.n8740 DVSS.n8739 0.00962857
R30090 DVSS.n8741 DVSS.n8740 0.00962857
R30091 DVSS.n8742 DVSS.n8741 0.00962857
R30092 DVSS.n8743 DVSS.n8742 0.00962857
R30093 DVSS.n8744 DVSS.n8743 0.00962857
R30094 DVSS.n8745 DVSS.n8744 0.00962857
R30095 DVSS.n8746 DVSS.n8745 0.00962857
R30096 DVSS.n8747 DVSS.n8746 0.00962857
R30097 DVSS.n8748 DVSS.n8747 0.00962857
R30098 DVSS.n8789 DVSS.n8788 0.00962857
R30099 DVSS.n11483 DVSS.n11465 0.00959676
R30100 DVSS.n11520 DVSS.n11502 0.00959676
R30101 DVSS.n11645 DVSS.n11627 0.00959676
R30102 DVSS.n11682 DVSS.n11664 0.00959676
R30103 DVSS.n11731 DVSS.n11713 0.00959676
R30104 DVSS.n20259 DVSS.n20258 0.00957614
R30105 DVSS.n20533 DVSS.n20532 0.00957614
R30106 DVSS.n19519 DVSS.n19518 0.00957614
R30107 DVSS.n19248 DVSS.n19247 0.00957614
R30108 DVSS.n20532 DVSS.n20531 0.00957614
R30109 DVSS.n20258 DVSS.n20257 0.00957614
R30110 DVSS.n2069 DVSS.n2067 0.00956429
R30111 DVSS.n1995 DVSS.n1994 0.00956429
R30112 DVSS.n172 DVSS.n171 0.00955887
R30113 DVSS.n17297 DVSS.n17296 0.00955028
R30114 DVSS.n17290 DVSS.n17288 0.00955028
R30115 DVSS.n16977 DVSS.n16975 0.00955028
R30116 DVSS.n16988 DVSS.n16987 0.00955028
R30117 DVSS.n12541 DVSS.n12540 0.00953846
R30118 DVSS.n12665 DVSS.n12664 0.00953846
R30119 DVSS.n12573 DVSS.n12572 0.00953846
R30120 DVSS.n12377 DVSS.n12376 0.00953846
R30121 DVSS.n12285 DVSS.n12284 0.00953846
R30122 DVSS.n12252 DVSS.n12251 0.00953846
R30123 DVSS.n3165 DVSS.n3164 0.00953846
R30124 DVSS.n3289 DVSS.n3288 0.00953846
R30125 DVSS.n3197 DVSS.n3196 0.00953846
R30126 DVSS.n3004 DVSS.n3003 0.00953846
R30127 DVSS.n2912 DVSS.n2911 0.00953846
R30128 DVSS.n2879 DVSS.n2878 0.00953846
R30129 DVSS.n3405 DVSS.n3404 0.00953846
R30130 DVSS.n5691 DVSS.n5690 0.00953543
R30131 DVSS.n10981 DVSS.n10980 0.00953543
R30132 DVSS.n16926 DVSS.n16925 0.00953543
R30133 DVSS.n4658 DVSS.n4657 0.00953543
R30134 DVSS.n9882 DVSS.n9881 0.00953543
R30135 DVSS.n17410 DVSS.n17409 0.00953543
R30136 DVSS.n4574 DVSS.n4573 0.00952778
R30137 DVSS.n4624 DVSS.n4623 0.00952778
R30138 DVSS.n17216 DVSS.n17215 0.0095
R30139 DVSS.n17228 DVSS.n17227 0.0095
R30140 DVSS.n15184 DVSS.n15183 0.0095
R30141 DVSS.n15147 DVSS.n15146 0.0095
R30142 DVSS.n15105 DVSS.n15104 0.0095
R30143 DVSS.n2351 DVSS.n2350 0.0095
R30144 DVSS.n2389 DVSS.n2388 0.0095
R30145 DVSS.n17694 DVSS.n17693 0.0095
R30146 DVSS.n5254 DVSS.n5253 0.00944366
R30147 DVSS.n5168 DVSS.n5167 0.00944366
R30148 DVSS.n5113 DVSS.n5112 0.00944366
R30149 DVSS.n10073 DVSS.n10072 0.00943572
R30150 DVSS.n10145 DVSS.n10144 0.00943572
R30151 DVSS.n10185 DVSS.n10184 0.00943572
R30152 DVSS.n8155 DVSS.n8154 0.00943572
R30153 DVSS.n8206 DVSS.n8205 0.00943572
R30154 DVSS.n8447 DVSS.n8446 0.00943572
R30155 DVSS.n8498 DVSS.n8497 0.00943572
R30156 DVSS.n8707 DVSS.n8706 0.00943572
R30157 DVSS.n8768 DVSS.n8767 0.00943572
R30158 DVSS.n19116 DVSS.n19107 0.00941892
R30159 DVSS.n19390 DVSS.n19379 0.00941892
R30160 DVSS.n20149 DVSS.n20148 0.00941892
R30161 DVSS.n20398 DVSS.n20384 0.00941892
R30162 DVSS.n16086 DVSS.n16085 0.00937324
R30163 DVSS.n15974 DVSS.n15973 0.00937324
R30164 DVSS.n4956 DVSS.n4955 0.00937143
R30165 DVSS.n4912 DVSS.n4911 0.00937143
R30166 DVSS.n6229 DVSS.n6228 0.00937143
R30167 DVSS.n6171 DVSS.n6170 0.00937143
R30168 DVSS.n21173 DVSS.n21172 0.0093706
R30169 DVSS.n5703 DVSS.n5702 0.00935827
R30170 DVSS.n10993 DVSS.n10992 0.00935827
R30171 DVSS.n16914 DVSS.n16913 0.00935827
R30172 DVSS.n9870 DVSS.n9869 0.00935827
R30173 DVSS.n17422 DVSS.n17421 0.00935827
R30174 DVSS.n12816 DVSS.n12800 0.00934615
R30175 DVSS.n3428 DVSS.n3412 0.00934615
R30176 DVSS.n12779 DVSS.n12778 0.00934615
R30177 DVSS.n935 DVSS.n934 0.00934615
R30178 DVSS.n21182 DVSS.n21168 0.00934615
R30179 DVSS.n931 DVSS.n930 0.00928172
R30180 DVSS.n15428 DVSS.n15427 0.009275
R30181 DVSS.n18284 DVSS.n18283 0.009275
R30182 DVSS.n18333 DVSS.n18332 0.009275
R30183 DVSS.n18342 DVSS.n18341 0.009275
R30184 DVSS.n10429 DVSS.n10428 0.00923239
R30185 DVSS.n10491 DVSS.n10490 0.00923239
R30186 DVSS.n6126 DVSS.n6125 0.00921251
R30187 DVSS.n5798 DVSS.n5797 0.0091811
R30188 DVSS.n5722 DVSS.n5721 0.0091811
R30189 DVSS.n9846 DVSS.n9845 0.0091811
R30190 DVSS.n11225 DVSS.n11224 0.0091811
R30191 DVSS.n12403 DVSS.n12402 0.0091811
R30192 DVSS.n12198 DVSS.n12197 0.0091811
R30193 DVSS.n17560 DVSS.n17559 0.0091811
R30194 DVSS.n17640 DVSS.n17639 0.0091811
R30195 DVSS.n3029 DVSS.n3028 0.0091811
R30196 DVSS.n2827 DVSS.n2826 0.0091811
R30197 DVSS.n11083 DVSS.n11082 0.0091811
R30198 DVSS.n11163 DVSS.n11162 0.0091811
R30199 DVSS.n16419 DVSS.n16418 0.0091811
R30200 DVSS.n16343 DVSS.n16342 0.0091811
R30201 DVSS.n6014 DVSS.n6013 0.00917063
R30202 DVSS.n6127 DVSS.n6126 0.00917063
R30203 DVSS.n17466 DVSS.n17465 0.00916197
R30204 DVSS.n16807 DVSS.n15873 0.00916197
R30205 DVSS.n12138 DVSS.n12137 0.00915385
R30206 DVSS.n12603 DVSS.n12602 0.00915385
R30207 DVSS.n12602 DVSS.n12601 0.00915385
R30208 DVSS.n12315 DVSS.n12314 0.00915385
R30209 DVSS.n12314 DVSS.n12313 0.00915385
R30210 DVSS.n12223 DVSS.n12222 0.00915385
R30211 DVSS.n2758 DVSS.n2757 0.00915385
R30212 DVSS.n3227 DVSS.n3226 0.00915385
R30213 DVSS.n3226 DVSS.n3225 0.00915385
R30214 DVSS.n2942 DVSS.n2941 0.00915385
R30215 DVSS.n2941 DVSS.n2940 0.00915385
R30216 DVSS.n877 DVSS.n876 0.00915385
R30217 DVSS.n14521 DVSS.n14520 0.00912168
R30218 DVSS.n16529 DVSS.n16528 0.00911913
R30219 DVSS.n18175 DVSS.n18174 0.00911913
R30220 DVSS.n14372 DVSS.n14371 0.00911913
R30221 DVSS.n14418 DVSS.n14417 0.00911913
R30222 DVSS.n14508 DVSS.n14507 0.00911913
R30223 DVSS.n19693 DVSS.n19692 0.00911913
R30224 DVSS.n19798 DVSS.n19797 0.00911913
R30225 DVSS.n19768 DVSS.n19767 0.00911913
R30226 DVSS.n149 DVSS.n148 0.00911913
R30227 DVSS.n239 DVSS.n238 0.00911913
R30228 DVSS.n209 DVSS.n208 0.00911913
R30229 DVSS.n182 DVSS.n181 0.00911913
R30230 DVSS.n14419 DVSS.n14418 0.00911913
R30231 DVSS.n18174 DVSS.n18173 0.00911913
R30232 DVSS.n16528 DVSS.n16527 0.00911913
R30233 DVSS.n14371 DVSS.n14370 0.00911913
R30234 DVSS.n16716 DVSS.n16715 0.00911913
R30235 DVSS.n15565 DVSS.n15564 0.00911913
R30236 DVSS.n14778 DVSS.n14777 0.00911913
R30237 DVSS.n14710 DVSS.n14709 0.00911913
R30238 DVSS.n14605 DVSS.n14604 0.00911913
R30239 DVSS.n19912 DVSS.n19911 0.00911913
R30240 DVSS.n20023 DVSS.n20022 0.00911913
R30241 DVSS.n19993 DVSS.n19992 0.00911913
R30242 DVSS.n309 DVSS.n308 0.00911913
R30243 DVSS.n447 DVSS.n446 0.00911913
R30244 DVSS.n417 DVSS.n416 0.00911913
R30245 DVSS.n391 DVSS.n390 0.00911913
R30246 DVSS.n14709 DVSS.n14708 0.00911913
R30247 DVSS.n15566 DVSS.n15565 0.00911913
R30248 DVSS.n16715 DVSS.n16714 0.00911913
R30249 DVSS.n14779 DVSS.n14778 0.00911913
R30250 DVSS.n19692 DVSS.n19691 0.00911913
R30251 DVSS.n19911 DVSS.n19910 0.00911913
R30252 DVSS.n14604 DVSS.n14603 0.00911913
R30253 DVSS.n14507 DVSS.n14506 0.00911913
R30254 DVSS.n20022 DVSS.n20021 0.00911913
R30255 DVSS.n19797 DVSS.n19796 0.00911913
R30256 DVSS.n19992 DVSS.n19991 0.00911913
R30257 DVSS.n19767 DVSS.n19766 0.00911913
R30258 DVSS.n310 DVSS.n309 0.00911913
R30259 DVSS.n150 DVSS.n149 0.00911913
R30260 DVSS.n390 DVSS.n389 0.00911913
R30261 DVSS.n446 DVSS.n445 0.00911913
R30262 DVSS.n238 DVSS.n237 0.00911913
R30263 DVSS.n416 DVSS.n415 0.00911913
R30264 DVSS.n208 DVSS.n207 0.00911913
R30265 DVSS.n183 DVSS.n182 0.00911913
R30266 DVSS.n14488 DVSS.n14487 0.00911702
R30267 DVSS.n14165 DVSS.n14163 0.00911702
R30268 DVSS.n14176 DVSS.n14174 0.00911702
R30269 DVSS.n14738 DVSS.n14736 0.00911702
R30270 DVSS.n14745 DVSS.n14743 0.00911702
R30271 DVSS.n4779 DVSS.n4778 0.00911429
R30272 DVSS.n4775 DVSS.n4774 0.00911429
R30273 DVSS.n8093 DVSS.n8092 0.00911429
R30274 DVSS.n8091 DVSS.n8090 0.00911429
R30275 DVSS.n11771 DVSS.n11770 0.00911429
R30276 DVSS.n11769 DVSS.n11768 0.00911429
R30277 DVSS.n8385 DVSS.n8384 0.00911429
R30278 DVSS.n8383 DVSS.n8382 0.00911429
R30279 DVSS.n8633 DVSS.n8632 0.00911429
R30280 DVSS.n8635 DVSS.n8634 0.00911429
R30281 DVSS.n5830 DVSS.n5827 0.00911111
R30282 DVSS.n5827 DVSS.n5825 0.00911111
R30283 DVSS.n5821 DVSS.n5818 0.00911111
R30284 DVSS.n5818 DVSS.n5816 0.00911111
R30285 DVSS.n5816 DVSS.n4583 0.00911111
R30286 DVSS.n5808 DVSS.n5806 0.00911111
R30287 DVSS.n5810 DVSS.n5808 0.00911111
R30288 DVSS.n17440 DVSS.n17438 0.00911111
R30289 DVSS.n17445 DVSS.n17440 0.00911111
R30290 DVSS.n17445 DVSS.n17444 0.00911111
R30291 DVSS.n16126 DVSS.n16124 0.00911111
R30292 DVSS.n17449 DVSS.n16126 0.00911111
R30293 DVSS.n17455 DVSS.n17453 0.00911111
R30294 DVSS.n17463 DVSS.n17461 0.00911111
R30295 DVSS.n17461 DVSS.n17459 0.00911111
R30296 DVSS.n17536 DVSS.n17534 0.00911111
R30297 DVSS.n17543 DVSS.n17541 0.00911111
R30298 DVSS.n17545 DVSS.n17543 0.00911111
R30299 DVSS.n17552 DVSS.n17549 0.00911111
R30300 DVSS.n16902 DVSS.n16899 0.00911111
R30301 DVSS.n16899 DVSS.n16897 0.00911111
R30302 DVSS.n16897 DVSS.n16894 0.00911111
R30303 DVSS.n16894 DVSS.n16892 0.00911111
R30304 DVSS.n11075 DVSS.n11072 0.00911111
R30305 DVSS.n11066 DVSS.n11063 0.00911111
R30306 DVSS.n11063 DVSS.n11061 0.00911111
R30307 DVSS.n11061 DVSS.n11058 0.00911111
R30308 DVSS.n11058 DVSS.n11056 0.00911111
R30309 DVSS.n11052 DVSS.n11049 0.00911111
R30310 DVSS.n11044 DVSS.n11041 0.00911111
R30311 DVSS.n11041 DVSS.n11039 0.00911111
R30312 DVSS.n11039 DVSS.n11036 0.00911111
R30313 DVSS.n11036 DVSS.n11034 0.00911111
R30314 DVSS.n2564 DVSS.n2562 0.00911111
R30315 DVSS.n2567 DVSS.n2564 0.00911111
R30316 DVSS.n2569 DVSS.n2567 0.00911111
R30317 DVSS.n4116 DVSS.n2569 0.00911111
R30318 DVSS.n4116 DVSS.n4115 0.00911111
R30319 DVSS.n4115 DVSS.n4113 0.00911111
R30320 DVSS.n4110 DVSS.n4107 0.00911111
R30321 DVSS.n4107 DVSS.n4105 0.00911111
R30322 DVSS.n4105 DVSS.n4102 0.00911111
R30323 DVSS.n4102 DVSS.n4100 0.00911111
R30324 DVSS.n4100 DVSS.n4097 0.00911111
R30325 DVSS.n4097 DVSS.n4095 0.00911111
R30326 DVSS.n7468 DVSS.n7466 0.00911111
R30327 DVSS.n18392 DVSS.n7468 0.00911111
R30328 DVSS.n18394 DVSS.n18392 0.00911111
R30329 DVSS.n18397 DVSS.n18394 0.00911111
R30330 DVSS.n18399 DVSS.n18397 0.00911111
R30331 DVSS.n18401 DVSS.n18399 0.00911111
R30332 DVSS.n18408 DVSS.n18406 0.00911111
R30333 DVSS.n18415 DVSS.n18408 0.00911111
R30334 DVSS.n18415 DVSS.n18414 0.00911111
R30335 DVSS.n18414 DVSS.n18412 0.00911111
R30336 DVSS.n15249 DVSS.n15248 0.00911111
R30337 DVSS.n15248 DVSS.n15246 0.00911111
R30338 DVSS.n15246 DVSS.n7710 0.00911111
R30339 DVSS.n14957 DVSS.n7710 0.00911111
R30340 DVSS.n14964 DVSS.n14962 0.00911111
R30341 DVSS.n14967 DVSS.n14964 0.00911111
R30342 DVSS.n14969 DVSS.n14967 0.00911111
R30343 DVSS.n14978 DVSS.n14969 0.00911111
R30344 DVSS.n14978 DVSS.n14977 0.00911111
R30345 DVSS.n14977 DVSS.n14975 0.00911111
R30346 DVSS.n9010 DVSS.n9008 0.00911111
R30347 DVSS.n9108 DVSS.n9010 0.00911111
R30348 DVSS.n9110 DVSS.n9108 0.00911111
R30349 DVSS.n9113 DVSS.n9110 0.00911111
R30350 DVSS.n9115 DVSS.n9113 0.00911111
R30351 DVSS.n9117 DVSS.n9115 0.00911111
R30352 DVSS.n9124 DVSS.n9122 0.00911111
R30353 DVSS.n9127 DVSS.n9124 0.00911111
R30354 DVSS.n9129 DVSS.n9127 0.00911111
R30355 DVSS.n9138 DVSS.n9129 0.00911111
R30356 DVSS.n9138 DVSS.n9137 0.00911111
R30357 DVSS.n9137 DVSS.n9135 0.00911111
R30358 DVSS.n2551 DVSS.n2549 0.00911111
R30359 DVSS.n2554 DVSS.n2551 0.00911111
R30360 DVSS.n2556 DVSS.n2554 0.00911111
R30361 DVSS.n4353 DVSS.n2556 0.00911111
R30362 DVSS.n4355 DVSS.n4353 0.00911111
R30363 DVSS.n4357 DVSS.n4355 0.00911111
R30364 DVSS.n4364 DVSS.n4362 0.00911111
R30365 DVSS.n4367 DVSS.n4364 0.00911111
R30366 DVSS.n4369 DVSS.n4367 0.00911111
R30367 DVSS.n4372 DVSS.n4369 0.00911111
R30368 DVSS.n4374 DVSS.n4372 0.00911111
R30369 DVSS.n4376 DVSS.n4374 0.00911111
R30370 DVSS.n7557 DVSS.n7555 0.00911111
R30371 DVSS.n18375 DVSS.n7557 0.00911111
R30372 DVSS.n18375 DVSS.n18374 0.00911111
R30373 DVSS.n18374 DVSS.n18372 0.00911111
R30374 DVSS.n18372 DVSS.n18371 0.00911111
R30375 DVSS.n18371 DVSS.n18369 0.00911111
R30376 DVSS.n18366 DVSS.n18365 0.00911111
R30377 DVSS.n18365 DVSS.n18363 0.00911111
R30378 DVSS.n18363 DVSS.n18362 0.00911111
R30379 DVSS.n18362 DVSS.n18360 0.00911111
R30380 DVSS.n7699 DVSS.n7697 0.00911111
R30381 DVSS.n15582 DVSS.n7699 0.00911111
R30382 DVSS.n15584 DVSS.n15582 0.00911111
R30383 DVSS.n15586 DVSS.n15584 0.00911111
R30384 DVSS.n15593 DVSS.n15591 0.00911111
R30385 DVSS.n15596 DVSS.n15593 0.00911111
R30386 DVSS.n15598 DVSS.n15596 0.00911111
R30387 DVSS.n15607 DVSS.n15598 0.00911111
R30388 DVSS.n15607 DVSS.n15606 0.00911111
R30389 DVSS.n15606 DVSS.n15604 0.00911111
R30390 DVSS.n8968 DVSS.n8966 0.00911111
R30391 DVSS.n9604 DVSS.n8968 0.00911111
R30392 DVSS.n9604 DVSS.n9603 0.00911111
R30393 DVSS.n9603 DVSS.n9601 0.00911111
R30394 DVSS.n9601 DVSS.n9600 0.00911111
R30395 DVSS.n9600 DVSS.n9598 0.00911111
R30396 DVSS.n9595 DVSS.n9594 0.00911111
R30397 DVSS.n9594 DVSS.n9592 0.00911111
R30398 DVSS.n9592 DVSS.n9591 0.00911111
R30399 DVSS.n9591 DVSS.n9589 0.00911111
R30400 DVSS.n9589 DVSS.n8985 0.00911111
R30401 DVSS.n8985 DVSS.n8983 0.00911111
R30402 DVSS.n6566 DVSS.n6556 0.00911111
R30403 DVSS.n6556 DVSS.n6554 0.00911111
R30404 DVSS.n6551 DVSS.n6548 0.00911111
R30405 DVSS.n6548 DVSS.n6546 0.00911111
R30406 DVSS.n6546 DVSS.n6543 0.00911111
R30407 DVSS.n6543 DVSS.n6541 0.00911111
R30408 DVSS.n6541 DVSS.n6538 0.00911111
R30409 DVSS.n6538 DVSS.n6536 0.00911111
R30410 DVSS.n16229 DVSS.n16227 0.00911111
R30411 DVSS.n16246 DVSS.n16229 0.00911111
R30412 DVSS.n16246 DVSS.n16245 0.00911111
R30413 DVSS.n16245 DVSS.n16243 0.00911111
R30414 DVSS.n16243 DVSS.n16242 0.00911111
R30415 DVSS.n16242 DVSS.n16240 0.00911111
R30416 DVSS.n16237 DVSS.n7614 0.00911111
R30417 DVSS.n18084 DVSS.n7614 0.00911111
R30418 DVSS.n18084 DVSS.n18083 0.00911111
R30419 DVSS.n18083 DVSS.n18081 0.00911111
R30420 DVSS.n7678 DVSS.n7676 0.00911111
R30421 DVSS.n15733 DVSS.n7678 0.00911111
R30422 DVSS.n15733 DVSS.n15732 0.00911111
R30423 DVSS.n15732 DVSS.n15730 0.00911111
R30424 DVSS.n15727 DVSS.n15726 0.00911111
R30425 DVSS.n15726 DVSS.n15724 0.00911111
R30426 DVSS.n15724 DVSS.n15723 0.00911111
R30427 DVSS.n15723 DVSS.n15721 0.00911111
R30428 DVSS.n15721 DVSS.n7693 0.00911111
R30429 DVSS.n7693 DVSS.n7691 0.00911111
R30430 DVSS.n8960 DVSS.n8958 0.00911111
R30431 DVSS.n9720 DVSS.n8960 0.00911111
R30432 DVSS.n9722 DVSS.n9720 0.00911111
R30433 DVSS.n9725 DVSS.n9722 0.00911111
R30434 DVSS.n9727 DVSS.n9725 0.00911111
R30435 DVSS.n9729 DVSS.n9727 0.00911111
R30436 DVSS.n9736 DVSS.n9734 0.00911111
R30437 DVSS.n9739 DVSS.n9736 0.00911111
R30438 DVSS.n9741 DVSS.n9739 0.00911111
R30439 DVSS.n9750 DVSS.n9741 0.00911111
R30440 DVSS.n9750 DVSS.n9749 0.00911111
R30441 DVSS.n9749 DVSS.n9747 0.00911111
R30442 DVSS.n6481 DVSS.n6479 0.00911111
R30443 DVSS.n6483 DVSS.n6481 0.00911111
R30444 DVSS.n6502 DVSS.n6501 0.00911111
R30445 DVSS.n6501 DVSS.n6499 0.00911111
R30446 DVSS.n6499 DVSS.n6498 0.00911111
R30447 DVSS.n6498 DVSS.n6496 0.00911111
R30448 DVSS.n6496 DVSS.n6495 0.00911111
R30449 DVSS.n6495 DVSS.n6493 0.00911111
R30450 DVSS.n16312 DVSS.n16310 0.00911111
R30451 DVSS.n16322 DVSS.n16312 0.00911111
R30452 DVSS.n16322 DVSS.n16319 0.00911111
R30453 DVSS.n16319 DVSS.n16317 0.00911111
R30454 DVSS.n16317 DVSS.n16314 0.00911111
R30455 DVSS.n16336 DVSS.n16333 0.00911111
R30456 DVSS.n16333 DVSS.n7634 0.00911111
R30457 DVSS.n7634 DVSS.n7633 0.00911111
R30458 DVSS.n7633 DVSS.n7631 0.00911111
R30459 DVSS.n17675 DVSS.n7653 0.00911111
R30460 DVSS.n7653 DVSS.n7651 0.00911111
R30461 DVSS.n7651 DVSS.n7650 0.00911111
R30462 DVSS.n17659 DVSS.n17656 0.00911111
R30463 DVSS.n17656 DVSS.n17654 0.00911111
R30464 DVSS.n17654 DVSS.n7664 0.00911111
R30465 DVSS.n7664 DVSS.n7662 0.00911111
R30466 DVSS.n7662 DVSS.n7661 0.00911111
R30467 DVSS.n9821 DVSS.n9819 0.00911111
R30468 DVSS.n9831 DVSS.n9821 0.00911111
R30469 DVSS.n9831 DVSS.n9830 0.00911111
R30470 DVSS.n9830 DVSS.n9828 0.00911111
R30471 DVSS.n9828 DVSS.n9827 0.00911111
R30472 DVSS.n11172 DVSS.n11170 0.00911111
R30473 DVSS.n11214 DVSS.n11172 0.00911111
R30474 DVSS.n11214 DVSS.n11211 0.00911111
R30475 DVSS.n11211 DVSS.n11209 0.00911111
R30476 DVSS.n11209 DVSS.n11208 0.00911111
R30477 DVSS.n11208 DVSS.n11206 0.00911111
R30478 DVSS.n6430 DVSS.n6420 0.00911111
R30479 DVSS.n6420 DVSS.n6418 0.00911111
R30480 DVSS.n6415 DVSS.n6412 0.00911111
R30481 DVSS.n6412 DVSS.n6410 0.00911111
R30482 DVSS.n6410 DVSS.n6407 0.00911111
R30483 DVSS.n6407 DVSS.n4477 0.00911111
R30484 DVSS.n4477 DVSS.n4474 0.00911111
R30485 DVSS.n4474 DVSS.n4472 0.00911111
R30486 DVSS.n16268 DVSS.n16266 0.00911111
R30487 DVSS.n16285 DVSS.n16268 0.00911111
R30488 DVSS.n16285 DVSS.n16284 0.00911111
R30489 DVSS.n16284 DVSS.n16282 0.00911111
R30490 DVSS.n16282 DVSS.n16281 0.00911111
R30491 DVSS.n16281 DVSS.n16279 0.00911111
R30492 DVSS.n16276 DVSS.n7622 0.00911111
R30493 DVSS.n17943 DVSS.n7622 0.00911111
R30494 DVSS.n17943 DVSS.n17942 0.00911111
R30495 DVSS.n17942 DVSS.n17940 0.00911111
R30496 DVSS.n7670 DVSS.n7668 0.00911111
R30497 DVSS.n15828 DVSS.n7670 0.00911111
R30498 DVSS.n15830 DVSS.n15828 0.00911111
R30499 DVSS.n15832 DVSS.n15830 0.00911111
R30500 DVSS.n15839 DVSS.n15837 0.00911111
R30501 DVSS.n15842 DVSS.n15839 0.00911111
R30502 DVSS.n15844 DVSS.n15842 0.00911111
R30503 DVSS.n15853 DVSS.n15844 0.00911111
R30504 DVSS.n15853 DVSS.n15852 0.00911111
R30505 DVSS.n15852 DVSS.n15850 0.00911111
R30506 DVSS.n8935 DVSS.n8933 0.00911111
R30507 DVSS.n9796 DVSS.n8935 0.00911111
R30508 DVSS.n9796 DVSS.n9795 0.00911111
R30509 DVSS.n9795 DVSS.n9793 0.00911111
R30510 DVSS.n9793 DVSS.n9792 0.00911111
R30511 DVSS.n9792 DVSS.n9790 0.00911111
R30512 DVSS.n9787 DVSS.n9786 0.00911111
R30513 DVSS.n9786 DVSS.n9784 0.00911111
R30514 DVSS.n9784 DVSS.n9783 0.00911111
R30515 DVSS.n9783 DVSS.n9781 0.00911111
R30516 DVSS.n9781 DVSS.n8952 0.00911111
R30517 DVSS.n8952 DVSS.n8950 0.00911111
R30518 DVSS.n2579 DVSS.n2577 0.00911111
R30519 DVSS.n4004 DVSS.n2579 0.00911111
R30520 DVSS.n4006 DVSS.n4004 0.00911111
R30521 DVSS.n4009 DVSS.n4006 0.00911111
R30522 DVSS.n4011 DVSS.n4009 0.00911111
R30523 DVSS.n4013 DVSS.n4011 0.00911111
R30524 DVSS.n4020 DVSS.n4018 0.00911111
R30525 DVSS.n4023 DVSS.n4020 0.00911111
R30526 DVSS.n4025 DVSS.n4023 0.00911111
R30527 DVSS.n4032 DVSS.n4025 0.00911111
R30528 DVSS.n4032 DVSS.n4031 0.00911111
R30529 DVSS.n4031 DVSS.n4029 0.00911111
R30530 DVSS.n7478 DVSS.n7476 0.00911111
R30531 DVSS.n7497 DVSS.n7478 0.00911111
R30532 DVSS.n7497 DVSS.n7496 0.00911111
R30533 DVSS.n7496 DVSS.n7494 0.00911111
R30534 DVSS.n7494 DVSS.n7493 0.00911111
R30535 DVSS.n7493 DVSS.n7491 0.00911111
R30536 DVSS.n7488 DVSS.n7487 0.00911111
R30537 DVSS.n7487 DVSS.n7458 0.00911111
R30538 DVSS.n7458 DVSS.n7457 0.00911111
R30539 DVSS.n7457 DVSS.n7455 0.00911111
R30540 DVSS.n15060 DVSS.n15059 0.00911111
R30541 DVSS.n15059 DVSS.n15057 0.00911111
R30542 DVSS.n15057 DVSS.n15056 0.00911111
R30543 DVSS.n15056 DVSS.n15054 0.00911111
R30544 DVSS.n15051 DVSS.n15050 0.00911111
R30545 DVSS.n15050 DVSS.n15048 0.00911111
R30546 DVSS.n15048 DVSS.n15047 0.00911111
R30547 DVSS.n15047 DVSS.n15045 0.00911111
R30548 DVSS.n15045 DVSS.n7783 0.00911111
R30549 DVSS.n7783 DVSS.n7781 0.00911111
R30550 DVSS.n9015 DVSS.n9013 0.00911111
R30551 DVSS.n9039 DVSS.n9015 0.00911111
R30552 DVSS.n9039 DVSS.n9038 0.00911111
R30553 DVSS.n9038 DVSS.n9036 0.00911111
R30554 DVSS.n9036 DVSS.n9035 0.00911111
R30555 DVSS.n9035 DVSS.n9033 0.00911111
R30556 DVSS.n9030 DVSS.n9029 0.00911111
R30557 DVSS.n9029 DVSS.n9027 0.00911111
R30558 DVSS.n9027 DVSS.n9026 0.00911111
R30559 DVSS.n9026 DVSS.n8059 0.00911111
R30560 DVSS.n8059 DVSS.n8058 0.00911111
R30561 DVSS.n8058 DVSS.n8056 0.00911111
R30562 DVSS.n5522 DVSS.n5520 0.00911111
R30563 DVSS.n5525 DVSS.n5522 0.00911111
R30564 DVSS.n5527 DVSS.n5525 0.00911111
R30565 DVSS.n5530 DVSS.n5527 0.00911111
R30566 DVSS.n5532 DVSS.n5530 0.00911111
R30567 DVSS.n5534 DVSS.n5532 0.00911111
R30568 DVSS.n5553 DVSS.n5551 0.00911111
R30569 DVSS.n5551 DVSS.n5549 0.00911111
R30570 DVSS.n5549 DVSS.n5548 0.00911111
R30571 DVSS.n5548 DVSS.n5546 0.00911111
R30572 DVSS.n5546 DVSS.n5545 0.00911111
R30573 DVSS.n5545 DVSS.n5543 0.00911111
R30574 DVSS.n16432 DVSS.n16430 0.00911111
R30575 DVSS.n16435 DVSS.n16432 0.00911111
R30576 DVSS.n16437 DVSS.n16435 0.00911111
R30577 DVSS.n16440 DVSS.n16437 0.00911111
R30578 DVSS.n16442 DVSS.n16440 0.00911111
R30579 DVSS.n17248 DVSS.n16442 0.00911111
R30580 DVSS.n17244 DVSS.n17243 0.00911111
R30581 DVSS.n17243 DVSS.n17241 0.00911111
R30582 DVSS.n17241 DVSS.n17238 0.00911111
R30583 DVSS.n17238 DVSS.n17236 0.00911111
R30584 DVSS.n16872 DVSS.n16870 0.00911111
R30585 DVSS.n17113 DVSS.n16872 0.00911111
R30586 DVSS.n17113 DVSS.n17110 0.00911111
R30587 DVSS.n17110 DVSS.n17108 0.00911111
R30588 DVSS.n17105 DVSS.n17104 0.00911111
R30589 DVSS.n17104 DVSS.n17102 0.00911111
R30590 DVSS.n17102 DVSS.n16888 0.00911111
R30591 DVSS.n16888 DVSS.n16886 0.00911111
R30592 DVSS.n16886 DVSS.n16883 0.00911111
R30593 DVSS.n16883 DVSS.n16881 0.00911111
R30594 DVSS.n9858 DVSS.n9856 0.00911111
R30595 DVSS.n9991 DVSS.n9858 0.00911111
R30596 DVSS.n9993 DVSS.n9991 0.00911111
R30597 DVSS.n9996 DVSS.n9993 0.00911111
R30598 DVSS.n9998 DVSS.n9996 0.00911111
R30599 DVSS.n10000 DVSS.n9998 0.00911111
R30600 DVSS.n10006 DVSS.n10004 0.00911111
R30601 DVSS.n10053 DVSS.n10006 0.00911111
R30602 DVSS.n10053 DVSS.n10052 0.00911111
R30603 DVSS.n10052 DVSS.n10050 0.00911111
R30604 DVSS.n10050 DVSS.n10047 0.00911111
R30605 DVSS.n10047 DVSS.n10045 0.00911111
R30606 DVSS.n16805 DVSS.n16804 0.0090896
R30607 DVSS.n7643 DVSS.n7642 0.0090896
R30608 DVSS.n19744 DVSS.n19743 0.00905176
R30609 DVSS.n19969 DVSS.n19968 0.00905176
R30610 DVSS.n7720 DVSS.n7719 0.00905
R30611 DVSS.n16051 DVSS.n16050 0.00905
R30612 DVSS.n5400 DVSS.n5398 0.00904749
R30613 DVSS.n10262 DVSS.n10261 0.00904749
R30614 DVSS.n5587 DVSS.n5586 0.00900394
R30615 DVSS.n10271 DVSS.n10270 0.00900394
R30616 DVSS.n17010 DVSS.n17009 0.00900394
R30617 DVSS.n10631 DVSS.n10630 0.00900394
R30618 DVSS.n5226 DVSS.n5225 0.00900394
R30619 DVSS.n9914 DVSS.n9913 0.00900394
R30620 DVSS.n17305 DVSS.n17304 0.00900394
R30621 DVSS.n5390 DVSS.n5389 0.00900394
R30622 DVSS.n18485 DVSS.n18484 0.0089507
R30623 DVSS.n15117 DVSS.n7711 0.0089507
R30624 DVSS.n6013 DVSS.n6012 0.00885505
R30625 DVSS.n6128 DVSS.n6127 0.00885505
R30626 DVSS.n5683 DVSS.n5682 0.00882677
R30627 DVSS.n5794 DVSS.n5793 0.00882677
R30628 DVSS.n10974 DVSS.n10973 0.00882677
R30629 DVSS.n9842 DVSS.n9841 0.00882677
R30630 DVSS.n16933 DVSS.n16932 0.00882677
R30631 DVSS.n17564 DVSS.n17563 0.00882677
R30632 DVSS.n10806 DVSS.n10805 0.00882677
R30633 DVSS.n4666 DVSS.n4665 0.00882677
R30634 DVSS.n9889 DVSS.n9888 0.00882677
R30635 DVSS.n11087 DVSS.n11086 0.00882677
R30636 DVSS.n17402 DVSS.n17401 0.00882677
R30637 DVSS.n16415 DVSS.n16414 0.00882677
R30638 DVSS.n5457 DVSS.n5456 0.00882677
R30639 DVSS.n16598 DVSS.n16597 0.008825
R30640 DVSS.n16605 DVSS.n16604 0.008825
R30641 DVSS.n18311 DVSS.n18310 0.008825
R30642 DVSS.n18318 DVSS.n18317 0.008825
R30643 DVSS.n14618 DVSS.n14617 0.00878984
R30644 DVSS.n6139 DVSS.n6138 0.0087865
R30645 DVSS.n6133 DVSS.n6132 0.0087865
R30646 DVSS.n6119 DVSS.n6118 0.0087865
R30647 DVSS.n6113 DVSS.n6112 0.0087865
R30648 DVSS.n12540 DVSS.n12539 0.00876923
R30649 DVSS.n12664 DVSS.n12663 0.00876923
R30650 DVSS.n12572 DVSS.n12571 0.00876923
R30651 DVSS.n12376 DVSS.n12375 0.00876923
R30652 DVSS.n12284 DVSS.n12283 0.00876923
R30653 DVSS.n12253 DVSS.n12252 0.00876923
R30654 DVSS.n3164 DVSS.n3163 0.00876923
R30655 DVSS.n3288 DVSS.n3287 0.00876923
R30656 DVSS.n3196 DVSS.n3195 0.00876923
R30657 DVSS.n3003 DVSS.n3002 0.00876923
R30658 DVSS.n2911 DVSS.n2910 0.00876923
R30659 DVSS.n2880 DVSS.n2879 0.00876923
R30660 DVSS.n5707 DVSS.n5706 0.00864961
R30661 DVSS.n10997 DVSS.n10996 0.00864961
R30662 DVSS.n12412 DVSS.n12411 0.00864961
R30663 DVSS.n16910 DVSS.n16909 0.00864961
R30664 DVSS.n3039 DVSS.n3038 0.00864961
R30665 DVSS.n9866 DVSS.n9865 0.00864961
R30666 DVSS.n17426 DVSS.n17425 0.00864961
R30667 DVSS.n7713 DVSS.n7712 0.0086
R30668 DVSS.n16095 DVSS.n16094 0.0086
R30669 DVSS.n16044 DVSS.n16043 0.0086
R30670 DVSS.n9964 DVSS.n9963 0.00857235
R30671 DVSS.n17368 DVSS.n17367 0.00857235
R30672 DVSS.n5377 DVSS.n5376 0.00854469
R30673 DVSS.n5373 DVSS.n5371 0.00854469
R30674 DVSS.n5594 DVSS.n5592 0.00854469
R30675 DVSS.n5597 DVSS.n5595 0.00854469
R30676 DVSS.n17312 DVSS.n17310 0.00854469
R30677 DVSS.n17315 DVSS.n17313 0.00854469
R30678 DVSS.n17017 DVSS.n17015 0.00854469
R30679 DVSS.n10227 DVSS.n10225 0.00854469
R30680 DVSS.n10233 DVSS.n10232 0.00854469
R30681 DVSS.n10278 DVSS.n10276 0.00854469
R30682 DVSS DVSS.n10589 0.00852817
R30683 DVSS.n10584 DVSS 0.00852817
R30684 DVSS.n979 DVSS.n978 0.00851368
R30685 DVSS.n20967 DVSS.n20966 0.00851368
R30686 DVSS.n14916 DVSS.n14883 0.0084922
R30687 DVSS.n6015 DVSS.n6014 0.00848752
R30688 DVSS.n21127 DVSS.n21126 0.00847244
R30689 DVSS.n798 DVSS.n797 0.00847244
R30690 DVSS.n2425 DVSS.n2424 0.00847143
R30691 DVSS.n10106 DVSS.n10105 0.00847143
R30692 DVSS.n10160 DVSS.n10159 0.00847143
R30693 DVSS.n10650 DVSS.n10649 0.00847143
R30694 DVSS.n8170 DVSS.n8169 0.00847143
R30695 DVSS.n8221 DVSS.n8220 0.00847143
R30696 DVSS.n11857 DVSS.n11856 0.00847143
R30697 DVSS.n11916 DVSS.n11915 0.00847143
R30698 DVSS.n8462 DVSS.n8461 0.00847143
R30699 DVSS.n8513 DVSS.n8512 0.00847143
R30700 DVSS.n8737 DVSS.n8736 0.00847143
R30701 DVSS.n8788 DVSS.n8787 0.00847143
R30702 DVSS.n8329 DVSS.n8328 0.00847143
R30703 DVSS.n12503 DVSS.n12502 0.00838462
R30704 DVSS.n12510 DVSS.n12509 0.00838462
R30705 DVSS.n12634 DVSS.n12633 0.00838462
R30706 DVSS.n12627 DVSS.n12626 0.00838462
R30707 DVSS.n12346 DVSS.n12345 0.00838462
R30708 DVSS.n12339 DVSS.n12338 0.00838462
R30709 DVSS.n21220 DVSS.n21219 0.00838462
R30710 DVSS.n3127 DVSS.n3126 0.00838462
R30711 DVSS.n3134 DVSS.n3133 0.00838462
R30712 DVSS.n3258 DVSS.n3257 0.00838462
R30713 DVSS.n3251 DVSS.n3250 0.00838462
R30714 DVSS.n2973 DVSS.n2972 0.00838462
R30715 DVSS.n2966 DVSS.n2965 0.00838462
R30716 DVSS.n901 DVSS.n900 0.00838462
R30717 DVSS.n908 DVSS.n907 0.00838462
R30718 DVSS.n3394 DVSS.n3393 0.00838462
R30719 DVSS.n3412 DVSS.n3411 0.00838462
R30720 DVSS.n12800 DVSS.n12792 0.00838462
R30721 DVSS.n12799 DVSS.n12798 0.00838462
R30722 DVSS.n15435 DVSS.n15434 0.008375
R30723 DVSS.n18277 DVSS.n18276 0.008375
R30724 DVSS.n18326 DVSS.n18325 0.008375
R30725 DVSS.n18349 DVSS.n18348 0.008375
R30726 DVSS.n18484 DVSS.n18483 0.0083169
R30727 DVSS.n15118 DVSS.n15117 0.0083169
R30728 DVSS.n3991 DVSS.n3990 0.00829908
R30729 DVSS.n20966 DVSS.n20965 0.00829908
R30730 DVSS.n20954 DVSS.n20953 0.00829908
R30731 DVSS.n9808 DVSS.n9807 0.00829908
R30732 DVSS.n9707 DVSS.n9706 0.00829908
R30733 DVSS.n9616 DVSS.n9615 0.00829908
R30734 DVSS.n9095 DVSS.n9094 0.00829908
R30735 DVSS.n9051 DVSS.n9050 0.00829908
R30736 DVSS.n16297 DVSS.n16296 0.00829908
R30737 DVSS.n16258 DVSS.n16257 0.00829908
R30738 DVSS.n16137 DVSS.n16136 0.00829908
R30739 DVSS.n18379 DVSS.n18378 0.00829908
R30740 DVSS.n7509 DVSS.n7508 0.00829908
R30741 DVSS.n11439 DVSS.n11438 0.00829528
R30742 DVSS.n6460 DVSS.n6459 0.00829528
R30743 DVSS.n17873 DVSS.n7620 0.00828229
R30744 DVSS.n18014 DVSS.n7612 0.00828229
R30745 DVSS.n18160 DVSS.n18159 0.00828229
R30746 DVSS.n7565 DVSS.n7459 0.00828229
R30747 DVSS.n15826 DVSS.n15825 0.00828229
R30748 DVSS.n15736 DVSS.n15735 0.00828229
R30749 DVSS.n15580 DVSS.n15579 0.00828229
R30750 DVSS.n15244 DVSS.n15243 0.00828229
R30751 DVSS.n18523 DVSS.n18522 0.00828229
R30752 DVSS.n7764 DVSS.n7763 0.00828229
R30753 DVSS.n6965 DVSS.n6964 0.00825207
R30754 DVSS.n7118 DVSS.n7117 0.00825207
R30755 DVSS.n7136 DVSS.n7135 0.00825207
R30756 DVSS.n13834 DVSS.n13833 0.00825207
R30757 DVSS.n13823 DVSS.n13822 0.00825207
R30758 DVSS.n13796 DVSS.n13795 0.00825207
R30759 DVSS.n13785 DVSS.n13784 0.00825207
R30760 DVSS.n13759 DVSS.n13758 0.00825207
R30761 DVSS.n13748 DVSS.n13747 0.00825207
R30762 DVSS.n13711 DVSS.n13710 0.00825207
R30763 DVSS.n13700 DVSS.n13699 0.00825207
R30764 DVSS.n13679 DVSS.n13678 0.00825207
R30765 DVSS.n13563 DVSS.n13562 0.00825207
R30766 DVSS.n13557 DVSS.n13556 0.00825207
R30767 DVSS.n13701 DVSS.n13700 0.00825207
R30768 DVSS.n13797 DVSS.n13796 0.00825207
R30769 DVSS.n13786 DVSS.n13785 0.00825207
R30770 DVSS.n13760 DVSS.n13759 0.00825207
R30771 DVSS.n13749 DVSS.n13748 0.00825207
R30772 DVSS.n13712 DVSS.n13711 0.00825207
R30773 DVSS.n13824 DVSS.n13823 0.00825207
R30774 DVSS.n13835 DVSS.n13834 0.00825207
R30775 DVSS.n7135 DVSS.n7134 0.00825207
R30776 DVSS.n13558 DVSS.n13557 0.00825207
R30777 DVSS.n7117 DVSS.n7116 0.00825207
R30778 DVSS.n13564 DVSS.n13563 0.00825207
R30779 DVSS.n6964 DVSS.n6963 0.00825207
R30780 DVSS.n13680 DVSS.n13679 0.00825207
R30781 DVSS.n13200 DVSS.n13199 0.00825207
R30782 DVSS.n13269 DVSS.n13268 0.00825207
R30783 DVSS.n13357 DVSS.n13356 0.00825207
R30784 DVSS.n13199 DVSS.n13192 0.00825207
R30785 DVSS.n13356 DVSS.n13355 0.00825207
R30786 DVSS.n13268 DVSS.n13267 0.00825207
R30787 DVSS.n18590 DVSS.n18589 0.00825207
R30788 DVSS.n18609 DVSS.n18608 0.00825207
R30789 DVSS.n18625 DVSS.n18624 0.00825207
R30790 DVSS.n18636 DVSS.n18635 0.00825207
R30791 DVSS.n18652 DVSS.n18651 0.00825207
R30792 DVSS.n18663 DVSS.n18662 0.00825207
R30793 DVSS.n18684 DVSS.n18683 0.00825207
R30794 DVSS.n18694 DVSS.n18693 0.00825207
R30795 DVSS.n18716 DVSS.n18715 0.00825207
R30796 DVSS.n18797 DVSS.n18796 0.00825207
R30797 DVSS.n18818 DVSS.n18817 0.00825207
R30798 DVSS.n18695 DVSS.n18694 0.00825207
R30799 DVSS.n18624 DVSS.n18623 0.00825207
R30800 DVSS.n18635 DVSS.n18634 0.00825207
R30801 DVSS.n18651 DVSS.n18650 0.00825207
R30802 DVSS.n18662 DVSS.n18661 0.00825207
R30803 DVSS.n18683 DVSS.n18682 0.00825207
R30804 DVSS.n18608 DVSS.n18607 0.00825207
R30805 DVSS.n18589 DVSS.n18584 0.00825207
R30806 DVSS.n18715 DVSS.n18710 0.00825207
R30807 DVSS.n18817 DVSS.n18816 0.00825207
R30808 DVSS.n18796 DVSS.n18795 0.00825207
R30809 DVSS.n10942 DVSS.n10941 0.00824041
R30810 DVSS.n17075 DVSS.n17074 0.00824041
R30811 DVSS.n4719 DVSS.n4718 0.00824041
R30812 DVSS.n5649 DVSS.n5648 0.0082404
R30813 DVSS.n20741 DVSS.n20740 0.00818173
R30814 DVSS.n1195 DVSS.n1194 0.00818173
R30815 DVSS.n10307 DVSS.n10306 0.00817606
R30816 DVSS.n14213 DVSS.n7451 0.00816024
R30817 DVSS.n7191 DVSS.n7189 0.00815957
R30818 DVSS.n7305 DVSS.n7304 0.00815957
R30819 DVSS.n18853 DVSS.n18851 0.00815957
R30820 DVSS.n7886 DVSS.n7884 0.00815957
R30821 DVSS.n13397 DVSS.n13395 0.00815957
R30822 DVSS.n7042 DVSS.n7040 0.00815957
R30823 DVSS.n7082 DVSS.n7080 0.00815957
R30824 DVSS.n7058 DVSS.n7057 0.00815957
R30825 DVSS.n7054 DVSS.n7052 0.00815957
R30826 DVSS.n13616 DVSS.n13613 0.00815957
R30827 DVSS.n13636 DVSS.n13633 0.00815957
R30828 DVSS.n13305 DVSS.n13303 0.00815957
R30829 DVSS.n13310 DVSS.n13309 0.00815957
R30830 DVSS.n17209 DVSS.n17208 0.00815
R30831 DVSS.n15154 DVSS.n15153 0.00815
R30832 DVSS.n15115 DVSS.n15111 0.00815
R30833 DVSS.n17687 DVSS.n17686 0.00815
R30834 DVSS.n12817 DVSS.n12777 0.00811811
R30835 DVSS.n3429 DVSS.n3389 0.00811811
R30836 DVSS.n10369 DVSS.n10368 0.00803521
R30837 DVSS.n11026 DVSS.n11024 0.008
R30838 DVSS.n6769 DVSS.n6764 0.008
R30839 DVSS.n11662 DVSS.n11660 0.008
R30840 DVSS.n11664 DVSS.n11662 0.008
R30841 DVSS.n6714 DVSS.n6709 0.008
R30842 DVSS.n11625 DVSS.n11623 0.008
R30843 DVSS.n11627 DVSS.n11625 0.008
R30844 DVSS.n6571 DVSS.n2541 0.008
R30845 DVSS.n11500 DVSS.n11498 0.008
R30846 DVSS.n11502 DVSS.n11500 0.008
R30847 DVSS.n11197 DVSS.n11195 0.008
R30848 DVSS.n6435 DVSS.n6402 0.008
R30849 DVSS.n11463 DVSS.n11461 0.008
R30850 DVSS.n11465 DVSS.n11463 0.008
R30851 DVSS.n12533 DVSS.n12532 0.008
R30852 DVSS.n12657 DVSS.n12656 0.008
R30853 DVSS.n12565 DVSS.n12564 0.008
R30854 DVSS.n12369 DVSS.n12368 0.008
R30855 DVSS.n12277 DVSS.n12276 0.008
R30856 DVSS.n12260 DVSS.n12259 0.008
R30857 DVSS.n6896 DVSS.n6891 0.008
R30858 DVSS.n11711 DVSS.n11709 0.008
R30859 DVSS.n11713 DVSS.n11711 0.008
R30860 DVSS.n10037 DVSS.n10035 0.008
R30861 DVSS.n3157 DVSS.n3156 0.008
R30862 DVSS.n3281 DVSS.n3280 0.008
R30863 DVSS.n3189 DVSS.n3188 0.008
R30864 DVSS.n2996 DVSS.n2995 0.008
R30865 DVSS.n2904 DVSS.n2903 0.008
R30866 DVSS.n2887 DVSS.n2886 0.008
R30867 DVSS.n10062 DVSS.n10061 0.00795714
R30868 DVSS.n12470 DVSS.n12469 0.00794094
R30869 DVSS.n3096 DVSS.n3095 0.00794094
R30870 DVSS.n15399 DVSS.n15398 0.007925
R30871 DVSS.n18292 DVSS.n18291 0.007925
R30872 DVSS.n18306 DVSS.n18305 0.007925
R30873 DVSS.n5241 DVSS.n5240 0.00789437
R30874 DVSS.n5158 DVSS.n5157 0.00789437
R30875 DVSS.n5104 DVSS.n5103 0.00789437
R30876 DVSS.n10320 DVSS.n10319 0.00789437
R30877 DVSS.n10352 DVSS.n10351 0.00789437
R30878 DVSS.n10360 DVSS.n10359 0.00789437
R30879 DVSS.n10419 DVSS.n10418 0.00789437
R30880 DVSS.n10478 DVSS.n10477 0.00789437
R30881 DVSS.n7214 DVSS.n7213 0.00786815
R30882 DVSS.n13517 DVSS.n13516 0.00786815
R30883 DVSS.n13419 DVSS.n13418 0.00786815
R30884 DVSS.n18874 DVSS.n18873 0.00786815
R30885 DVSS.n4579 DVSS.n4577 0.00786111
R30886 DVSS.n6764 DVSS.n6762 0.00786111
R30887 DVSS.n6709 DVSS.n6707 0.00786111
R30888 DVSS.n2541 DVSS.n2539 0.00786111
R30889 DVSS.n4525 DVSS.n4523 0.00786111
R30890 DVSS.n6402 DVSS.n6400 0.00786111
R30891 DVSS.n6891 DVSS.n6889 0.00786111
R30892 DVSS.n5509 DVSS.n5507 0.00786111
R30893 DVSS.n1710 VSS 0.00782857
R30894 DVSS.n2238 VSS 0.00782857
R30895 VSS DVSS.n2239 0.00782857
R30896 VSS DVSS.n1711 0.00782857
R30897 DVSS DVSS.n10715 0.00782857
R30898 DVSS.n10714 DVSS 0.00782857
R30899 DVSS DVSS.n8312 0.00782857
R30900 DVSS.n8311 DVSS 0.00782857
R30901 DVSS.n12973 DVSS 0.00782857
R30902 DVSS.n12974 DVSS 0.00782857
R30903 DVSS.n11307 DVSS 0.00782857
R30904 DVSS.n11308 DVSS 0.00782857
R30905 DVSS.n8887 DVSS 0.00782857
R30906 DVSS DVSS.n8888 0.00782857
R30907 DVSS.n10198 DVSS.n10197 0.00781054
R30908 DVSS.n10915 DVSS.n10914 0.00781054
R30909 DVSS.n10928 DVSS.n10927 0.00781054
R30910 DVSS.n11285 DVSS.n11284 0.00781054
R30911 DVSS.n11271 DVSS.n11270 0.00781054
R30912 DVSS.n9517 DVSS.n9516 0.00781054
R30913 DVSS.n9546 DVSS.n9545 0.00781054
R30914 DVSS.n9573 DVSS.n9572 0.00781054
R30915 DVSS.n8998 DVSS.n8997 0.00781054
R30916 DVSS.n13130 DVSS.n13129 0.00781054
R30917 DVSS.n12953 DVSS.n12952 0.00781054
R30918 DVSS.n12928 DVSS.n12927 0.00781054
R30919 DVSS.n12892 DVSS.n12891 0.00781054
R30920 DVSS.n12862 DVSS.n12861 0.00781054
R30921 DVSS.n11284 DVSS.n11283 0.00781054
R30922 DVSS.n12929 DVSS.n12928 0.00781054
R30923 DVSS.n9547 DVSS.n9546 0.00781054
R30924 DVSS.n9516 DVSS.n9515 0.00781054
R30925 DVSS.n9572 DVSS.n9571 0.00781054
R30926 DVSS.n8999 DVSS.n8998 0.00781054
R30927 DVSS.n13129 DVSS.n13128 0.00781054
R30928 DVSS.n10916 DVSS.n10915 0.00781054
R30929 DVSS.n10929 DVSS.n10928 0.00781054
R30930 DVSS.n10197 DVSS.n10196 0.00781054
R30931 DVSS.n12952 DVSS.n12951 0.00781054
R30932 DVSS.n11272 DVSS.n11271 0.00781054
R30933 DVSS.n16943 DVSS.n16942 0.00781054
R30934 DVSS.n17048 DVSS.n17047 0.00781054
R30935 DVSS.n17061 DVSS.n17060 0.00781054
R30936 DVSS.n17580 DVSS.n17579 0.00781054
R30937 DVSS.n17594 DVSS.n17593 0.00781054
R30938 DVSS.n15680 DVSS.n15679 0.00781054
R30939 DVSS.n15651 DVSS.n15650 0.00781054
R30940 DVSS.n15624 DVSS.n15623 0.00781054
R30941 DVSS.n14996 DVSS.n14995 0.00781054
R30942 DVSS.n15024 DVSS.n15023 0.00781054
R30943 DVSS.n13665 DVSS.n13664 0.00781054
R30944 DVSS.n13577 DVSS.n13576 0.00781054
R30945 DVSS.n20187 DVSS.n20186 0.00781054
R30946 DVSS.n20303 DVSS.n20302 0.00781054
R30947 DVSS.n20273 DVSS.n20272 0.00781054
R30948 DVSS.n20843 DVSS.n20842 0.00781054
R30949 DVSS.n20809 DVSS.n20808 0.00781054
R30950 DVSS.n20779 DVSS.n20778 0.00781054
R30951 DVSS.n20753 DVSS.n20752 0.00781054
R30952 DVSS.n17581 DVSS.n17580 0.00781054
R30953 DVSS.n13578 DVSS.n13577 0.00781054
R30954 DVSS.n15650 DVSS.n15649 0.00781054
R30955 DVSS.n15681 DVSS.n15680 0.00781054
R30956 DVSS.n15625 DVSS.n15624 0.00781054
R30957 DVSS.n14997 DVSS.n14996 0.00781054
R30958 DVSS.n15025 DVSS.n15024 0.00781054
R30959 DVSS.n17049 DVSS.n17048 0.00781054
R30960 DVSS.n17062 DVSS.n17061 0.00781054
R30961 DVSS.n16942 DVSS.n16941 0.00781054
R30962 DVSS.n17593 DVSS.n17592 0.00781054
R30963 DVSS.n13666 DVSS.n13665 0.00781054
R30964 DVSS.n10602 DVSS.n10601 0.00781054
R30965 DVSS.n10847 DVSS.n10846 0.00781054
R30966 DVSS.n10834 DVSS.n10833 0.00781054
R30967 DVSS.n11377 DVSS.n11376 0.00781054
R30968 DVSS.n11391 DVSS.n11390 0.00781054
R30969 DVSS.n11555 DVSS.n11554 0.00781054
R30970 DVSS.n11584 DVSS.n11583 0.00781054
R30971 DVSS.n11611 DVSS.n11610 0.00781054
R30972 DVSS.n11694 DVSS.n11693 0.00781054
R30973 DVSS.n13071 DVSS.n13070 0.00781054
R30974 DVSS.n13039 DVSS.n13038 0.00781054
R30975 DVSS.n12044 DVSS.n12043 0.00781054
R30976 DVSS.n12077 DVSS.n12076 0.00781054
R30977 DVSS.n34 DVSS.n33 0.00781054
R30978 DVSS.n59 DVSS.n58 0.00781054
R30979 DVSS.n21541 DVSS.n21540 0.00781054
R30980 DVSS.n21511 DVSS.n21510 0.00781054
R30981 DVSS.n21485 DVSS.n21484 0.00781054
R30982 DVSS.n21453 DVSS.n21452 0.00781054
R30983 DVSS.n21423 DVSS.n21422 0.00781054
R30984 DVSS.n21398 DVSS.n21397 0.00781054
R30985 DVSS.n11378 DVSS.n11377 0.00781054
R30986 DVSS.n12043 DVSS.n12042 0.00781054
R30987 DVSS.n13040 DVSS.n13039 0.00781054
R30988 DVSS.n11585 DVSS.n11584 0.00781054
R30989 DVSS.n11554 DVSS.n11553 0.00781054
R30990 DVSS.n11610 DVSS.n11609 0.00781054
R30991 DVSS.n11693 DVSS.n11692 0.00781054
R30992 DVSS.n13072 DVSS.n13071 0.00781054
R30993 DVSS.n10846 DVSS.n10845 0.00781054
R30994 DVSS.n10833 DVSS.n10832 0.00781054
R30995 DVSS.n10601 DVSS.n10600 0.00781054
R30996 DVSS.n11390 DVSS.n11389 0.00781054
R30997 DVSS.n9899 DVSS.n9898 0.00781054
R30998 DVSS.n9937 DVSS.n9936 0.00781054
R30999 DVSS.n9950 DVSS.n9949 0.00781054
R31000 DVSS.n11103 DVSS.n11102 0.00781054
R31001 DVSS.n11117 DVSS.n11116 0.00781054
R31002 DVSS.n9677 DVSS.n9676 0.00781054
R31003 DVSS.n9648 DVSS.n9647 0.00781054
R31004 DVSS.n9621 DVSS.n9620 0.00781054
R31005 DVSS.n9088 DVSS.n9087 0.00781054
R31006 DVSS.n9060 DVSS.n9059 0.00781054
R31007 DVSS.n13210 DVSS.n13209 0.00781054
R31008 DVSS.n13255 DVSS.n13254 0.00781054
R31009 DVSS.n20458 DVSS.n20457 0.00781054
R31010 DVSS.n20577 DVSS.n20576 0.00781054
R31011 DVSS.n20547 DVSS.n20546 0.00781054
R31012 DVSS.n21069 DVSS.n21068 0.00781054
R31013 DVSS.n21035 DVSS.n21034 0.00781054
R31014 DVSS.n21005 DVSS.n21004 0.00781054
R31015 DVSS.n20979 DVSS.n20978 0.00781054
R31016 DVSS.n11104 DVSS.n11103 0.00781054
R31017 DVSS.n13254 DVSS.n13253 0.00781054
R31018 DVSS.n9647 DVSS.n9646 0.00781054
R31019 DVSS.n9678 DVSS.n9677 0.00781054
R31020 DVSS.n9622 DVSS.n9621 0.00781054
R31021 DVSS.n9089 DVSS.n9088 0.00781054
R31022 DVSS.n9061 DVSS.n9060 0.00781054
R31023 DVSS.n9938 DVSS.n9937 0.00781054
R31024 DVSS.n9951 DVSS.n9950 0.00781054
R31025 DVSS.n9898 DVSS.n9897 0.00781054
R31026 DVSS.n11116 DVSS.n11115 0.00781054
R31027 DVSS.n13209 DVSS.n13208 0.00781054
R31028 DVSS.n60 DVSS.n59 0.00781054
R31029 DVSS.n20186 DVSS.n20185 0.00781054
R31030 DVSS.n20457 DVSS.n20456 0.00781054
R31031 DVSS.n12863 DVSS.n12862 0.00781054
R31032 DVSS.n33 DVSS.n32 0.00781054
R31033 DVSS.n12893 DVSS.n12892 0.00781054
R31034 DVSS.n12078 DVSS.n12077 0.00781054
R31035 DVSS.n20400 DVSS.n20399 0.00781054
R31036 DVSS.n20117 DVSS.n20116 0.00781054
R31037 DVSS.n21542 DVSS.n21541 0.00781054
R31038 DVSS.n20576 DVSS.n20575 0.00781054
R31039 DVSS.n20302 DVSS.n20301 0.00781054
R31040 DVSS.n21512 DVSS.n21511 0.00781054
R31041 DVSS.n20546 DVSS.n20545 0.00781054
R31042 DVSS.n20272 DVSS.n20271 0.00781054
R31043 DVSS.n21486 DVSS.n21485 0.00781054
R31044 DVSS.n21070 DVSS.n21069 0.00781054
R31045 DVSS.n20844 DVSS.n20843 0.00781054
R31046 DVSS.n20752 DVSS.n20751 0.00781054
R31047 DVSS.n21454 DVSS.n21453 0.00781054
R31048 DVSS.n21034 DVSS.n21033 0.00781054
R31049 DVSS.n20808 DVSS.n20807 0.00781054
R31050 DVSS.n21424 DVSS.n21423 0.00781054
R31051 DVSS.n21004 DVSS.n21003 0.00781054
R31052 DVSS.n20778 DVSS.n20777 0.00781054
R31053 DVSS.n20978 DVSS.n20977 0.00781054
R31054 DVSS.n21397 DVSS.n21396 0.00781054
R31055 DVSS.n20248 DVSS.n20247 0.00780945
R31056 DVSS.n20522 DVSS.n20521 0.00780945
R31057 DVSS.n19509 DVSS.n19508 0.00780945
R31058 DVSS.n19643 DVSS.n19641 0.0077973
R31059 DVSS.n19681 DVSS.n19678 0.0077973
R31060 DVSS.n19900 DVSS.n19899 0.0077973
R31061 DVSS.n19875 DVSS.n19874 0.0077973
R31062 DVSS.n2361 DVSS.n2360 0.00779557
R31063 DVSS.n2405 DVSS.n2404 0.00779557
R31064 DVSS.n2393 DVSS.n2392 0.0077955
R31065 DVSS.n2372 DVSS.n2371 0.0077955
R31066 DVSS.n2346 DVSS.n2345 0.00779539
R31067 DVSS.n2376 DVSS.n2375 0.00779449
R31068 DVSS.n2365 DVSS.n2364 0.00779416
R31069 DVSS.n2401 DVSS.n2400 0.00779416
R31070 DVSS.n2357 DVSS.n2356 0.00779335
R31071 DVSS.n2342 DVSS.n2341 0.00779236
R31072 DVSS.n6137 DVSS.n6136 0.0077918
R31073 DVSS.n6131 DVSS.n6130 0.0077918
R31074 DVSS.n6123 DVSS.n6122 0.0077918
R31075 DVSS.n6117 DVSS.n6116 0.0077918
R31076 DVSS.n6111 DVSS.n6110 0.0077918
R31077 DVSS.n5712 DVSS.n5711 0.00776378
R31078 DVSS.n11002 DVSS.n11001 0.00776378
R31079 DVSS.n16905 DVSS.n16904 0.00776378
R31080 DVSS.n9861 DVSS.n9840 0.00776378
R31081 DVSS.n17431 DVSS.n17430 0.00776378
R31082 DVSS.n17220 DVSS.n17219 0.0077
R31083 DVSS.n17224 DVSS.n17223 0.0077
R31084 DVSS.n15188 DVSS.n15187 0.0077
R31085 DVSS.n15143 DVSS.n15142 0.0077
R31086 DVSS.n17698 DVSS.n17697 0.0077
R31087 DVSS.n17778 DVSS.n17777 0.0076831
R31088 DVSS.n15885 DVSS.n15884 0.0076831
R31089 DVSS.n14399 DVSS.n14398 0.0076451
R31090 DVSS.n14400 DVSS.n14399 0.0076451
R31091 DVSS.n14728 DVSS.n14727 0.0076451
R31092 DVSS.n14729 DVSS.n14728 0.0076451
R31093 DVSS.n12146 DVSS.n12145 0.00761538
R31094 DVSS.n12610 DVSS.n12609 0.00761538
R31095 DVSS.n12595 DVSS.n12594 0.00761538
R31096 DVSS.n12322 DVSS.n12321 0.00761538
R31097 DVSS.n12307 DVSS.n12306 0.00761538
R31098 DVSS.n12230 DVSS.n12229 0.00761538
R31099 DVSS.n2766 DVSS.n2765 0.00761538
R31100 DVSS.n3234 DVSS.n3233 0.00761538
R31101 DVSS.n3219 DVSS.n3218 0.00761538
R31102 DVSS.n2949 DVSS.n2948 0.00761538
R31103 DVSS.n2934 DVSS.n2933 0.00761538
R31104 DVSS.n2857 DVSS.n2856 0.00761538
R31105 DVSS.n884 DVSS.n883 0.00761538
R31106 DVSS.n2051 DVSS.n2050 0.00757143
R31107 DVSS.n1723 DVSS.n1722 0.00757143
R31108 DVSS.n8065 DVSS.n8064 0.00750714
R31109 DVSS.n11742 DVSS.n11741 0.00750714
R31110 DVSS.n8357 DVSS.n8356 0.00750714
R31111 DVSS.n19238 DVSS.n19237 0.00747736
R31112 DVSS.n15424 DVSS.n15423 0.007475
R31113 DVSS.n18288 DVSS.n18287 0.007475
R31114 DVSS.n18337 DVSS.n18336 0.007475
R31115 DVSS.n18338 DVSS.n18337 0.007475
R31116 DVSS.n12705 DVSS.n12704 0.00740945
R31117 DVSS.n10795 DVSS.n10794 0.00740945
R31118 DVSS.n3328 DVSS.n3327 0.00740945
R31119 DVSS.n5469 DVSS.n5468 0.00740945
R31120 DVSS.n8120 DVSS.n8118 0.00737857
R31121 DVSS.n11799 DVSS.n11797 0.00737857
R31122 DVSS.n8412 DVSS.n8410 0.00737857
R31123 DVSS.n12829 DVSS.n12828 0.00735992
R31124 DVSS.n21139 DVSS.n21138 0.00735992
R31125 DVSS.n21136 DVSS.n21135 0.00735992
R31126 DVSS.n3789 DVSS.n3788 0.00735992
R31127 DVSS.n13850 DVSS.n13849 0.00733971
R31128 DVSS.n12942 DVSS.n8049 0.00733971
R31129 DVSS.n13182 DVSS.n13181 0.00733971
R31130 DVSS.n18574 DVSS.n18573 0.00733971
R31131 DVSS.n6953 DVSS.n6952 0.00733971
R31132 DVSS.n2012 DVSS.n2011 0.00731429
R31133 DVSS.n2458 DVSS.n2457 0.00731429
R31134 DVSS.n7724 DVSS.n7723 0.00725
R31135 DVSS.n2004 DVSS.n2003 0.00725
R31136 DVSS.n2332 DVSS.n2331 0.00725
R31137 DVSS.n16055 DVSS.n16054 0.00725
R31138 DVSS.n17683 DVSS.n17682 0.00725
R31139 DVSS.n4968 DVSS.n4967 0.00725
R31140 DVSS.n4924 DVSS.n4923 0.00725
R31141 DVSS.n4864 DVSS.n4863 0.00725
R31142 DVSS.n4794 DVSS.n4793 0.00725
R31143 DVSS.n10103 DVSS.n10102 0.00725
R31144 DVSS.n10148 DVSS.n10147 0.00725
R31145 DVSS.n4813 DVSS.n4812 0.00725
R31146 DVSS.n3909 DVSS.n3908 0.00725
R31147 DVSS.n3863 DVSS.n3862 0.00725
R31148 DVSS.n8076 DVSS.n8075 0.00725
R31149 DVSS.n8104 DVSS.n8103 0.00725
R31150 DVSS.n8112 DVSS.n8111 0.00725
R31151 DVSS.n8163 DVSS.n8162 0.00725
R31152 DVSS.n8214 DVSS.n8213 0.00725
R31153 DVSS.n2703 DVSS.n2702 0.00725
R31154 DVSS.n2649 DVSS.n2648 0.00725
R31155 DVSS.n11755 DVSS.n11754 0.00725
R31156 DVSS.n11781 DVSS.n11780 0.00725
R31157 DVSS.n11789 DVSS.n11788 0.00725
R31158 DVSS.n11848 DVSS.n11847 0.00725
R31159 DVSS.n11907 DVSS.n11906 0.00725
R31160 DVSS.n5987 DVSS.n5986 0.00725
R31161 DVSS.n5941 DVSS.n5940 0.00725
R31162 DVSS.n8368 DVSS.n8367 0.00725
R31163 DVSS.n8396 DVSS.n8395 0.00725
R31164 DVSS.n8404 DVSS.n8403 0.00725
R31165 DVSS.n8455 DVSS.n8454 0.00725
R31166 DVSS.n8506 DVSS.n8505 0.00725
R31167 DVSS.n8601 DVSS.n8600 0.00725
R31168 DVSS.n6240 DVSS.n6239 0.00725
R31169 DVSS.n6182 DVSS.n6181 0.00725
R31170 DVSS.n8616 DVSS.n8615 0.00725
R31171 DVSS.n8646 DVSS.n8645 0.00725
R31172 DVSS.n8717 DVSS.n8716 0.00725
R31173 DVSS.n8778 DVSS.n8777 0.00725
R31174 DVSS.n12706 DVSS.n12705 0.00723228
R31175 DVSS.n3329 DVSS.n3328 0.00723228
R31176 DVSS.n12548 DVSS.n12547 0.00723077
R31177 DVSS.n12672 DVSS.n12671 0.00723077
R31178 DVSS.n12580 DVSS.n12579 0.00723077
R31179 DVSS.n12384 DVSS.n12383 0.00723077
R31180 DVSS.n12292 DVSS.n12291 0.00723077
R31181 DVSS.n12245 DVSS.n12244 0.00723077
R31182 DVSS.n3172 DVSS.n3171 0.00723077
R31183 DVSS.n3296 DVSS.n3295 0.00723077
R31184 DVSS.n3204 DVSS.n3203 0.00723077
R31185 DVSS.n3011 DVSS.n3010 0.00723077
R31186 DVSS.n2919 DVSS.n2918 0.00723077
R31187 DVSS.n2872 DVSS.n2871 0.00723077
R31188 DVSS.n14468 DVSS.n14467 0.00722377
R31189 DVSS.n14467 DVSS.n14466 0.00722377
R31190 DVSS.n14654 DVSS.n14653 0.00722377
R31191 DVSS.n14655 DVSS.n14654 0.00722377
R31192 DVSS.n6514 DVSS.n6513 0.00722225
R31193 DVSS.n9772 DVSS.n9771 0.00722225
R31194 DVSS.n9760 DVSS.n9759 0.00722225
R31195 DVSS.n9580 DVSS.n9579 0.00722225
R31196 DVSS.n9148 DVSS.n9147 0.00722225
R31197 DVSS.n15863 DVSS.n15862 0.00722225
R31198 DVSS.n15712 DVSS.n15711 0.00722225
R31199 DVSS.n15617 DVSS.n15616 0.00722225
R31200 DVSS.n14982 DVSS.n14981 0.00722225
R31201 DVSS.n13141 DVSS.n13140 0.00722225
R31202 DVSS.n15036 DVSS.n15035 0.00722225
R31203 DVSS.n4042 DVSS.n4041 0.00722225
R31204 DVSS.n4344 DVSS.n4343 0.00722225
R31205 DVSS.n4126 DVSS.n4125 0.00722225
R31206 DVSS.n5249 DVSS.n5248 0.00719014
R31207 DVSS.n5166 DVSS.n5165 0.00719014
R31208 DVSS.n5114 DVSS.n5111 0.00719014
R31209 DVSS.n6521 DVSS.n6520 0.00716351
R31210 DVSS.n6534 DVSS.n6533 0.00716351
R31211 DVSS.n4379 DVSS.n4378 0.00716351
R31212 DVSS.n4093 DVSS.n4092 0.00716351
R31213 DVSS.n4035 DVSS.n4034 0.00716351
R31214 DVSS.n9779 DVSS.n9778 0.00716351
R31215 DVSS.n9753 DVSS.n9752 0.00716351
R31216 DVSS.n9587 DVSS.n9586 0.00716351
R31217 DVSS.n9141 DVSS.n9140 0.00716351
R31218 DVSS.n13148 DVSS.n13147 0.00716351
R31219 DVSS.n15856 DVSS.n15855 0.00716351
R31220 DVSS.n15719 DVSS.n15718 0.00716351
R31221 DVSS.n15610 DVSS.n15609 0.00716351
R31222 DVSS.n14989 DVSS.n14988 0.00716351
R31223 DVSS.n15043 DVSS.n15042 0.00716351
R31224 DVSS.n4351 DVSS.n4350 0.00716351
R31225 DVSS.n4119 DVSS.n4118 0.00716351
R31226 DVSS.n4000 DVSS.n3999 0.00716351
R31227 DVSS.n9799 DVSS.n9798 0.00716351
R31228 DVSS.n9716 DVSS.n9715 0.00716351
R31229 DVSS.n9607 DVSS.n9606 0.00716351
R31230 DVSS.n9104 DVSS.n9103 0.00716351
R31231 DVSS.n9042 DVSS.n9041 0.00716351
R31232 DVSS.n16288 DVSS.n16287 0.00716351
R31233 DVSS.n16249 DVSS.n16248 0.00716351
R31234 DVSS.n16128 DVSS.n7548 0.00716351
R31235 DVSS.n18388 DVSS.n18387 0.00716351
R31236 DVSS.n7500 DVSS.n7499 0.00716351
R31237 DVSS.n16610 DVSS.n16609 0.00706915
R31238 DVSS.n16614 DVSS.n16613 0.00706915
R31239 DVSS.n16618 DVSS.n16617 0.00706915
R31240 DVSS.n16622 DVSS.n16621 0.00706915
R31241 DVSS.n16781 DVSS.n16780 0.00706915
R31242 DVSS.n16785 DVSS.n16784 0.00706915
R31243 DVSS.n16628 DVSS.n16627 0.00706915
R31244 DVSS.n16790 DVSS.n16789 0.00706915
R31245 DVSS.n16794 DVSS.n16793 0.00706915
R31246 DVSS.n16710 DVSS.n16709 0.00706915
R31247 DVSS.n17191 DVSS.n17190 0.00706915
R31248 DVSS.n17194 DVSS.n17193 0.00706915
R31249 DVSS.n17197 DVSS.n17196 0.00706915
R31250 DVSS.n17200 DVSS.n17199 0.00706915
R31251 DVSS.n17203 DVSS.n17202 0.00706915
R31252 DVSS.n17206 DVSS.n17205 0.00706915
R31253 DVSS.n17222 DVSS.n17221 0.00706915
R31254 DVSS.n17223 DVSS.n17222 0.00706915
R31255 DVSS.n17207 DVSS.n17206 0.00706915
R31256 DVSS.n17204 DVSS.n17203 0.00706915
R31257 DVSS.n17201 DVSS.n17200 0.00706915
R31258 DVSS.n17198 DVSS.n17197 0.00706915
R31259 DVSS.n17195 DVSS.n17194 0.00706915
R31260 DVSS.n17192 DVSS.n17191 0.00706915
R31261 DVSS.n17189 DVSS.n16710 0.00706915
R31262 DVSS.n16795 DVSS.n16794 0.00706915
R31263 DVSS.n16791 DVSS.n16790 0.00706915
R31264 DVSS.n16629 DVSS.n16628 0.00706915
R31265 DVSS.n16786 DVSS.n16785 0.00706915
R31266 DVSS.n16782 DVSS.n16781 0.00706915
R31267 DVSS.n16623 DVSS.n16622 0.00706915
R31268 DVSS.n16619 DVSS.n16618 0.00706915
R31269 DVSS.n16615 DVSS.n16614 0.00706915
R31270 DVSS.n16611 DVSS.n16610 0.00706915
R31271 DVSS.n15189 DVSS.n15188 0.00706915
R31272 DVSS.n15155 DVSS.n15154 0.00706915
R31273 DVSS.n7725 DVSS.n7724 0.00706915
R31274 DVSS.n15103 DVSS.n15102 0.00706915
R31275 DVSS.n15100 DVSS.n15099 0.00706915
R31276 DVSS.n15097 DVSS.n15096 0.00706915
R31277 DVSS.n15094 DVSS.n15093 0.00706915
R31278 DVSS.n15091 DVSS.n15090 0.00706915
R31279 DVSS.n15088 DVSS.n15087 0.00706915
R31280 DVSS.n15085 DVSS.n15084 0.00706915
R31281 DVSS.n15082 DVSS.n15081 0.00706915
R31282 DVSS.n15079 DVSS.n15078 0.00706915
R31283 DVSS.n15076 DVSS.n15075 0.00706915
R31284 DVSS.n15073 DVSS.n15072 0.00706915
R31285 DVSS.n15072 DVSS.n15068 0.00706915
R31286 DVSS.n15075 DVSS.n15074 0.00706915
R31287 DVSS.n15078 DVSS.n15077 0.00706915
R31288 DVSS.n15081 DVSS.n15080 0.00706915
R31289 DVSS.n15084 DVSS.n15083 0.00706915
R31290 DVSS.n15087 DVSS.n15086 0.00706915
R31291 DVSS.n15090 DVSS.n15089 0.00706915
R31292 DVSS.n15093 DVSS.n15092 0.00706915
R31293 DVSS.n15096 DVSS.n15095 0.00706915
R31294 DVSS.n15099 DVSS.n15098 0.00706915
R31295 DVSS.n15102 DVSS.n15101 0.00706915
R31296 DVSS.n15116 DVSS.n7725 0.00706915
R31297 DVSS.n15156 DVSS.n15155 0.00706915
R31298 DVSS.n15190 DVSS.n15189 0.00706915
R31299 DVSS.n15180 DVSS.n15179 0.00706915
R31300 DVSS.n15207 DVSS.n15206 0.00706915
R31301 DVSS.n16096 DVSS.n16095 0.00706915
R31302 DVSS.n16083 DVSS.n16082 0.00706915
R31303 DVSS.n16056 DVSS.n16055 0.00706915
R31304 DVSS.n16040 DVSS.n16039 0.00706915
R31305 DVSS.n16036 DVSS.n16035 0.00706915
R31306 DVSS.n16032 DVSS.n16031 0.00706915
R31307 DVSS.n16028 DVSS.n16027 0.00706915
R31308 DVSS.n16024 DVSS.n16023 0.00706915
R31309 DVSS.n16020 DVSS.n16019 0.00706915
R31310 DVSS.n16016 DVSS.n16015 0.00706915
R31311 DVSS.n7646 DVSS.n7645 0.00706915
R31312 DVSS.n17719 DVSS.n17718 0.00706915
R31313 DVSS.n17716 DVSS.n17715 0.00706915
R31314 DVSS.n17713 DVSS.n17712 0.00706915
R31315 DVSS.n17710 DVSS.n17709 0.00706915
R31316 DVSS.n17707 DVSS.n17706 0.00706915
R31317 DVSS.n17704 DVSS.n17703 0.00706915
R31318 DVSS.n17701 DVSS.n17700 0.00706915
R31319 DVSS.n17686 DVSS.n17685 0.00706915
R31320 DVSS.n17685 DVSS.n17684 0.00706915
R31321 DVSS.n17700 DVSS.n17699 0.00706915
R31322 DVSS.n17703 DVSS.n17702 0.00706915
R31323 DVSS.n17706 DVSS.n17705 0.00706915
R31324 DVSS.n17709 DVSS.n17708 0.00706915
R31325 DVSS.n17712 DVSS.n17711 0.00706915
R31326 DVSS.n17715 DVSS.n17714 0.00706915
R31327 DVSS.n17718 DVSS.n17717 0.00706915
R31328 DVSS.n17720 DVSS.n7646 0.00706915
R31329 DVSS.n16017 DVSS.n16016 0.00706915
R31330 DVSS.n16021 DVSS.n16020 0.00706915
R31331 DVSS.n16025 DVSS.n16024 0.00706915
R31332 DVSS.n16029 DVSS.n16028 0.00706915
R31333 DVSS.n16033 DVSS.n16032 0.00706915
R31334 DVSS.n16037 DVSS.n16036 0.00706915
R31335 DVSS.n16041 DVSS.n16040 0.00706915
R31336 DVSS.n16057 DVSS.n16056 0.00706915
R31337 DVSS.n16084 DVSS.n16083 0.00706915
R31338 DVSS.n16097 DVSS.n16096 0.00706915
R31339 DVSS.n17493 DVSS.n17492 0.00706915
R31340 DVSS.n17496 DVSS.n17495 0.00706915
R31341 DVSS.n17499 DVSS.n17498 0.00706915
R31342 DVSS.n17502 DVSS.n17501 0.00706915
R31343 DVSS.n17505 DVSS.n17504 0.00706915
R31344 DVSS.n17508 DVSS.n17507 0.00706915
R31345 DVSS.n17511 DVSS.n17510 0.00706915
R31346 DVSS.n17514 DVSS.n17513 0.00706915
R31347 DVSS.n17517 DVSS.n17516 0.00706915
R31348 DVSS.n17520 DVSS.n17519 0.00706915
R31349 DVSS.n17523 DVSS.n17522 0.00706915
R31350 DVSS.n17524 DVSS.n17523 0.00706915
R31351 DVSS.n17518 DVSS.n17517 0.00706915
R31352 DVSS.n17512 DVSS.n17511 0.00706915
R31353 DVSS.n17509 DVSS.n17508 0.00706915
R31354 DVSS.n17506 DVSS.n17505 0.00706915
R31355 DVSS.n17503 DVSS.n17502 0.00706915
R31356 DVSS.n17500 DVSS.n17499 0.00706915
R31357 DVSS.n17497 DVSS.n17496 0.00706915
R31358 DVSS.n17494 DVSS.n17493 0.00706915
R31359 DVSS.n16490 DVSS.n16489 0.00706915
R31360 DVSS.n16486 DVSS.n16485 0.00706915
R31361 DVSS.n16482 DVSS.n16481 0.00706915
R31362 DVSS.n16478 DVSS.n16477 0.00706915
R31363 DVSS.n16474 DVSS.n16473 0.00706915
R31364 DVSS.n16470 DVSS.n16469 0.00706915
R31365 DVSS.n16466 DVSS.n16465 0.00706915
R31366 DVSS.n16462 DVSS.n16461 0.00706915
R31367 DVSS.n16458 DVSS.n16457 0.00706915
R31368 DVSS.n16454 DVSS.n16453 0.00706915
R31369 DVSS.n16450 DVSS.n16449 0.00706915
R31370 DVSS.n16446 DVSS.n16445 0.00706915
R31371 DVSS.n16004 DVSS.n16003 0.00706915
R31372 DVSS.n17515 DVSS.n17514 0.00706915
R31373 DVSS.n17521 DVSS.n17520 0.00706915
R31374 DVSS.n15299 DVSS.n15298 0.00706915
R31375 DVSS.n15296 DVSS.n15295 0.00706915
R31376 DVSS.n15293 DVSS.n15292 0.00706915
R31377 DVSS.n15290 DVSS.n15289 0.00706915
R31378 DVSS.n15287 DVSS.n15286 0.00706915
R31379 DVSS.n15284 DVSS.n15283 0.00706915
R31380 DVSS.n15281 DVSS.n15280 0.00706915
R31381 DVSS.n15278 DVSS.n15277 0.00706915
R31382 DVSS.n15275 DVSS.n15274 0.00706915
R31383 DVSS.n15272 DVSS.n15271 0.00706915
R31384 DVSS.n15269 DVSS.n15268 0.00706915
R31385 DVSS.n15268 DVSS.n15267 0.00706915
R31386 DVSS.n15274 DVSS.n15273 0.00706915
R31387 DVSS.n15277 DVSS.n15276 0.00706915
R31388 DVSS.n15280 DVSS.n15279 0.00706915
R31389 DVSS.n15283 DVSS.n15282 0.00706915
R31390 DVSS.n15286 DVSS.n15285 0.00706915
R31391 DVSS.n15289 DVSS.n15288 0.00706915
R31392 DVSS.n15292 DVSS.n15291 0.00706915
R31393 DVSS.n15295 DVSS.n15294 0.00706915
R31394 DVSS.n15298 DVSS.n15297 0.00706915
R31395 DVSS.n15357 DVSS.n15356 0.00706915
R31396 DVSS.n15353 DVSS.n15352 0.00706915
R31397 DVSS.n15349 DVSS.n15348 0.00706915
R31398 DVSS.n15345 DVSS.n15344 0.00706915
R31399 DVSS.n15341 DVSS.n15340 0.00706915
R31400 DVSS.n15337 DVSS.n15336 0.00706915
R31401 DVSS.n15333 DVSS.n15332 0.00706915
R31402 DVSS.n15329 DVSS.n15328 0.00706915
R31403 DVSS.n15325 DVSS.n15324 0.00706915
R31404 DVSS.n15321 DVSS.n15320 0.00706915
R31405 DVSS.n15317 DVSS.n15316 0.00706915
R31406 DVSS.n15313 DVSS.n15312 0.00706915
R31407 DVSS.n7704 DVSS.n7703 0.00706915
R31408 DVSS.n15271 DVSS.n15270 0.00706915
R31409 DVSS.n15400 DVSS.n15399 0.00706915
R31410 DVSS.n15436 DVSS.n15435 0.00706915
R31411 DVSS.n18289 DVSS.n18288 0.00706915
R31412 DVSS.n18323 DVSS.n18322 0.00706915
R31413 DVSS.n18324 DVSS.n18323 0.00706915
R31414 DVSS.n18290 DVSS.n18289 0.00706915
R31415 DVSS.n15437 DVSS.n15436 0.00706915
R31416 DVSS.n15401 DVSS.n15400 0.00706915
R31417 DVSS.n15391 DVSS.n15390 0.00706915
R31418 DVSS.n18041 DVSS.n18040 0.00706915
R31419 DVSS.n18044 DVSS.n18043 0.00706915
R31420 DVSS.n18047 DVSS.n18046 0.00706915
R31421 DVSS.n18050 DVSS.n18049 0.00706915
R31422 DVSS.n18053 DVSS.n18052 0.00706915
R31423 DVSS.n18056 DVSS.n18055 0.00706915
R31424 DVSS.n18059 DVSS.n18058 0.00706915
R31425 DVSS.n18062 DVSS.n18061 0.00706915
R31426 DVSS.n18065 DVSS.n18064 0.00706915
R31427 DVSS.n18068 DVSS.n18067 0.00706915
R31428 DVSS.n18071 DVSS.n18070 0.00706915
R31429 DVSS.n18072 DVSS.n18071 0.00706915
R31430 DVSS.n18069 DVSS.n18068 0.00706915
R31431 DVSS.n18066 DVSS.n18065 0.00706915
R31432 DVSS.n18063 DVSS.n18062 0.00706915
R31433 DVSS.n18060 DVSS.n18059 0.00706915
R31434 DVSS.n18057 DVSS.n18056 0.00706915
R31435 DVSS.n18054 DVSS.n18053 0.00706915
R31436 DVSS.n18051 DVSS.n18050 0.00706915
R31437 DVSS.n18048 DVSS.n18047 0.00706915
R31438 DVSS.n18045 DVSS.n18044 0.00706915
R31439 DVSS.n18042 DVSS.n18041 0.00706915
R31440 DVSS.n17957 DVSS.n17956 0.00706915
R31441 DVSS.n17961 DVSS.n17960 0.00706915
R31442 DVSS.n17965 DVSS.n17964 0.00706915
R31443 DVSS.n17969 DVSS.n17968 0.00706915
R31444 DVSS.n17973 DVSS.n17972 0.00706915
R31445 DVSS.n17977 DVSS.n17976 0.00706915
R31446 DVSS.n17981 DVSS.n17980 0.00706915
R31447 DVSS.n17985 DVSS.n17984 0.00706915
R31448 DVSS.n17989 DVSS.n17988 0.00706915
R31449 DVSS.n17993 DVSS.n17992 0.00706915
R31450 DVSS.n17997 DVSS.n17996 0.00706915
R31451 DVSS.n18001 DVSS.n18000 0.00706915
R31452 DVSS.n7619 DVSS.n7618 0.00706915
R31453 DVSS.n17900 DVSS.n17899 0.00706915
R31454 DVSS.n17903 DVSS.n17902 0.00706915
R31455 DVSS.n17906 DVSS.n17905 0.00706915
R31456 DVSS.n17909 DVSS.n17908 0.00706915
R31457 DVSS.n17912 DVSS.n17911 0.00706915
R31458 DVSS.n17915 DVSS.n17914 0.00706915
R31459 DVSS.n17918 DVSS.n17917 0.00706915
R31460 DVSS.n17921 DVSS.n17920 0.00706915
R31461 DVSS.n17924 DVSS.n17923 0.00706915
R31462 DVSS.n17927 DVSS.n17926 0.00706915
R31463 DVSS.n17930 DVSS.n17929 0.00706915
R31464 DVSS.n17931 DVSS.n17930 0.00706915
R31465 DVSS.n17928 DVSS.n17927 0.00706915
R31466 DVSS.n17925 DVSS.n17924 0.00706915
R31467 DVSS.n17922 DVSS.n17921 0.00706915
R31468 DVSS.n17919 DVSS.n17918 0.00706915
R31469 DVSS.n17916 DVSS.n17915 0.00706915
R31470 DVSS.n17913 DVSS.n17912 0.00706915
R31471 DVSS.n17910 DVSS.n17909 0.00706915
R31472 DVSS.n17907 DVSS.n17906 0.00706915
R31473 DVSS.n17904 DVSS.n17903 0.00706915
R31474 DVSS.n17901 DVSS.n17900 0.00706915
R31475 DVSS.n17816 DVSS.n17815 0.00706915
R31476 DVSS.n17820 DVSS.n17819 0.00706915
R31477 DVSS.n17824 DVSS.n17823 0.00706915
R31478 DVSS.n17828 DVSS.n17827 0.00706915
R31479 DVSS.n17832 DVSS.n17831 0.00706915
R31480 DVSS.n17836 DVSS.n17835 0.00706915
R31481 DVSS.n17840 DVSS.n17839 0.00706915
R31482 DVSS.n17844 DVSS.n17843 0.00706915
R31483 DVSS.n17848 DVSS.n17847 0.00706915
R31484 DVSS.n17852 DVSS.n17851 0.00706915
R31485 DVSS.n17856 DVSS.n17855 0.00706915
R31486 DVSS.n17860 DVSS.n17859 0.00706915
R31487 DVSS.n7627 DVSS.n7626 0.00706915
R31488 DVSS.n13862 DVSS.n13861 0.00706915
R31489 DVSS.n13866 DVSS.n13865 0.00706915
R31490 DVSS.n13870 DVSS.n13869 0.00706915
R31491 DVSS.n13874 DVSS.n13873 0.00706915
R31492 DVSS.n13878 DVSS.n13877 0.00706915
R31493 DVSS.n13882 DVSS.n13881 0.00706915
R31494 DVSS.n13886 DVSS.n13885 0.00706915
R31495 DVSS.n13890 DVSS.n13889 0.00706915
R31496 DVSS.n13894 DVSS.n13893 0.00706915
R31497 DVSS.n13898 DVSS.n13897 0.00706915
R31498 DVSS.n13902 DVSS.n13901 0.00706915
R31499 DVSS.n13906 DVSS.n13905 0.00706915
R31500 DVSS.n13910 DVSS.n13909 0.00706915
R31501 DVSS.n13936 DVSS.n13935 0.00706915
R31502 DVSS.n13939 DVSS.n13938 0.00706915
R31503 DVSS.n13942 DVSS.n13941 0.00706915
R31504 DVSS.n13945 DVSS.n13944 0.00706915
R31505 DVSS.n13948 DVSS.n13947 0.00706915
R31506 DVSS.n13951 DVSS.n13950 0.00706915
R31507 DVSS.n13954 DVSS.n13953 0.00706915
R31508 DVSS.n13958 DVSS.n13957 0.00706915
R31509 DVSS.n13960 DVSS.n13959 0.00706915
R31510 DVSS.n13964 DVSS.n13963 0.00706915
R31511 DVSS.n13969 DVSS.n13965 0.00706915
R31512 DVSS.n13911 DVSS.n13910 0.00706915
R31513 DVSS.n13907 DVSS.n13906 0.00706915
R31514 DVSS.n13903 DVSS.n13902 0.00706915
R31515 DVSS.n13899 DVSS.n13898 0.00706915
R31516 DVSS.n13895 DVSS.n13894 0.00706915
R31517 DVSS.n13891 DVSS.n13890 0.00706915
R31518 DVSS.n13887 DVSS.n13886 0.00706915
R31519 DVSS.n13883 DVSS.n13882 0.00706915
R31520 DVSS.n13879 DVSS.n13878 0.00706915
R31521 DVSS.n13875 DVSS.n13874 0.00706915
R31522 DVSS.n13871 DVSS.n13870 0.00706915
R31523 DVSS.n13867 DVSS.n13866 0.00706915
R31524 DVSS.n13863 DVSS.n13862 0.00706915
R31525 DVSS.n13853 DVSS.n13852 0.00706915
R31526 DVSS.n13937 DVSS.n13936 0.00706915
R31527 DVSS.n13940 DVSS.n13939 0.00706915
R31528 DVSS.n13943 DVSS.n13942 0.00706915
R31529 DVSS.n13946 DVSS.n13945 0.00706915
R31530 DVSS.n13949 DVSS.n13948 0.00706915
R31531 DVSS.n13952 DVSS.n13951 0.00706915
R31532 DVSS.n13957 DVSS.n13956 0.00706915
R31533 DVSS.n13955 DVSS.n13954 0.00706915
R31534 DVSS.n13961 DVSS.n13960 0.00706915
R31535 DVSS.n13963 DVSS.n13962 0.00706915
R31536 DVSS.n13970 DVSS.n13969 0.00706915
R31537 DVSS.n6112 DVSS.n6111 0.00706681
R31538 DVSS.n6124 DVSS.n6123 0.00706681
R31539 DVSS.n6132 DVSS.n6131 0.00706681
R31540 DVSS.n6138 DVSS.n6137 0.00706681
R31541 DVSS.n6118 DVSS.n6117 0.00706681
R31542 DVSS.n17470 DVSS.n17469 0.0070493
R31543 DVSS.n18179 DVSS.n18178 0.0070493
R31544 DVSS.n16811 DVSS.n16810 0.0070493
R31545 DVSS.n15561 DVSS.n15560 0.0070493
R31546 DVSS.n16594 DVSS.n16593 0.007025
R31547 DVSS.n16609 DVSS.n16608 0.007025
R31548 DVSS.n18307 DVSS.n18306 0.007025
R31549 DVSS.n18322 DVSS.n18321 0.007025
R31550 DVSS.n4744 DVSS.n4743 0.00699286
R31551 DVSS.n8666 DVSS.n8664 0.00699286
R31552 DVSS.n3439 DVSS.n3438 0.0069488
R31553 DVSS.n10427 DVSS.n10426 0.00690845
R31554 DVSS.n10486 DVSS.n10485 0.00690845
R31555 DVSS.n10583 DVSS.n10581 0.00690845
R31556 DVSS.n6527 DVSS.n6526 0.00689005
R31557 DVSS.n4386 DVSS.n4385 0.00689005
R31558 DVSS.n4086 DVSS.n4085 0.00689005
R31559 DVSS.n10759 DVSS.n10758 0.00687795
R31560 DVSS.n5485 DVSS.n4528 0.00687795
R31561 DVSS.n3813 DVSS.n3812 0.00686429
R31562 DVSS.n3916 DVSS.n3914 0.00686429
R31563 DVSS.n3870 DVSS.n3868 0.00686429
R31564 DVSS.n2586 DVSS.n2585 0.00686429
R31565 DVSS.n5994 DVSS.n5992 0.00686429
R31566 DVSS.n5948 DVSS.n5946 0.00686429
R31567 DVSS.n12736 DVSS.n12735 0.00684615
R31568 DVSS.n12518 DVSS.n12517 0.00684615
R31569 DVSS.n12642 DVSS.n12641 0.00684615
R31570 DVSS.n12619 DVSS.n12618 0.00684615
R31571 DVSS.n12354 DVSS.n12353 0.00684615
R31572 DVSS.n12331 DVSS.n12330 0.00684615
R31573 DVSS.n2774 DVSS.n2773 0.00684615
R31574 DVSS.n3142 DVSS.n3141 0.00684615
R31575 DVSS.n3266 DVSS.n3265 0.00684615
R31576 DVSS.n3243 DVSS.n3242 0.00684615
R31577 DVSS.n2981 DVSS.n2980 0.00684615
R31578 DVSS.n2958 DVSS.n2957 0.00684615
R31579 DVSS.n893 DVSS.n892 0.00684615
R31580 DVSS.n3409 DVSS.n3408 0.00684615
R31581 DVSS.n12783 DVSS.n12782 0.00684615
R31582 DVSS.n2380 DVSS.n2379 0.0068424
R31583 DVSS.n2379 DVSS.n2378 0.0068424
R31584 DVSS.n16082 DVSS.n16081 0.0068
R31585 DVSS.n5403 DVSS.n5397 0.00678492
R31586 DVSS.n1372 DVSS.n1371 0.00678492
R31587 DVSS.n6886 DVSS.n6885 0.00668725
R31588 DVSS.n6759 DVSS.n6758 0.00668725
R31589 DVSS.n6704 DVSS.n6703 0.00668725
R31590 DVSS.n2536 DVSS.n2535 0.00668725
R31591 DVSS.n6397 DVSS.n6396 0.00668725
R31592 DVSS.n2043 DVSS.n2042 0.00667143
R31593 DVSS.n2415 DVSS.n2414 0.00667143
R31594 DVSS.n8171 DVSS.n8168 0.00667143
R31595 DVSS.n8222 DVSS.n8219 0.00667143
R31596 DVSS.n8306 DVSS.n8304 0.00667143
R31597 DVSS.n12981 DVSS.n12980 0.00667143
R31598 DVSS.n8463 DVSS.n8460 0.00667143
R31599 DVSS.n8514 DVSS.n8511 0.00667143
R31600 DVSS.n11315 DVSS.n11314 0.00667143
R31601 DVSS.n18226 DVSS.n18225 0.00662676
R31602 DVSS.n15514 DVSS.n15513 0.00662676
R31603 DVSS.n2368 DVSS.n2367 0.00661798
R31604 DVSS.n2397 DVSS.n2396 0.00661798
R31605 DVSS.n2398 DVSS.n2397 0.00661798
R31606 DVSS.n2712 DVSS.n2710 0.00660714
R31607 DVSS.n2658 DVSS.n2656 0.00660714
R31608 DVSS.n7088 DVSS.n7087 0.0065738
R31609 DVSS.n13595 DVSS.n13594 0.0065738
R31610 DVSS.n7087 DVSS.n7086 0.0065738
R31611 DVSS.n13596 DVSS.n13595 0.0065738
R31612 DVSS.n13237 DVSS.n13236 0.0065738
R31613 DVSS.n13236 DVSS.n13235 0.0065738
R31614 DVSS.n18767 DVSS.n18766 0.0065738
R31615 DVSS.n18766 DVSS.n18765 0.0065738
R31616 DVSS.n933 DVSS.n932 0.00656106
R31617 DVSS.n941 DVSS.n940 0.00656106
R31618 DVSS.n942 DVSS.n941 0.00656106
R31619 DVSS.n21166 DVSS.n21165 0.00656106
R31620 DVSS.n21167 DVSS.n21166 0.00656106
R31621 DVSS.n21181 DVSS.n21180 0.00656106
R31622 DVSS.n5735 DVSS.n5734 0.00652362
R31623 DVSS.n11238 DVSS.n11237 0.00652362
R31624 DVSS.n17627 DVSS.n17626 0.00652362
R31625 DVSS.n11426 DVSS.n11425 0.00652362
R31626 DVSS.n11150 DVSS.n11149 0.00652362
R31627 DVSS.n16356 DVSS.n16355 0.00652362
R31628 DVSS.n6348 DVSS.n6347 0.00652362
R31629 DVSS.n12525 DVSS.n12524 0.00646154
R31630 DVSS.n12649 DVSS.n12648 0.00646154
R31631 DVSS.n12361 DVSS.n12360 0.00646154
R31632 DVSS.n12269 DVSS.n12268 0.00646154
R31633 DVSS.n12268 DVSS.n12267 0.00646154
R31634 DVSS.n3149 DVSS.n3148 0.00646154
R31635 DVSS.n3273 DVSS.n3272 0.00646154
R31636 DVSS.n2988 DVSS.n2987 0.00646154
R31637 DVSS.n2896 DVSS.n2895 0.00646154
R31638 DVSS.n2895 DVSS.n2894 0.00646154
R31639 DVSS.n16863 DVSS.n16862 0.00641549
R31640 DVSS.n2356 DVSS.n2355 0.00639353
R31641 DVSS.n6559 DVSS.n6558 0.00639353
R31642 DVSS.n6423 DVSS.n6422 0.00639353
R31643 DVSS.n11858 DVSS.n11855 0.00635
R31644 DVSS.n11917 DVSS.n11914 0.00635
R31645 DVSS.n11438 DVSS.n11437 0.00634646
R31646 DVSS.n6461 DVSS.n6460 0.00634646
R31647 DVSS.n6443 DVSS.n6442 0.00628209
R31648 DVSS.n6354 DVSS.n6353 0.00628209
R31649 DVSS.n6659 DVSS.n6658 0.00628209
R31650 DVSS.n6720 DVSS.n6719 0.00628209
R31651 DVSS.n6841 DVSS.n6840 0.00628209
R31652 DVSS.n11686 DVSS.n11685 0.0062233
R31653 DVSS.n11649 DVSS.n11648 0.0062233
R31654 DVSS.n11524 DVSS.n11523 0.0062233
R31655 DVSS.n11487 DVSS.n11486 0.0062233
R31656 DVSS.n13055 DVSS.n13054 0.0062233
R31657 DVSS.n6438 DVSS.n6437 0.0062233
R31658 DVSS.n6349 DVSS.n1402 0.0062233
R31659 DVSS.n6664 DVSS.n6663 0.0062233
R31660 DVSS.n6725 DVSS.n6724 0.0062233
R31661 DVSS.n6846 DVSS.n6845 0.0062233
R31662 DVSS.n7155 DVSS.n7154 0.00622032
R31663 DVSS.n13538 DVSS.n13537 0.00622032
R31664 DVSS.n7154 DVSS.n7153 0.00622032
R31665 DVSS.n13539 DVSS.n13538 0.00622032
R31666 DVSS.n13379 DVSS.n13378 0.00622032
R31667 DVSS.n13378 DVSS.n13374 0.00622032
R31668 DVSS.n18837 DVSS.n18836 0.00622032
R31669 DVSS.n18836 DVSS.n18835 0.00622032
R31670 DVSS.n19704 DVSS.n19703 0.00620423
R31671 DVSS.n19783 DVSS.n19782 0.00620423
R31672 DVSS.n135 DVSS.n134 0.00620423
R31673 DVSS.n224 DVSS.n223 0.00620423
R31674 DVSS.n197 DVSS.n196 0.00620423
R31675 DVSS.n19923 DVSS.n19922 0.00620423
R31676 DVSS.n20008 DVSS.n20007 0.00620423
R31677 DVSS.n295 DVSS.n294 0.00620423
R31678 DVSS.n432 DVSS.n431 0.00620423
R31679 DVSS.n405 DVSS.n404 0.00620423
R31680 DVSS.n19167 DVSS.n19166 0.00617568
R31681 DVSS.n19111 DVSS.n19110 0.00617568
R31682 DVSS.n19438 DVSS.n19436 0.00617568
R31683 DVSS.n19386 DVSS.n19385 0.00617568
R31684 DVSS.n20175 DVSS.n20174 0.00617568
R31685 DVSS.n20143 DVSS.n20142 0.00617568
R31686 DVSS.n20446 DVSS.n20444 0.00617568
R31687 DVSS.n20394 DVSS.n20393 0.00617568
R31688 DVSS.n8145 DVSS.n8144 0.00615714
R31689 DVSS.n8196 DVSS.n8195 0.00615714
R31690 DVSS.n8231 DVSS.n8230 0.00615714
R31691 DVSS.n8315 DVSS.n8314 0.00615714
R31692 DVSS.n11926 DVSS.n11925 0.00615714
R31693 DVSS.n12971 DVSS.n12970 0.00615714
R31694 DVSS.n8437 DVSS.n8436 0.00615714
R31695 DVSS.n8488 DVSS.n8487 0.00615714
R31696 DVSS.n8523 DVSS.n8522 0.00615714
R31697 DVSS.n16595 DVSS.n16594 0.006125
R31698 DVSS.n16608 DVSS.n16607 0.006125
R31699 DVSS.n18308 DVSS.n18307 0.006125
R31700 DVSS.n18321 DVSS.n18320 0.006125
R31701 DVSS.n12737 DVSS.n12736 0.00607692
R31702 DVSS.n12618 DVSS.n12617 0.00607692
R31703 DVSS.n12587 DVSS.n12586 0.00607692
R31704 DVSS.n12330 DVSS.n12329 0.00607692
R31705 DVSS.n12299 DVSS.n12298 0.00607692
R31706 DVSS.n12238 DVSS.n12237 0.00607692
R31707 DVSS.n21333 DVSS.n21332 0.00607692
R31708 DVSS.n2775 DVSS.n2774 0.00607692
R31709 DVSS.n3242 DVSS.n3241 0.00607692
R31710 DVSS.n3211 DVSS.n3210 0.00607692
R31711 DVSS.n2957 DVSS.n2956 0.00607692
R31712 DVSS.n2926 DVSS.n2925 0.00607692
R31713 DVSS.n2865 DVSS.n2864 0.00607692
R31714 DVSS.n892 DVSS.n891 0.00607692
R31715 DVSS.n3408 DVSS.n3407 0.00607692
R31716 DVSS.n12782 DVSS.n12781 0.00607692
R31717 DVSS.n5378 DVSS.n5377 0.00603073
R31718 DVSS.n5371 DVSS.n5370 0.00603073
R31719 DVSS.n17030 DVSS.n17024 0.00603073
R31720 DVSS.n10225 DVSS.n10224 0.00603073
R31721 DVSS.n10236 DVSS.n10233 0.00603073
R31722 DVSS.n10291 DVSS.n10285 0.00603073
R31723 DVSS.n10627 DVSS.n10624 0.00603073
R31724 DVSS.n8031 DVSS.n8029 0.00603073
R31725 DVSS.n8032 DVSS.n8031 0.00601993
R31726 DVSS.n16098 DVSS.n16090 0.00599296
R31727 DVSS.n18229 DVSS.n18228 0.00599296
R31728 DVSS.n18459 DVSS.n18458 0.00599296
R31729 DVSS.n19651 DVSS.n19650 0.00599296
R31730 DVSS.n19707 DVSS.n19706 0.00599296
R31731 DVSS.n19724 DVSS.n19723 0.00599296
R31732 DVSS.n19786 DVSS.n19785 0.00599296
R31733 DVSS.n138 DVSS.n137 0.00599296
R31734 DVSS.n227 DVSS.n226 0.00599296
R31735 DVSS.n194 DVSS.n193 0.00599296
R31736 DVSS.n178 DVSS.n177 0.00599296
R31737 DVSS.n15979 DVSS.n15978 0.00599296
R31738 DVSS.n15511 DVSS.n15510 0.00599296
R31739 DVSS.n15158 DVSS.n15157 0.00599296
R31740 DVSS.n19860 DVSS.n19859 0.00599296
R31741 DVSS.n19926 DVSS.n19925 0.00599296
R31742 DVSS.n19943 DVSS.n19942 0.00599296
R31743 DVSS.n20011 DVSS.n20010 0.00599296
R31744 DVSS.n298 DVSS.n297 0.00599296
R31745 DVSS.n435 DVSS.n434 0.00599296
R31746 DVSS.n402 DVSS.n401 0.00599296
R31747 DVSS.n386 DVSS.n385 0.00599296
R31748 DVSS.n5708 DVSS.n5707 0.00599213
R31749 DVSS.n10998 DVSS.n10997 0.00599213
R31750 DVSS.n21235 DVSS.n21234 0.00599213
R31751 DVSS.n16909 DVSS.n16908 0.00599213
R31752 DVSS.n766 DVSS.n765 0.00599213
R31753 DVSS.n9865 DVSS.n9864 0.00599213
R31754 DVSS.n17427 DVSS.n17426 0.00599213
R31755 DVSS.n6803 DVSS.n6802 0.00596429
R31756 DVSS.n3925 DVSS.n3924 0.00596429
R31757 DVSS.n3895 DVSS.n3894 0.00596429
R31758 DVSS.n3849 DVSS.n3848 0.00596429
R31759 DVSS.n3619 DVSS.n3618 0.00596429
R31760 DVSS.n2721 DVSS.n2720 0.00596429
R31761 DVSS.n5973 DVSS.n5972 0.00596429
R31762 DVSS.n5927 DVSS.n5926 0.00596429
R31763 DVSS.n11456 DVSS.n11455 0.00594972
R31764 DVSS.n11493 DVSS.n11492 0.00594972
R31765 DVSS.n11618 DVSS.n11617 0.00594972
R31766 DVSS.n11655 DVSS.n11654 0.00594972
R31767 DVSS.n13060 DVSS.n13059 0.00594972
R31768 DVSS.n17526 DVSS.n17525 0.00594611
R31769 DVSS.n17527 DVSS.n17526 0.00594611
R31770 DVSS.n15266 DVSS.n15265 0.00594611
R31771 DVSS.n15265 DVSS.n15264 0.00594611
R31772 DVSS.n18354 DVSS.n18353 0.00594611
R31773 DVSS.n18353 DVSS.n18349 0.00594611
R31774 DVSS.n18074 DVSS.n18073 0.00594611
R31775 DVSS.n18075 DVSS.n18074 0.00594611
R31776 DVSS.n17933 DVSS.n17932 0.00594611
R31777 DVSS.n17934 DVSS.n17933 0.00594611
R31778 DVSS.n2400 DVSS.n2399 0.00594456
R31779 DVSS.n949 DVSS.n948 0.00594375
R31780 DVSS.n10316 DVSS.n10315 0.00592254
R31781 DVSS.n10358 DVSS.n10357 0.00592254
R31782 DVSS.n7723 DVSS.n7722 0.0059
R31783 DVSS.n16054 DVSS.n16053 0.0059
R31784 DVSS.n4977 DVSS.n4976 0.0059
R31785 DVSS.n4933 DVSS.n4932 0.0059
R31786 DVSS.n4873 DVSS.n4872 0.0059
R31787 DVSS.n6248 DVSS.n6247 0.0059
R31788 DVSS.n6191 DVSS.n6189 0.0059
R31789 DVSS.n10976 DVSS.n10975 0.00587205
R31790 DVSS.n21163 DVSS.n21162 0.00584085
R31791 DVSS.n16592 DVSS.n16591 0.00583379
R31792 DVSS.n16593 DVSS.n16592 0.00583379
R31793 DVSS.n15213 DVSS.n15212 0.00583379
R31794 DVSS.n15214 DVSS.n15213 0.00583379
R31795 DVSS.n16496 DVSS.n16495 0.00583379
R31796 DVSS.n16497 DVSS.n16496 0.00583379
R31797 DVSS.n15363 DVSS.n15362 0.00583379
R31798 DVSS.n15364 DVSS.n15363 0.00583379
R31799 DVSS.n18093 DVSS.n18092 0.00583379
R31800 DVSS.n18094 DVSS.n18093 0.00583379
R31801 DVSS.n17952 DVSS.n17951 0.00583379
R31802 DVSS.n17953 DVSS.n17952 0.00583379
R31803 DVSS.n17811 DVSS.n17810 0.00583379
R31804 DVSS.n17812 DVSS.n17811 0.00583379
R31805 DVSS.n21168 DVSS.n21167 0.00581245
R31806 DVSS.n21180 DVSS.n21173 0.00581245
R31807 DVSS.n932 DVSS.n931 0.00581245
R31808 DVSS.n940 DVSS.n935 0.00581245
R31809 DVSS.n21165 DVSS.n21164 0.00581245
R31810 DVSS.n943 DVSS.n942 0.00581245
R31811 DVSS.n16550 DVSS.n16549 0.00578169
R31812 DVSS.n16565 DVSS.n16564 0.00578169
R31813 DVSS.n16588 DVSS.n16587 0.00578169
R31814 DVSS.n17768 DVSS.n17767 0.00578169
R31815 DVSS.n18116 DVSS.n18115 0.00578169
R31816 DVSS.n18230 DVSS.n18229 0.00578169
R31817 DVSS.n19761 DVSS.n19760 0.00578169
R31818 DVSS.n165 DVSS.n164 0.00578169
R31819 DVSS.n16737 DVSS.n16736 0.00578169
R31820 DVSS.n16752 DVSS.n16751 0.00578169
R31821 DVSS.n16775 DVSS.n16774 0.00578169
R31822 DVSS.n15895 DVSS.n15894 0.00578169
R31823 DVSS.n15406 DVSS.n15405 0.00578169
R31824 DVSS.n15510 DVSS.n15509 0.00578169
R31825 DVSS.n19986 DVSS.n19985 0.00578169
R31826 DVSS.n325 DVSS.n324 0.00578169
R31827 DVSS.n7186 DVSS.n7181 0.00576596
R31828 DVSS.n7307 DVSS.n7305 0.00576596
R31829 DVSS.n7883 DVSS.n7874 0.00576596
R31830 DVSS.n7962 DVSS.n7961 0.00576596
R31831 DVSS.n7040 DVSS.n7039 0.00576596
R31832 DVSS.n7080 DVSS.n7079 0.00576596
R31833 DVSS.n7052 DVSS.n7051 0.00576596
R31834 DVSS.n13613 DVSS.n13612 0.00576596
R31835 DVSS.n13633 DVSS.n13632 0.00576596
R31836 DVSS.n13303 DVSS.n13302 0.00576596
R31837 DVSS.n2339 DVSS.n2338 0.00572004
R31838 DVSS.n2377 DVSS.n2376 0.00572004
R31839 DVSS.n6028 DVSS.n6026 0.00570714
R31840 DVSS.n15425 DVSS.n15424 0.005675
R31841 DVSS.n18287 DVSS.n18286 0.005675
R31842 DVSS.n18336 DVSS.n18335 0.005675
R31843 DVSS.n18339 DVSS.n18338 0.005675
R31844 DVSS.n10090 DVSS.n10089 0.00564286
R31845 DVSS.n10157 DVSS.n10156 0.00564286
R31846 DVSS.n10710 DVSS.n10707 0.00564286
R31847 DVSS.n8725 DVSS.n8724 0.00564286
R31848 DVSS.n8786 DVSS.n8785 0.00564286
R31849 DVSS.n8882 DVSS.n8880 0.00564286
R31850 DVSS.n10395 DVSS.n10394 0.00564085
R31851 DVSS.n10454 DVSS.n10453 0.00564085
R31852 DVSS.n10497 DVSS.n10496 0.00564085
R31853 DVSS.n16518 DVSS.n16517 0.00560681
R31854 DVSS.n6022 DVSS.n6006 0.00557857
R31855 DVSS.n18253 DVSS.n18252 0.00557042
R31856 DVSS.n18479 DVSS.n18478 0.00557042
R31857 DVSS.n15487 DVSS.n15486 0.00557042
R31858 DVSS.n15123 DVSS.n15122 0.00557042
R31859 DVSS.n10263 DVSS.n10262 0.00552793
R31860 DVSS.n11220 DVSS.n11219 0.00551772
R31861 DVSS.n17649 DVSS.n17648 0.00551772
R31862 DVSS.n9837 DVSS.n9836 0.00551772
R31863 DVSS.n17219 DVSS.n17218 0.00545
R31864 DVSS.n17225 DVSS.n17224 0.00545
R31865 DVSS.n17230 DVSS.n17229 0.00545
R31866 DVSS.n15187 DVSS.n15186 0.00545
R31867 DVSS.n15144 DVSS.n15143 0.00545
R31868 DVSS.n2385 DVSS.n2384 0.00545
R31869 DVSS.n2061 DVSS.n2044 0.00545
R31870 DVSS.n2002 DVSS.n2001 0.00545
R31871 DVSS.n17697 DVSS.n17696 0.00545
R31872 DVSS.n6798 DVSS.n6797 0.00545
R31873 DVSS.n3826 DVSS.n3825 0.00545
R31874 DVSS.n3906 DVSS.n3905 0.00545
R31875 DVSS.n3860 DVSS.n3859 0.00545
R31876 DVSS.n8072 DVSS.n8071 0.00545
R31877 DVSS.n8110 DVSS.n8109 0.00545
R31878 DVSS.n8161 DVSS.n8160 0.00545
R31879 DVSS.n8212 DVSS.n8211 0.00545
R31880 DVSS.n8297 DVSS.n8296 0.00545
R31881 DVSS.n13097 DVSS.n13096 0.00545
R31882 DVSS.n3605 DVSS.n3604 0.00545
R31883 DVSS.n2594 DVSS.n2593 0.00545
R31884 DVSS.n11751 DVSS.n11750 0.00545
R31885 DVSS.n11787 DVSS.n11786 0.00545
R31886 DVSS.n12989 DVSS.n12988 0.00545
R31887 DVSS.n13014 DVSS.n13013 0.00545
R31888 DVSS.n5984 DVSS.n5983 0.00545
R31889 DVSS.n5938 DVSS.n5937 0.00545
R31890 DVSS.n8364 DVSS.n8363 0.00545
R31891 DVSS.n8402 DVSS.n8401 0.00545
R31892 DVSS.n8453 DVSS.n8452 0.00545
R31893 DVSS.n8504 DVSS.n8503 0.00545
R31894 DVSS.n11323 DVSS.n11322 0.00545
R31895 DVSS.n2054 DVSS.n2052 0.00543435
R31896 DVSS.n19167 DVSS.n19158 0.00536486
R31897 DVSS.n19110 DVSS.n19108 0.00536486
R31898 DVSS.n19438 DVSS.n19430 0.00536486
R31899 DVSS.n19385 DVSS.n19383 0.00536486
R31900 DVSS.n20175 DVSS.n20167 0.00536486
R31901 DVSS.n20142 DVSS.n20140 0.00536486
R31902 DVSS.n20446 DVSS.n20438 0.00536486
R31903 DVSS.n20393 DVSS.n20390 0.00536486
R31904 DVSS.n5177 DVSS.n5176 0.00535915
R31905 DVSS.n5139 DVSS.n5138 0.00535915
R31906 DVSS.n5085 DVSS.n5084 0.00535915
R31907 DVSS.n10592 DVSS.n10591 0.00535915
R31908 DVSS.n18118 DVSS.n18117 0.00535915
R31909 DVSS.n18153 DVSS.n18152 0.00535915
R31910 DVSS.n18201 DVSS.n18200 0.00535915
R31911 DVSS.n18434 DVSS.n18433 0.00535915
R31912 DVSS.n15408 DVSS.n15407 0.00535915
R31913 DVSS.n15458 DVSS.n15457 0.00535915
R31914 DVSS.n15539 DVSS.n15538 0.00535915
R31915 DVSS.n15195 DVSS.n15194 0.00535915
R31916 DVSS.n11251 DVSS.n11250 0.00534055
R31917 DVSS.n17614 DVSS.n17613 0.00534055
R31918 DVSS.n11137 DVSS.n11136 0.00534055
R31919 DVSS.n17799 DVSS.n17798 0.00532561
R31920 DVSS.n17773 DVSS.n17772 0.00532561
R31921 DVSS.n17766 DVSS.n17765 0.00532561
R31922 DVSS.n15897 DVSS.n15896 0.00532561
R31923 DVSS.n12772 DVSS.n12771 0.00530769
R31924 DVSS.n12742 DVSS.n12737 0.00530769
R31925 DVSS.n12617 DVSS.n12616 0.00530769
R31926 DVSS.n12592 DVSS.n12587 0.00530769
R31927 DVSS.n12329 DVSS.n12328 0.00530769
R31928 DVSS.n12304 DVSS.n12299 0.00530769
R31929 DVSS.n12237 DVSS.n12236 0.00530769
R31930 DVSS.n21340 DVSS.n21333 0.00530769
R31931 DVSS.n21183 DVSS.n21182 0.00530769
R31932 DVSS.n3384 DVSS.n3383 0.00530769
R31933 DVSS.n2780 DVSS.n2775 0.00530769
R31934 DVSS.n3241 DVSS.n3240 0.00530769
R31935 DVSS.n3216 DVSS.n3211 0.00530769
R31936 DVSS.n2956 DVSS.n2955 0.00530769
R31937 DVSS.n2931 DVSS.n2926 0.00530769
R31938 DVSS.n2864 DVSS.n2863 0.00530769
R31939 DVSS.n891 DVSS.n890 0.00530769
R31940 DVSS.n934 DVSS.n927 0.00530769
R31941 DVSS.n3407 DVSS.n3406 0.00530769
R31942 DVSS.n12781 DVSS.n12780 0.00530769
R31943 DVSS.n4430 DVSS.n4429 0.00528346
R31944 DVSS.n4406 DVSS.n4405 0.00528346
R31945 DVSS.n19187 DVSS.n19186 0.00528346
R31946 DVSS.n19274 DVSS.n19273 0.00528346
R31947 DVSS.n846 DVSS.n845 0.00528346
R31948 DVSS.n1029 DVSS.n1028 0.00528346
R31949 DVSS.n1005 DVSS.n1004 0.00528346
R31950 DVSS.n9531 DVSS.n9530 0.00528346
R31951 DVSS.n9558 DVSS.n9557 0.00528346
R31952 DVSS.n12878 DVSS.n12877 0.00528346
R31953 DVSS.n12851 DVSS.n12850 0.00528346
R31954 DVSS.n12674 DVSS.n12497 0.00528346
R31955 DVSS.n15666 DVSS.n15665 0.00528346
R31956 DVSS.n15639 DVSS.n15638 0.00528346
R31957 DVSS.n20198 DVSS.n20197 0.00528346
R31958 DVSS.n20288 DVSS.n20287 0.00528346
R31959 DVSS.n20829 DVSS.n20828 0.00528346
R31960 DVSS.n20794 DVSS.n20793 0.00528346
R31961 DVSS.n20767 DVSS.n20766 0.00528346
R31962 DVSS.n11569 DVSS.n11568 0.00528346
R31963 DVSS.n11596 DVSS.n11595 0.00528346
R31964 DVSS.n18 DVSS.n17 0.00528346
R31965 DVSS.n45 DVSS.n44 0.00528346
R31966 DVSS.n21527 DVSS.n21526 0.00528346
R31967 DVSS.n21500 DVSS.n21499 0.00528346
R31968 DVSS.n21439 DVSS.n21438 0.00528346
R31969 DVSS.n21412 DVSS.n21411 0.00528346
R31970 DVSS.n4300 DVSS.n4299 0.00528346
R31971 DVSS.n4324 DVSS.n4323 0.00528346
R31972 DVSS.n3487 DVSS.n3486 0.00528346
R31973 DVSS.n3463 DVSS.n3462 0.00528346
R31974 DVSS.n3298 DVSS.n3121 0.00528346
R31975 DVSS.n9663 DVSS.n9662 0.00528346
R31976 DVSS.n9636 DVSS.n9635 0.00528346
R31977 DVSS.n20469 DVSS.n20468 0.00528346
R31978 DVSS.n20562 DVSS.n20561 0.00528346
R31979 DVSS.n21055 DVSS.n21054 0.00528346
R31980 DVSS.n21020 DVSS.n21019 0.00528346
R31981 DVSS.n20993 DVSS.n20992 0.00528346
R31982 DVSS.n16180 DVSS.n16179 0.00528346
R31983 DVSS.n16155 DVSS.n16154 0.00528346
R31984 DVSS.n19458 DVSS.n19457 0.00528346
R31985 DVSS.n19545 DVSS.n19544 0.00528346
R31986 DVSS.n1133 DVSS.n1132 0.00528346
R31987 DVSS.n1244 DVSS.n1243 0.00528346
R31988 DVSS.n1220 DVSS.n1219 0.00528346
R31989 DVSS.n6614 DVSS.n6613 0.00528346
R31990 DVSS.n6639 DVSS.n6638 0.00528346
R31991 DVSS.n3549 DVSS.n3548 0.00528346
R31992 DVSS.n18946 DVSS.n18945 0.00528346
R31993 DVSS.n18993 DVSS.n18992 0.00528346
R31994 DVSS.n524 DVSS.n523 0.00528346
R31995 DVSS.n595 DVSS.n594 0.00528346
R31996 DVSS.n571 DVSS.n570 0.00528346
R31997 DVSS.n948 DVSS.n943 0.00527824
R31998 DVSS.n11760 DVSS.n11759 0.00525714
R31999 DVSS.n16072 DVSS.n16071 0.0052251
R32000 DVSS.n15964 DVSS.n15963 0.0052251
R32001 DVSS.n15398 DVSS.n15397 0.005225
R32002 DVSS.n18293 DVSS.n18292 0.005225
R32003 DVSS.n4580 DVSS.n4579 0.00522222
R32004 DVSS.n11027 DVSS.n11026 0.00522222
R32005 DVSS.n4526 DVSS.n4525 0.00522222
R32006 DVSS.n11198 DVSS.n11197 0.00522222
R32007 DVSS.n5510 DVSS.n5509 0.00522222
R32008 DVSS.n10038 DVSS.n10037 0.00522222
R32009 DVSS.n5185 DVSS.n5184 0.00521831
R32010 DVSS.n5147 DVSS.n5146 0.00521831
R32011 DVSS.n5093 DVSS.n5092 0.00521831
R32012 DVSS.n10885 DVSS.n10884 0.00521831
R32013 DVSS.n11430 DVSS.n11429 0.00520602
R32014 DVSS.n11824 DVSS.n11823 0.00519286
R32015 DVSS.n11883 DVSS.n11882 0.00519286
R32016 DVSS.n21164 DVSS.n21163 0.0051892
R32017 DVSS.n17875 DVSS.n17874 0.00518499
R32018 DVSS.n18016 DVSS.n18015 0.00518499
R32019 DVSS.n18162 DVSS.n18161 0.00518499
R32020 DVSS.n7567 DVSS.n7566 0.00518499
R32021 DVSS.n14446 DVSS.n14445 0.00518499
R32022 DVSS.n15824 DVSS.n15823 0.00518499
R32023 DVSS.n15738 DVSS.n15737 0.00518499
R32024 DVSS.n15578 DVSS.n15577 0.00518499
R32025 DVSS.n15242 DVSS.n15241 0.00518499
R32026 DVSS.n18521 DVSS.n18520 0.00518499
R32027 DVSS.n7762 DVSS.n7761 0.00518499
R32028 DVSS.n10408 DVSS.n10407 0.00514789
R32029 DVSS.n10467 DVSS.n10466 0.00514789
R32030 DVSS.n10899 DVSS.n10898 0.00514789
R32031 DVSS.n16559 DVSS.n16558 0.00514789
R32032 DVSS.n16560 DVSS.n16559 0.00514789
R32033 DVSS.n16564 DVSS.n16563 0.00514789
R32034 DVSS.n16658 DVSS.n16657 0.00514789
R32035 DVSS.n16670 DVSS.n16669 0.00514789
R32036 DVSS.n17730 DVSS.n17729 0.00514789
R32037 DVSS.n18443 DVSS.n18442 0.00514789
R32038 DVSS.n14395 DVSS.n14394 0.00514789
R32039 DVSS.n19721 DVSS.n19720 0.00514789
R32040 DVSS.n16746 DVSS.n16745 0.00514789
R32041 DVSS.n16747 DVSS.n16746 0.00514789
R32042 DVSS.n16751 DVSS.n16750 0.00514789
R32043 DVSS.n17165 DVSS.n17164 0.00514789
R32044 DVSS.n17153 DVSS.n17152 0.00514789
R32045 DVSS.n15933 DVSS.n15932 0.00514789
R32046 DVSS.n15174 DVSS.n15173 0.00514789
R32047 DVSS.n14755 DVSS.n14754 0.00514789
R32048 DVSS.n19940 DVSS.n19939 0.00514789
R32049 DVSS.n11779 DVSS.n11778 0.00512857
R32050 DVSS.n16654 DVSS.n16653 0.0051193
R32051 DVSS.n17169 DVSS.n17168 0.0051193
R32052 DVSS.n18149 DVSS.n18148 0.00511916
R32053 DVSS.n15454 DVSS.n15453 0.00511916
R32054 DVSS.n4433 DVSS.n4432 0.0051063
R32055 DVSS.n4403 DVSS.n4402 0.0051063
R32056 DVSS.n19128 DVSS.n19127 0.0051063
R32057 DVSS.n19190 DVSS.n19189 0.0051063
R32058 DVSS.n19277 DVSS.n19276 0.0051063
R32059 DVSS.n849 DVSS.n848 0.0051063
R32060 DVSS.n1032 DVSS.n1031 0.0051063
R32061 DVSS.n1002 DVSS.n1001 0.0051063
R32062 DVSS.n985 DVSS.n984 0.0051063
R32063 DVSS.n9528 DVSS.n9527 0.0051063
R32064 DVSS.n9561 DVSS.n9560 0.0051063
R32065 DVSS.n12881 DVSS.n12880 0.0051063
R32066 DVSS.n12848 DVSS.n12847 0.0051063
R32067 DVSS.n15669 DVSS.n15668 0.0051063
R32068 DVSS.n15636 DVSS.n15635 0.0051063
R32069 DVSS.n20128 DVSS.n20127 0.0051063
R32070 DVSS.n20201 DVSS.n20200 0.0051063
R32071 DVSS.n20291 DVSS.n20290 0.0051063
R32072 DVSS.n20832 DVSS.n20831 0.0051063
R32073 DVSS.n20797 DVSS.n20796 0.0051063
R32074 DVSS.n20764 DVSS.n20763 0.0051063
R32075 DVSS.n20747 DVSS.n20746 0.0051063
R32076 DVSS.n11566 DVSS.n11565 0.0051063
R32077 DVSS.n11599 DVSS.n11598 0.0051063
R32078 DVSS.n12066 DVSS.n12065 0.0051063
R32079 DVSS.n48 DVSS.n47 0.0051063
R32080 DVSS.n21530 DVSS.n21529 0.0051063
R32081 DVSS.n21497 DVSS.n21496 0.0051063
R32082 DVSS.n21442 DVSS.n21441 0.0051063
R32083 DVSS.n21409 DVSS.n21408 0.0051063
R32084 DVSS.n4297 DVSS.n4296 0.0051063
R32085 DVSS.n4327 DVSS.n4326 0.0051063
R32086 DVSS.n3490 DVSS.n3489 0.0051063
R32087 DVSS.n3460 DVSS.n3459 0.0051063
R32088 DVSS.n9666 DVSS.n9665 0.0051063
R32089 DVSS.n9633 DVSS.n9632 0.0051063
R32090 DVSS.n20411 DVSS.n20410 0.0051063
R32091 DVSS.n20472 DVSS.n20471 0.0051063
R32092 DVSS.n20565 DVSS.n20564 0.0051063
R32093 DVSS.n21058 DVSS.n21057 0.0051063
R32094 DVSS.n21023 DVSS.n21022 0.0051063
R32095 DVSS.n20990 DVSS.n20989 0.0051063
R32096 DVSS.n20973 DVSS.n20972 0.0051063
R32097 DVSS.n16183 DVSS.n16182 0.0051063
R32098 DVSS.n16152 DVSS.n16151 0.0051063
R32099 DVSS.n19402 DVSS.n19401 0.0051063
R32100 DVSS.n19461 DVSS.n19460 0.0051063
R32101 DVSS.n19548 DVSS.n19547 0.0051063
R32102 DVSS.n1136 DVSS.n1135 0.0051063
R32103 DVSS.n1247 DVSS.n1246 0.0051063
R32104 DVSS.n1217 DVSS.n1216 0.0051063
R32105 DVSS.n1201 DVSS.n1200 0.0051063
R32106 DVSS.n6611 DVSS.n6610 0.0051063
R32107 DVSS.n6642 DVSS.n6641 0.0051063
R32108 DVSS.n3552 DVSS.n3551 0.0051063
R32109 DVSS.n18949 DVSS.n18948 0.0051063
R32110 DVSS.n18996 DVSS.n18995 0.0051063
R32111 DVSS.n527 DVSS.n526 0.0051063
R32112 DVSS.n598 DVSS.n597 0.0051063
R32113 DVSS.n568 DVSS.n567 0.0051063
R32114 DVSS.n5265 DVSS.n5264 0.00507746
R32115 DVSS.n5260 DVSS.n5259 0.00507746
R32116 DVSS.n6807 DVSS.n6806 0.00506429
R32117 DVSS.n3929 DVSS.n3928 0.00506429
R32118 DVSS.n3899 DVSS.n3898 0.00506429
R32119 DVSS.n3853 DVSS.n3852 0.00506429
R32120 DVSS.n3625 DVSS.n3614 0.00506429
R32121 DVSS.n2756 DVSS.n2606 0.00506429
R32122 DVSS.n5977 DVSS.n5976 0.00506429
R32123 DVSS.n5931 DVSS.n5930 0.00506429
R32124 DVSS.n16804 DVSS.n16800 0.0050448
R32125 DVSS.n7642 DVSS.n7638 0.0050448
R32126 DVSS.n16012 DVSS.n16011 0.0050448
R32127 DVSS.n15309 DVSS.n15308 0.0050448
R32128 DVSS.n18011 DVSS.n18010 0.0050448
R32129 DVSS.n17870 DVSS.n17869 0.0050448
R32130 DVSS.n17465 DVSS.n17464 0.00504436
R32131 DVSS.n14443 DVSS.n14433 0.00504436
R32132 DVSS.n17878 DVSS.n17877 0.00504436
R32133 DVSS.n18019 DVSS.n18018 0.00504436
R32134 DVSS.n18165 DVSS.n18164 0.00504436
R32135 DVSS.n7570 DVSS.n7569 0.00504436
R32136 DVSS.n17539 DVSS.n15873 0.00504436
R32137 DVSS.n15821 DVSS.n15820 0.00504436
R32138 DVSS.n15741 DVSS.n15740 0.00504436
R32139 DVSS.n15575 DVSS.n15574 0.00504436
R32140 DVSS.n15239 DVSS.n15238 0.00504436
R32141 DVSS.n15884 DVSS.n15883 0.00504436
R32142 DVSS.n14694 DVSS.n14693 0.00504436
R32143 DVSS.n7759 DVSS.n7758 0.00504436
R32144 DVSS.n18518 DVSS.n18517 0.00504436
R32145 DVSS.n17114 DVSS.n16868 0.00504436
R32146 DVSS.n16708 DVSS.n16523 0.00504436
R32147 DVSS.n17298 DVSS.n17297 0.00502514
R32148 DVSS.n17288 DVSS.n17287 0.00502514
R32149 DVSS.n16975 DVSS.n16974 0.00502514
R32150 DVSS.n16990 DVSS.n16988 0.00502514
R32151 DVSS.n10628 DVSS.n10627 0.00502514
R32152 DVSS.n17210 DVSS.n17209 0.005
R32153 DVSS.n15153 DVSS.n15152 0.005
R32154 DVSS.n15111 DVSS.n15110 0.005
R32155 DVSS.n17688 DVSS.n17687 0.005
R32156 DVSS.n8153 DVSS.n8152 0.005
R32157 DVSS.n8204 DVSS.n8203 0.005
R32158 DVSS.n13114 DVSS.n13113 0.005
R32159 DVSS.n13087 DVSS.n13086 0.005
R32160 DVSS.n12968 DVSS.n12967 0.005
R32161 DVSS.n13024 DVSS.n13023 0.005
R32162 DVSS.n8445 DVSS.n8444 0.005
R32163 DVSS.n8496 DVSS.n8495 0.005
R32164 DVSS.n11300 DVSS.n11299 0.005
R32165 DVSS.n14911 DVSS.n14910 0.005
R32166 DVSS.n5306 DVSS.n5305 0.00494444
R32167 DVSS.n5305 DVSS.n5304 0.00494444
R32168 DVSS.n5304 DVSS.n5303 0.00494444
R32169 DVSS.n5303 DVSS.n5302 0.00494444
R32170 DVSS.n5302 DVSS.n5301 0.00494444
R32171 DVSS.n5301 DVSS.n5300 0.00494444
R32172 DVSS.n5300 DVSS.n5299 0.00494444
R32173 DVSS.n5299 DVSS.n5298 0.00494444
R32174 DVSS.n5298 DVSS.n5297 0.00494444
R32175 DVSS.n5297 DVSS.n5296 0.00494444
R32176 DVSS.n5296 DVSS.n5295 0.00494444
R32177 DVSS.n5295 DVSS.n5294 0.00494444
R32178 DVSS.n5294 DVSS.n5293 0.00494444
R32179 DVSS.n5293 DVSS.n5292 0.00494444
R32180 DVSS.n5292 DVSS.n5291 0.00494444
R32181 DVSS.n5291 DVSS.n5290 0.00494444
R32182 DVSS.n5290 DVSS.n5289 0.00494444
R32183 DVSS.n5289 DVSS.n5288 0.00494444
R32184 DVSS.n5288 DVSS.n5287 0.00494444
R32185 DVSS.n5287 DVSS.n5286 0.00494444
R32186 DVSS.n5286 DVSS.n5285 0.00494444
R32187 DVSS.n5285 DVSS.n5284 0.00494444
R32188 DVSS.n5284 DVSS.n5283 0.00494444
R32189 DVSS.n5283 DVSS.n5282 0.00494444
R32190 DVSS.n5282 DVSS.n5281 0.00494444
R32191 DVSS.n5281 DVSS.n5280 0.00494444
R32192 DVSS.n5280 DVSS.n5279 0.00494444
R32193 DVSS.n5279 DVSS.n5278 0.00494444
R32194 DVSS.n5278 DVSS.n5277 0.00494444
R32195 DVSS.n5277 DVSS.n5276 0.00494444
R32196 DVSS.n5276 DVSS.n5275 0.00494444
R32197 DVSS.n5275 DVSS.n5274 0.00494444
R32198 DVSS.n5274 DVSS.n5273 0.00494444
R32199 DVSS.n5273 DVSS.n5272 0.00494444
R32200 DVSS.n5272 DVSS.n5271 0.00494444
R32201 DVSS.n10505 DVSS.n10504 0.00494444
R32202 DVSS.n10506 DVSS.n10505 0.00494444
R32203 DVSS.n10507 DVSS.n10506 0.00494444
R32204 DVSS.n10508 DVSS.n10507 0.00494444
R32205 DVSS.n10509 DVSS.n10508 0.00494444
R32206 DVSS.n10510 DVSS.n10509 0.00494444
R32207 DVSS.n10511 DVSS.n10510 0.00494444
R32208 DVSS.n10512 DVSS.n10511 0.00494444
R32209 DVSS.n10513 DVSS.n10512 0.00494444
R32210 DVSS.n10514 DVSS.n10513 0.00494444
R32211 DVSS.n10515 DVSS.n10514 0.00494444
R32212 DVSS.n10516 DVSS.n10515 0.00494444
R32213 DVSS.n10517 DVSS.n10516 0.00494444
R32214 DVSS.n10518 DVSS.n10517 0.00494444
R32215 DVSS.n10519 DVSS.n10518 0.00494444
R32216 DVSS.n10520 DVSS.n10519 0.00494444
R32217 DVSS.n10521 DVSS.n10520 0.00494444
R32218 DVSS.n10522 DVSS.n10521 0.00494444
R32219 DVSS.n10523 DVSS.n10522 0.00494444
R32220 DVSS.n10524 DVSS.n10523 0.00494444
R32221 DVSS.n10525 DVSS.n10524 0.00494444
R32222 DVSS.n10526 DVSS.n10525 0.00494444
R32223 DVSS.n10527 DVSS.n10526 0.00494444
R32224 DVSS.n10528 DVSS.n10527 0.00494444
R32225 DVSS.n10529 DVSS.n10528 0.00494444
R32226 DVSS.n10530 DVSS.n10529 0.00494444
R32227 DVSS.n10531 DVSS.n10530 0.00494444
R32228 DVSS.n10532 DVSS.n10531 0.00494444
R32229 DVSS.n10533 DVSS.n10532 0.00494444
R32230 DVSS.n10534 DVSS.n10533 0.00494444
R32231 DVSS.n10535 DVSS.n10534 0.00494444
R32232 DVSS.n10536 DVSS.n10535 0.00494444
R32233 DVSS.n10537 DVSS.n10536 0.00494444
R32234 DVSS.n10538 DVSS.n10537 0.00494444
R32235 DVSS.n10539 DVSS.n10538 0.00494444
R32236 DVSS.n10540 DVSS.n10539 0.00494444
R32237 DVSS.n10541 DVSS.n10540 0.00494444
R32238 DVSS.n10542 DVSS.n10541 0.00494444
R32239 DVSS.n10543 DVSS.n10542 0.00494444
R32240 DVSS.n10544 DVSS.n10543 0.00494444
R32241 DVSS.n10545 DVSS.n10544 0.00494444
R32242 DVSS.n10546 DVSS.n10545 0.00494444
R32243 DVSS.n10547 DVSS.n10546 0.00494444
R32244 DVSS.n10548 DVSS.n10547 0.00494444
R32245 DVSS.n10549 DVSS.n10548 0.00494444
R32246 DVSS.n10550 DVSS.n10549 0.00494444
R32247 DVSS.n10551 DVSS.n10550 0.00494444
R32248 DVSS.n10552 DVSS.n10551 0.00494444
R32249 DVSS.n10553 DVSS.n10552 0.00494444
R32250 DVSS.n10554 DVSS.n10553 0.00494444
R32251 DVSS.n10555 DVSS.n10554 0.00494444
R32252 DVSS.n10556 DVSS.n10555 0.00494444
R32253 DVSS.n10557 DVSS.n10556 0.00494444
R32254 DVSS.n10558 DVSS.n10557 0.00494444
R32255 DVSS.n10895 DVSS.n10894 0.00494444
R32256 DVSS.n10894 DVSS.n10893 0.00494444
R32257 DVSS.n10893 DVSS.n10892 0.00494444
R32258 DVSS.n10892 DVSS.n10891 0.00494444
R32259 DVSS.n10891 DVSS.n10890 0.00494444
R32260 DVSS.n10890 DVSS.n10889 0.00494444
R32261 DVSS.n10878 DVSS.n10877 0.00494444
R32262 DVSS.n16548 DVSS.n16547 0.00493662
R32263 DVSS.n16078 DVSS.n16077 0.00493662
R32264 DVSS.n17785 DVSS.n17784 0.00493662
R32265 DVSS.n18106 DVSS.n18105 0.00493662
R32266 DVSS.n18270 DVSS.n18269 0.00493662
R32267 DVSS.n18256 DVSS.n18255 0.00493662
R32268 DVSS.n16735 DVSS.n16734 0.00493662
R32269 DVSS.n15970 DVSS.n15969 0.00493662
R32270 DVSS.n15878 DVSS.n15877 0.00493662
R32271 DVSS.n15384 DVSS.n15383 0.00493662
R32272 DVSS.n15470 DVSS.n15469 0.00493662
R32273 DVSS.n15484 DVSS.n15483 0.00493662
R32274 DVSS.n10718 DVSS.n10717 0.00493571
R32275 DVSS.n8152 DVSS.n8151 0.00493571
R32276 DVSS.n8203 DVSS.n8202 0.00493571
R32277 DVSS.n13114 DVSS.n8288 0.00493571
R32278 DVSS.n13086 DVSS.n8322 0.00493571
R32279 DVSS.n2683 DVSS.n2682 0.00493571
R32280 DVSS.n2629 DVSS.n2628 0.00493571
R32281 DVSS.n12967 DVSS.n11983 0.00493571
R32282 DVSS.n13024 DVSS.n13004 0.00493571
R32283 DVSS.n8444 DVSS.n8443 0.00493571
R32284 DVSS.n8495 DVSS.n8494 0.00493571
R32285 DVSS.n11299 DVSS.n8585 0.00493571
R32286 DVSS.n11305 DVSS.n11304 0.00493571
R32287 DVSS.n8891 DVSS.n8890 0.00493571
R32288 DVSS.n5601 DVSS.n5591 0.00492913
R32289 DVSS.n5647 DVSS.n5646 0.00492913
R32290 DVSS.n5717 DVSS.n5716 0.00492913
R32291 DVSS.n4459 DVSS.n4458 0.00492913
R32292 DVSS.n19255 DVSS.n19254 0.00492913
R32293 DVSS.n874 DVSS.n873 0.00492913
R32294 DVSS.n10284 DVSS.n10275 0.00492913
R32295 DVSS.n10940 DVSS.n10939 0.00492913
R32296 DVSS.n9500 DVSS.n9499 0.00492913
R32297 DVSS.n12909 DVSS.n12908 0.00492913
R32298 DVSS.n12773 DVSS.n12764 0.00492913
R32299 DVSS.n12734 DVSS.n12733 0.00492913
R32300 DVSS.n12443 DVSS.n12442 0.00492913
R32301 DVSS.n12419 DVSS.n12418 0.00492913
R32302 DVSS.n12169 DVSS.n12168 0.00492913
R32303 DVSS.n21231 DVSS.n21230 0.00492913
R32304 DVSS.n21195 DVSS.n21194 0.00492913
R32305 DVSS.n21330 DVSS.n21329 0.00492913
R32306 DVSS.n17023 DVSS.n17014 0.00492913
R32307 DVSS.n17073 DVSS.n17072 0.00492913
R32308 DVSS.n15697 DVSS.n15696 0.00492913
R32309 DVSS.n20266 DVSS.n20265 0.00492913
R32310 DVSS.n20859 DVSS.n20858 0.00492913
R32311 DVSS.n10636 DVSS.n10635 0.00492913
R32312 DVSS.n10822 DVSS.n10821 0.00492913
R32313 DVSS.n11538 DVSS.n11537 0.00492913
R32314 DVSS.n12063 DVSS.n12062 0.00492913
R32315 DVSS.n75 DVSS.n74 0.00492913
R32316 DVSS.n21470 DVSS.n21469 0.00492913
R32317 DVSS.n5231 DVSS.n5230 0.00492913
R32318 DVSS.n4717 DVSS.n4716 0.00492913
R32319 DVSS.n4271 DVSS.n4270 0.00492913
R32320 DVSS.n3733 DVSS.n3732 0.00492913
R32321 DVSS.n3385 DVSS.n3376 0.00492913
R32322 DVSS.n3356 DVSS.n3355 0.00492913
R32323 DVSS.n3070 DVSS.n3069 0.00492913
R32324 DVSS.n3046 DVSS.n3045 0.00492913
R32325 DVSS.n2797 DVSS.n2796 0.00492913
R32326 DVSS.n761 DVSS.n760 0.00492913
R32327 DVSS.n802 DVSS.n801 0.00492913
R32328 DVSS.n728 DVSS.n727 0.00492913
R32329 DVSS.n9919 DVSS.n9918 0.00492913
R32330 DVSS.n9962 DVSS.n9961 0.00492913
R32331 DVSS.n9694 DVSS.n9693 0.00492913
R32332 DVSS.n20540 DVSS.n20539 0.00492913
R32333 DVSS.n21085 DVSS.n21084 0.00492913
R32334 DVSS.n17319 DVSS.n17309 0.00492913
R32335 DVSS.n17366 DVSS.n17365 0.00492913
R32336 DVSS.n16329 DVSS.n16328 0.00492913
R32337 DVSS.n16209 DVSS.n16208 0.00492913
R32338 DVSS.n19526 DVSS.n19525 0.00492913
R32339 DVSS.n1161 DVSS.n1160 0.00492913
R32340 DVSS.n5395 DVSS.n5394 0.00492913
R32341 DVSS.n5442 DVSS.n5441 0.00492913
R32342 DVSS.n6470 DVSS.n6469 0.00492913
R32343 DVSS.n6585 DVSS.n6584 0.00492913
R32344 DVSS.n3658 DVSS.n3657 0.00492913
R32345 DVSS.n18974 DVSS.n18973 0.00492913
R32346 DVSS.n552 DVSS.n551 0.00492913
R32347 DVSS.n12530 DVSS.n12525 0.00492308
R32348 DVSS.n12654 DVSS.n12649 0.00492308
R32349 DVSS.n12366 DVSS.n12361 0.00492308
R32350 DVSS.n12274 DVSS.n12269 0.00492308
R32351 DVSS.n12267 DVSS.n12266 0.00492308
R32352 DVSS.n3154 DVSS.n3149 0.00492308
R32353 DVSS.n3278 DVSS.n3273 0.00492308
R32354 DVSS.n2993 DVSS.n2988 0.00492308
R32355 DVSS.n2901 DVSS.n2896 0.00492308
R32356 DVSS.n2894 DVSS.n2893 0.00492308
R32357 DVSS.n6120 DVSS.n6119 0.00489325
R32358 DVSS.n6114 DVSS.n6113 0.00489325
R32359 DVSS.n6134 DVSS.n6133 0.00489325
R32360 DVSS.n6140 DVSS.n6139 0.00489325
R32361 DVSS.n5069 DVSS.n5068 0.0048662
R32362 DVSS.n2384 DVSS.n2383 0.00482175
R32363 DVSS.n2345 DVSS.n2344 0.00482175
R32364 DVSS.n2383 DVSS.n2382 0.00482175
R32365 DVSS.n14490 DVSS.n14488 0.00480851
R32366 DVSS.n14472 DVSS.n14469 0.00480851
R32367 DVSS.n14081 DVSS.n14080 0.00480851
R32368 DVSS.n14650 DVSS.n14645 0.00480851
R32369 DVSS.n14163 DVSS.n14162 0.00480851
R32370 DVSS.n14743 DVSS.n14742 0.00480851
R32371 DVSS.n10723 DVSS.n10644 0.00480714
R32372 DVSS.n6806 DVSS.n6805 0.00480714
R32373 DVSS.n3928 DVSS.n3927 0.00480714
R32374 DVSS.n3898 DVSS.n3897 0.00480714
R32375 DVSS.n3852 DVSS.n3851 0.00480714
R32376 DVSS.n3625 DVSS.n3624 0.00480714
R32377 DVSS.n2756 DVSS.n2755 0.00480714
R32378 DVSS.n2691 DVSS.n2690 0.00480714
R32379 DVSS.n2637 DVSS.n2636 0.00480714
R32380 DVSS.n5976 DVSS.n5975 0.00480714
R32381 DVSS.n5930 DVSS.n5929 0.00480714
R32382 DVSS.n11339 DVSS.n11338 0.00480714
R32383 DVSS.n8901 DVSS.n8900 0.00480714
R32384 DVSS.n10870 DVSS.n10869 0.00479577
R32385 DVSS.n16093 DVSS.n16092 0.004775
R32386 DVSS.n15434 DVSS.n15433 0.004775
R32387 DVSS.n18278 DVSS.n18277 0.004775
R32388 DVSS.n18327 DVSS.n18326 0.004775
R32389 DVSS.n18348 DVSS.n18347 0.004775
R32390 DVSS.n5349 DVSS.n5348 0.00477374
R32391 DVSS.n4136 DVSS.n4135 0.00476
R32392 DVSS.n4197 DVSS.n4196 0.00476
R32393 DVSS.n4193 DVSS.n4192 0.00476
R32394 DVSS.n4189 DVSS.n4188 0.00476
R32395 DVSS.n4183 DVSS.n4182 0.00476
R32396 DVSS.n9236 DVSS.n9235 0.00476
R32397 DVSS.n9299 DVSS.n9298 0.00476
R32398 DVSS.n9300 DVSS.n9299 0.00476
R32399 DVSS.n4133 DVSS.n4131 0.00476
R32400 DVSS.n4134 DVSS.n4133 0.00476
R32401 DVSS.n4137 DVSS.n4134 0.00476
R32402 DVSS.n4233 DVSS.n4231 0.00476
R32403 DVSS.n4231 DVSS.n4229 0.00476
R32404 DVSS.n4229 DVSS.n4227 0.00476
R32405 DVSS.n4227 DVSS.n4225 0.00476
R32406 DVSS.n4202 DVSS.n4200 0.00476
R32407 DVSS.n4200 DVSS.n4198 0.00476
R32408 DVSS.n4198 DVSS.n4195 0.00476
R32409 DVSS.n4195 DVSS.n4194 0.00476
R32410 DVSS.n4194 DVSS.n4191 0.00476
R32411 DVSS.n4191 DVSS.n4190 0.00476
R32412 DVSS.n4190 DVSS.n4187 0.00476
R32413 DVSS.n4187 DVSS.n4186 0.00476
R32414 DVSS.n4186 DVSS.n4184 0.00476
R32415 DVSS.n4184 DVSS.n4181 0.00476
R32416 DVSS.n4181 DVSS.n4180 0.00476
R32417 DVSS.n4180 DVSS.n4178 0.00476
R32418 DVSS.n4156 DVSS.n4154 0.00476
R32419 DVSS.n4154 DVSS.n4152 0.00476
R32420 DVSS.n4152 DVSS.n4150 0.00476
R32421 DVSS.n4150 DVSS.n4148 0.00476
R32422 DVSS.n9155 DVSS.n9153 0.00476
R32423 DVSS.n9157 DVSS.n9155 0.00476
R32424 DVSS.n9159 DVSS.n9157 0.00476
R32425 DVSS.n9161 DVSS.n9159 0.00476
R32426 DVSS.n9163 DVSS.n9161 0.00476
R32427 DVSS.n9165 DVSS.n9163 0.00476
R32428 DVSS.n9167 DVSS.n9165 0.00476
R32429 DVSS.n9229 DVSS.n9227 0.00476
R32430 DVSS.n9231 DVSS.n9229 0.00476
R32431 DVSS.n9233 DVSS.n9231 0.00476
R32432 DVSS.n9234 DVSS.n9233 0.00476
R32433 DVSS.n9237 DVSS.n9234 0.00476
R32434 DVSS.n9239 DVSS.n9237 0.00476
R32435 DVSS.n9241 DVSS.n9239 0.00476
R32436 DVSS.n9243 DVSS.n9241 0.00476
R32437 DVSS.n9245 DVSS.n9243 0.00476
R32438 DVSS.n9247 DVSS.n9245 0.00476
R32439 DVSS.n9249 DVSS.n9247 0.00476
R32440 DVSS.n9251 DVSS.n9249 0.00476
R32441 DVSS.n9281 DVSS.n9279 0.00476
R32442 DVSS.n9283 DVSS.n9281 0.00476
R32443 DVSS.n9285 DVSS.n9283 0.00476
R32444 DVSS.n9287 DVSS.n9285 0.00476
R32445 DVSS.n9289 DVSS.n9287 0.00476
R32446 DVSS.n9291 DVSS.n9289 0.00476
R32447 DVSS.n9293 DVSS.n9291 0.00476
R32448 DVSS.n9295 DVSS.n9293 0.00476
R32449 DVSS.n9296 DVSS.n9295 0.00476
R32450 DVSS.n9297 DVSS.n9296 0.00476
R32451 DVSS.n9301 DVSS.n9297 0.00476
R32452 DVSS.n9303 DVSS.n9301 0.00476
R32453 DVSS.n9333 DVSS.n9331 0.00476
R32454 DVSS.n9335 DVSS.n9333 0.00476
R32455 DVSS.n9337 DVSS.n9335 0.00476
R32456 DVSS.n9339 DVSS.n9337 0.00476
R32457 DVSS.n9463 DVSS.n9461 0.00476
R32458 DVSS.n9465 DVSS.n9463 0.00476
R32459 DVSS.n9475 DVSS.n9465 0.00476
R32460 DVSS.n12112 DVSS.n12111 0.00476
R32461 DVSS.n12114 DVSS.n12113 0.00476
R32462 DVSS.n12113 DVSS.n12014 0.00476
R32463 DVSS.n5789 DVSS.n5788 0.00475197
R32464 DVSS.n5749 DVSS.n5748 0.00475197
R32465 DVSS.n4063 DVSS.n4062 0.00475197
R32466 DVSS.n11296 DVSS.n11295 0.00475197
R32467 DVSS.n13118 DVSS.n13117 0.00475197
R32468 DVSS.n12940 DVSS.n12939 0.00475197
R32469 DVSS.n12466 DVSS.n12465 0.00475197
R32470 DVSS.n12195 DVSS.n12194 0.00475197
R32471 DVSS.n12188 DVSS.n12187 0.00475197
R32472 DVSS.n21232 DVSS.n21231 0.00475197
R32473 DVSS.n21236 DVSS.n21235 0.00475197
R32474 DVSS.n17569 DVSS.n17568 0.00475197
R32475 DVSS.n15013 DVSS.n15012 0.00475197
R32476 DVSS.n10800 DVSS.n10799 0.00475197
R32477 DVSS.n10747 DVSS.n10746 0.00475197
R32478 DVSS.n11366 DVSS.n11365 0.00475197
R32479 DVSS.n13083 DVSS.n13082 0.00475197
R32480 DVSS.n12032 DVSS.n12031 0.00475197
R32481 DVSS.n3972 DVSS.n3971 0.00475197
R32482 DVSS.n3762 DVSS.n3761 0.00475197
R32483 DVSS.n3092 DVSS.n3091 0.00475197
R32484 DVSS.n2824 DVSS.n2823 0.00475197
R32485 DVSS.n2817 DVSS.n2816 0.00475197
R32486 DVSS.n762 DVSS.n761 0.00475197
R32487 DVSS.n767 DVSS.n766 0.00475197
R32488 DVSS.n11092 DVSS.n11091 0.00475197
R32489 DVSS.n9072 DVSS.n9071 0.00475197
R32490 DVSS.n16410 DVSS.n16409 0.00475197
R32491 DVSS.n16370 DVSS.n16369 0.00475197
R32492 DVSS.n7528 DVSS.n7527 0.00475197
R32493 DVSS.n5464 DVSS.n5463 0.00475197
R32494 DVSS.n5847 DVSS.n5846 0.00475197
R32495 DVSS.n6053 DVSS.n6052 0.00475197
R32496 DVSS.n6820 DVSS.n6819 0.00475197
R32497 DVSS.n3629 DVSS.n3628 0.00475197
R32498 DVSS.n11837 DVSS.n11836 0.00474286
R32499 DVSS.n11896 DVSS.n11895 0.00474286
R32500 DVSS.n17611 DVSS.n17610 0.00473539
R32501 DVSS.n17620 DVSS.n17619 0.00473539
R32502 DVSS.n11134 DVSS.n11133 0.00473539
R32503 DVSS.n11143 DVSS.n11142 0.00473539
R32504 DVSS.n16372 DVSS.n16371 0.00473539
R32505 DVSS.n16363 DVSS.n16362 0.00473539
R32506 DVSS.n16642 DVSS.n16641 0.00472535
R32507 DVSS.n16113 DVSS.n16112 0.00472535
R32508 DVSS.n17746 DVSS.n17745 0.00472535
R32509 DVSS.n17756 DVSS.n17755 0.00472535
R32510 DVSS.n18457 DVSS.n18456 0.00472535
R32511 DVSS.n18489 DVSS.n18488 0.00472535
R32512 DVSS.n18490 DVSS.n18489 0.00472535
R32513 DVSS.n14383 DVSS.n14382 0.00472535
R32514 DVSS.n19751 DVSS.n19750 0.00472535
R32515 DVSS.n17181 DVSS.n17180 0.00472535
R32516 DVSS.n15994 DVSS.n15993 0.00472535
R32517 DVSS.n15917 DVSS.n15916 0.00472535
R32518 DVSS.n15907 DVSS.n15906 0.00472535
R32519 DVSS.n15160 DVSS.n15159 0.00472535
R32520 DVSS.n7730 DVSS.n7729 0.00472535
R32521 DVSS.n7731 DVSS.n7730 0.00472535
R32522 DVSS.n14767 DVSS.n14766 0.00472535
R32523 DVSS.n19976 DVSS.n19975 0.00472535
R32524 DVSS.n5057 DVSS.n5056 0.00467857
R32525 DVSS.n4987 DVSS.n4986 0.00467857
R32526 DVSS.n6042 DVSS.n6041 0.00467857
R32527 DVSS.n6037 DVSS.n6036 0.00467857
R32528 DVSS.n6325 DVSS.n6324 0.00467857
R32529 DVSS.n6285 DVSS.n6284 0.00467857
R32530 DVSS.n9262 DVSS.n9261 0.00467
R32531 DVSS.n9315 DVSS.n9314 0.00467
R32532 DVSS.n17791 DVSS.n17790 0.00465899
R32533 DVSS.n15890 DVSS.n15889 0.00465899
R32534 DVSS.n17665 DVSS.n17664 0.00465899
R32535 DVSS.n17672 DVSS.n7654 0.00465899
R32536 DVSS.n4163 DVSS.n4162 0.00464
R32537 DVSS.n5731 DVSS.n5730 0.00461744
R32538 DVSS.n6519 DVSS.n6518 0.00461744
R32539 DVSS.n9777 DVSS.n9776 0.00461744
R32540 DVSS.n9755 DVSS.n9754 0.00461744
R32541 DVSS.n9585 DVSS.n9584 0.00461744
R32542 DVSS.n9143 DVSS.n9142 0.00461744
R32543 DVSS.n15858 DVSS.n15857 0.00461744
R32544 DVSS.n15717 DVSS.n15716 0.00461744
R32545 DVSS.n15612 DVSS.n15611 0.00461744
R32546 DVSS.n14987 DVSS.n14986 0.00461744
R32547 DVSS.n7134 DVSS.n7133 0.00461744
R32548 DVSS.n10755 DVSS.n10754 0.00461744
R32549 DVSS.n4037 DVSS.n4036 0.00461744
R32550 DVSS.n15041 DVSS.n15040 0.00461744
R32551 DVSS.n13146 DVSS.n13145 0.00461744
R32552 DVSS.n4349 DVSS.n4348 0.00461744
R32553 DVSS.n4121 DVSS.n4120 0.00461744
R32554 DVSS.n3998 DVSS.n3997 0.00461744
R32555 DVSS.n9801 DVSS.n9800 0.00461744
R32556 DVSS.n9714 DVSS.n9713 0.00461744
R32557 DVSS.n9609 DVSS.n9608 0.00461744
R32558 DVSS.n9102 DVSS.n9101 0.00461744
R32559 DVSS.n9044 DVSS.n9043 0.00461744
R32560 DVSS.n13355 DVSS.n13354 0.00461744
R32561 DVSS.n16290 DVSS.n16289 0.00461744
R32562 DVSS.n16251 DVSS.n16250 0.00461744
R32563 DVSS.n16130 DVSS.n16129 0.00461744
R32564 DVSS.n18386 DVSS.n18385 0.00461744
R32565 DVSS.n7502 DVSS.n7501 0.00461744
R32566 DVSS.n4802 DVSS.n4801 0.00461429
R32567 DVSS.n8610 DVSS.n8609 0.00461429
R32568 DVSS.n18428 DVSS.n18427 0.00459139
R32569 DVSS.n15201 DVSS.n15200 0.00459139
R32570 DVSS DVSS.n21360 0.00458
R32571 DVSS.n21365 DVSS 0.00458
R32572 DVSS.n16931 DVSS.n16930 0.00457827
R32573 DVSS.n9887 DVSS.n9886 0.00457827
R32574 DVSS.n5615 DVSS.n5614 0.0045748
R32575 DVSS.n10904 DVSS.n10903 0.0045748
R32576 DVSS.n12698 DVSS.n12697 0.0045748
R32577 DVSS.n12477 DVSS.n12476 0.0045748
R32578 DVSS.n12196 DVSS.n12195 0.0045748
R32579 DVSS.n17037 DVSS.n17036 0.0045748
R32580 DVSS.n10858 DVSS.n10857 0.0045748
R32581 DVSS.n5205 DVSS.n5204 0.0045748
R32582 DVSS.n3321 DVSS.n3320 0.0045748
R32583 DVSS.n3103 DVSS.n3102 0.0045748
R32584 DVSS.n2825 DVSS.n2824 0.0045748
R32585 DVSS.n9926 DVSS.n9925 0.0045748
R32586 DVSS.n17334 DVSS.n17333 0.0045748
R32587 DVSS.n5410 DVSS.n5409 0.0045748
R32588 DVSS.n6322 DVSS.n6321 0.00455714
R32589 DVSS.n6321 DVSS.n6320 0.00455714
R32590 DVSS.n6320 DVSS.n6319 0.00455714
R32591 DVSS.n6319 DVSS.n6318 0.00455714
R32592 DVSS.n6318 DVSS.n6317 0.00455714
R32593 DVSS.n6317 DVSS.n6316 0.00455714
R32594 DVSS.n6316 DVSS.n6315 0.00455714
R32595 DVSS.n6315 DVSS.n6314 0.00455714
R32596 DVSS.n6314 DVSS.n6313 0.00455714
R32597 DVSS.n6313 DVSS.n6312 0.00455714
R32598 DVSS.n6312 DVSS.n6311 0.00455714
R32599 DVSS.n6311 DVSS.n6310 0.00455714
R32600 DVSS.n6310 DVSS.n6309 0.00455714
R32601 DVSS.n6309 DVSS.n6308 0.00455714
R32602 DVSS.n6308 DVSS.n6307 0.00455714
R32603 DVSS.n6307 DVSS.n6306 0.00455714
R32604 DVSS.n6306 DVSS.n6305 0.00455714
R32605 DVSS.n6305 DVSS.n6304 0.00455714
R32606 DVSS.n6304 DVSS.n6303 0.00455714
R32607 DVSS.n6303 DVSS.n6302 0.00455714
R32608 DVSS.n6302 DVSS.n6301 0.00455714
R32609 DVSS.n6301 DVSS.n6300 0.00455714
R32610 DVSS.n6300 DVSS.n6299 0.00455714
R32611 DVSS.n6299 DVSS.n6298 0.00455714
R32612 DVSS.n6298 DVSS.n6297 0.00455714
R32613 DVSS.n6297 DVSS.n6296 0.00455714
R32614 DVSS.n6296 DVSS.n6295 0.00455714
R32615 DVSS.n6295 DVSS.n6294 0.00455714
R32616 DVSS.n6294 DVSS.n6293 0.00455714
R32617 DVSS.n6293 DVSS.n6292 0.00455714
R32618 DVSS.n6292 DVSS.n6291 0.00455714
R32619 DVSS.n6291 DVSS.n6290 0.00455714
R32620 DVSS.n6290 DVSS.n6289 0.00455714
R32621 DVSS.n6289 DVSS.n6288 0.00455714
R32622 DVSS.n8805 DVSS.n8804 0.00455714
R32623 DVSS.n8806 DVSS.n8805 0.00455714
R32624 DVSS.n8807 DVSS.n8806 0.00455714
R32625 DVSS.n8808 DVSS.n8807 0.00455714
R32626 DVSS.n8809 DVSS.n8808 0.00455714
R32627 DVSS.n8810 DVSS.n8809 0.00455714
R32628 DVSS.n8811 DVSS.n8810 0.00455714
R32629 DVSS.n8812 DVSS.n8811 0.00455714
R32630 DVSS.n8813 DVSS.n8812 0.00455714
R32631 DVSS.n8814 DVSS.n8813 0.00455714
R32632 DVSS.n8815 DVSS.n8814 0.00455714
R32633 DVSS.n8816 DVSS.n8815 0.00455714
R32634 DVSS.n8817 DVSS.n8816 0.00455714
R32635 DVSS.n8818 DVSS.n8817 0.00455714
R32636 DVSS.n8819 DVSS.n8818 0.00455714
R32637 DVSS.n8820 DVSS.n8819 0.00455714
R32638 DVSS.n8821 DVSS.n8820 0.00455714
R32639 DVSS.n8822 DVSS.n8821 0.00455714
R32640 DVSS.n8823 DVSS.n8822 0.00455714
R32641 DVSS.n8824 DVSS.n8823 0.00455714
R32642 DVSS.n8825 DVSS.n8824 0.00455714
R32643 DVSS.n8826 DVSS.n8825 0.00455714
R32644 DVSS.n8827 DVSS.n8826 0.00455714
R32645 DVSS.n8828 DVSS.n8827 0.00455714
R32646 DVSS.n8829 DVSS.n8828 0.00455714
R32647 DVSS.n8830 DVSS.n8829 0.00455714
R32648 DVSS.n8831 DVSS.n8830 0.00455714
R32649 DVSS.n8832 DVSS.n8831 0.00455714
R32650 DVSS.n8833 DVSS.n8832 0.00455714
R32651 DVSS.n8834 DVSS.n8833 0.00455714
R32652 DVSS.n8835 DVSS.n8834 0.00455714
R32653 DVSS.n8836 DVSS.n8835 0.00455714
R32654 DVSS.n8837 DVSS.n8836 0.00455714
R32655 DVSS.n8838 DVSS.n8837 0.00455714
R32656 DVSS.n8839 DVSS.n8838 0.00455714
R32657 DVSS.n8840 DVSS.n8839 0.00455714
R32658 DVSS.n8841 DVSS.n8840 0.00455714
R32659 DVSS.n8842 DVSS.n8841 0.00455714
R32660 DVSS.n8843 DVSS.n8842 0.00455714
R32661 DVSS.n8844 DVSS.n8843 0.00455714
R32662 DVSS.n8845 DVSS.n8844 0.00455714
R32663 DVSS.n8846 DVSS.n8845 0.00455714
R32664 DVSS.n8847 DVSS.n8846 0.00455714
R32665 DVSS.n8848 DVSS.n8847 0.00455714
R32666 DVSS.n8849 DVSS.n8848 0.00455714
R32667 DVSS.n8850 DVSS.n8849 0.00455714
R32668 DVSS.n8851 DVSS.n8850 0.00455714
R32669 DVSS.n8852 DVSS.n8851 0.00455714
R32670 DVSS.n8853 DVSS.n8852 0.00455714
R32671 DVSS.n8854 DVSS.n8853 0.00455714
R32672 DVSS.n8855 DVSS.n8854 0.00455714
R32673 DVSS.n8856 DVSS.n8855 0.00455714
R32674 DVSS.n8857 DVSS.n8856 0.00455714
R32675 DVSS.n8858 DVSS.n8857 0.00455714
R32676 DVSS.n8918 DVSS.n8917 0.00455714
R32677 DVSS.n8917 DVSS.n8916 0.00455714
R32678 DVSS.n8916 DVSS.n8915 0.00455714
R32679 DVSS.n8915 DVSS.n8914 0.00455714
R32680 DVSS.n8914 DVSS.n8913 0.00455714
R32681 DVSS.n8913 DVSS.n8912 0.00455714
R32682 DVSS.n8911 DVSS.n8910 0.00455714
R32683 DVSS.n2455 DVSS.n2454 0.00455714
R32684 DVSS.n2454 DVSS.n2453 0.00455714
R32685 DVSS.n2453 DVSS.n2452 0.00455714
R32686 DVSS.n2452 DVSS.n2451 0.00455714
R32687 DVSS.n2451 DVSS.n2450 0.00455714
R32688 DVSS.n2450 DVSS.n2449 0.00455714
R32689 DVSS.n2449 DVSS.n2448 0.00455714
R32690 DVSS.n2448 DVSS.n2447 0.00455714
R32691 DVSS.n2447 DVSS.n2446 0.00455714
R32692 DVSS.n2446 DVSS.n2445 0.00455714
R32693 DVSS.n2445 DVSS.n2444 0.00455714
R32694 DVSS.n2444 DVSS.n2443 0.00455714
R32695 DVSS.n2443 DVSS.n2442 0.00455714
R32696 DVSS.n2442 DVSS.n2441 0.00455714
R32697 DVSS.n2441 DVSS.n2440 0.00455714
R32698 DVSS.n2440 DVSS.n2439 0.00455714
R32699 DVSS.n2439 DVSS.n2438 0.00455714
R32700 DVSS.n2438 DVSS.n2437 0.00455714
R32701 DVSS.n2437 DVSS.n2436 0.00455714
R32702 DVSS.n1555 DVSS.n1554 0.00455714
R32703 DVSS.n1556 DVSS.n1555 0.00455714
R32704 DVSS.n1557 DVSS.n1556 0.00455714
R32705 DVSS.n1558 DVSS.n1557 0.00455714
R32706 DVSS.n1559 DVSS.n1558 0.00455714
R32707 DVSS.n1560 DVSS.n1559 0.00455714
R32708 DVSS.n1561 DVSS.n1560 0.00455714
R32709 DVSS.n1562 DVSS.n1561 0.00455714
R32710 DVSS.n1563 DVSS.n1562 0.00455714
R32711 DVSS.n1564 DVSS.n1563 0.00455714
R32712 DVSS.n1565 DVSS.n1564 0.00455714
R32713 DVSS.n1566 DVSS.n1565 0.00455714
R32714 DVSS.n1567 DVSS.n1566 0.00455714
R32715 DVSS.n1568 DVSS.n1567 0.00455714
R32716 DVSS.n1569 DVSS.n1568 0.00455714
R32717 DVSS.n1570 DVSS.n1569 0.00455714
R32718 DVSS.n1571 DVSS.n1570 0.00455714
R32719 DVSS.n1572 DVSS.n1571 0.00455714
R32720 DVSS.n1574 DVSS.n1572 0.00455714
R32721 DVSS.n1576 DVSS.n1574 0.00455714
R32722 DVSS.n1578 DVSS.n1576 0.00455714
R32723 DVSS.n1580 DVSS.n1578 0.00455714
R32724 DVSS.n1582 DVSS.n1580 0.00455714
R32725 DVSS.n1584 DVSS.n1582 0.00455714
R32726 DVSS.n1586 DVSS.n1584 0.00455714
R32727 DVSS.n1588 DVSS.n1586 0.00455714
R32728 DVSS.n1590 DVSS.n1588 0.00455714
R32729 DVSS.n1592 DVSS.n1590 0.00455714
R32730 DVSS.n1594 DVSS.n1592 0.00455714
R32731 DVSS.n1596 DVSS.n1594 0.00455714
R32732 DVSS.n1598 DVSS.n1596 0.00455714
R32733 DVSS.n1600 DVSS.n1598 0.00455714
R32734 DVSS.n1602 DVSS.n1600 0.00455714
R32735 DVSS.n1604 DVSS.n1602 0.00455714
R32736 DVSS.n1606 DVSS.n1604 0.00455714
R32737 DVSS.n1608 DVSS.n1606 0.00455714
R32738 DVSS.n1610 DVSS.n1608 0.00455714
R32739 DVSS.n1612 DVSS.n1610 0.00455714
R32740 DVSS.n1614 DVSS.n1612 0.00455714
R32741 DVSS.n1616 DVSS.n1614 0.00455714
R32742 DVSS.n1618 DVSS.n1616 0.00455714
R32743 DVSS.n1620 DVSS.n1618 0.00455714
R32744 DVSS.n1622 DVSS.n1620 0.00455714
R32745 DVSS.n1624 DVSS.n1622 0.00455714
R32746 DVSS.n1626 DVSS.n1624 0.00455714
R32747 DVSS.n1628 DVSS.n1626 0.00455714
R32748 DVSS.n1630 DVSS.n1628 0.00455714
R32749 DVSS.n1632 DVSS.n1630 0.00455714
R32750 DVSS.n1634 DVSS.n1632 0.00455714
R32751 DVSS.n1636 DVSS.n1634 0.00455714
R32752 DVSS.n1638 DVSS.n1636 0.00455714
R32753 DVSS.n1640 DVSS.n1638 0.00455714
R32754 DVSS.n1642 DVSS.n1640 0.00455714
R32755 DVSS.n1645 DVSS.n1642 0.00455714
R32756 DVSS.n1648 DVSS.n1645 0.00455714
R32757 DVSS.n1651 DVSS.n1648 0.00455714
R32758 DVSS.n1654 DVSS.n1651 0.00455714
R32759 DVSS.n1657 DVSS.n1654 0.00455714
R32760 DVSS.n1660 DVSS.n1657 0.00455714
R32761 DVSS.n1663 DVSS.n1660 0.00455714
R32762 DVSS.n1666 DVSS.n1663 0.00455714
R32763 DVSS.n1669 DVSS.n1666 0.00455714
R32764 DVSS.n1672 DVSS.n1669 0.00455714
R32765 DVSS.n1675 DVSS.n1672 0.00455714
R32766 DVSS.n1678 DVSS.n1675 0.00455714
R32767 DVSS.n1681 DVSS.n1678 0.00455714
R32768 DVSS.n1684 DVSS.n1681 0.00455714
R32769 DVSS.n1687 DVSS.n1684 0.00455714
R32770 DVSS.n1690 DVSS.n1687 0.00455714
R32771 DVSS.n1693 DVSS.n1690 0.00455714
R32772 DVSS.n1696 DVSS.n1693 0.00455714
R32773 DVSS.n1699 DVSS.n1696 0.00455714
R32774 DVSS.n1702 DVSS.n1699 0.00455714
R32775 DVSS.n1705 DVSS.n1702 0.00455714
R32776 DVSS.n1708 DVSS.n1705 0.00455714
R32777 DVSS.n1709 DVSS.n1708 0.00455714
R32778 DVSS.n1718 DVSS.n1709 0.00455714
R32779 DVSS.n1720 DVSS.n1719 0.00455714
R32780 DVSS.n2018 DVSS.n2017 0.00455714
R32781 DVSS.n2017 DVSS.n2016 0.00455714
R32782 DVSS.n2016 DVSS.n2015 0.00455714
R32783 DVSS.n2015 DVSS.n2014 0.00455714
R32784 DVSS.n2014 DVSS.n2013 0.00455714
R32785 DVSS.n2039 DVSS.n2038 0.00455714
R32786 DVSS.n2040 DVSS.n2039 0.00455714
R32787 DVSS.n2330 DVSS.n2329 0.00455714
R32788 DVSS.n2329 DVSS.n2328 0.00455714
R32789 DVSS.n2328 DVSS.n2327 0.00455714
R32790 DVSS.n2327 DVSS.n2326 0.00455714
R32791 DVSS.n2326 DVSS.n2325 0.00455714
R32792 DVSS.n2325 DVSS.n2324 0.00455714
R32793 DVSS.n2324 DVSS.n2323 0.00455714
R32794 DVSS.n2323 DVSS.n2322 0.00455714
R32795 DVSS.n2322 DVSS.n2321 0.00455714
R32796 DVSS.n2321 DVSS.n2320 0.00455714
R32797 DVSS.n2320 DVSS.n2319 0.00455714
R32798 DVSS.n2319 DVSS.n2318 0.00455714
R32799 DVSS.n2318 DVSS.n2317 0.00455714
R32800 DVSS.n2317 DVSS.n2316 0.00455714
R32801 DVSS.n2316 DVSS.n2315 0.00455714
R32802 DVSS.n2315 DVSS.n2314 0.00455714
R32803 DVSS.n2314 DVSS.n2313 0.00455714
R32804 DVSS.n2313 DVSS.n2312 0.00455714
R32805 DVSS.n2312 DVSS.n2311 0.00455714
R32806 DVSS.n2311 DVSS.n2310 0.00455714
R32807 DVSS.n2310 DVSS.n2309 0.00455714
R32808 DVSS.n2309 DVSS.n2308 0.00455714
R32809 DVSS.n2308 DVSS.n2307 0.00455714
R32810 DVSS.n2307 DVSS.n2306 0.00455714
R32811 DVSS.n2306 DVSS.n2305 0.00455714
R32812 DVSS.n2305 DVSS.n2304 0.00455714
R32813 DVSS.n2304 DVSS.n2303 0.00455714
R32814 DVSS.n2303 DVSS.n2302 0.00455714
R32815 DVSS.n2302 DVSS.n2301 0.00455714
R32816 DVSS.n2301 DVSS.n2300 0.00455714
R32817 DVSS.n2300 DVSS.n2299 0.00455714
R32818 DVSS.n2299 DVSS.n2298 0.00455714
R32819 DVSS.n2298 DVSS.n2297 0.00455714
R32820 DVSS.n2297 DVSS.n2296 0.00455714
R32821 DVSS.n2296 DVSS.n2295 0.00455714
R32822 DVSS.n2295 DVSS.n2294 0.00455714
R32823 DVSS.n2294 DVSS.n2293 0.00455714
R32824 DVSS.n2293 DVSS.n2292 0.00455714
R32825 DVSS.n2292 DVSS.n2291 0.00455714
R32826 DVSS.n2291 DVSS.n2290 0.00455714
R32827 DVSS.n2290 DVSS.n2289 0.00455714
R32828 DVSS.n2289 DVSS.n2288 0.00455714
R32829 DVSS.n2288 DVSS.n2287 0.00455714
R32830 DVSS.n2287 DVSS.n2286 0.00455714
R32831 DVSS.n2286 DVSS.n2285 0.00455714
R32832 DVSS.n2285 DVSS.n2284 0.00455714
R32833 DVSS.n2284 DVSS.n2283 0.00455714
R32834 DVSS.n2283 DVSS.n2282 0.00455714
R32835 DVSS.n2282 DVSS.n2281 0.00455714
R32836 DVSS.n2281 DVSS.n2280 0.00455714
R32837 DVSS.n2280 DVSS.n2279 0.00455714
R32838 DVSS.n2279 DVSS.n2278 0.00455714
R32839 DVSS.n2278 DVSS.n2277 0.00455714
R32840 DVSS.n2277 DVSS.n2276 0.00455714
R32841 DVSS.n2276 DVSS.n2275 0.00455714
R32842 DVSS.n2275 DVSS.n2274 0.00455714
R32843 DVSS.n2274 DVSS.n2273 0.00455714
R32844 DVSS.n2273 DVSS.n2272 0.00455714
R32845 DVSS.n2272 DVSS.n2271 0.00455714
R32846 DVSS.n2271 DVSS.n2270 0.00455714
R32847 DVSS.n2270 DVSS.n2269 0.00455714
R32848 DVSS.n2269 DVSS.n2268 0.00455714
R32849 DVSS.n2268 DVSS.n2267 0.00455714
R32850 DVSS.n2267 DVSS.n2266 0.00455714
R32851 DVSS.n2266 DVSS.n2265 0.00455714
R32852 DVSS.n2265 DVSS.n2264 0.00455714
R32853 DVSS.n2264 DVSS.n2263 0.00455714
R32854 DVSS.n2263 DVSS.n2262 0.00455714
R32855 DVSS.n2262 DVSS.n2261 0.00455714
R32856 DVSS.n2261 DVSS.n2260 0.00455714
R32857 DVSS.n2260 DVSS.n2259 0.00455714
R32858 DVSS.n2259 DVSS.n2258 0.00455714
R32859 DVSS.n2258 DVSS.n2257 0.00455714
R32860 DVSS.n2257 DVSS.n2256 0.00455714
R32861 DVSS.n2256 DVSS.n2255 0.00455714
R32862 DVSS.n2255 DVSS.n2254 0.00455714
R32863 DVSS.n2254 DVSS.n2253 0.00455714
R32864 DVSS.n2253 DVSS.n2252 0.00455714
R32865 DVSS.n2252 DVSS.n2251 0.00455714
R32866 DVSS.n2251 DVSS.n2250 0.00455714
R32867 DVSS.n2250 DVSS.n2249 0.00455714
R32868 DVSS.n2249 DVSS.n2248 0.00455714
R32869 DVSS.n2248 DVSS.n2247 0.00455714
R32870 DVSS.n2247 DVSS.n2246 0.00455714
R32871 DVSS.n2246 DVSS.n2245 0.00455714
R32872 DVSS.n2245 DVSS.n2244 0.00455714
R32873 DVSS.n2244 DVSS.n2243 0.00455714
R32874 DVSS.n2243 DVSS.n2242 0.00455714
R32875 DVSS.n2242 DVSS.n2060 0.00455714
R32876 DVSS.n2060 DVSS.n2057 0.00455714
R32877 DVSS.n4642 DVSS.n4641 0.00455714
R32878 DVSS.n5054 DVSS.n5053 0.00455714
R32879 DVSS.n5053 DVSS.n5052 0.00455714
R32880 DVSS.n5052 DVSS.n5051 0.00455714
R32881 DVSS.n5051 DVSS.n5050 0.00455714
R32882 DVSS.n5050 DVSS.n5049 0.00455714
R32883 DVSS.n5049 DVSS.n5048 0.00455714
R32884 DVSS.n5048 DVSS.n5047 0.00455714
R32885 DVSS.n5047 DVSS.n5046 0.00455714
R32886 DVSS.n5046 DVSS.n5045 0.00455714
R32887 DVSS.n5045 DVSS.n5044 0.00455714
R32888 DVSS.n5044 DVSS.n5043 0.00455714
R32889 DVSS.n5043 DVSS.n5042 0.00455714
R32890 DVSS.n5042 DVSS.n5041 0.00455714
R32891 DVSS.n5041 DVSS.n5040 0.00455714
R32892 DVSS.n5040 DVSS.n5039 0.00455714
R32893 DVSS.n5039 DVSS.n5038 0.00455714
R32894 DVSS.n5038 DVSS.n5037 0.00455714
R32895 DVSS.n5037 DVSS.n5036 0.00455714
R32896 DVSS.n5036 DVSS.n5035 0.00455714
R32897 DVSS.n5035 DVSS.n5034 0.00455714
R32898 DVSS.n5034 DVSS.n5033 0.00455714
R32899 DVSS.n5033 DVSS.n5032 0.00455714
R32900 DVSS.n5032 DVSS.n5031 0.00455714
R32901 DVSS.n5031 DVSS.n5030 0.00455714
R32902 DVSS.n5030 DVSS.n5029 0.00455714
R32903 DVSS.n5029 DVSS.n5028 0.00455714
R32904 DVSS.n5028 DVSS.n5027 0.00455714
R32905 DVSS.n5027 DVSS.n5026 0.00455714
R32906 DVSS.n5026 DVSS.n5025 0.00455714
R32907 DVSS.n5025 DVSS.n5024 0.00455714
R32908 DVSS.n5024 DVSS.n5023 0.00455714
R32909 DVSS.n5023 DVSS.n5022 0.00455714
R32910 DVSS.n5022 DVSS.n5021 0.00455714
R32911 DVSS.n5021 DVSS.n5020 0.00455714
R32912 DVSS.n5020 DVSS.n5019 0.00455714
R32913 DVSS.n5019 DVSS.n5018 0.00455714
R32914 DVSS.n5018 DVSS.n5017 0.00455714
R32915 DVSS.n5017 DVSS.n5016 0.00455714
R32916 DVSS.n5016 DVSS.n5015 0.00455714
R32917 DVSS.n5015 DVSS.n5014 0.00455714
R32918 DVSS.n5014 DVSS.n5013 0.00455714
R32919 DVSS.n5013 DVSS.n5012 0.00455714
R32920 DVSS.n5012 DVSS.n5011 0.00455714
R32921 DVSS.n5011 DVSS.n5010 0.00455714
R32922 DVSS.n5010 DVSS.n5009 0.00455714
R32923 DVSS.n5009 DVSS.n5008 0.00455714
R32924 DVSS.n5008 DVSS.n5007 0.00455714
R32925 DVSS.n5007 DVSS.n5006 0.00455714
R32926 DVSS.n5006 DVSS.n5005 0.00455714
R32927 DVSS.n5005 DVSS.n5004 0.00455714
R32928 DVSS.n5004 DVSS.n5003 0.00455714
R32929 DVSS.n5003 DVSS.n5002 0.00455714
R32930 DVSS.n5002 DVSS.n5001 0.00455714
R32931 DVSS.n5001 DVSS.n5000 0.00455714
R32932 DVSS.n5000 DVSS.n4999 0.00455714
R32933 DVSS.n4999 DVSS.n4998 0.00455714
R32934 DVSS.n4998 DVSS.n4997 0.00455714
R32935 DVSS.n4997 DVSS.n4996 0.00455714
R32936 DVSS.n4996 DVSS.n4995 0.00455714
R32937 DVSS.n4995 DVSS.n4994 0.00455714
R32938 DVSS.n4994 DVSS.n4993 0.00455714
R32939 DVSS.n4993 DVSS.n4992 0.00455714
R32940 DVSS.n4992 DVSS.n4991 0.00455714
R32941 DVSS.n4991 DVSS.n4990 0.00455714
R32942 DVSS.n10662 DVSS.n10661 0.00455714
R32943 DVSS.n10663 DVSS.n10662 0.00455714
R32944 DVSS.n10664 DVSS.n10663 0.00455714
R32945 DVSS.n10665 DVSS.n10664 0.00455714
R32946 DVSS.n10666 DVSS.n10665 0.00455714
R32947 DVSS.n10667 DVSS.n10666 0.00455714
R32948 DVSS.n10668 DVSS.n10667 0.00455714
R32949 DVSS.n10669 DVSS.n10668 0.00455714
R32950 DVSS.n10670 DVSS.n10669 0.00455714
R32951 DVSS.n10671 DVSS.n10670 0.00455714
R32952 DVSS.n10672 DVSS.n10671 0.00455714
R32953 DVSS.n10673 DVSS.n10672 0.00455714
R32954 DVSS.n10674 DVSS.n10673 0.00455714
R32955 DVSS.n10675 DVSS.n10674 0.00455714
R32956 DVSS.n10676 DVSS.n10675 0.00455714
R32957 DVSS.n10677 DVSS.n10676 0.00455714
R32958 DVSS.n10678 DVSS.n10677 0.00455714
R32959 DVSS.n10679 DVSS.n10678 0.00455714
R32960 DVSS.n10680 DVSS.n10679 0.00455714
R32961 DVSS.n10681 DVSS.n10680 0.00455714
R32962 DVSS.n10682 DVSS.n10681 0.00455714
R32963 DVSS.n10683 DVSS.n10682 0.00455714
R32964 DVSS.n10684 DVSS.n10683 0.00455714
R32965 DVSS.n10685 DVSS.n10684 0.00455714
R32966 DVSS.n10686 DVSS.n10685 0.00455714
R32967 DVSS.n10687 DVSS.n10686 0.00455714
R32968 DVSS.n10688 DVSS.n10687 0.00455714
R32969 DVSS.n10689 DVSS.n10688 0.00455714
R32970 DVSS.n10690 DVSS.n10689 0.00455714
R32971 DVSS.n10691 DVSS.n10690 0.00455714
R32972 DVSS.n10692 DVSS.n10691 0.00455714
R32973 DVSS.n10726 DVSS.n10692 0.00455714
R32974 DVSS.n10728 DVSS.n10727 0.00455714
R32975 DVSS.n6812 DVSS.n6811 0.00455714
R32976 DVSS.n6811 DVSS.n6810 0.00455714
R32977 DVSS.n3818 DVSS.n3817 0.00455714
R32978 DVSS.n3819 DVSS.n3818 0.00455714
R32979 DVSS.n3820 DVSS.n3819 0.00455714
R32980 DVSS.n3821 DVSS.n3820 0.00455714
R32981 DVSS.n3964 DVSS.n3963 0.00455714
R32982 DVSS.n3963 DVSS.n3962 0.00455714
R32983 DVSS.n3962 DVSS.n3961 0.00455714
R32984 DVSS.n3961 DVSS.n3960 0.00455714
R32985 DVSS.n3960 DVSS.n3959 0.00455714
R32986 DVSS.n3959 DVSS.n3958 0.00455714
R32987 DVSS.n3958 DVSS.n3957 0.00455714
R32988 DVSS.n3957 DVSS.n3956 0.00455714
R32989 DVSS.n3956 DVSS.n3955 0.00455714
R32990 DVSS.n3955 DVSS.n3954 0.00455714
R32991 DVSS.n3954 DVSS.n3953 0.00455714
R32992 DVSS.n3953 DVSS.n3952 0.00455714
R32993 DVSS.n3952 DVSS.n3951 0.00455714
R32994 DVSS.n3951 DVSS.n3950 0.00455714
R32995 DVSS.n3950 DVSS.n3949 0.00455714
R32996 DVSS.n3949 DVSS.n3948 0.00455714
R32997 DVSS.n3948 DVSS.n3947 0.00455714
R32998 DVSS.n3947 DVSS.n3946 0.00455714
R32999 DVSS.n3946 DVSS.n3945 0.00455714
R33000 DVSS.n3945 DVSS.n3944 0.00455714
R33001 DVSS.n3944 DVSS.n3943 0.00455714
R33002 DVSS.n3943 DVSS.n3942 0.00455714
R33003 DVSS.n3942 DVSS.n3941 0.00455714
R33004 DVSS.n3941 DVSS.n3940 0.00455714
R33005 DVSS.n3940 DVSS.n3939 0.00455714
R33006 DVSS.n3939 DVSS.n3938 0.00455714
R33007 DVSS.n3938 DVSS.n3937 0.00455714
R33008 DVSS.n3937 DVSS.n3936 0.00455714
R33009 DVSS.n3936 DVSS.n3935 0.00455714
R33010 DVSS.n3935 DVSS.n3934 0.00455714
R33011 DVSS.n3934 DVSS.n3933 0.00455714
R33012 DVSS.n3933 DVSS.n3932 0.00455714
R33013 DVSS.n8237 DVSS.n8236 0.00455714
R33014 DVSS.n8238 DVSS.n8237 0.00455714
R33015 DVSS.n8239 DVSS.n8238 0.00455714
R33016 DVSS.n8240 DVSS.n8239 0.00455714
R33017 DVSS.n8241 DVSS.n8240 0.00455714
R33018 DVSS.n8242 DVSS.n8241 0.00455714
R33019 DVSS.n8243 DVSS.n8242 0.00455714
R33020 DVSS.n8244 DVSS.n8243 0.00455714
R33021 DVSS.n8245 DVSS.n8244 0.00455714
R33022 DVSS.n8246 DVSS.n8245 0.00455714
R33023 DVSS.n8247 DVSS.n8246 0.00455714
R33024 DVSS.n8248 DVSS.n8247 0.00455714
R33025 DVSS.n8249 DVSS.n8248 0.00455714
R33026 DVSS.n8250 DVSS.n8249 0.00455714
R33027 DVSS.n8251 DVSS.n8250 0.00455714
R33028 DVSS.n8252 DVSS.n8251 0.00455714
R33029 DVSS.n8253 DVSS.n8252 0.00455714
R33030 DVSS.n8254 DVSS.n8253 0.00455714
R33031 DVSS.n8255 DVSS.n8254 0.00455714
R33032 DVSS.n8256 DVSS.n8255 0.00455714
R33033 DVSS.n8257 DVSS.n8256 0.00455714
R33034 DVSS.n8258 DVSS.n8257 0.00455714
R33035 DVSS.n8259 DVSS.n8258 0.00455714
R33036 DVSS.n8260 DVSS.n8259 0.00455714
R33037 DVSS.n8261 DVSS.n8260 0.00455714
R33038 DVSS.n8262 DVSS.n8261 0.00455714
R33039 DVSS.n8263 DVSS.n8262 0.00455714
R33040 DVSS.n8264 DVSS.n8263 0.00455714
R33041 DVSS.n8265 DVSS.n8264 0.00455714
R33042 DVSS.n8266 DVSS.n8265 0.00455714
R33043 DVSS.n8267 DVSS.n8266 0.00455714
R33044 DVSS.n8268 DVSS.n8267 0.00455714
R33045 DVSS.n8269 DVSS.n8268 0.00455714
R33046 DVSS.n8270 DVSS.n8269 0.00455714
R33047 DVSS.n8271 DVSS.n8270 0.00455714
R33048 DVSS.n8272 DVSS.n8271 0.00455714
R33049 DVSS.n8273 DVSS.n8272 0.00455714
R33050 DVSS.n8274 DVSS.n8273 0.00455714
R33051 DVSS.n8275 DVSS.n8274 0.00455714
R33052 DVSS.n8276 DVSS.n8275 0.00455714
R33053 DVSS.n8277 DVSS.n8276 0.00455714
R33054 DVSS.n8278 DVSS.n8277 0.00455714
R33055 DVSS.n8279 DVSS.n8278 0.00455714
R33056 DVSS.n8280 DVSS.n8279 0.00455714
R33057 DVSS.n8281 DVSS.n8280 0.00455714
R33058 DVSS.n8282 DVSS.n8281 0.00455714
R33059 DVSS.n8283 DVSS.n8282 0.00455714
R33060 DVSS.n8284 DVSS.n8283 0.00455714
R33061 DVSS.n8285 DVSS.n8284 0.00455714
R33062 DVSS.n13110 DVSS.n13109 0.00455714
R33063 DVSS.n13109 DVSS.n13108 0.00455714
R33064 DVSS.n13108 DVSS.n13107 0.00455714
R33065 DVSS.n13107 DVSS.n13106 0.00455714
R33066 DVSS.n13106 DVSS.n13105 0.00455714
R33067 DVSS.n13105 DVSS.n13104 0.00455714
R33068 DVSS.n13104 DVSS.n13103 0.00455714
R33069 DVSS.n13102 DVSS.n8292 0.00455714
R33070 DVSS.n3610 DVSS.n3609 0.00455714
R33071 DVSS.n3622 DVSS.n3621 0.00455714
R33072 DVSS.n3621 DVSS.n3620 0.00455714
R33073 DVSS.n2600 DVSS.n2599 0.00455714
R33074 DVSS.n2601 DVSS.n2600 0.00455714
R33075 DVSS.n2602 DVSS.n2601 0.00455714
R33076 DVSS.n2603 DVSS.n2602 0.00455714
R33077 DVSS.n2753 DVSS.n2752 0.00455714
R33078 DVSS.n2752 DVSS.n2751 0.00455714
R33079 DVSS.n2751 DVSS.n2750 0.00455714
R33080 DVSS.n2750 DVSS.n2749 0.00455714
R33081 DVSS.n2749 DVSS.n2748 0.00455714
R33082 DVSS.n2748 DVSS.n2747 0.00455714
R33083 DVSS.n2747 DVSS.n2746 0.00455714
R33084 DVSS.n2746 DVSS.n2745 0.00455714
R33085 DVSS.n2745 DVSS.n2744 0.00455714
R33086 DVSS.n2744 DVSS.n2743 0.00455714
R33087 DVSS.n2743 DVSS.n2742 0.00455714
R33088 DVSS.n2742 DVSS.n2741 0.00455714
R33089 DVSS.n2741 DVSS.n2740 0.00455714
R33090 DVSS.n2740 DVSS.n2739 0.00455714
R33091 DVSS.n2739 DVSS.n2738 0.00455714
R33092 DVSS.n2738 DVSS.n2737 0.00455714
R33093 DVSS.n2737 DVSS.n2736 0.00455714
R33094 DVSS.n2736 DVSS.n2735 0.00455714
R33095 DVSS.n2735 DVSS.n2734 0.00455714
R33096 DVSS.n2734 DVSS.n2733 0.00455714
R33097 DVSS.n2733 DVSS.n2732 0.00455714
R33098 DVSS.n2732 DVSS.n2731 0.00455714
R33099 DVSS.n2731 DVSS.n2730 0.00455714
R33100 DVSS.n2730 DVSS.n2729 0.00455714
R33101 DVSS.n2729 DVSS.n2728 0.00455714
R33102 DVSS.n2728 DVSS.n2727 0.00455714
R33103 DVSS.n2727 DVSS.n2726 0.00455714
R33104 DVSS.n2726 DVSS.n2725 0.00455714
R33105 DVSS.n2725 DVSS.n2724 0.00455714
R33106 DVSS.n2724 DVSS.n2723 0.00455714
R33107 DVSS.n2723 DVSS.n2722 0.00455714
R33108 DVSS.n11932 DVSS.n11931 0.00455714
R33109 DVSS.n11933 DVSS.n11932 0.00455714
R33110 DVSS.n11934 DVSS.n11933 0.00455714
R33111 DVSS.n11935 DVSS.n11934 0.00455714
R33112 DVSS.n11936 DVSS.n11935 0.00455714
R33113 DVSS.n11937 DVSS.n11936 0.00455714
R33114 DVSS.n11938 DVSS.n11937 0.00455714
R33115 DVSS.n11939 DVSS.n11938 0.00455714
R33116 DVSS.n11940 DVSS.n11939 0.00455714
R33117 DVSS.n11941 DVSS.n11940 0.00455714
R33118 DVSS.n11942 DVSS.n11941 0.00455714
R33119 DVSS.n11943 DVSS.n11942 0.00455714
R33120 DVSS.n11944 DVSS.n11943 0.00455714
R33121 DVSS.n11945 DVSS.n11944 0.00455714
R33122 DVSS.n11946 DVSS.n11945 0.00455714
R33123 DVSS.n11947 DVSS.n11946 0.00455714
R33124 DVSS.n11948 DVSS.n11947 0.00455714
R33125 DVSS.n11949 DVSS.n11948 0.00455714
R33126 DVSS.n11950 DVSS.n11949 0.00455714
R33127 DVSS.n11951 DVSS.n11950 0.00455714
R33128 DVSS.n11952 DVSS.n11951 0.00455714
R33129 DVSS.n11953 DVSS.n11952 0.00455714
R33130 DVSS.n11954 DVSS.n11953 0.00455714
R33131 DVSS.n11955 DVSS.n11954 0.00455714
R33132 DVSS.n11956 DVSS.n11955 0.00455714
R33133 DVSS.n11957 DVSS.n11956 0.00455714
R33134 DVSS.n11958 DVSS.n11957 0.00455714
R33135 DVSS.n11959 DVSS.n11958 0.00455714
R33136 DVSS.n11960 DVSS.n11959 0.00455714
R33137 DVSS.n11961 DVSS.n11960 0.00455714
R33138 DVSS.n11962 DVSS.n11961 0.00455714
R33139 DVSS.n11963 DVSS.n11962 0.00455714
R33140 DVSS.n11964 DVSS.n11963 0.00455714
R33141 DVSS.n11965 DVSS.n11964 0.00455714
R33142 DVSS.n11966 DVSS.n11965 0.00455714
R33143 DVSS.n11967 DVSS.n11966 0.00455714
R33144 DVSS.n11968 DVSS.n11967 0.00455714
R33145 DVSS.n11969 DVSS.n11968 0.00455714
R33146 DVSS.n11970 DVSS.n11969 0.00455714
R33147 DVSS.n11971 DVSS.n11970 0.00455714
R33148 DVSS.n11972 DVSS.n11971 0.00455714
R33149 DVSS.n11973 DVSS.n11972 0.00455714
R33150 DVSS.n11974 DVSS.n11973 0.00455714
R33151 DVSS.n11975 DVSS.n11974 0.00455714
R33152 DVSS.n11976 DVSS.n11975 0.00455714
R33153 DVSS.n11977 DVSS.n11976 0.00455714
R33154 DVSS.n11978 DVSS.n11977 0.00455714
R33155 DVSS.n11979 DVSS.n11978 0.00455714
R33156 DVSS.n11980 DVSS.n11979 0.00455714
R33157 DVSS.n12995 DVSS.n12994 0.00455714
R33158 DVSS.n12996 DVSS.n12995 0.00455714
R33159 DVSS.n12997 DVSS.n12996 0.00455714
R33160 DVSS.n12998 DVSS.n12997 0.00455714
R33161 DVSS.n12999 DVSS.n12998 0.00455714
R33162 DVSS.n13001 DVSS.n13000 0.00455714
R33163 DVSS.n13020 DVSS.n13019 0.00455714
R33164 DVSS.n5909 DVSS.n5908 0.00455714
R33165 DVSS.n5908 DVSS.n5907 0.00455714
R33166 DVSS.n5907 DVSS.n5906 0.00455714
R33167 DVSS.n5906 DVSS.n5905 0.00455714
R33168 DVSS.n5905 DVSS.n5904 0.00455714
R33169 DVSS.n5904 DVSS.n5903 0.00455714
R33170 DVSS.n5903 DVSS.n5902 0.00455714
R33171 DVSS.n5902 DVSS.n5901 0.00455714
R33172 DVSS.n5901 DVSS.n5900 0.00455714
R33173 DVSS.n5900 DVSS.n5899 0.00455714
R33174 DVSS.n5899 DVSS.n5898 0.00455714
R33175 DVSS.n5898 DVSS.n5897 0.00455714
R33176 DVSS.n5897 DVSS.n5896 0.00455714
R33177 DVSS.n5896 DVSS.n5895 0.00455714
R33178 DVSS.n5895 DVSS.n5894 0.00455714
R33179 DVSS.n5894 DVSS.n5893 0.00455714
R33180 DVSS.n5893 DVSS.n5892 0.00455714
R33181 DVSS.n5892 DVSS.n5891 0.00455714
R33182 DVSS.n5891 DVSS.n5890 0.00455714
R33183 DVSS.n5890 DVSS.n5889 0.00455714
R33184 DVSS.n5889 DVSS.n5888 0.00455714
R33185 DVSS.n5888 DVSS.n5887 0.00455714
R33186 DVSS.n5887 DVSS.n5886 0.00455714
R33187 DVSS.n5886 DVSS.n5885 0.00455714
R33188 DVSS.n5885 DVSS.n5884 0.00455714
R33189 DVSS.n5884 DVSS.n5883 0.00455714
R33190 DVSS.n5883 DVSS.n5882 0.00455714
R33191 DVSS.n5882 DVSS.n5881 0.00455714
R33192 DVSS.n5881 DVSS.n5880 0.00455714
R33193 DVSS.n5880 DVSS.n5879 0.00455714
R33194 DVSS.n5879 DVSS.n5878 0.00455714
R33195 DVSS.n5878 DVSS.n5877 0.00455714
R33196 DVSS.n5877 DVSS.n5876 0.00455714
R33197 DVSS.n5876 DVSS.n5875 0.00455714
R33198 DVSS.n5875 DVSS.n5874 0.00455714
R33199 DVSS.n8529 DVSS.n8528 0.00455714
R33200 DVSS.n8530 DVSS.n8529 0.00455714
R33201 DVSS.n8531 DVSS.n8530 0.00455714
R33202 DVSS.n8532 DVSS.n8531 0.00455714
R33203 DVSS.n8533 DVSS.n8532 0.00455714
R33204 DVSS.n8534 DVSS.n8533 0.00455714
R33205 DVSS.n8535 DVSS.n8534 0.00455714
R33206 DVSS.n8536 DVSS.n8535 0.00455714
R33207 DVSS.n8537 DVSS.n8536 0.00455714
R33208 DVSS.n8538 DVSS.n8537 0.00455714
R33209 DVSS.n8539 DVSS.n8538 0.00455714
R33210 DVSS.n8540 DVSS.n8539 0.00455714
R33211 DVSS.n8541 DVSS.n8540 0.00455714
R33212 DVSS.n8542 DVSS.n8541 0.00455714
R33213 DVSS.n8543 DVSS.n8542 0.00455714
R33214 DVSS.n8544 DVSS.n8543 0.00455714
R33215 DVSS.n8545 DVSS.n8544 0.00455714
R33216 DVSS.n8546 DVSS.n8545 0.00455714
R33217 DVSS.n8547 DVSS.n8546 0.00455714
R33218 DVSS.n8548 DVSS.n8547 0.00455714
R33219 DVSS.n8549 DVSS.n8548 0.00455714
R33220 DVSS.n8550 DVSS.n8549 0.00455714
R33221 DVSS.n8551 DVSS.n8550 0.00455714
R33222 DVSS.n8552 DVSS.n8551 0.00455714
R33223 DVSS.n8553 DVSS.n8552 0.00455714
R33224 DVSS.n8554 DVSS.n8553 0.00455714
R33225 DVSS.n8555 DVSS.n8554 0.00455714
R33226 DVSS.n8556 DVSS.n8555 0.00455714
R33227 DVSS.n8557 DVSS.n8556 0.00455714
R33228 DVSS.n8558 DVSS.n8557 0.00455714
R33229 DVSS.n8559 DVSS.n8558 0.00455714
R33230 DVSS.n8560 DVSS.n8559 0.00455714
R33231 DVSS.n8561 DVSS.n8560 0.00455714
R33232 DVSS.n8562 DVSS.n8561 0.00455714
R33233 DVSS.n8563 DVSS.n8562 0.00455714
R33234 DVSS.n8564 DVSS.n8563 0.00455714
R33235 DVSS.n8565 DVSS.n8564 0.00455714
R33236 DVSS.n8566 DVSS.n8565 0.00455714
R33237 DVSS.n8567 DVSS.n8566 0.00455714
R33238 DVSS.n8568 DVSS.n8567 0.00455714
R33239 DVSS.n8569 DVSS.n8568 0.00455714
R33240 DVSS.n8570 DVSS.n8569 0.00455714
R33241 DVSS.n8571 DVSS.n8570 0.00455714
R33242 DVSS.n8572 DVSS.n8571 0.00455714
R33243 DVSS.n8573 DVSS.n8572 0.00455714
R33244 DVSS.n8574 DVSS.n8573 0.00455714
R33245 DVSS.n8575 DVSS.n8574 0.00455714
R33246 DVSS.n8576 DVSS.n8575 0.00455714
R33247 DVSS.n8577 DVSS.n8576 0.00455714
R33248 DVSS.n8578 DVSS.n8577 0.00455714
R33249 DVSS.n8579 DVSS.n8578 0.00455714
R33250 DVSS.n8580 DVSS.n8579 0.00455714
R33251 DVSS.n8581 DVSS.n8580 0.00455714
R33252 DVSS.n8582 DVSS.n8581 0.00455714
R33253 DVSS.n11329 DVSS.n11328 0.00455714
R33254 DVSS.n11330 DVSS.n11329 0.00455714
R33255 DVSS.n11331 DVSS.n11330 0.00455714
R33256 DVSS.n11332 DVSS.n11331 0.00455714
R33257 DVSS.n11333 DVSS.n11332 0.00455714
R33258 DVSS.n11334 DVSS.n11333 0.00455714
R33259 DVSS.n11357 DVSS.n11356 0.00455714
R33260 DVSS.n7714 DVSS.n7713 0.00455
R33261 DVSS.n16045 DVSS.n16044 0.00455
R33262 DVSS.n6024 DVSS.n6022 0.00455
R33263 DVSS.n10209 DVSS.n10208 0.0045432
R33264 DVSS.n16954 DVSS.n16953 0.0045432
R33265 DVSS.n9910 DVSS.n9909 0.0045432
R33266 DVSS.n12517 DVSS.n12516 0.00453846
R33267 DVSS.n12641 DVSS.n12640 0.00453846
R33268 DVSS.n12624 DVSS.n12619 0.00453846
R33269 DVSS.n12353 DVSS.n12352 0.00453846
R33270 DVSS.n12336 DVSS.n12331 0.00453846
R33271 DVSS.n21323 DVSS.n21318 0.00453846
R33272 DVSS.n21183 DVSS.n21161 0.00453846
R33273 DVSS.n3141 DVSS.n3140 0.00453846
R33274 DVSS.n3265 DVSS.n3264 0.00453846
R33275 DVSS.n3248 DVSS.n3243 0.00453846
R33276 DVSS.n2980 DVSS.n2979 0.00453846
R33277 DVSS.n2963 DVSS.n2958 0.00453846
R33278 DVSS.n898 DVSS.n893 0.00453846
R33279 DVSS.n927 DVSS.n926 0.00453846
R33280 DVSS.n3410 DVSS.n3409 0.00453846
R33281 DVSS.n12791 DVSS.n12783 0.00453846
R33282 DVSS.n9198 DVSS.n9197 0.00452
R33283 DVSS.n9196 DVSS.n9195 0.00452
R33284 DVSS.n14258 DVSS.n14257 0.00451837
R33285 DVSS.n14283 DVSS.n14282 0.00451837
R33286 DVSS.n14312 DVSS.n14311 0.00451837
R33287 DVSS.n17456 DVSS.n16121 0.00451837
R33288 DVSS.n14398 DVSS.n14397 0.00451837
R33289 DVSS.n14857 DVSS.n14856 0.00451837
R33290 DVSS.n14840 DVSS.n14839 0.00451837
R33291 DVSS.n14823 DVSS.n14822 0.00451837
R33292 DVSS.n14752 DVSS.n14729 0.00451837
R33293 DVSS.n17537 DVSS.n16002 0.00451837
R33294 DVSS.n15881 DVSS.n15880 0.00451837
R33295 DVSS.n14691 DVSS.n14675 0.00451837
R33296 DVSS.n16508 DVSS.n16507 0.00451408
R33297 DVSS.n16106 DVSS.n16105 0.00451408
R33298 DVSS.n16103 DVSS.n16102 0.00451408
R33299 DVSS.n16060 DVSS.n16059 0.00451408
R33300 DVSS.n18129 DVSS.n18128 0.00451408
R33301 DVSS.n18132 DVSS.n18131 0.00451408
R33302 DVSS.n18137 DVSS.n18136 0.00451408
R33303 DVSS.n18220 DVSS.n18219 0.00451408
R33304 DVSS.n18187 DVSS.n18186 0.00451408
R33305 DVSS.n18432 DVSS.n18431 0.00451408
R33306 DVSS.n18480 DVSS.n18479 0.00451408
R33307 DVSS.n14519 DVSS.n14518 0.00451408
R33308 DVSS.n19809 DVSS.n19808 0.00451408
R33309 DVSS.n250 DVSS.n249 0.00451408
R33310 DVSS.n16854 DVSS.n16853 0.00451408
R33311 DVSS.n15987 DVSS.n15986 0.00451408
R33312 DVSS.n15984 DVSS.n15983 0.00451408
R33313 DVSS.n15952 DVSS.n15951 0.00451408
R33314 DVSS.n15419 DVSS.n15418 0.00451408
R33315 DVSS.n15422 DVSS.n15421 0.00451408
R33316 DVSS.n15442 DVSS.n15441 0.00451408
R33317 DVSS.n15520 DVSS.n15519 0.00451408
R33318 DVSS.n15553 DVSS.n15552 0.00451408
R33319 DVSS.n15197 DVSS.n15196 0.00451408
R33320 DVSS.n15122 DVSS.n15121 0.00451408
R33321 DVSS.n14616 DVSS.n14615 0.00451408
R33322 DVSS.n20034 DVSS.n20033 0.00451408
R33323 DVSS.n458 DVSS.n457 0.00451408
R33324 DVSS.n1719 VSS 0.0045
R33325 DVSS.n5813 DVSS.n5712 0.00449949
R33326 DVSS.n6529 DVSS.n6528 0.00449949
R33327 DVSS.n4384 DVSS.n4383 0.00449949
R33328 DVSS.n4088 DVSS.n4087 0.00449949
R33329 DVSS.n6516 DVSS.n6515 0.00449949
R33330 DVSS.n11045 DVSS.n11002 0.00449949
R33331 DVSS.n9774 DVSS.n9773 0.00449949
R33332 DVSS.n9758 DVSS.n9757 0.00449949
R33333 DVSS.n9582 DVSS.n9581 0.00449949
R33334 DVSS.n9146 DVSS.n9145 0.00449949
R33335 DVSS.n11237 DVSS.n11236 0.00449949
R33336 DVSS.n16904 DVSS.n16903 0.00449949
R33337 DVSS.n15861 DVSS.n15860 0.00449949
R33338 DVSS.n15714 DVSS.n15713 0.00449949
R33339 DVSS.n15615 DVSS.n15614 0.00449949
R33340 DVSS.n14984 DVSS.n14983 0.00449949
R33341 DVSS.n17628 DVSS.n17627 0.00449949
R33342 DVSS.n7131 DVSS.n7118 0.00449949
R33343 DVSS.n4040 DVSS.n4039 0.00449949
R33344 DVSS.n15038 DVSS.n15037 0.00449949
R33345 DVSS.n13143 DVSS.n13142 0.00449949
R33346 DVSS.n5678 DVSS.n5677 0.00449949
R33347 DVSS.n10969 DVSS.n10968 0.00449949
R33348 DVSS.n17101 DVSS.n16937 0.00449949
R33349 DVSS.n4346 DVSS.n4345 0.00449949
R33350 DVSS.n4124 DVSS.n4123 0.00449949
R33351 DVSS.n3995 DVSS.n3994 0.00449949
R33352 DVSS.n11067 DVSS.n9840 0.00449949
R33353 DVSS.n9804 DVSS.n9803 0.00449949
R33354 DVSS.n9711 DVSS.n9710 0.00449949
R33355 DVSS.n9612 DVSS.n9611 0.00449949
R33356 DVSS.n9099 DVSS.n9098 0.00449949
R33357 DVSS.n9047 DVSS.n9046 0.00449949
R33358 DVSS.n11151 DVSS.n11150 0.00449949
R33359 DVSS.n9990 DVSS.n9893 0.00449949
R33360 DVSS.n13352 DVSS.n13269 0.00449949
R33361 DVSS.n16293 DVSS.n16292 0.00449949
R33362 DVSS.n16254 DVSS.n16253 0.00449949
R33363 DVSS.n16133 DVSS.n16132 0.00449949
R33364 DVSS.n18383 DVSS.n18382 0.00449949
R33365 DVSS.n7505 DVSS.n7504 0.00449949
R33366 DVSS.n16355 DVSS.n16354 0.00449949
R33367 DVSS.n18647 DVSS.n18636 0.00449949
R33368 DVSS.n18679 DVSS.n18663 0.00449949
R33369 DVSS.n18620 DVSS.n18609 0.00449949
R33370 DVSS.n17397 DVSS.n17396 0.00449949
R33371 DVSS.n17446 DVSS.n17431 0.00449949
R33372 DVSS.n6471 DVSS.n6348 0.00449949
R33373 DVSS.n5836 DVSS.n4528 0.00449949
R33374 DVSS.n19655 DVSS.n19654 0.00448591
R33375 DVSS.n19864 DVSS.n19863 0.00448591
R33376 DVSS.n4634 DVSS.n4633 0.00448571
R33377 DVSS.n4755 DVSS.n4754 0.00448571
R33378 DVSS.n10055 DVSS.n10054 0.00448571
R33379 DVSS.n10120 DVSS.n10119 0.00448571
R33380 DVSS.n10168 DVSS.n10167 0.00448571
R33381 DVSS.n5870 DVSS.n5869 0.00448571
R33382 DVSS.n6097 DVSS.n6096 0.00448571
R33383 DVSS.n8655 DVSS.n8654 0.00448571
R33384 DVSS.n8691 DVSS.n8690 0.00448571
R33385 DVSS.n8752 DVSS.n8751 0.00448571
R33386 DVSS.n8797 DVSS.n8796 0.00448571
R33387 DVSS DVSS.n13102 0.00447143
R33388 DVSS.n5239 DVSS.n5238 0.00444366
R33389 DVSS.n5156 DVSS.n5155 0.00444366
R33390 DVSS.n5102 DVSS.n5101 0.00444366
R33391 DVSS.n10325 DVSS.n10324 0.00444366
R33392 DVSS.n10654 DVSS.n10653 0.00442143
R33393 DVSS.n6026 DVSS.n6024 0.00442143
R33394 DVSS.n11349 DVSS.n11348 0.00442143
R33395 DVSS.n8334 DVSS.n8333 0.00442143
R33396 DVSS.n6995 DVSS.n6994 0.00439764
R33397 DVSS.n19204 DVSS.n19203 0.00439764
R33398 DVSS.n21312 DVSS.n21311 0.00439764
R33399 DVSS.n21279 DVSS.n21278 0.00439764
R33400 DVSS.n21184 DVSS.n21144 0.00439764
R33401 DVSS.n13643 DVSS.n13642 0.00439764
R33402 DVSS.n20215 DVSS.n20214 0.00439764
R33403 DVSS.n782 DVSS.n781 0.00439764
R33404 DVSS.n656 DVSS.n655 0.00439764
R33405 DVSS.n698 DVSS.n697 0.00439764
R33406 DVSS.n13232 DVSS.n13231 0.00439764
R33407 DVSS.n20486 DVSS.n20485 0.00439764
R33408 DVSS.n18762 DVSS.n18761 0.00439764
R33409 DVSS.n19475 DVSS.n19474 0.00439764
R33410 DVSS.n16542 DVSS.n16541 0.00437965
R33411 DVSS.n16729 DVSS.n16728 0.00437965
R33412 DVSS.n14255 DVSS.n14246 0.00437774
R33413 DVSS.n14280 DVSS.n14271 0.00437774
R33414 DVSS.n14309 DVSS.n14296 0.00437774
R33415 DVSS.n14860 DVSS.n14859 0.00437774
R33416 DVSS.n14843 DVSS.n14842 0.00437774
R33417 DVSS.n14826 DVSS.n14825 0.00437774
R33418 DVSS.n10417 DVSS.n10416 0.00437324
R33419 DVSS.n10476 DVSS.n10475 0.00437324
R33420 DVSS.n10572 DVSS.n10571 0.00437324
R33421 DVSS.n2360 DVSS.n2359 0.00437247
R33422 DVSS.n2406 DVSS.n2405 0.00437247
R33423 DVSS.n16599 DVSS.n16598 0.004325
R33424 DVSS.n16604 DVSS.n16603 0.004325
R33425 DVSS.n18312 DVSS.n18311 0.004325
R33426 DVSS.n18317 DVSS.n18316 0.004325
R33427 DVSS.n16679 DVSS.n16678 0.00430282
R33428 DVSS.n16693 DVSS.n16692 0.00430282
R33429 DVSS.n18122 DVSS.n18121 0.00430282
R33430 DVSS.n18204 DVSS.n18203 0.00430282
R33431 DVSS.n19700 DVSS.n19699 0.00430282
R33432 DVSS.n19779 DVSS.n19778 0.00430282
R33433 DVSS.n131 DVSS.n130 0.00430282
R33434 DVSS.n220 DVSS.n219 0.00430282
R33435 DVSS.n201 DVSS.n200 0.00430282
R33436 DVSS.n17144 DVSS.n17143 0.00430282
R33437 DVSS.n17130 DVSS.n17129 0.00430282
R33438 DVSS.n15412 DVSS.n15411 0.00430282
R33439 DVSS.n15536 DVSS.n15535 0.00430282
R33440 DVSS.n19919 DVSS.n19918 0.00430282
R33441 DVSS.n20004 DVSS.n20003 0.00430282
R33442 DVSS.n291 DVSS.n290 0.00430282
R33443 DVSS.n428 DVSS.n427 0.00430282
R33444 DVSS.n409 DVSS.n408 0.00430282
R33445 DVSS.n10965 DVSS.n10964 0.00427756
R33446 DVSS.n17098 DVSS.n17097 0.00427756
R33447 DVSS.n9987 DVSS.n9986 0.00427756
R33448 DVSS.n10640 DVSS.n10638 0.00426578
R33449 DVSS.n8036 DVSS.n8034 0.00426578
R33450 DVSS.n10350 DVSS.n10349 0.00423239
R33451 DVSS.n4943 DVSS.n4942 0.00422857
R33452 DVSS.n4899 DVSS.n4898 0.00422857
R33453 DVSS.n4839 DVSS.n4838 0.00422857
R33454 DVSS.n6216 DVSS.n6215 0.00422857
R33455 DVSS.n6158 DVSS.n6157 0.00422857
R33456 DVSS.n5590 DVSS.n5589 0.00422047
R33457 DVSS.n5728 DVSS.n5727 0.00422047
R33458 DVSS.n10274 DVSS.n10273 0.00422047
R33459 DVSS.n12713 DVSS.n12712 0.00422047
R33460 DVSS.n12712 DVSS.n12711 0.00422047
R33461 DVSS.n12214 DVSS.n12213 0.00422047
R33462 DVSS.n12187 DVSS.n12186 0.00422047
R33463 DVSS.n21281 DVSS.n21280 0.00422047
R33464 DVSS.n17013 DVSS.n17012 0.00422047
R33465 DVSS.n10634 DVSS.n10633 0.00422047
R33466 DVSS.n10762 DVSS.n10761 0.00422047
R33467 DVSS.n11432 DVSS.n11431 0.00422047
R33468 DVSS.n5229 DVSS.n5228 0.00422047
R33469 DVSS.n3336 DVSS.n3335 0.00422047
R33470 DVSS.n3335 DVSS.n3334 0.00422047
R33471 DVSS.n2844 DVSS.n2843 0.00422047
R33472 DVSS.n2816 DVSS.n2815 0.00422047
R33473 DVSS.n658 DVSS.n657 0.00422047
R33474 DVSS.n9917 DVSS.n9916 0.00422047
R33475 DVSS.n17308 DVSS.n17307 0.00422047
R33476 DVSS.n16349 DVSS.n16348 0.00422047
R33477 DVSS.n5393 DVSS.n5392 0.00422047
R33478 DVSS.n5488 DVSS.n5487 0.00422047
R33479 DVSS.n6467 DVSS.n6466 0.00422047
R33480 DVSS.n9438 DVSS.n9437 0.00422
R33481 DVSS.n18487 DVSS.n18486 0.00416802
R33482 DVSS.n7728 DVSS.n7727 0.00416802
R33483 DVSS.n18228 DVSS.n18227 0.00416734
R33484 DVSS.n15512 DVSS.n15511 0.00416734
R33485 DVSS.n6805 DVSS.n6803 0.00416429
R33486 DVSS.n3927 DVSS.n3925 0.00416429
R33487 DVSS.n3897 DVSS.n3895 0.00416429
R33488 DVSS.n3851 DVSS.n3849 0.00416429
R33489 DVSS.n3624 DVSS.n3619 0.00416429
R33490 DVSS.n2755 DVSS.n2721 0.00416429
R33491 DVSS.n5975 DVSS.n5973 0.00416429
R33492 DVSS.n5929 DVSS.n5927 0.00416429
R33493 DVSS.n12547 DVSS.n12546 0.00415385
R33494 DVSS.n12671 DVSS.n12670 0.00415385
R33495 DVSS.n12579 DVSS.n12578 0.00415385
R33496 DVSS.n12383 DVSS.n12382 0.00415385
R33497 DVSS.n12291 DVSS.n12290 0.00415385
R33498 DVSS.n12250 DVSS.n12245 0.00415385
R33499 DVSS.n3171 DVSS.n3170 0.00415385
R33500 DVSS.n3295 DVSS.n3294 0.00415385
R33501 DVSS.n3203 DVSS.n3202 0.00415385
R33502 DVSS.n3010 DVSS.n3009 0.00415385
R33503 DVSS.n2918 DVSS.n2917 0.00415385
R33504 DVSS.n2877 DVSS.n2872 0.00415385
R33505 DVSS.n1367 DVSS.n1366 0.00414027
R33506 DVSS.n1368 DVSS.n1367 0.00414027
R33507 DVSS.n7719 DVSS.n7718 0.0041
R33508 DVSS.n15066 DVSS.n15065 0.0041
R33509 DVSS.n16050 DVSS.n16049 0.0041
R33510 DVSS.n17529 DVSS.n17528 0.0041
R33511 DVSS.n15263 DVSS.n15262 0.0041
R33512 DVSS.n18356 DVSS.n18355 0.0041
R33513 DVSS.n18077 DVSS.n18076 0.0041
R33514 DVSS.n17936 DVSS.n17935 0.0041
R33515 DVSS.n8081 DVSS.n8080 0.0041
R33516 DVSS.n2700 DVSS.n2699 0.0041
R33517 DVSS.n2646 DVSS.n2645 0.0041
R33518 DVSS.n11335 DVSS 0.0041
R33519 DVSS.n8373 DVSS.n8372 0.0041
R33520 DVSS.n13973 DVSS.n13972 0.0041
R33521 DVSS.n5347 DVSS.n5346 0.00409785
R33522 DVSS.n1365 DVSS.n1364 0.00409785
R33523 DVSS.n16573 DVSS.n16572 0.00409155
R33524 DVSS.n16676 DVSS.n16675 0.00409155
R33525 DVSS.n16076 DVSS.n16075 0.00409155
R33526 DVSS.n18272 DVSS.n18271 0.00409155
R33527 DVSS.n18246 DVSS.n18245 0.00409155
R33528 DVSS.n18237 DVSS.n18236 0.00409155
R33529 DVSS.n18185 DVSS.n18184 0.00409155
R33530 DVSS.n18449 DVSS.n18448 0.00409155
R33531 DVSS.n19647 DVSS.n19646 0.00409155
R33532 DVSS.n19711 DVSS.n19710 0.00409155
R33533 DVSS.n19790 DVSS.n19789 0.00409155
R33534 DVSS.n142 DVSS.n141 0.00409155
R33535 DVSS.n231 DVSS.n230 0.00409155
R33536 DVSS.n190 DVSS.n189 0.00409155
R33537 DVSS.n16760 DVSS.n16759 0.00409155
R33538 DVSS.n17147 DVSS.n17146 0.00409155
R33539 DVSS.n15968 DVSS.n15967 0.00409155
R33540 DVSS.n15468 DVSS.n15467 0.00409155
R33541 DVSS.n15494 DVSS.n15493 0.00409155
R33542 DVSS.n15503 DVSS.n15502 0.00409155
R33543 DVSS.n15555 DVSS.n15554 0.00409155
R33544 DVSS.n15168 DVSS.n15167 0.00409155
R33545 DVSS.n19856 DVSS.n19855 0.00409155
R33546 DVSS.n19930 DVSS.n19929 0.00409155
R33547 DVSS.n20015 DVSS.n20014 0.00409155
R33548 DVSS.n302 DVSS.n301 0.00409155
R33549 DVSS.n439 DVSS.n438 0.00409155
R33550 DVSS.n398 DVSS.n397 0.00409155
R33551 DVSS.n5751 DVSS.n5750 0.00406877
R33552 DVSS.n5742 DVSS.n5741 0.00406877
R33553 DVSS.n5720 DVSS.n5719 0.00406877
R33554 DVSS.n6504 DVSS.n6503 0.00406877
R33555 DVSS.n11254 DVSS.n11253 0.00406877
R33556 DVSS.n11215 DVSS.n8926 0.00406877
R33557 DVSS.n11245 DVSS.n11244 0.00406877
R33558 DVSS.n11223 DVSS.n11222 0.00406877
R33559 DVSS.n17646 DVSS.n17645 0.00406877
R33560 DVSS.n17653 DVSS.n15871 0.00406877
R33561 DVSS.n11164 DVSS.n9839 0.00406877
R33562 DVSS.n9832 DVSS.n9814 0.00406877
R33563 DVSS.n16341 DVSS.n16331 0.00406877
R33564 DVSS.n16323 DVSS.n16304 0.00406877
R33565 DVSS.n18494 DVSS.n18493 0.00406336
R33566 DVSS.n14479 DVSS.n14478 0.00406336
R33567 DVSS.n7735 DVSS.n7734 0.00406336
R33568 DVSS.n14637 DVSS.n14636 0.00406336
R33569 DVSS.n18234 DVSS.n18233 0.00406318
R33570 DVSS.n15506 DVSS.n15505 0.00406318
R33571 DVSS.n5795 DVSS.n5794 0.00404331
R33572 DVSS.n5757 DVSS.n5756 0.00404331
R33573 DVSS.n4068 DVSS.n4067 0.00404331
R33574 DVSS.n6984 DVSS.n6983 0.00404331
R33575 DVSS.n9843 DVSS.n9842 0.00404331
R33576 DVSS.n11260 DVSS.n11259 0.00404331
R33577 DVSS.n8987 DVSS.n8986 0.00404331
R33578 DVSS.n12964 DVSS.n12963 0.00404331
R33579 DVSS.n12821 DVSS.n12820 0.00404331
R33580 DVSS.n12758 DVSS.n12757 0.00404331
R33581 DVSS.n21298 DVSS.n21297 0.00404331
R33582 DVSS.n17563 DVSS.n17562 0.00404331
R33583 DVSS.n17605 DVSS.n17604 0.00404331
R33584 DVSS.n15008 DVSS.n15007 0.00404331
R33585 DVSS.n13654 DVSS.n13653 0.00404331
R33586 DVSS.n11402 DVSS.n11401 0.00404331
R33587 DVSS.n11705 DVSS.n11704 0.00404331
R33588 DVSS.n13028 DVSS.n13027 0.00404331
R33589 DVSS.n3805 DVSS.n3804 0.00404331
R33590 DVSS.n3767 DVSS.n3766 0.00404331
R33591 DVSS.n3433 DVSS.n3432 0.00404331
R33592 DVSS.n3371 DVSS.n3370 0.00404331
R33593 DVSS.n708 DVSS.n707 0.00404331
R33594 DVSS.n11086 DVSS.n11085 0.00404331
R33595 DVSS.n11128 DVSS.n11127 0.00404331
R33596 DVSS.n9077 DVSS.n9076 0.00404331
R33597 DVSS.n13221 DVSS.n13220 0.00404331
R33598 DVSS.n16416 DVSS.n16415 0.00404331
R33599 DVSS.n16378 DVSS.n16377 0.00404331
R33600 DVSS.n7533 DVSS.n7532 0.00404331
R33601 DVSS.n18751 DVSS.n18750 0.00404331
R33602 DVSS.n5449 DVSS.n5448 0.00404331
R33603 DVSS.n6085 DVSS.n6084 0.00404331
R33604 DVSS.n6786 DVSS.n6785 0.00404331
R33605 DVSS.n3594 DVSS.n3593 0.00404331
R33606 DVSS.n4791 DVSS.n4790 0.00403571
R33607 DVSS.n11846 DVSS.n11845 0.00403571
R33608 DVSS.n11905 DVSS.n11904 0.00403571
R33609 DVSS.n8621 DVSS.n8620 0.00403571
R33610 DVSS.n14474 DVSS.n14473 0.0040341
R33611 DVSS.n14652 DVSS.n14651 0.0040341
R33612 DVSS.n5383 DVSS.n5382 0.00401955
R33613 DVSS.n5366 DVSS.n5365 0.00401955
R33614 DVSS.n5608 DVSS.n5607 0.00401955
R33615 DVSS.n5576 DVSS.n5572 0.00401955
R33616 DVSS.n17327 DVSS.n17325 0.00401955
R33617 DVSS.n17303 DVSS.n17277 0.00401955
R33618 DVSS.n16998 DVSS.n16997 0.00401955
R33619 DVSS.n17008 DVSS.n17005 0.00401955
R33620 DVSS.n10218 DVSS.n10217 0.00401955
R33621 DVSS.n10242 DVSS.n10240 0.00401955
R33622 DVSS.n10250 DVSS.n10249 0.00401955
R33623 DVSS.n10269 DVSS.n10257 0.00401955
R33624 DVSS.n5685 DVSS.n5684 0.00397904
R33625 DVSS.n4664 DVSS.n4663 0.00397904
R33626 DVSS.n17404 DVSS.n17403 0.00397904
R33627 DVSS.n4575 DVSS.n4574 0.00397222
R33628 DVSS.n5505 DVSS.n4624 0.00397222
R33629 DVSS.n6274 DVSS.n6273 0.00397143
R33630 DVSS.n19691 DVSS.n19690 0.0039558
R33631 DVSS.n19769 DVSS.n19768 0.0039558
R33632 DVSS.n210 DVSS.n209 0.0039558
R33633 DVSS.n19910 DVSS.n19909 0.0039558
R33634 DVSS.n19994 DVSS.n19993 0.0039558
R33635 DVSS.n418 DVSS.n417 0.0039558
R33636 DVSS.n19690 DVSS.n19689 0.0039558
R33637 DVSS.n19909 DVSS.n19908 0.0039558
R33638 DVSS.n19770 DVSS.n19769 0.0039558
R33639 DVSS.n19995 DVSS.n19994 0.0039558
R33640 DVSS.n211 DVSS.n210 0.0039558
R33641 DVSS.n419 DVSS.n418 0.0039558
R33642 DVSS.n5811 DVSS.n5803 0.00395082
R33643 DVSS.n7086 DVSS.n7085 0.00395082
R33644 DVSS.n6532 DVSS.n6531 0.00395082
R33645 DVSS.n4381 DVSS.n4380 0.00395082
R33646 DVSS.n4091 DVSS.n4090 0.00395082
R33647 DVSS.n11047 DVSS.n9851 0.00395082
R33648 DVSS.n11234 DVSS.n11233 0.00395082
R33649 DVSS.n17554 DVSS.n17553 0.00395082
R33650 DVSS.n13819 DVSS.n13797 0.00395082
R33651 DVSS.n13781 DVSS.n13760 0.00395082
R33652 DVSS.n13744 DVSS.n13712 0.00395082
R33653 DVSS.n17631 DVSS.n17630 0.00395082
R33654 DVSS.n13640 DVSS.n13596 0.00395082
R33655 DVSS.n11077 DVSS.n11076 0.00395082
R33656 DVSS.n11154 DVSS.n11153 0.00395082
R33657 DVSS.n16352 DVSS.n16351 0.00395082
R33658 DVSS.n18623 DVSS.n18622 0.00395082
R33659 DVSS.n18650 DVSS.n18649 0.00395082
R33660 DVSS.n18682 DVSS.n18681 0.00395082
R33661 DVSS.n17448 DVSS.n16424 0.00395082
R33662 DVSS.n18816 DVSS.n18815 0.00395082
R33663 DVSS.n5264 DVSS.n5262 0.0039507
R33664 DVSS.n9766 DVSS.n9765 0.00392323
R33665 DVSS.n15869 DVSS.n15868 0.00392323
R33666 DVSS.n9812 DVSS.n9811 0.00392323
R33667 DVSS.n2362 DVSS.n2361 0.0039231
R33668 DVSS.n2404 DVSS.n2403 0.0039231
R33669 DVSS DVSS.n9476 0.00392
R33670 DVSS.n9475 DVSS 0.00392
R33671 DVSS.n12111 DVSS 0.00392
R33672 DVSS DVSS.n12014 0.00392
R33673 DVSS.n10889 DVSS 0.00391158
R33674 DVSS.n4965 DVSS.n4964 0.00390714
R33675 DVSS.n4921 DVSS.n4920 0.00390714
R33676 DVSS.n4861 DVSS.n4860 0.00390714
R33677 DVSS.n4766 DVSS.n4765 0.00390714
R33678 DVSS.n8102 DVSS.n8101 0.00390714
R33679 DVSS.n8394 DVSS.n8393 0.00390714
R33680 DVSS.n6237 DVSS.n6236 0.00390714
R33681 DVSS.n6179 DVSS.n6178 0.00390714
R33682 DVSS.n8644 DVSS.n8643 0.00390714
R33683 DVSS.n12439 DVSS.n12438 0.00389055
R33684 DVSS.n16668 DVSS.n16667 0.00388028
R33685 DVSS.n17477 DVSS.n17476 0.00388028
R33686 DVSS.n16068 DVSS.n16067 0.00388028
R33687 DVSS.n17775 DVSS.n17774 0.00388028
R33688 DVSS.n17884 DVSS.n17883 0.00388028
R33689 DVSS.n18025 DVSS.n18024 0.00388028
R33690 DVSS.n18264 DVSS.n18263 0.00388028
R33691 DVSS.n18180 DVSS.n18179 0.00388028
R33692 DVSS.n7576 DVSS.n7575 0.00388028
R33693 DVSS.n18472 DVSS.n18471 0.00388028
R33694 DVSS.n18512 DVSS.n18511 0.00388028
R33695 DVSS.n18557 DVSS.n18556 0.00388028
R33696 DVSS.n19757 DVSS.n19756 0.00388028
R33697 DVSS.n161 DVSS.n160 0.00388028
R33698 DVSS.n17155 DVSS.n17154 0.00388028
R33699 DVSS.n16818 DVSS.n16817 0.00388028
R33700 DVSS.n15960 DVSS.n15959 0.00388028
R33701 DVSS.n15888 DVSS.n15887 0.00388028
R33702 DVSS.n15815 DVSS.n15814 0.00388028
R33703 DVSS.n15747 DVSS.n15746 0.00388028
R33704 DVSS.n15476 DVSS.n15475 0.00388028
R33705 DVSS.n15560 DVSS.n15559 0.00388028
R33706 DVSS.n15233 DVSS.n15232 0.00388028
R33707 DVSS.n15130 DVSS.n15129 0.00388028
R33708 DVSS.n7753 DVSS.n7752 0.00388028
R33709 DVSS.n13919 DVSS.n13851 0.00388028
R33710 DVSS.n19982 DVSS.n19981 0.00388028
R33711 DVSS.n321 DVSS.n320 0.00388028
R33712 DVSS.n16590 DVSS.n16589 0.003875
R33713 DVSS.n15211 DVSS.n15210 0.003875
R33714 DVSS.n16494 DVSS.n16493 0.003875
R33715 DVSS.n15361 DVSS.n15360 0.003875
R33716 DVSS.n18091 DVSS.n18090 0.003875
R33717 DVSS.n15429 DVSS.n15428 0.003875
R33718 DVSS.n18283 DVSS.n18282 0.003875
R33719 DVSS.n18332 DVSS.n18331 0.003875
R33720 DVSS.n18343 DVSS.n18342 0.003875
R33721 DVSS.n17950 DVSS.n17949 0.003875
R33722 DVSS.n17809 DVSS.n17808 0.003875
R33723 DVSS.n13859 DVSS.n13858 0.003875
R33724 DVSS.n5697 DVSS.n5696 0.00386614
R33725 DVSS.n4454 DVSS.n4453 0.00386614
R33726 DVSS.n7212 DVSS.n7211 0.00386614
R33727 DVSS.n19298 DVSS.n19297 0.00386614
R33728 DVSS.n1053 DVSS.n1052 0.00386614
R33729 DVSS.n9505 DVSS.n9504 0.00386614
R33730 DVSS.n12904 DVSS.n12903 0.00386614
R33731 DVSS.n12831 DVSS.n12830 0.00386614
R33732 DVSS.n12405 DVSS.n12404 0.00386614
R33733 DVSS.n12212 DVSS.n12211 0.00386614
R33734 DVSS.n21311 DVSS.n21310 0.00386614
R33735 DVSS.n21302 DVSS.n21301 0.00386614
R33736 DVSS.n15692 DVSS.n15691 0.00386614
R33737 DVSS.n13515 DVSS.n13514 0.00386614
R33738 DVSS.n20314 DVSS.n20313 0.00386614
R33739 DVSS.n20820 DVSS.n20819 0.00386614
R33740 DVSS.n10812 DVSS.n10811 0.00386614
R33741 DVSS.n10792 DVSS.n10791 0.00386614
R33742 DVSS.n10739 DVSS.n10738 0.00386614
R33743 DVSS.n11543 DVSS.n11542 0.00386614
R33744 DVSS.n12089 DVSS.n12088 0.00386614
R33745 DVSS.n21553 DVSS.n21552 0.00386614
R33746 DVSS.n21465 DVSS.n21464 0.00386614
R33747 DVSS.n4652 DVSS.n4651 0.00386614
R33748 DVSS.n4276 DVSS.n4275 0.00386614
R33749 DVSS.n3511 DVSS.n3510 0.00386614
R33750 DVSS.n3443 DVSS.n3442 0.00386614
R33751 DVSS.n3031 DVSS.n3030 0.00386614
R33752 DVSS.n2842 DVSS.n2841 0.00386614
R33753 DVSS.n781 DVSS.n780 0.00386614
R33754 DVSS.n665 DVSS.n664 0.00386614
R33755 DVSS.n9689 DVSS.n9688 0.00386614
R33756 DVSS.n13417 DVSS.n13416 0.00386614
R33757 DVSS.n20588 DVSS.n20587 0.00386614
R33758 DVSS.n21046 DVSS.n21045 0.00386614
R33759 DVSS.n17416 DVSS.n17415 0.00386614
R33760 DVSS.n16204 DVSS.n16203 0.00386614
R33761 DVSS.n18872 DVSS.n18871 0.00386614
R33762 DVSS.n19569 DVSS.n19568 0.00386614
R33763 DVSS.n1268 DVSS.n1267 0.00386614
R33764 DVSS.n5451 DVSS.n5450 0.00386614
R33765 DVSS.n5472 DVSS.n5471 0.00386614
R33766 DVSS.n5854 DVSS.n5853 0.00386614
R33767 DVSS.n6590 DVSS.n6589 0.00386614
R33768 DVSS.n3573 DVSS.n3572 0.00386614
R33769 DVSS.n19017 DVSS.n19016 0.00386614
R33770 DVSS.n619 DVSS.n618 0.00386614
R33771 DVSS.n7164 DVSS.n7163 0.00385106
R33772 DVSS.n1314 DVSS.n1311 0.00385106
R33773 DVSS.n7299 DVSS.n7298 0.00385106
R33774 DVSS.n7313 DVSS.n7310 0.00385106
R33775 DVSS.n7868 DVSS.n7867 0.00385106
R33776 DVSS.n7878 DVSS.n7877 0.00385106
R33777 DVSS.n7956 DVSS.n7955 0.00385106
R33778 DVSS.n7973 DVSS.n7965 0.00385106
R33779 DVSS.n7033 DVSS.n7032 0.00385106
R33780 DVSS.n7074 DVSS.n7073 0.00385106
R33781 DVSS.n7065 DVSS.n7064 0.00385106
R33782 DVSS.n14154 DVSS.n14152 0.00385106
R33783 DVSS.n13604 DVSS.n13603 0.00385106
R33784 DVSS.n13624 DVSS.n13623 0.00385106
R33785 DVSS.n13319 DVSS.n13317 0.00385106
R33786 DVSS.n16686 DVSS.n16685 0.00385031
R33787 DVSS.n18173 DVSS.n18172 0.00385031
R33788 DVSS.n14509 DVSS.n14508 0.00385031
R33789 DVSS.n19799 DVSS.n19798 0.00385031
R33790 DVSS.n152 DVSS.n151 0.00385031
R33791 DVSS.n240 DVSS.n239 0.00385031
R33792 DVSS.n18461 DVSS.n18460 0.00385031
R33793 DVSS.n18172 DVSS.n18171 0.00385031
R33794 DVSS.n17136 DVSS.n17135 0.00385031
R33795 DVSS.n15567 DVSS.n15566 0.00385031
R33796 DVSS.n14606 DVSS.n14605 0.00385031
R33797 DVSS.n20024 DVSS.n20023 0.00385031
R33798 DVSS.n312 DVSS.n311 0.00385031
R33799 DVSS.n448 DVSS.n447 0.00385031
R33800 DVSS.n15141 DVSS.n15140 0.00385031
R33801 DVSS.n15568 DVSS.n15567 0.00385031
R33802 DVSS.n17137 DVSS.n17136 0.00385031
R33803 DVSS.n16687 DVSS.n16686 0.00385031
R33804 DVSS.n14510 DVSS.n14509 0.00385031
R33805 DVSS.n14607 DVSS.n14606 0.00385031
R33806 DVSS.n19800 DVSS.n19799 0.00385031
R33807 DVSS.n20025 DVSS.n20024 0.00385031
R33808 DVSS.n311 DVSS.n310 0.00385031
R33809 DVSS.n151 DVSS.n150 0.00385031
R33810 DVSS.n241 DVSS.n240 0.00385031
R33811 DVSS.n449 DVSS.n448 0.00385031
R33812 DVSS.n10082 DVSS.n10081 0.00384286
R33813 DVSS.n10143 DVSS.n10142 0.00384286
R33814 DVSS.n10697 DVSS.n10696 0.00384286
R33815 DVSS.n6262 DVSS.n6261 0.00384286
R33816 DVSS.n8715 DVSS.n8714 0.00384286
R33817 DVSS.n8776 DVSS.n8775 0.00384286
R33818 DVSS.n8871 DVSS.n8870 0.00384286
R33819 DVSS.n5734 DVSS.n5733 0.00383286
R33820 DVSS.n13822 DVSS.n13821 0.00383286
R33821 DVSS.n13784 DVSS.n13783 0.00383286
R33822 DVSS.n13747 DVSS.n13746 0.00383286
R33823 DVSS.n4671 DVSS.n4670 0.00383286
R33824 DVSS.n18813 DVSS.n18797 0.00383286
R33825 DVSS.n12408 DVSS.n12407 0.00380239
R33826 DVSS.n3016 DVSS.n3015 0.00380234
R33827 DVSS.n9168 DVSS.n9167 0.00377
R33828 DVSS.n12144 DVSS.n12143 0.00376923
R33829 DVSS.n12151 DVSS.n12146 0.00376923
R33830 DVSS.n12609 DVSS.n12608 0.00376923
R33831 DVSS.n12600 DVSS.n12595 0.00376923
R33832 DVSS.n12321 DVSS.n12320 0.00376923
R33833 DVSS.n12312 DVSS.n12307 0.00376923
R33834 DVSS.n12229 DVSS.n12228 0.00376923
R33835 DVSS.n21205 DVSS.n21202 0.00376923
R33836 DVSS.n2764 DVSS.n2763 0.00376923
R33837 DVSS.n2771 DVSS.n2766 0.00376923
R33838 DVSS.n3233 DVSS.n3232 0.00376923
R33839 DVSS.n3224 DVSS.n3219 0.00376923
R33840 DVSS.n2948 DVSS.n2947 0.00376923
R33841 DVSS.n2939 DVSS.n2934 0.00376923
R33842 DVSS.n2856 DVSS.n2855 0.00376923
R33843 DVSS.n883 DVSS.n882 0.00376923
R33844 DVSS.n11242 DVSS.n11241 0.00374606
R33845 DVSS.n17623 DVSS.n17622 0.00374606
R33846 DVSS.n11146 DVSS.n11145 0.00374606
R33847 DVSS.n19142 DVSS.n19136 0.00374577
R33848 DVSS.n20153 DVSS.n20135 0.00374577
R33849 DVSS.n20424 DVSS.n20418 0.00374577
R33850 DVSS.n19416 DVSS.n19410 0.00374577
R33851 DVSS.n17468 DVSS.n17467 0.0037448
R33852 DVSS.n17794 DVSS.n17793 0.0037448
R33853 DVSS.n14374 DVSS.n14373 0.0037448
R33854 DVSS.n180 DVSS.n179 0.0037448
R33855 DVSS.n17469 DVSS.n17468 0.0037448
R33856 DVSS.n18227 DVSS.n18226 0.0037448
R33857 DVSS.n17795 DVSS.n17794 0.0037448
R33858 DVSS.n14373 DVSS.n14372 0.0037448
R33859 DVSS.n16809 DVSS.n16808 0.0037448
R33860 DVSS.n17668 DVSS.n17667 0.0037448
R33861 DVSS.n15513 DVSS.n15512 0.0037448
R33862 DVSS.n14777 DVSS.n14776 0.0037448
R33863 DVSS.n388 DVSS.n387 0.0037448
R33864 DVSS.n16810 DVSS.n16809 0.0037448
R33865 DVSS.n17669 DVSS.n17668 0.0037448
R33866 DVSS.n14776 DVSS.n14775 0.0037448
R33867 DVSS.n389 DVSS.n388 0.0037448
R33868 DVSS.n181 DVSS.n180 0.0037448
R33869 DVSS.n19643 DVSS.n19636 0.00374324
R33870 DVSS.n19681 DVSS.n19679 0.00374324
R33871 DVSS.n19900 DVSS.n19893 0.00374324
R33872 DVSS.n19874 DVSS.n19872 0.00374324
R33873 DVSS.n9227 DVSS.n9225 0.00371
R33874 DVSS.n2373 DVSS.n2372 0.00369838
R33875 DVSS.n2392 DVSS.n2391 0.00369838
R33876 DVSS.n5660 DVSS.n5659 0.00368898
R33877 DVSS.n5674 DVSS.n5673 0.00368898
R33878 DVSS.n4426 DVSS.n4425 0.00368898
R33879 DVSS.n4410 DVSS.n4409 0.00368898
R33880 DVSS.n19183 DVSS.n19182 0.00368898
R33881 DVSS.n19270 DVSS.n19269 0.00368898
R33882 DVSS.n842 DVSS.n841 0.00368898
R33883 DVSS.n1025 DVSS.n1024 0.00368898
R33884 DVSS.n1009 DVSS.n1008 0.00368898
R33885 DVSS.n10953 DVSS.n10952 0.00368898
R33886 DVSS.n9535 DVSS.n9534 0.00368898
R33887 DVSS.n9554 DVSS.n9553 0.00368898
R33888 DVSS.n12874 DVSS.n12873 0.00368898
R33889 DVSS.n12855 DVSS.n12854 0.00368898
R33890 DVSS.n12823 DVSS.n12822 0.00368898
R33891 DVSS.n12699 DVSS.n12698 0.00368898
R33892 DVSS.n12426 DVSS.n12425 0.00368898
R33893 DVSS.n21287 DVSS.n21286 0.00368898
R33894 DVSS.n21197 DVSS.n21196 0.00368898
R33895 DVSS.n17086 DVSS.n17085 0.00368898
R33896 DVSS.n15662 DVSS.n15661 0.00368898
R33897 DVSS.n15643 DVSS.n15642 0.00368898
R33898 DVSS.n20194 DVSS.n20193 0.00368898
R33899 DVSS.n20284 DVSS.n20283 0.00368898
R33900 DVSS.n20825 DVSS.n20824 0.00368898
R33901 DVSS.n20790 DVSS.n20789 0.00368898
R33902 DVSS.n20771 DVSS.n20770 0.00368898
R33903 DVSS.n11419 DVSS.n11418 0.00368898
R33904 DVSS.n11445 DVSS.n11444 0.00368898
R33905 DVSS.n11446 DVSS.n11445 0.00368898
R33906 DVSS.n11573 DVSS.n11572 0.00368898
R33907 DVSS.n11592 DVSS.n11591 0.00368898
R33908 DVSS.n22 DVSS.n21 0.00368898
R33909 DVSS.n41 DVSS.n40 0.00368898
R33910 DVSS.n21523 DVSS.n21522 0.00368898
R33911 DVSS.n21504 DVSS.n21503 0.00368898
R33912 DVSS.n21435 DVSS.n21434 0.00368898
R33913 DVSS.n21416 DVSS.n21415 0.00368898
R33914 DVSS.n4689 DVSS.n4688 0.00368898
R33915 DVSS.n4675 DVSS.n4674 0.00368898
R33916 DVSS.n4304 DVSS.n4303 0.00368898
R33917 DVSS.n4320 DVSS.n4319 0.00368898
R33918 DVSS.n3483 DVSS.n3482 0.00368898
R33919 DVSS.n3467 DVSS.n3466 0.00368898
R33920 DVSS.n3435 DVSS.n3434 0.00368898
R33921 DVSS.n3322 DVSS.n3321 0.00368898
R33922 DVSS.n3052 DVSS.n3051 0.00368898
R33923 DVSS.n737 DVSS.n736 0.00368898
R33924 DVSS.n804 DVSS.n803 0.00368898
R33925 DVSS.n9975 DVSS.n9974 0.00368898
R33926 DVSS.n9659 DVSS.n9658 0.00368898
R33927 DVSS.n9640 DVSS.n9639 0.00368898
R33928 DVSS.n20465 DVSS.n20464 0.00368898
R33929 DVSS.n20558 DVSS.n20557 0.00368898
R33930 DVSS.n21051 DVSS.n21050 0.00368898
R33931 DVSS.n21016 DVSS.n21015 0.00368898
R33932 DVSS.n20997 DVSS.n20996 0.00368898
R33933 DVSS.n17379 DVSS.n17378 0.00368898
R33934 DVSS.n17393 DVSS.n17392 0.00368898
R33935 DVSS.n16176 DVSS.n16175 0.00368898
R33936 DVSS.n16159 DVSS.n16158 0.00368898
R33937 DVSS.n19454 DVSS.n19453 0.00368898
R33938 DVSS.n19541 DVSS.n19540 0.00368898
R33939 DVSS.n1129 DVSS.n1128 0.00368898
R33940 DVSS.n1240 DVSS.n1239 0.00368898
R33941 DVSS.n1224 DVSS.n1223 0.00368898
R33942 DVSS.n6341 DVSS.n6340 0.00368898
R33943 DVSS.n6454 DVSS.n6453 0.00368898
R33944 DVSS.n6453 DVSS.n6452 0.00368898
R33945 DVSS.n6618 DVSS.n6617 0.00368898
R33946 DVSS.n6635 DVSS.n6634 0.00368898
R33947 DVSS.n3545 DVSS.n3544 0.00368898
R33948 DVSS.n18942 DVSS.n18941 0.00368898
R33949 DVSS.n18989 DVSS.n18988 0.00368898
R33950 DVSS.n520 DVSS.n519 0.00368898
R33951 DVSS.n591 DVSS.n590 0.00368898
R33952 DVSS.n575 DVSS.n574 0.00368898
R33953 DVSS.n5348 DVSS.n5347 0.00368083
R33954 DVSS.n1366 DVSS.n1365 0.00368083
R33955 DVSS.n5268 DVSS.n5267 0.00366901
R33956 DVSS.n5181 DVSS.n5179 0.00366901
R33957 DVSS.n5143 DVSS.n5141 0.00366901
R33958 DVSS.n5089 DVSS.n5087 0.00366901
R33959 DVSS.n10405 DVSS.n10404 0.00366901
R33960 DVSS.n10464 DVSS.n10463 0.00366901
R33961 DVSS.n10562 DVSS.n10561 0.00366901
R33962 DVSS.n16557 DVSS.n16556 0.00366901
R33963 DVSS.n16502 DVSS.n16501 0.00366901
R33964 DVSS.n16121 DVSS.n16120 0.00366901
R33965 DVSS.n16089 DVSS.n16088 0.00366901
R33966 DVSS.n17806 DVSS.n17805 0.00366901
R33967 DVSS.n17947 DVSS.n17946 0.00366901
R33968 DVSS.n18088 DVSS.n18087 0.00366901
R33969 DVSS.n18123 DVSS.n18122 0.00366901
R33970 DVSS.n18146 DVSS.n18145 0.00366901
R33971 DVSS.n18147 DVSS.n18146 0.00366901
R33972 DVSS.n18211 DVSS.n18210 0.00366901
R33973 DVSS.n7606 DVSS.n7605 0.00366901
R33974 DVSS.n18419 DVSS.n18418 0.00366901
R33975 DVSS.n18474 DVSS.n18473 0.00366901
R33976 DVSS.n18527 DVSS.n18526 0.00366901
R33977 DVSS.n14411 DVSS.n14410 0.00366901
R33978 DVSS.n16744 DVSS.n16743 0.00366901
R33979 DVSS.n16848 DVSS.n16847 0.00366901
R33980 DVSS.n16002 DVSS.n16001 0.00366901
R33981 DVSS.n15977 DVSS.n15976 0.00366901
R33982 DVSS.n15785 DVSS.n15784 0.00366901
R33983 DVSS.n15777 DVSS.n15776 0.00366901
R33984 DVSS.n15372 DVSS.n15371 0.00366901
R33985 DVSS.n15413 DVSS.n15412 0.00366901
R33986 DVSS.n15451 DVSS.n15450 0.00366901
R33987 DVSS.n15452 DVSS.n15451 0.00366901
R33988 DVSS.n15529 DVSS.n15528 0.00366901
R33989 DVSS.n15369 DVSS.n15368 0.00366901
R33990 DVSS.n15219 DVSS.n15218 0.00366901
R33991 DVSS.n15128 DVSS.n15127 0.00366901
R33992 DVSS.n13856 DVSS.n13855 0.00366901
R33993 DVSS.n14717 DVSS.n14716 0.00366901
R33994 DVSS.n17215 DVSS.n17214 0.00365
R33995 DVSS.n15183 DVSS.n15182 0.00365
R33996 DVSS.n15148 DVSS.n15147 0.00365
R33997 DVSS.n2338 DVSS.n2337 0.00365
R33998 DVSS.n17693 DVSS.n17692 0.00365
R33999 DVSS.n17682 DVSS.n17681 0.00365
R34000 DVSS.n17680 DVSS.n17679 0.00365
R34001 DVSS.n5056 DVSS.n4989 0.00365
R34002 DVSS.n6041 DVSS.n6039 0.00365
R34003 DVSS.n6324 DVSS.n6287 0.00365
R34004 DVSS.n13000 DVSS 0.00364286
R34005 DVSS.n18223 DVSS.n18222 0.00364043
R34006 DVSS.n15517 DVSS.n15516 0.00364043
R34007 DVSS.n18482 DVSS.n18481 0.00363995
R34008 DVSS.n15120 DVSS.n15119 0.00363995
R34009 DVSS.n16530 DVSS.n16529 0.0036393
R34010 DVSS.n17782 DVSS.n17781 0.0036393
R34011 DVSS.n14264 DVSS.n14263 0.0036393
R34012 DVSS.n14289 DVSS.n14288 0.0036393
R34013 DVSS.n14318 DVSS.n14317 0.0036393
R34014 DVSS.n14421 DVSS.n14420 0.0036393
R34015 DVSS.n14452 DVSS.n14451 0.0036393
R34016 DVSS.n14420 DVSS.n14419 0.0036393
R34017 DVSS.n14317 DVSS.n14316 0.0036393
R34018 DVSS.n14288 DVSS.n14287 0.0036393
R34019 DVSS.n14263 DVSS.n14262 0.0036393
R34020 DVSS.n18248 DVSS.n18247 0.0036393
R34021 DVSS.n17781 DVSS.n17780 0.0036393
R34022 DVSS.n16531 DVSS.n16530 0.0036393
R34023 DVSS.n14451 DVSS.n14450 0.0036393
R34024 DVSS.n16718 DVSS.n16717 0.0036393
R34025 DVSS.n14851 DVSS.n14850 0.0036393
R34026 DVSS.n14834 DVSS.n14833 0.0036393
R34027 DVSS.n14817 DVSS.n14816 0.0036393
R34028 DVSS.n14707 DVSS.n14706 0.0036393
R34029 DVSS.n14670 DVSS.n14669 0.0036393
R34030 DVSS.n14708 DVSS.n14707 0.0036393
R34031 DVSS.n15492 DVSS.n15491 0.0036393
R34032 DVSS.n14852 DVSS.n14851 0.0036393
R34033 DVSS.n14835 DVSS.n14834 0.0036393
R34034 DVSS.n14818 DVSS.n14817 0.0036393
R34035 DVSS.n16717 DVSS.n16716 0.0036393
R34036 DVSS.n14671 DVSS.n14670 0.0036393
R34037 DVSS.n7060 DVSS.n7059 0.00363144
R34038 DVSS.n13313 DVSS.n13311 0.00363144
R34039 DVSS.n13311 DVSS.n13310 0.00363144
R34040 DVSS.n7059 DVSS.n7058 0.00363144
R34041 DVSS.n10616 DVSS.n10615 0.00362543
R34042 DVSS.n10882 DVSS.n10881 0.00359859
R34043 DVSS.n11019 DVSS.n11015 0.00355556
R34044 DVSS.n11679 DVSS.n11675 0.00355556
R34045 DVSS.n11642 DVSS.n11638 0.00355556
R34046 DVSS.n11517 DVSS.n11513 0.00355556
R34047 DVSS.n11189 DVSS.n11185 0.00355556
R34048 DVSS.n11480 DVSS.n11476 0.00355556
R34049 DVSS.n11728 DVSS.n11724 0.00355556
R34050 DVSS.n10029 DVSS.n10025 0.00355556
R34051 DVSS.n18475 DVSS.n18474 0.0035352
R34052 DVSS.n15127 DVSS.n15126 0.0035352
R34053 DVSS.n16585 DVSS.n16584 0.00353378
R34054 DVSS.n16689 DVSS.n16688 0.00353378
R34055 DVSS.n16699 DVSS.n16698 0.00353378
R34056 DVSS.n16515 DVSS.n16514 0.00353378
R34057 DVSS.n16506 DVSS.n16505 0.00353378
R34058 DVSS.n17780 DVSS.n17779 0.00353378
R34059 DVSS.n14242 DVSS.n14241 0.00353378
R34060 DVSS.n14267 DVSS.n14266 0.00353378
R34061 DVSS.n14292 DVSS.n14291 0.00353378
R34062 DVSS.n14429 DVSS.n14428 0.00353378
R34063 DVSS.n176 DVSS.n175 0.00353378
R34064 DVSS.n18198 DVSS.n18197 0.00353378
R34065 DVSS.n14241 DVSS.n14240 0.00353378
R34066 DVSS.n14266 DVSS.n14265 0.00353378
R34067 DVSS.n14291 DVSS.n14290 0.00353378
R34068 DVSS.n17779 DVSS.n17778 0.00353378
R34069 DVSS.n16584 DVSS.n16583 0.00353378
R34070 DVSS.n14428 DVSS.n14427 0.00353378
R34071 DVSS.n16772 DVSS.n16771 0.00353378
R34072 DVSS.n17134 DVSS.n17133 0.00353378
R34073 DVSS.n17124 DVSS.n17123 0.00353378
R34074 DVSS.n16861 DVSS.n16860 0.00353378
R34075 DVSS.n16852 DVSS.n16851 0.00353378
R34076 DVSS.n14865 DVSS.n14864 0.00353378
R34077 DVSS.n14848 DVSS.n14847 0.00353378
R34078 DVSS.n14831 DVSS.n14830 0.00353378
R34079 DVSS.n14699 DVSS.n14698 0.00353378
R34080 DVSS.n384 DVSS.n383 0.00353378
R34081 DVSS.n14700 DVSS.n14699 0.00353378
R34082 DVSS.n15542 DVSS.n15541 0.00353378
R34083 DVSS.n14866 DVSS.n14865 0.00353378
R34084 DVSS.n14849 DVSS.n14848 0.00353378
R34085 DVSS.n14832 DVSS.n14831 0.00353378
R34086 DVSS.n16771 DVSS.n16770 0.00353378
R34087 DVSS.n16862 DVSS.n16861 0.00353378
R34088 DVSS.n16516 DVSS.n16515 0.00353378
R34089 DVSS.n16698 DVSS.n16697 0.00353378
R34090 DVSS.n17135 DVSS.n17134 0.00353378
R34091 DVSS.n16688 DVSS.n16687 0.00353378
R34092 DVSS.n17125 DVSS.n17124 0.00353378
R34093 DVSS.n16853 DVSS.n16852 0.00353378
R34094 DVSS.n16507 DVSS.n16506 0.00353378
R34095 DVSS.n385 DVSS.n384 0.00353378
R34096 DVSS.n177 DVSS.n176 0.00353378
R34097 DVSS.n5182 DVSS.n5181 0.00352817
R34098 DVSS.n5144 DVSS.n5143 0.00352817
R34099 DVSS.n5090 DVSS.n5089 0.00352817
R34100 DVSS.n5384 DVSS.n5383 0.00351676
R34101 DVSS.n5365 DVSS.n5364 0.00351676
R34102 DVSS.n5608 DVSS.n5602 0.00351676
R34103 DVSS.n5576 DVSS.n5573 0.00351676
R34104 DVSS.n17327 DVSS.n17322 0.00351676
R34105 DVSS.n17303 DVSS.n17302 0.00351676
R34106 DVSS.n16998 DVSS.n16994 0.00351676
R34107 DVSS.n17008 DVSS.n17006 0.00351676
R34108 DVSS.n10217 DVSS.n10214 0.00351676
R34109 DVSS.n10243 DVSS.n10242 0.00351676
R34110 DVSS.n10250 DVSS.n10246 0.00351676
R34111 DVSS.n10269 DVSS.n10267 0.00351676
R34112 DVSS.n4437 DVSS.n4436 0.00351181
R34113 DVSS.n4399 DVSS.n4398 0.00351181
R34114 DVSS.n19124 DVSS.n19123 0.00351181
R34115 DVSS.n19194 DVSS.n19193 0.00351181
R34116 DVSS.n19281 DVSS.n19280 0.00351181
R34117 DVSS.n853 DVSS.n852 0.00351181
R34118 DVSS.n1036 DVSS.n1035 0.00351181
R34119 DVSS.n998 DVSS.n997 0.00351181
R34120 DVSS.n9524 DVSS.n9523 0.00351181
R34121 DVSS.n9565 DVSS.n9564 0.00351181
R34122 DVSS.n12885 DVSS.n12884 0.00351181
R34123 DVSS.n12844 DVSS.n12843 0.00351181
R34124 DVSS.n12749 DVSS.n12748 0.00351181
R34125 DVSS.n12691 DVSS.n12690 0.00351181
R34126 DVSS.n12464 DVSS.n12463 0.00351181
R34127 DVSS.n12435 DVSS.n12434 0.00351181
R34128 DVSS.n12417 DVSS.n12416 0.00351181
R34129 DVSS.n21306 DVSS.n21305 0.00351181
R34130 DVSS.n21201 DVSS.n21200 0.00351181
R34131 DVSS.n15673 DVSS.n15672 0.00351181
R34132 DVSS.n15632 DVSS.n15631 0.00351181
R34133 DVSS.n20124 DVSS.n20123 0.00351181
R34134 DVSS.n20205 DVSS.n20204 0.00351181
R34135 DVSS.n20295 DVSS.n20294 0.00351181
R34136 DVSS.n20836 DVSS.n20835 0.00351181
R34137 DVSS.n20801 DVSS.n20800 0.00351181
R34138 DVSS.n20760 DVSS.n20759 0.00351181
R34139 DVSS.n11562 DVSS.n11561 0.00351181
R34140 DVSS.n11603 DVSS.n11602 0.00351181
R34141 DVSS.n12070 DVSS.n12069 0.00351181
R34142 DVSS.n52 DVSS.n51 0.00351181
R34143 DVSS.n21534 DVSS.n21533 0.00351181
R34144 DVSS.n21493 DVSS.n21492 0.00351181
R34145 DVSS.n21446 DVSS.n21445 0.00351181
R34146 DVSS.n21405 DVSS.n21404 0.00351181
R34147 DVSS.n4293 DVSS.n4292 0.00351181
R34148 DVSS.n4331 DVSS.n4330 0.00351181
R34149 DVSS.n3494 DVSS.n3493 0.00351181
R34150 DVSS.n3456 DVSS.n3455 0.00351181
R34151 DVSS.n3362 DVSS.n3361 0.00351181
R34152 DVSS.n3314 DVSS.n3313 0.00351181
R34153 DVSS.n3090 DVSS.n3089 0.00351181
R34154 DVSS.n3061 DVSS.n3060 0.00351181
R34155 DVSS.n3044 DVSS.n3043 0.00351181
R34156 DVSS.n670 DVSS.n669 0.00351181
R34157 DVSS.n786 DVSS.n785 0.00351181
R34158 DVSS.n9670 DVSS.n9669 0.00351181
R34159 DVSS.n9629 DVSS.n9628 0.00351181
R34160 DVSS.n20407 DVSS.n20406 0.00351181
R34161 DVSS.n20476 DVSS.n20475 0.00351181
R34162 DVSS.n20569 DVSS.n20568 0.00351181
R34163 DVSS.n21062 DVSS.n21061 0.00351181
R34164 DVSS.n21027 DVSS.n21026 0.00351181
R34165 DVSS.n20986 DVSS.n20985 0.00351181
R34166 DVSS.n16187 DVSS.n16186 0.00351181
R34167 DVSS.n16148 DVSS.n16147 0.00351181
R34168 DVSS.n19398 DVSS.n19397 0.00351181
R34169 DVSS.n19465 DVSS.n19464 0.00351181
R34170 DVSS.n19552 DVSS.n19551 0.00351181
R34171 DVSS.n1140 DVSS.n1139 0.00351181
R34172 DVSS.n1251 DVSS.n1250 0.00351181
R34173 DVSS.n1213 DVSS.n1212 0.00351181
R34174 DVSS.n6607 DVSS.n6606 0.00351181
R34175 DVSS.n6646 DVSS.n6645 0.00351181
R34176 DVSS.n3556 DVSS.n3555 0.00351181
R34177 DVSS.n18953 DVSS.n18952 0.00351181
R34178 DVSS.n19000 DVSS.n18999 0.00351181
R34179 DVSS.n531 DVSS.n530 0.00351181
R34180 DVSS.n602 DVSS.n601 0.00351181
R34181 DVSS.n564 DVSS.n563 0.00351181
R34182 DVSS.n8033 DVSS.n8032 0.00350954
R34183 DVSS.n4418 DVSS.n4417 0.00347895
R34184 DVSS.n9545 DVSS.n9544 0.00347895
R34185 DVSS.n12864 DVSS.n12863 0.00347895
R34186 DVSS.n9544 DVSS.n9543 0.00347895
R34187 DVSS.n15652 DVSS.n15651 0.00347895
R34188 DVSS.n20185 DVSS.n20184 0.00347895
R34189 DVSS.n20274 DVSS.n20273 0.00347895
R34190 DVSS.n20780 DVSS.n20779 0.00347895
R34191 DVSS.n15653 DVSS.n15652 0.00347895
R34192 DVSS.n11583 DVSS.n11582 0.00347895
R34193 DVSS.n32 DVSS.n31 0.00347895
R34194 DVSS.n21513 DVSS.n21512 0.00347895
R34195 DVSS.n21425 DVSS.n21424 0.00347895
R34196 DVSS.n11582 DVSS.n11581 0.00347895
R34197 DVSS.n4312 DVSS.n4311 0.00347895
R34198 DVSS.n9649 DVSS.n9648 0.00347895
R34199 DVSS.n20456 DVSS.n20455 0.00347895
R34200 DVSS.n20548 DVSS.n20547 0.00347895
R34201 DVSS.n21006 DVSS.n21005 0.00347895
R34202 DVSS.n9650 DVSS.n9649 0.00347895
R34203 DVSS.n16167 DVSS.n16166 0.00347895
R34204 DVSS.n16168 DVSS.n16167 0.00347895
R34205 DVSS.n6627 DVSS.n6626 0.00347895
R34206 DVSS.n6626 DVSS.n6625 0.00347895
R34207 DVSS.n3537 DVSS.n3536 0.00347895
R34208 DVSS.n3475 DVSS.n3474 0.00347895
R34209 DVSS.n19175 DVSS.n19174 0.00347895
R34210 DVSS.n20455 DVSS.n20454 0.00347895
R34211 DVSS.n12865 DVSS.n12864 0.00347895
R34212 DVSS.n31 DVSS.n30 0.00347895
R34213 DVSS.n19446 DVSS.n19445 0.00347895
R34214 DVSS.n20184 DVSS.n20183 0.00347895
R34215 DVSS.n18981 DVSS.n18980 0.00347895
R34216 DVSS.n19533 DVSS.n19532 0.00347895
R34217 DVSS.n21514 DVSS.n21513 0.00347895
R34218 DVSS.n19262 DVSS.n19261 0.00347895
R34219 DVSS.n20549 DVSS.n20548 0.00347895
R34220 DVSS.n20275 DVSS.n20274 0.00347895
R34221 DVSS.n583 DVSS.n582 0.00347895
R34222 DVSS.n1232 DVSS.n1231 0.00347895
R34223 DVSS.n21426 DVSS.n21425 0.00347895
R34224 DVSS.n1017 DVSS.n1016 0.00347895
R34225 DVSS.n21007 DVSS.n21006 0.00347895
R34226 DVSS.n20781 DVSS.n20780 0.00347895
R34227 DVSS.n2347 DVSS.n2346 0.00347364
R34228 DVSS.n4138 DVSS.n4137 0.00347
R34229 DVSS.n4225 DVSS.n4223 0.00347
R34230 DVSS.n4178 DVSS.n4176 0.00347
R34231 DVSS.n16581 DVSS.n16580 0.00345775
R34232 DVSS.n16651 DVSS.n16650 0.00345775
R34233 DVSS.n17758 DVSS.n17757 0.00345775
R34234 DVSS.n17760 DVSS.n17759 0.00345775
R34235 DVSS.n18101 DVSS.n18100 0.00345775
R34236 DVSS.n18214 DVSS.n18213 0.00345775
R34237 DVSS.n18425 DVSS.n18424 0.00345775
R34238 DVSS.n18442 DVSS.n18441 0.00345775
R34239 DVSS.n18498 DVSS.n18497 0.00345775
R34240 DVSS.n16768 DVSS.n16767 0.00345775
R34241 DVSS.n17172 DVSS.n17171 0.00345775
R34242 DVSS.n15905 DVSS.n15904 0.00345775
R34243 DVSS.n15903 DVSS.n15902 0.00345775
R34244 DVSS.n15379 DVSS.n15378 0.00345775
R34245 DVSS.n15526 DVSS.n15525 0.00345775
R34246 DVSS.n15204 DVSS.n15203 0.00345775
R34247 DVSS.n15175 DVSS.n15174 0.00345775
R34248 DVSS.n7739 DVSS.n7738 0.00345775
R34249 DVSS.n3349 DVSS.n3348 0.00344838
R34250 DVSS.n16520 DVSS.n16519 0.00342827
R34251 DVSS.n16865 DVSS.n16864 0.00342827
R34252 DVSS.n16521 DVSS.n16520 0.00342827
R34253 DVSS.n16866 DVSS.n16865 0.00342827
R34254 DVSS DVSS.n17189 0.003425
R34255 DVSS.n15106 DVSS 0.003425
R34256 DVSS.n17720 DVSS 0.003425
R34257 DVSS DVSS.n17491 0.003425
R34258 DVSS.n15300 DVSS 0.003425
R34259 DVSS.n15393 DVSS.n15392 0.003425
R34260 DVSS.n15394 DVSS.n15393 0.003425
R34261 DVSS.n18300 DVSS.n18299 0.003425
R34262 DVSS.n18301 DVSS.n18300 0.003425
R34263 DVSS DVSS.n18304 0.003425
R34264 DVSS DVSS.n18039 0.003425
R34265 DVSS DVSS.n17898 0.003425
R34266 DVSS DVSS.n13933 0.003425
R34267 DVSS.n11481 DVSS.n11480 0.00340612
R34268 DVSS.n11518 DVSS.n11517 0.00340612
R34269 DVSS.n11643 DVSS.n11642 0.00340612
R34270 DVSS.n11680 DVSS.n11679 0.00340612
R34271 DVSS.n11729 DVSS.n11728 0.00340612
R34272 DVSS.n4646 DVSS.n4645 0.00339286
R34273 DVSS.n2687 DVSS.n2685 0.00339286
R34274 DVSS.n2633 DVSS.n2631 0.00339286
R34275 DVSS.n11834 DVSS.n11833 0.00339286
R34276 DVSS.n11893 DVSS.n11892 0.00339286
R34277 DVSS.n6045 DVSS.n6044 0.00339286
R34278 DVSS.n6108 DVSS.n6107 0.00339286
R34279 DVSS.n7197 DVSS.n7196 0.00339173
R34280 DVSS.n13523 DVSS.n13522 0.00339173
R34281 DVSS.n13401 DVSS.n13400 0.00339173
R34282 DVSS.n18857 DVSS.n18856 0.00339173
R34283 DVSS.n20256 DVSS.n20255 0.00339144
R34284 DVSS.n20530 DVSS.n20529 0.00339144
R34285 DVSS.n20219 DVSS.n20218 0.00339064
R34286 DVSS.n20490 DVSS.n20489 0.00339064
R34287 DVSS.n5654 DVSS.n5653 0.00339046
R34288 DVSS.n4391 DVSS.n4390 0.00339046
R34289 DVSS.n861 DVSS.n860 0.00339046
R34290 DVSS.n4445 DVSS.n4444 0.00339046
R34291 DVSS.n5653 DVSS.n5652 0.00339046
R34292 DVSS.n10947 DVSS.n10946 0.00339046
R34293 DVSS.n9515 DVSS.n9514 0.00339046
R34294 DVSS.n9574 DVSS.n9573 0.00339046
R34295 DVSS.n12894 DVSS.n12893 0.00339046
R34296 DVSS.n9575 DVSS.n9574 0.00339046
R34297 DVSS.n9514 DVSS.n9513 0.00339046
R34298 DVSS.n10946 DVSS.n10945 0.00339046
R34299 DVSS.n17080 DVSS.n17079 0.00339046
R34300 DVSS.n15682 DVSS.n15681 0.00339046
R34301 DVSS.n15623 DVSS.n15622 0.00339046
R34302 DVSS.n13505 DVSS.n13504 0.00339046
R34303 DVSS.n20304 DVSS.n20303 0.00339046
R34304 DVSS.n20846 DVSS.n20845 0.00339046
R34305 DVSS.n20810 DVSS.n20809 0.00339046
R34306 DVSS.n15683 DVSS.n15682 0.00339046
R34307 DVSS.n15622 DVSS.n15621 0.00339046
R34308 DVSS.n17079 DVSS.n17078 0.00339046
R34309 DVSS.n11553 DVSS.n11552 0.00339046
R34310 DVSS.n11612 DVSS.n11611 0.00339046
R34311 DVSS.n12079 DVSS.n12078 0.00339046
R34312 DVSS.n62 DVSS.n61 0.00339046
R34313 DVSS.n21543 DVSS.n21542 0.00339046
R34314 DVSS.n21483 DVSS.n21482 0.00339046
R34315 DVSS.n21455 DVSS.n21454 0.00339046
R34316 DVSS.n21396 DVSS.n21395 0.00339046
R34317 DVSS.n11613 DVSS.n11612 0.00339046
R34318 DVSS.n11552 DVSS.n11551 0.00339046
R34319 DVSS.n5686 DVSS.n5685 0.00339046
R34320 DVSS.n4695 DVSS.n4694 0.00339046
R34321 DVSS.n4663 DVSS.n4662 0.00339046
R34322 DVSS.n4696 DVSS.n4695 0.00339046
R34323 DVSS.n4339 DVSS.n4338 0.00339046
R34324 DVSS.n4285 DVSS.n4284 0.00339046
R34325 DVSS.n9969 DVSS.n9968 0.00339046
R34326 DVSS.n9679 DVSS.n9678 0.00339046
R34327 DVSS.n9620 DVSS.n9619 0.00339046
R34328 DVSS.n13407 DVSS.n13406 0.00339046
R34329 DVSS.n20578 DVSS.n20577 0.00339046
R34330 DVSS.n21072 DVSS.n21071 0.00339046
R34331 DVSS.n21036 DVSS.n21035 0.00339046
R34332 DVSS.n9680 DVSS.n9679 0.00339046
R34333 DVSS.n9619 DVSS.n9618 0.00339046
R34334 DVSS.n9968 DVSS.n9967 0.00339046
R34335 DVSS.n17373 DVSS.n17372 0.00339046
R34336 DVSS.n17405 DVSS.n17404 0.00339046
R34337 DVSS.n16140 DVSS.n16139 0.00339046
R34338 DVSS.n1148 DVSS.n1147 0.00339046
R34339 DVSS.n16195 DVSS.n16194 0.00339046
R34340 DVSS.n17372 DVSS.n17371 0.00339046
R34341 DVSS.n6654 DVSS.n6653 0.00339046
R34342 DVSS.n18961 DVSS.n18960 0.00339046
R34343 DVSS.n539 DVSS.n538 0.00339046
R34344 DVSS.n556 DVSS.n555 0.00339046
R34345 DVSS.n6599 DVSS.n6598 0.00339046
R34346 DVSS.n3564 DVSS.n3563 0.00339046
R34347 DVSS.n61 DVSS.n60 0.00339046
R34348 DVSS.n12080 DVSS.n12079 0.00339046
R34349 DVSS.n3502 DVSS.n3501 0.00339046
R34350 DVSS.n12895 DVSS.n12894 0.00339046
R34351 DVSS.n18863 DVSS.n18862 0.00339046
R34352 DVSS.n7203 DVSS.n7202 0.00339046
R34353 DVSS.n13408 DVSS.n13407 0.00339046
R34354 DVSS.n13506 DVSS.n13505 0.00339046
R34355 DVSS.n19008 DVSS.n19007 0.00339046
R34356 DVSS.n19560 DVSS.n19559 0.00339046
R34357 DVSS.n21544 DVSS.n21543 0.00339046
R34358 DVSS.n19289 DVSS.n19288 0.00339046
R34359 DVSS.n21484 DVSS.n21483 0.00339046
R34360 DVSS.n21071 DVSS.n21070 0.00339046
R34361 DVSS.n20845 DVSS.n20844 0.00339046
R34362 DVSS.n20579 DVSS.n20578 0.00339046
R34363 DVSS.n20305 DVSS.n20304 0.00339046
R34364 DVSS.n610 DVSS.n609 0.00339046
R34365 DVSS.n1259 DVSS.n1258 0.00339046
R34366 DVSS.n21456 DVSS.n21455 0.00339046
R34367 DVSS.n1044 DVSS.n1043 0.00339046
R34368 DVSS.n21037 DVSS.n21036 0.00339046
R34369 DVSS.n20811 DVSS.n20810 0.00339046
R34370 DVSS.n21395 DVSS.n21394 0.00339046
R34371 DVSS.n12538 DVSS.n12533 0.00338462
R34372 DVSS.n12662 DVSS.n12657 0.00338462
R34373 DVSS.n12570 DVSS.n12565 0.00338462
R34374 DVSS.n12374 DVSS.n12369 0.00338462
R34375 DVSS.n12282 DVSS.n12277 0.00338462
R34376 DVSS.n12259 DVSS.n12258 0.00338462
R34377 DVSS.n3162 DVSS.n3157 0.00338462
R34378 DVSS.n3286 DVSS.n3281 0.00338462
R34379 DVSS.n3194 DVSS.n3189 0.00338462
R34380 DVSS.n3001 DVSS.n2996 0.00338462
R34381 DVSS.n2909 DVSS.n2904 0.00338462
R34382 DVSS.n2886 DVSS.n2885 0.00338462
R34383 DVSS.n9279 DVSS.n9277 0.00338
R34384 DVSS.n9331 DVSS.n9329 0.00338
R34385 DVSS.n9461 DVSS.n9459 0.00338
R34386 DVSS.n16932 DVSS.n16931 0.00337808
R34387 DVSS.n9888 DVSS.n9887 0.00337808
R34388 DVSS.n7163 DVSS.n7161 0.00337234
R34389 DVSS.n1314 DVSS.n1312 0.00337234
R34390 DVSS.n7298 DVSS.n7296 0.00337234
R34391 DVSS.n7313 DVSS.n7311 0.00337234
R34392 DVSS.n7867 DVSS.n7865 0.00337234
R34393 DVSS.n7877 DVSS.n7875 0.00337234
R34394 DVSS.n7955 DVSS.n7953 0.00337234
R34395 DVSS.n7973 DVSS.n7971 0.00337234
R34396 DVSS.n13295 DVSS.n13293 0.00337234
R34397 DVSS.n12182 DVSS.n12181 0.00335984
R34398 DVSS.n5568 DVSS.n5567 0.00333465
R34399 DVSS.n5643 DVSS.n5642 0.00333465
R34400 DVSS.n6507 DVSS.n6506 0.00333465
R34401 DVSS.n4463 DVSS.n4462 0.00333465
R34402 DVSS.n19251 DVSS.n19250 0.00333465
R34403 DVSS.n870 DVSS.n869 0.00333465
R34404 DVSS.n10936 DVSS.n10935 0.00333465
R34405 DVSS.n9496 DVSS.n9495 0.00333465
R34406 DVSS.n12913 DVSS.n12912 0.00333465
R34407 DVSS.n12775 DVSS.n12774 0.00333465
R34408 DVSS.n12484 DVSS.n12483 0.00333465
R34409 DVSS.n12445 DVSS.n12444 0.00333465
R34410 DVSS.n12208 DVSS.n12207 0.00333465
R34411 DVSS.n12171 DVSS.n12170 0.00333465
R34412 DVSS.n12160 DVSS.n12159 0.00333465
R34413 DVSS.n21186 DVSS.n21185 0.00333465
R34414 DVSS.n17069 DVSS.n17068 0.00333465
R34415 DVSS.n15701 DVSS.n15700 0.00333465
R34416 DVSS.n20262 DVSS.n20261 0.00333465
R34417 DVSS.n20855 DVSS.n20854 0.00333465
R34418 DVSS.n10826 DVSS.n10825 0.00333465
R34419 DVSS.n10748 DVSS.n10747 0.00333465
R34420 DVSS.n11534 DVSS.n11533 0.00333465
R34421 DVSS.n12059 DVSS.n12058 0.00333465
R34422 DVSS.n71 DVSS.n70 0.00333465
R34423 DVSS.n21474 DVSS.n21473 0.00333465
R34424 DVSS.n5221 DVSS.n5220 0.00333465
R34425 DVSS.n4713 DVSS.n4712 0.00333465
R34426 DVSS.n4267 DVSS.n4266 0.00333465
R34427 DVSS.n3737 DVSS.n3736 0.00333465
R34428 DVSS.n3387 DVSS.n3386 0.00333465
R34429 DVSS.n3109 DVSS.n3108 0.00333465
R34430 DVSS.n3072 DVSS.n3071 0.00333465
R34431 DVSS.n2838 DVSS.n2837 0.00333465
R34432 DVSS.n2799 DVSS.n2798 0.00333465
R34433 DVSS.n2788 DVSS.n2787 0.00333465
R34434 DVSS.n700 DVSS.n699 0.00333465
R34435 DVSS.n9958 DVSS.n9957 0.00333465
R34436 DVSS.n9698 DVSS.n9697 0.00333465
R34437 DVSS.n20536 DVSS.n20535 0.00333465
R34438 DVSS.n21081 DVSS.n21080 0.00333465
R34439 DVSS.n17263 DVSS.n17262 0.00333465
R34440 DVSS.n17362 DVSS.n17361 0.00333465
R34441 DVSS.n16302 DVSS.n16301 0.00333465
R34442 DVSS.n16213 DVSS.n16212 0.00333465
R34443 DVSS.n19522 DVSS.n19521 0.00333465
R34444 DVSS.n1157 DVSS.n1156 0.00333465
R34445 DVSS.n5438 DVSS.n5437 0.00333465
R34446 DVSS.n5846 DVSS.n5845 0.00333465
R34447 DVSS.n6581 DVSS.n6580 0.00333465
R34448 DVSS.n3654 DVSS.n3653 0.00333465
R34449 DVSS.n18970 DVSS.n18969 0.00333465
R34450 DVSS.n548 DVSS.n547 0.00333465
R34451 DVSS.n4954 DVSS.n4953 0.00332857
R34452 DVSS.n4910 DVSS.n4909 0.00332857
R34453 DVSS.n4851 DVSS.n4850 0.00332857
R34454 DVSS.n10732 DVSS.n10731 0.00332857
R34455 DVSS.n11361 DVSS.n11360 0.00332857
R34456 DVSS.n6227 DVSS.n6226 0.00332857
R34457 DVSS.n6169 DVSS.n6168 0.00332857
R34458 DVSS.n8904 DVSS.n8903 0.00332857
R34459 DVSS.n16526 DVSS.n16525 0.00332274
R34460 DVSS.n16527 DVSS.n16526 0.00332274
R34461 DVSS.n16713 DVSS.n16712 0.00332274
R34462 DVSS.n16714 DVSS.n16713 0.00332274
R34463 DVSS.n14417 DVSS.n14416 0.00332274
R34464 DVSS.n14416 DVSS.n14415 0.00332274
R34465 DVSS.n14711 DVSS.n14710 0.00332274
R34466 DVSS.n14712 DVSS.n14711 0.00332274
R34467 DVSS.n3699 DVSS.n3698 0.00332
R34468 DVSS.n19085 DVSS.n19084 0.00332
R34469 DVSS.n822 DVSS.n821 0.00332
R34470 DVSS.n823 DVSS.n820 0.00332
R34471 DVSS.n19086 DVSS.n19083 0.00332
R34472 DVSS.n3700 DVSS.n3697 0.00332
R34473 DVSS.n16517 DVSS.n16516 0.00330302
R34474 DVSS.n5710 DVSS.n5709 0.00330197
R34475 DVSS.n5766 DVSS.n5765 0.00330197
R34476 DVSS.n4077 DVSS.n4076 0.00330197
R34477 DVSS.n989 DVSS.n988 0.00330197
R34478 DVSS.n5709 DVSS.n5708 0.00330197
R34479 DVSS.n5635 DVSS.n5634 0.00330197
R34480 DVSS.n6975 DVSS.n6974 0.00330197
R34481 DVSS.n10927 DVSS.n10926 0.00330197
R34482 DVSS.n11000 DVSS.n10999 0.00330197
R34483 DVSS.n11270 DVSS.n11269 0.00330197
R34484 DVSS.n8996 DVSS.n8995 0.00330197
R34485 DVSS.n12955 DVSS.n12954 0.00330197
R34486 DVSS.n12676 DVSS.n12675 0.00330197
R34487 DVSS.n12438 DVSS.n12437 0.00330197
R34488 DVSS.n12164 DVSS.n12163 0.00330197
R34489 DVSS.n10999 DVSS.n10998 0.00330197
R34490 DVSS.n8997 DVSS.n8996 0.00330197
R34491 DVSS.n10926 DVSS.n10925 0.00330197
R34492 DVSS.n12954 DVSS.n12953 0.00330197
R34493 DVSS.n11269 DVSS.n11268 0.00330197
R34494 DVSS.n17060 DVSS.n17059 0.00330197
R34495 DVSS.n16907 DVSS.n16906 0.00330197
R34496 DVSS.n17595 DVSS.n17594 0.00330197
R34497 DVSS.n14999 DVSS.n14998 0.00330197
R34498 DVSS.n13664 DVSS.n13663 0.00330197
R34499 DVSS.n20750 DVSS.n20749 0.00330197
R34500 DVSS.n16908 DVSS.n16907 0.00330197
R34501 DVSS.n14998 DVSS.n14997 0.00330197
R34502 DVSS.n17059 DVSS.n17058 0.00330197
R34503 DVSS.n17596 DVSS.n17595 0.00330197
R34504 DVSS.n13663 DVSS.n13662 0.00330197
R34505 DVSS.n10835 DVSS.n10834 0.00330197
R34506 DVSS.n11392 DVSS.n11391 0.00330197
R34507 DVSS.n11696 DVSS.n11695 0.00330197
R34508 DVSS.n13037 DVSS.n13036 0.00330197
R34509 DVSS.n11695 DVSS.n11694 0.00330197
R34510 DVSS.n10836 DVSS.n10835 0.00330197
R34511 DVSS.n11393 DVSS.n11392 0.00330197
R34512 DVSS.n13038 DVSS.n13037 0.00330197
R34513 DVSS.n4705 DVSS.n4704 0.00330197
R34514 DVSS.n3796 DVSS.n3795 0.00330197
R34515 DVSS.n3776 DVSS.n3775 0.00330197
R34516 DVSS.n3300 DVSS.n3299 0.00330197
R34517 DVSS.n3064 DVSS.n3063 0.00330197
R34518 DVSS.n2792 DVSS.n2791 0.00330197
R34519 DVSS.n9949 DVSS.n9948 0.00330197
R34520 DVSS.n9863 DVSS.n9862 0.00330197
R34521 DVSS.n11118 DVSS.n11117 0.00330197
R34522 DVSS.n9086 DVSS.n9085 0.00330197
R34523 DVSS.n13211 DVSS.n13210 0.00330197
R34524 DVSS.n20976 DVSS.n20975 0.00330197
R34525 DVSS.n9864 DVSS.n9863 0.00330197
R34526 DVSS.n9087 DVSS.n9086 0.00330197
R34527 DVSS.n9948 DVSS.n9947 0.00330197
R34528 DVSS.n11119 DVSS.n11118 0.00330197
R34529 DVSS.n13212 DVSS.n13211 0.00330197
R34530 DVSS.n17429 DVSS.n17428 0.00330197
R34531 DVSS.n7542 DVSS.n7541 0.00330197
R34532 DVSS.n18742 DVSS.n18741 0.00330197
R34533 DVSS.n1205 DVSS.n1204 0.00330197
R34534 DVSS.n17428 DVSS.n17427 0.00330197
R34535 DVSS.n17354 DVSS.n17353 0.00330197
R34536 DVSS.n16387 DVSS.n16386 0.00330197
R34537 DVSS.n6076 DVSS.n6075 0.00330197
R34538 DVSS.n6777 DVSS.n6776 0.00330197
R34539 DVSS.n3585 DVSS.n3584 0.00330197
R34540 DVSS.n5430 DVSS.n5429 0.00330197
R34541 DVSS.n3301 DVSS.n3300 0.00330197
R34542 DVSS.n12677 DVSS.n12676 0.00330197
R34543 DVSS.n3065 DVSS.n3064 0.00330197
R34544 DVSS.n20977 DVSS.n20976 0.00330197
R34545 DVSS.n20751 DVSS.n20750 0.00330197
R34546 DVSS.n2793 DVSS.n2792 0.00330197
R34547 DVSS.n12165 DVSS.n12164 0.00330197
R34548 DVSS.n990 DVSS.n989 0.00330197
R34549 DVSS.n5835 DVSS.n4580 0.00327778
R34550 DVSS.n11028 DVSS.n11027 0.00327778
R34551 DVSS.n6472 DVSS.n4526 0.00327778
R34552 DVSS.n11201 DVSS.n11198 0.00327778
R34553 DVSS.n5512 DVSS.n5510 0.00327778
R34554 DVSS.n10039 DVSS.n10038 0.00327778
R34555 DVSS.n3077 DVSS.n3076 0.00327131
R34556 DVSS.n3115 DVSS.n3114 0.00327102
R34557 DVSS.n10071 DVSS.n10070 0.00326429
R34558 DVSS.n10135 DVSS.n10134 0.00326429
R34559 DVSS.n10183 DVSS.n10182 0.00326429
R34560 DVSS.n2688 DVSS.n2687 0.00326429
R34561 DVSS.n2634 DVSS.n2633 0.00326429
R34562 DVSS.n8703 DVSS.n8702 0.00326429
R34563 DVSS.n8766 DVSS.n8765 0.00326429
R34564 DVSS.n8923 DVSS.n8922 0.00326429
R34565 DVSS.n16539 DVSS.n16538 0.00324648
R34566 DVSS.n16652 DVSS.n16651 0.00324648
R34567 DVSS.n17738 DVSS.n17737 0.00324648
R34568 DVSS.n17741 DVSS.n17740 0.00324648
R34569 DVSS.n17743 DVSS.n17742 0.00324648
R34570 DVSS.n18098 DVSS.n18097 0.00324648
R34571 DVSS.n18261 DVSS.n18260 0.00324648
R34572 DVSS.n18221 DVSS.n18220 0.00324648
R34573 DVSS.n14466 DVSS.n14465 0.00324648
R34574 DVSS.n14499 DVSS.n14498 0.00324648
R34575 DVSS.n16726 DVSS.n16725 0.00324648
R34576 DVSS.n17171 DVSS.n17170 0.00324648
R34577 DVSS.n15925 DVSS.n15924 0.00324648
R34578 DVSS.n15922 DVSS.n15921 0.00324648
R34579 DVSS.n15920 DVSS.n15919 0.00324648
R34580 DVSS.n15376 DVSS.n15375 0.00324648
R34581 DVSS.n15479 DVSS.n15478 0.00324648
R34582 DVSS.n15519 DVSS.n15518 0.00324648
R34583 DVSS.n14656 DVSS.n14655 0.00324648
R34584 DVSS.n14623 DVSS.n14622 0.00324648
R34585 DVSS.n16661 DVSS.n16660 0.00321722
R34586 DVSS.n17472 DVSS.n17471 0.00321722
R34587 DVSS.n17735 DVSS.n17734 0.00321722
R34588 DVSS.n17788 DVSS.n17787 0.00321722
R34589 DVSS.n14369 DVSS.n14368 0.00321722
R34590 DVSS.n14455 DVSS.n14454 0.00321722
R34591 DVSS.n156 DVSS.n155 0.00321722
R34592 DVSS.n18209 DVSS.n18208 0.00321722
R34593 DVSS.n17734 DVSS.n17733 0.00321722
R34594 DVSS.n17473 DVSS.n17472 0.00321722
R34595 DVSS.n16660 DVSS.n16659 0.00321722
R34596 DVSS.n17787 DVSS.n17786 0.00321722
R34597 DVSS.n14370 DVSS.n14369 0.00321722
R34598 DVSS.n14475 DVSS.n14474 0.00321722
R34599 DVSS.n17162 DVSS.n17161 0.00321722
R34600 DVSS.n16813 DVSS.n16812 0.00321722
R34601 DVSS.n15928 DVSS.n15927 0.00321722
R34602 DVSS.n15875 DVSS.n15874 0.00321722
R34603 DVSS.n14781 DVSS.n14780 0.00321722
R34604 DVSS.n14667 DVSS.n14666 0.00321722
R34605 DVSS.n316 DVSS.n315 0.00321722
R34606 DVSS.n14651 DVSS.n14644 0.00321722
R34607 DVSS.n15531 DVSS.n15530 0.00321722
R34608 DVSS.n16814 DVSS.n16813 0.00321722
R34609 DVSS.n17163 DVSS.n17162 0.00321722
R34610 DVSS.n15929 DVSS.n15928 0.00321722
R34611 DVSS.n15876 DVSS.n15875 0.00321722
R34612 DVSS.n14780 DVSS.n14779 0.00321722
R34613 DVSS.n14668 DVSS.n14667 0.00321722
R34614 DVSS.n14454 DVSS.n14453 0.00321722
R34615 DVSS.n315 DVSS.n314 0.00321722
R34616 DVSS.n155 DVSS.n154 0.00321722
R34617 DVSS.n5777 DVSS.n5776 0.00321348
R34618 DVSS.n5559 DVSS.n5558 0.00321348
R34619 DVSS.n13132 DVSS.n13131 0.00321348
R34620 DVSS.n13131 DVSS.n13130 0.00321348
R34621 DVSS.n13069 DVSS.n13068 0.00321348
R34622 DVSS.n13070 DVSS.n13069 0.00321348
R34623 DVSS.n9058 DVSS.n9057 0.00321348
R34624 DVSS.n9059 DVSS.n9058 0.00321348
R34625 DVSS.n4051 DVSS.n4050 0.00321348
R34626 DVSS.n7106 DVSS.n7105 0.00321348
R34627 DVSS.n7140 DVSS.n7139 0.00321348
R34628 DVSS.n19208 DVSS.n19207 0.00321348
R34629 DVSS.n10199 DVSS.n10198 0.00321348
R34630 DVSS.n11282 DVSS.n11281 0.00321348
R34631 DVSS.n12926 DVSS.n12925 0.00321348
R34632 DVSS.n11283 DVSS.n11282 0.00321348
R34633 DVSS.n12927 DVSS.n12926 0.00321348
R34634 DVSS.n10200 DVSS.n10199 0.00321348
R34635 DVSS.n16944 DVSS.n16943 0.00321348
R34636 DVSS.n17583 DVSS.n17582 0.00321348
R34637 DVSS.n15027 DVSS.n15026 0.00321348
R34638 DVSS.n13792 DVSS.n13791 0.00321348
R34639 DVSS.n13755 DVSS.n13754 0.00321348
R34640 DVSS.n13707 DVSS.n13706 0.00321348
R34641 DVSS.n13575 DVSS.n13574 0.00321348
R34642 DVSS.n13559 DVSS.n13558 0.00321348
R34643 DVSS.n13553 DVSS.n13552 0.00321348
R34644 DVSS.n17582 DVSS.n17581 0.00321348
R34645 DVSS.n13576 DVSS.n13575 0.00321348
R34646 DVSS.n15026 DVSS.n15025 0.00321348
R34647 DVSS.n13708 DVSS.n13707 0.00321348
R34648 DVSS.n13756 DVSS.n13755 0.00321348
R34649 DVSS.n13793 DVSS.n13792 0.00321348
R34650 DVSS.n16945 DVSS.n16944 0.00321348
R34651 DVSS.n13554 DVSS.n13553 0.00321348
R34652 DVSS.n7139 DVSS.n7138 0.00321348
R34653 DVSS.n13560 DVSS.n13559 0.00321348
R34654 DVSS.n10603 DVSS.n10602 0.00321348
R34655 DVSS.n11380 DVSS.n11379 0.00321348
R34656 DVSS.n12046 DVSS.n12045 0.00321348
R34657 DVSS.n11684 DVSS.n11683 0.00321348
R34658 DVSS.n11647 DVSS.n11646 0.00321348
R34659 DVSS.n11522 DVSS.n11521 0.00321348
R34660 DVSS.n11485 DVSS.n11484 0.00321348
R34661 DVSS.n11379 DVSS.n11378 0.00321348
R34662 DVSS.n12045 DVSS.n12044 0.00321348
R34663 DVSS.n10604 DVSS.n10603 0.00321348
R34664 DVSS.n13057 DVSS.n13056 0.00321348
R34665 DVSS.n5212 DVSS.n5211 0.00321348
R34666 DVSS.n3984 DVSS.n3983 0.00321348
R34667 DVSS.n3750 DVSS.n3749 0.00321348
R34668 DVSS.n9900 DVSS.n9899 0.00321348
R34669 DVSS.n11106 DVSS.n11105 0.00321348
R34670 DVSS.n13235 DVSS.n13234 0.00321348
R34671 DVSS.n13257 DVSS.n13256 0.00321348
R34672 DVSS.n13361 DVSS.n13360 0.00321348
R34673 DVSS.n11105 DVSS.n11104 0.00321348
R34674 DVSS.n13256 DVSS.n13255 0.00321348
R34675 DVSS.n9901 DVSS.n9900 0.00321348
R34676 DVSS.n13234 DVSS.n13233 0.00321348
R34677 DVSS.n13360 DVSS.n13359 0.00321348
R34678 DVSS.n7516 DVSS.n7515 0.00321348
R34679 DVSS.n18629 DVSS.n18628 0.00321348
R34680 DVSS.n18656 DVSS.n18655 0.00321348
R34681 DVSS.n18688 DVSS.n18687 0.00321348
R34682 DVSS.n18765 DVSS.n18764 0.00321348
R34683 DVSS.n18785 DVSS.n18784 0.00321348
R34684 DVSS.n18822 DVSS.n18821 0.00321348
R34685 DVSS.n19479 DVSS.n19478 0.00321348
R34686 DVSS.n18628 DVSS.n18627 0.00321348
R34687 DVSS.n18655 DVSS.n18654 0.00321348
R34688 DVSS.n18687 DVSS.n18686 0.00321348
R34689 DVSS.n18821 DVSS.n18820 0.00321348
R34690 DVSS.n18764 DVSS.n18763 0.00321348
R34691 DVSS.n16398 DVSS.n16397 0.00321348
R34692 DVSS.n17254 DVSS.n17253 0.00321348
R34693 DVSS.n5317 DVSS.n5316 0.00321348
R34694 DVSS.n5839 DVSS.n5838 0.00321348
R34695 DVSS.n6065 DVSS.n6064 0.00321348
R34696 DVSS.n6832 DVSS.n6831 0.00321348
R34697 DVSS.n3641 DVSS.n3640 0.00321348
R34698 DVSS.n5838 DVSS.n5837 0.00321348
R34699 DVSS.n20489 DVSS.n20488 0.00321348
R34700 DVSS.n20218 DVSS.n20217 0.00321348
R34701 DVSS.n19478 DVSS.n19477 0.00321348
R34702 DVSS.n19207 DVSS.n19206 0.00321348
R34703 DVSS.n17214 DVSS.n17213 0.0032
R34704 DVSS.n15182 DVSS.n15181 0.0032
R34705 DVSS.n15149 DVSS.n15148 0.0032
R34706 DVSS.n15107 DVSS.n15106 0.0032
R34707 DVSS.n17692 DVSS.n17691 0.0032
R34708 DVSS.n17681 DVSS.n17680 0.0032
R34709 DVSS.n10066 DVSS.n10065 0.0032
R34710 DVSS.n10130 DVSS.n10129 0.0032
R34711 DVSS.n10178 DVSS.n10177 0.0032
R34712 DVSS.n8698 DVSS.n8697 0.0032
R34713 DVSS.n8761 DVSS.n8760 0.0032
R34714 DVSS.n8862 DVSS.n8861 0.0032
R34715 DVSS.n10803 DVSS.n10802 0.0031825
R34716 DVSS.n19594 DVSS.n1302 0.00316667
R34717 DVSS.n20673 DVSS.n80 0.00316667
R34718 DVSS.n19594 DVSS.n18919 0.00316667
R34719 DVSS.n20079 DVSS.n81 0.00316667
R34720 DVSS.n20079 DVSS.n504 0.00316667
R34721 DVSS.n21107 DVSS.n20673 0.00316667
R34722 DVSS.n17798 DVSS.n17797 0.00316244
R34723 DVSS.n17765 DVSS.n17764 0.00316244
R34724 DVSS.n17772 DVSS.n17771 0.00316244
R34725 DVSS.n15898 DVSS.n15897 0.00316244
R34726 DVSS.n5803 DVSS.n5802 0.00315748
R34727 DVSS.n5785 DVSS.n5784 0.00315748
R34728 DVSS.n5740 DVSS.n5739 0.00315748
R34729 DVSS.n4059 DVSS.n4058 0.00315748
R34730 DVSS.n7098 DVSS.n7097 0.00315748
R34731 DVSS.n9851 DVSS.n9850 0.00315748
R34732 DVSS.n11292 DVSS.n11291 0.00315748
R34733 DVSS.n13122 DVSS.n13121 0.00315748
R34734 DVSS.n12936 DVSS.n12935 0.00315748
R34735 DVSS.n12689 DVSS.n12688 0.00315748
R34736 DVSS.n12476 DVSS.n12475 0.00315748
R34737 DVSS.n12395 DVSS.n12394 0.00315748
R34738 DVSS.n12204 DVSS.n12203 0.00315748
R34739 DVSS.n21290 DVSS.n21289 0.00315748
R34740 DVSS.n21243 DVSS.n21242 0.00315748
R34741 DVSS.n21316 DVSS.n21315 0.00315748
R34742 DVSS.n17555 DVSS.n17554 0.00315748
R34743 DVSS.n17573 DVSS.n17572 0.00315748
R34744 DVSS.n15017 DVSS.n15016 0.00315748
R34745 DVSS.n13585 DVSS.n13584 0.00315748
R34746 DVSS.n10764 DVSS.n10763 0.00315748
R34747 DVSS.n10754 DVSS.n10753 0.00315748
R34748 DVSS.n10737 DVSS.n10736 0.00315748
R34749 DVSS.n11370 DVSS.n11369 0.00315748
R34750 DVSS.n11421 DVSS.n11420 0.00315748
R34751 DVSS.n13079 DVSS.n13078 0.00315748
R34752 DVSS.n12036 DVSS.n12035 0.00315748
R34753 DVSS.n3976 DVSS.n3975 0.00315748
R34754 DVSS.n3758 DVSS.n3757 0.00315748
R34755 DVSS.n3312 DVSS.n3311 0.00315748
R34756 DVSS.n3102 DVSS.n3101 0.00315748
R34757 DVSS.n3021 DVSS.n3020 0.00315748
R34758 DVSS.n2834 DVSS.n2833 0.00315748
R34759 DVSS.n740 DVSS.n739 0.00315748
R34760 DVSS.n774 DVSS.n773 0.00315748
R34761 DVSS.n674 DVSS.n673 0.00315748
R34762 DVSS.n11078 DVSS.n11077 0.00315748
R34763 DVSS.n11096 DVSS.n11095 0.00315748
R34764 DVSS.n9068 DVSS.n9067 0.00315748
R34765 DVSS.n13247 DVSS.n13246 0.00315748
R34766 DVSS.n16424 DVSS.n16423 0.00315748
R34767 DVSS.n16406 DVSS.n16405 0.00315748
R34768 DVSS.n16361 DVSS.n16360 0.00315748
R34769 DVSS.n7524 DVSS.n7523 0.00315748
R34770 DVSS.n18777 DVSS.n18776 0.00315748
R34771 DVSS.n5490 DVSS.n5489 0.00315748
R34772 DVSS.n5840 DVSS.n5839 0.00315748
R34773 DVSS.n5856 DVSS.n5855 0.00315748
R34774 DVSS.n6057 DVSS.n6056 0.00315748
R34775 DVSS.n6343 DVSS.n6342 0.00315748
R34776 DVSS.n6824 DVSS.n6823 0.00315748
R34777 DVSS.n3633 DVSS.n3632 0.00315748
R34778 DVSS.n14174 DVSS.n14173 0.00315322
R34779 DVSS.n14736 DVSS.n14735 0.00315322
R34780 DVSS.n14173 DVSS.n14172 0.00315322
R34781 DVSS.n14735 DVSS.n14734 0.00315322
R34782 DVSS.n9252 DVSS.n9251 0.00314
R34783 DVSS.n9304 DVSS.n9303 0.00314
R34784 DVSS.n9340 DVSS.n9339 0.00314
R34785 DVSS.n9474 DVSS.n9473 0.00314
R34786 DVSS.n21363 DVSS.n21362 0.00314
R34787 DVSS.n5627 DVSS.n5626 0.00312498
R34788 DVSS.n5656 DVSS.n5655 0.00312498
R34789 DVSS.n5667 DVSS.n5666 0.00312498
R34790 DVSS.n5687 DVSS.n5686 0.00312498
R34791 DVSS.n5699 DVSS.n5698 0.00312498
R34792 DVSS.n7114 DVSS.n7113 0.00312498
R34793 DVSS.n983 DVSS.n982 0.00312498
R34794 DVSS.n10918 DVSS.n10917 0.00312498
R34795 DVSS.n10949 DVSS.n10948 0.00312498
R34796 DVSS.n10959 DVSS.n10958 0.00312498
R34797 DVSS.n10978 DVSS.n10977 0.00312498
R34798 DVSS.n10989 DVSS.n10988 0.00312498
R34799 DVSS.n12746 DVSS.n12745 0.00312498
R34800 DVSS.n10917 DVSS.n10916 0.00312498
R34801 DVSS.n17051 DVSS.n17050 0.00312498
R34802 DVSS.n17082 DVSS.n17081 0.00312498
R34803 DVSS.n17092 DVSS.n17091 0.00312498
R34804 DVSS.n16929 DVSS.n16928 0.00312498
R34805 DVSS.n16918 DVSS.n16917 0.00312498
R34806 DVSS.n13827 DVSS.n13826 0.00312498
R34807 DVSS.n13789 DVSS.n13788 0.00312498
R34808 DVSS.n13752 DVSS.n13751 0.00312498
R34809 DVSS.n13567 DVSS.n13566 0.00312498
R34810 DVSS.n13561 DVSS.n13560 0.00312498
R34811 DVSS.n20745 DVSS.n20744 0.00312498
R34812 DVSS.n13828 DVSS.n13827 0.00312498
R34813 DVSS.n13790 DVSS.n13789 0.00312498
R34814 DVSS.n13753 DVSS.n13752 0.00312498
R34815 DVSS.n17050 DVSS.n17049 0.00312498
R34816 DVSS.n13562 DVSS.n13561 0.00312498
R34817 DVSS.n13568 DVSS.n13567 0.00312498
R34818 DVSS.n7113 DVSS.n7112 0.00312498
R34819 DVSS.n10844 DVSS.n10843 0.00312498
R34820 DVSS.n10757 DVSS.n10756 0.00312498
R34821 DVSS.n11428 DVSS.n11427 0.00312498
R34822 DVSS.n11484 DVSS.n11457 0.00312498
R34823 DVSS.n11521 DVSS.n11494 0.00312498
R34824 DVSS.n11646 DVSS.n11619 0.00312498
R34825 DVSS.n11683 DVSS.n11656 0.00312498
R34826 DVSS.n11427 DVSS.n11426 0.00312498
R34827 DVSS.n10758 DVSS.n10757 0.00312498
R34828 DVSS.n10845 DVSS.n10844 0.00312498
R34829 DVSS.n13058 DVSS.n13057 0.00312498
R34830 DVSS.n5698 DVSS.n5697 0.00312498
R34831 DVSS.n16930 DVSS.n16929 0.00312498
R34832 DVSS.n5666 DVSS.n5665 0.00312498
R34833 DVSS.n10958 DVSS.n10957 0.00312498
R34834 DVSS.n10988 DVSS.n10987 0.00312498
R34835 DVSS.n10977 DVSS.n10976 0.00312498
R34836 DVSS.n10948 DVSS.n10947 0.00312498
R34837 DVSS.n5655 DVSS.n5654 0.00312498
R34838 DVSS.n17081 DVSS.n17080 0.00312498
R34839 DVSS.n17091 DVSS.n17090 0.00312498
R34840 DVSS.n5688 DVSS.n5687 0.00312498
R34841 DVSS.n16919 DVSS.n16918 0.00312498
R34842 DVSS.n5193 DVSS.n5192 0.00312498
R34843 DVSS.n4693 DVSS.n4692 0.00312498
R34844 DVSS.n4682 DVSS.n4681 0.00312498
R34845 DVSS.n4662 DVSS.n4661 0.00312498
R34846 DVSS.n4650 DVSS.n4649 0.00312498
R34847 DVSS.n4651 DVSS.n4650 0.00312498
R34848 DVSS.n4683 DVSS.n4682 0.00312498
R34849 DVSS.n4694 DVSS.n4693 0.00312498
R34850 DVSS.n4661 DVSS.n4660 0.00312498
R34851 DVSS.n3359 DVSS.n3358 0.00312498
R34852 DVSS.n735 DVSS.n732 0.00312498
R34853 DVSS.n9940 DVSS.n9939 0.00312498
R34854 DVSS.n9971 DVSS.n9970 0.00312498
R34855 DVSS.n9981 DVSS.n9980 0.00312498
R34856 DVSS.n9885 DVSS.n9884 0.00312498
R34857 DVSS.n9874 DVSS.n9873 0.00312498
R34858 DVSS.n13265 DVSS.n13264 0.00312498
R34859 DVSS.n20971 DVSS.n20970 0.00312498
R34860 DVSS.n13264 DVSS.n13263 0.00312498
R34861 DVSS.n9980 DVSS.n9979 0.00312498
R34862 DVSS.n9939 DVSS.n9938 0.00312498
R34863 DVSS.n9970 DVSS.n9969 0.00312498
R34864 DVSS.n9875 DVSS.n9874 0.00312498
R34865 DVSS.n9886 DVSS.n9885 0.00312498
R34866 DVSS.n17375 DVSS.n17374 0.00312498
R34867 DVSS.n17386 DVSS.n17385 0.00312498
R34868 DVSS.n17407 DVSS.n17406 0.00312498
R34869 DVSS.n17418 DVSS.n17417 0.00312498
R34870 DVSS.n18605 DVSS.n18604 0.00312498
R34871 DVSS.n18632 DVSS.n18631 0.00312498
R34872 DVSS.n18659 DVSS.n18658 0.00312498
R34873 DVSS.n18793 DVSS.n18792 0.00312498
R34874 DVSS.n1200 DVSS.n1199 0.00312498
R34875 DVSS.n18792 DVSS.n18791 0.00312498
R34876 DVSS.n18604 DVSS.n18603 0.00312498
R34877 DVSS.n18631 DVSS.n18630 0.00312498
R34878 DVSS.n18658 DVSS.n18657 0.00312498
R34879 DVSS.n17417 DVSS.n17416 0.00312498
R34880 DVSS.n17406 DVSS.n17405 0.00312498
R34881 DVSS.n17385 DVSS.n17384 0.00312498
R34882 DVSS.n17374 DVSS.n17373 0.00312498
R34883 DVSS.n17346 DVSS.n17345 0.00312498
R34884 DVSS.n1199 DVSS.n1198 0.00312498
R34885 DVSS.n5422 DVSS.n5421 0.00312498
R34886 DVSS.n6441 DVSS.n6440 0.00312498
R34887 DVSS.n6352 DVSS.n6351 0.00312498
R34888 DVSS.n6661 DVSS.n6660 0.00312498
R34889 DVSS.n6722 DVSS.n6721 0.00312498
R34890 DVSS.n6843 DVSS.n6842 0.00312498
R34891 DVSS.n3360 DVSS.n3359 0.00312498
R34892 DVSS.n12747 DVSS.n12746 0.00312498
R34893 DVSS.n735 DVSS.n734 0.00312498
R34894 DVSS.n20972 DVSS.n20971 0.00312498
R34895 DVSS.n20746 DVSS.n20745 0.00312498
R34896 DVSS.n21252 DVSS.n21251 0.00312498
R34897 DVSS.n984 DVSS.n983 0.00312498
R34898 DVSS.n14722 DVSS.n14721 0.00311264
R34899 DVSS.n14406 DVSS.n14405 0.00311264
R34900 DVSS.n18440 DVSS.n18439 0.00311219
R34901 DVSS.n15177 DVSS.n15176 0.00311219
R34902 DVSS.n18156 DVSS.n18155 0.00311168
R34903 DVSS.n18176 DVSS.n18175 0.00311168
R34904 DVSS.n14218 DVSS.n14217 0.00311168
R34905 DVSS.n14505 DVSS.n14504 0.00311168
R34906 DVSS.n19717 DVSS.n19716 0.00311168
R34907 DVSS.n19795 DVSS.n19794 0.00311168
R34908 DVSS.n148 DVSS.n147 0.00311168
R34909 DVSS.n236 DVSS.n235 0.00311168
R34910 DVSS.n185 DVSS.n184 0.00311168
R34911 DVSS.n14217 DVSS.n14216 0.00311168
R34912 DVSS.n18177 DVSS.n18176 0.00311168
R34913 DVSS.n18259 DVSS.n18258 0.00311168
R34914 DVSS.n18155 DVSS.n18154 0.00311168
R34915 DVSS.n18486 DVSS.n18485 0.00311168
R34916 DVSS.n15461 DVSS.n15460 0.00311168
R34917 DVSS.n15481 DVSS.n15480 0.00311168
R34918 DVSS.n15564 DVSS.n15563 0.00311168
R34919 DVSS.n7727 DVSS.n7711 0.00311168
R34920 DVSS.n14879 DVSS.n14878 0.00311168
R34921 DVSS.n14602 DVSS.n14601 0.00311168
R34922 DVSS.n19936 DVSS.n19935 0.00311168
R34923 DVSS.n20020 DVSS.n20019 0.00311168
R34924 DVSS.n308 DVSS.n307 0.00311168
R34925 DVSS.n444 DVSS.n443 0.00311168
R34926 DVSS.n393 DVSS.n392 0.00311168
R34927 DVSS.n15460 DVSS.n15459 0.00311168
R34928 DVSS.n15563 DVSS.n15562 0.00311168
R34929 DVSS.n14880 DVSS.n14879 0.00311168
R34930 DVSS.n19716 DVSS.n19715 0.00311168
R34931 DVSS.n14603 DVSS.n14602 0.00311168
R34932 DVSS.n14506 DVSS.n14505 0.00311168
R34933 DVSS.n19935 DVSS.n19934 0.00311168
R34934 DVSS.n147 DVSS.n146 0.00311168
R34935 DVSS.n307 DVSS.n306 0.00311168
R34936 DVSS.n20021 DVSS.n20020 0.00311168
R34937 DVSS.n19796 DVSS.n19795 0.00311168
R34938 DVSS.n445 DVSS.n444 0.00311168
R34939 DVSS.n237 DVSS.n236 0.00311168
R34940 DVSS.n184 DVSS.n183 0.00311168
R34941 DVSS.n392 DVSS.n391 0.00311168
R34942 DVSS.n3308 DVSS.n3307 0.00309404
R34943 DVSS.n17876 DVSS.n17875 0.00309215
R34944 DVSS.n18017 DVSS.n18016 0.00309215
R34945 DVSS.n18163 DVSS.n18162 0.00309215
R34946 DVSS.n7568 DVSS.n7567 0.00309215
R34947 DVSS.n14445 DVSS.n14444 0.00309215
R34948 DVSS.n15739 DVSS.n15738 0.00309215
R34949 DVSS.n15823 DVSS.n15822 0.00309215
R34950 DVSS.n15241 DVSS.n15240 0.00309215
R34951 DVSS.n15577 DVSS.n15576 0.00309215
R34952 DVSS.n18520 DVSS.n18519 0.00309215
R34953 DVSS.n7761 DVSS.n7760 0.00309215
R34954 DVSS.n4949 DVSS.n4948 0.00307143
R34955 DVSS.n4905 DVSS.n4904 0.00307143
R34956 DVSS.n4846 DVSS.n4845 0.00307143
R34957 DVSS.n6222 DVSS.n6221 0.00307143
R34958 DVSS.n6164 DVSS.n6163 0.00307143
R34959 DVSS.n1391 DVSS.n1390 0.00305
R34960 DVSS.n4234 DVSS.n4233 0.00305
R34961 DVSS.n4203 DVSS.n4202 0.00305
R34962 DVSS.n4157 DVSS.n4156 0.00305
R34963 DVSS.n3672 DVSS.n3671 0.00305
R34964 DVSS.n19025 DVSS.n19024 0.00305
R34965 DVSS.n634 DVSS.n633 0.00305
R34966 DVSS.n5682 DVSS.n5681 0.00303648
R34967 DVSS.n5624 DVSS.n5623 0.00303648
R34968 DVSS.n10914 DVSS.n10913 0.00303648
R34969 DVSS.n10913 DVSS.n10912 0.00303648
R34970 DVSS.n17047 DVSS.n17046 0.00303648
R34971 DVSS.n16934 DVSS.n16933 0.00303648
R34972 DVSS.n17046 DVSS.n17045 0.00303648
R34973 DVSS.n10848 DVSS.n10847 0.00303648
R34974 DVSS.n10796 DVSS.n10795 0.00303648
R34975 DVSS.n10849 DVSS.n10848 0.00303648
R34976 DVSS.n5681 DVSS.n5680 0.00303648
R34977 DVSS.n16935 DVSS.n16934 0.00303648
R34978 DVSS.n10797 DVSS.n10796 0.00303648
R34979 DVSS.n5196 DVSS.n5195 0.00303648
R34980 DVSS.n9936 DVSS.n9935 0.00303648
R34981 DVSS.n9935 DVSS.n9934 0.00303648
R34982 DVSS.n17401 DVSS.n17400 0.00303648
R34983 DVSS.n17400 DVSS.n17399 0.00303648
R34984 DVSS.n17343 DVSS.n17342 0.00303648
R34985 DVSS.n5468 DVSS.n5467 0.00303648
R34986 DVSS.n5419 DVSS.n5418 0.00303648
R34987 DVSS.n5467 DVSS.n5466 0.00303648
R34988 DVSS.n10973 DVSS.n10972 0.00303648
R34989 DVSS.n10972 DVSS.n10971 0.00303648
R34990 DVSS.n4667 DVSS.n4666 0.00303648
R34991 DVSS.n4668 DVSS.n4667 0.00303648
R34992 DVSS.n9890 DVSS.n9889 0.00303648
R34993 DVSS.n9891 DVSS.n9890 0.00303648
R34994 DVSS.n16576 DVSS.n16575 0.00303521
R34995 DVSS.n16650 DVSS.n16649 0.00303521
R34996 DVSS.n16090 DVSS.n16089 0.00303521
R34997 DVSS.n17740 DVSS.n17739 0.00303521
R34998 DVSS.n17759 DVSS.n17758 0.00303521
R34999 DVSS.n17774 DVSS.n17773 0.00303521
R35000 DVSS.n18196 DVSS.n18195 0.00303521
R35001 DVSS.n18193 DVSS.n18192 0.00303521
R35002 DVSS.n18424 DVSS.n18423 0.00303521
R35003 DVSS.n18452 DVSS.n18451 0.00303521
R35004 DVSS.n18495 DVSS.n18494 0.00303521
R35005 DVSS.n18497 DVSS.n18496 0.00303521
R35006 DVSS.n14385 DVSS.n14384 0.00303521
R35007 DVSS.n14426 DVSS.n14425 0.00303521
R35008 DVSS.n14500 DVSS.n14499 0.00303521
R35009 DVSS.n16763 DVSS.n16762 0.00303521
R35010 DVSS.n17173 DVSS.n17172 0.00303521
R35011 DVSS.n15978 DVSS.n15977 0.00303521
R35012 DVSS.n15923 DVSS.n15922 0.00303521
R35013 DVSS.n15904 DVSS.n15903 0.00303521
R35014 DVSS.n15889 DVSS.n15888 0.00303521
R35015 DVSS.n15544 DVSS.n15543 0.00303521
R35016 DVSS.n15547 DVSS.n15546 0.00303521
R35017 DVSS.n15205 DVSS.n15204 0.00303521
R35018 DVSS.n15165 DVSS.n15164 0.00303521
R35019 DVSS.n7736 DVSS.n7735 0.00303521
R35020 DVSS.n7738 DVSS.n7737 0.00303521
R35021 DVSS.n14765 DVSS.n14764 0.00303521
R35022 DVSS.n14702 DVSS.n14701 0.00303521
R35023 DVSS.n14622 DVSS.n14621 0.00303521
R35024 DVSS.n17877 DVSS.n17876 0.00302184
R35025 DVSS.n18018 DVSS.n18017 0.00302184
R35026 DVSS.n18164 DVSS.n18163 0.00302184
R35027 DVSS.n7569 DVSS.n7568 0.00302184
R35028 DVSS.n15883 DVSS.n15882 0.00302184
R35029 DVSS.n14693 DVSS.n14692 0.00302184
R35030 DVSS.n15822 DVSS.n15821 0.00302184
R35031 DVSS.n15740 DVSS.n15739 0.00302184
R35032 DVSS.n15576 DVSS.n15575 0.00302184
R35033 DVSS.n15240 DVSS.n15239 0.00302184
R35034 DVSS.n18519 DVSS.n18518 0.00302184
R35035 DVSS.n7760 DVSS.n7759 0.00302184
R35036 DVSS.n16708 DVSS.n16707 0.00302184
R35037 DVSS.n17115 DVSS.n17114 0.00302184
R35038 DVSS.n17464 DVSS.n17457 0.00302184
R35039 DVSS.n14444 DVSS.n14443 0.00302184
R35040 DVSS.n17539 DVSS.n17538 0.00302184
R35041 DVSS.n18184 DVSS.n18183 0.00300702
R35042 DVSS.n15556 DVSS.n15555 0.00300702
R35043 DVSS.n16705 DVSS.n16704 0.00300615
R35044 DVSS.n16510 DVSS.n16509 0.00300615
R35045 DVSS.n19687 DVSS.n19686 0.00300615
R35046 DVSS.n19695 DVSS.n19694 0.00300615
R35047 DVSS.n19773 DVSS.n19772 0.00300615
R35048 DVSS.n19765 DVSS.n19764 0.00300615
R35049 DVSS.n214 DVSS.n213 0.00300615
R35050 DVSS.n206 DVSS.n205 0.00300615
R35051 DVSS.n18135 DVSS.n18134 0.00300615
R35052 DVSS.n18454 DVSS.n18453 0.00300615
R35053 DVSS.n18483 DVSS.n18482 0.00300615
R35054 DVSS.n16704 DVSS.n16703 0.00300615
R35055 DVSS.n16511 DVSS.n16510 0.00300615
R35056 DVSS.n17118 DVSS.n17117 0.00300615
R35057 DVSS.n16856 DVSS.n16855 0.00300615
R35058 DVSS.n15163 DVSS.n15162 0.00300615
R35059 DVSS.n15119 DVSS.n15118 0.00300615
R35060 DVSS.n19906 DVSS.n19905 0.00300615
R35061 DVSS.n19914 DVSS.n19913 0.00300615
R35062 DVSS.n19998 DVSS.n19997 0.00300615
R35063 DVSS.n19990 DVSS.n19989 0.00300615
R35064 DVSS.n422 DVSS.n421 0.00300615
R35065 DVSS.n414 DVSS.n413 0.00300615
R35066 DVSS.n15440 DVSS.n15439 0.00300615
R35067 DVSS.n17119 DVSS.n17118 0.00300615
R35068 DVSS.n16857 DVSS.n16856 0.00300615
R35069 DVSS.n19686 DVSS.n19685 0.00300615
R35070 DVSS.n19913 DVSS.n19912 0.00300615
R35071 DVSS.n19694 DVSS.n19693 0.00300615
R35072 DVSS.n19905 DVSS.n19904 0.00300615
R35073 DVSS.n19774 DVSS.n19773 0.00300615
R35074 DVSS.n19999 DVSS.n19998 0.00300615
R35075 DVSS.n19991 DVSS.n19990 0.00300615
R35076 DVSS.n19766 DVSS.n19765 0.00300615
R35077 DVSS.n215 DVSS.n214 0.00300615
R35078 DVSS.n423 DVSS.n422 0.00300615
R35079 DVSS.n415 DVSS.n414 0.00300615
R35080 DVSS.n207 DVSS.n206 0.00300615
R35081 DVSS.n6336 DVSS.n6335 0.00300558
R35082 DVSS.n11022 DVSS.n11021 0.003
R35083 DVSS.n11020 DVSS.n11019 0.003
R35084 DVSS.n11192 DVSS.n11191 0.003
R35085 DVSS.n11190 DVSS.n11189 0.003
R35086 DVSS.n12508 DVSS.n12503 0.003
R35087 DVSS.n12509 DVSS.n12508 0.003
R35088 DVSS.n12633 DVSS.n12632 0.003
R35089 DVSS.n12632 DVSS.n12627 0.003
R35090 DVSS.n12345 DVSS.n12344 0.003
R35091 DVSS.n12344 DVSS.n12339 0.003
R35092 DVSS.n21218 DVSS.n21213 0.003
R35093 DVSS.n21220 DVSS.n21218 0.003
R35094 DVSS.n10032 DVSS.n10031 0.003
R35095 DVSS.n10030 DVSS.n10029 0.003
R35096 DVSS.n3132 DVSS.n3127 0.003
R35097 DVSS.n3133 DVSS.n3132 0.003
R35098 DVSS.n3257 DVSS.n3256 0.003
R35099 DVSS.n3256 DVSS.n3251 0.003
R35100 DVSS.n2972 DVSS.n2971 0.003
R35101 DVSS.n2971 DVSS.n2966 0.003
R35102 DVSS.n906 DVSS.n901 0.003
R35103 DVSS.n907 DVSS.n906 0.003
R35104 DVSS.n3392 DVSS.n3391 0.003
R35105 DVSS.n3393 DVSS.n3392 0.003
R35106 DVSS.n12798 DVSS.n12797 0.003
R35107 DVSS.n12797 DVSS.n12796 0.003
R35108 DVSS.n5619 DVSS.n5618 0.00298032
R35109 DVSS.n10908 DVSS.n10907 0.00298032
R35110 DVSS.n17041 DVSS.n17040 0.00298032
R35111 DVSS.n10854 DVSS.n10853 0.00298032
R35112 DVSS.n5201 DVSS.n5200 0.00298032
R35113 DVSS.n9930 DVSS.n9929 0.00298032
R35114 DVSS.n17338 DVSS.n17337 0.00298032
R35115 DVSS.n5414 DVSS.n5413 0.00298032
R35116 DVSS.n16591 DVSS.n16590 0.002975
R35117 DVSS.n15212 DVSS.n15211 0.002975
R35118 DVSS.n16495 DVSS.n16494 0.002975
R35119 DVSS.n15362 DVSS.n15361 0.002975
R35120 DVSS.n18092 DVSS.n18091 0.002975
R35121 DVSS.n15430 DVSS.n15429 0.002975
R35122 DVSS.n18282 DVSS.n18281 0.002975
R35123 DVSS.n18331 DVSS.n18330 0.002975
R35124 DVSS.n18344 DVSS.n18343 0.002975
R35125 DVSS.n17951 DVSS.n17950 0.002975
R35126 DVSS.n17810 DVSS.n17809 0.002975
R35127 DVSS.n13860 DVSS.n13859 0.002975
R35128 DVSS.n5556 DVSS.n5555 0.00294798
R35129 DVSS.n5780 DVSS.n5779 0.00294798
R35130 DVSS.n7103 DVSS.n7102 0.00294798
R35131 DVSS.n4054 DVSS.n4053 0.00294798
R35132 DVSS.n10196 DVSS.n10195 0.00294798
R35133 DVSS.n11286 DVSS.n11285 0.00294798
R35134 DVSS.n13128 DVSS.n13127 0.00294798
R35135 DVSS.n12930 DVSS.n12929 0.00294798
R35136 DVSS.n12931 DVSS.n12930 0.00294798
R35137 DVSS.n13127 DVSS.n13126 0.00294798
R35138 DVSS.n10195 DVSS.n10194 0.00294798
R35139 DVSS.n11287 DVSS.n11286 0.00294798
R35140 DVSS.n16941 DVSS.n16940 0.00294798
R35141 DVSS.n17579 DVSS.n17578 0.00294798
R35142 DVSS.n15023 DVSS.n15022 0.00294798
R35143 DVSS.n13579 DVSS.n13578 0.00294798
R35144 DVSS.n13580 DVSS.n13579 0.00294798
R35145 DVSS.n15022 DVSS.n15021 0.00294798
R35146 DVSS.n16940 DVSS.n16939 0.00294798
R35147 DVSS.n17578 DVSS.n17577 0.00294798
R35148 DVSS.n10600 DVSS.n10599 0.00294798
R35149 DVSS.n11376 DVSS.n11375 0.00294798
R35150 DVSS.n13073 DVSS.n13072 0.00294798
R35151 DVSS.n12042 DVSS.n12041 0.00294798
R35152 DVSS.n12041 DVSS.n12040 0.00294798
R35153 DVSS.n13074 DVSS.n13073 0.00294798
R35154 DVSS.n11375 DVSS.n11374 0.00294798
R35155 DVSS.n10599 DVSS.n10598 0.00294798
R35156 DVSS.n5209 DVSS.n5208 0.00294798
R35157 DVSS.n3753 DVSS.n3752 0.00294798
R35158 DVSS.n3981 DVSS.n3980 0.00294798
R35159 DVSS.n9897 DVSS.n9896 0.00294798
R35160 DVSS.n11102 DVSS.n11101 0.00294798
R35161 DVSS.n9062 DVSS.n9061 0.00294798
R35162 DVSS.n13253 DVSS.n13252 0.00294798
R35163 DVSS.n13252 DVSS.n13251 0.00294798
R35164 DVSS.n9063 DVSS.n9062 0.00294798
R35165 DVSS.n9896 DVSS.n9895 0.00294798
R35166 DVSS.n11101 DVSS.n11100 0.00294798
R35167 DVSS.n7519 DVSS.n7518 0.00294798
R35168 DVSS.n18782 DVSS.n18781 0.00294798
R35169 DVSS.n16401 DVSS.n16400 0.00294798
R35170 DVSS.n17251 DVSS.n17250 0.00294798
R35171 DVSS.n6062 DVSS.n6061 0.00294798
R35172 DVSS.n6829 DVSS.n6828 0.00294798
R35173 DVSS.n3638 DVSS.n3637 0.00294798
R35174 DVSS.n5314 DVSS.n5313 0.00294798
R35175 DVSS DVSS.n10726 0.00292857
R35176 DVSS.n14461 DVSS.n14460 0.00290105
R35177 DVSS.n14661 DVSS.n14660 0.00290105
R35178 DVSS.n16697 DVSS.n16696 0.00290061
R35179 DVSS.n18142 DVSS.n18141 0.00290061
R35180 DVSS.n14513 DVSS.n14512 0.00290061
R35181 DVSS.n19803 DVSS.n19802 0.00290061
R35182 DVSS.n244 DVSS.n243 0.00290061
R35183 DVSS.n18141 DVSS.n18140 0.00290061
R35184 DVSS.n18126 DVSS.n18125 0.00290061
R35185 DVSS.n16696 DVSS.n16695 0.00290061
R35186 DVSS.n17127 DVSS.n17126 0.00290061
R35187 DVSS.n15447 DVSS.n15446 0.00290061
R35188 DVSS.n14610 DVSS.n14609 0.00290061
R35189 DVSS.n20028 DVSS.n20027 0.00290061
R35190 DVSS.n452 DVSS.n451 0.00290061
R35191 DVSS.n15416 DVSS.n15415 0.00290061
R35192 DVSS.n15446 DVSS.n15445 0.00290061
R35193 DVSS.n17126 DVSS.n17125 0.00290061
R35194 DVSS.n14514 DVSS.n14513 0.00290061
R35195 DVSS.n14611 DVSS.n14610 0.00290061
R35196 DVSS.n19804 DVSS.n19803 0.00290061
R35197 DVSS.n20029 DVSS.n20028 0.00290061
R35198 DVSS.n245 DVSS.n244 0.00290061
R35199 DVSS.n453 DVSS.n452 0.00290061
R35200 DVSS.n17619 DVSS.n17618 0.00286739
R35201 DVSS.n17610 DVSS.n17609 0.00286739
R35202 DVSS.n11133 DVSS.n11132 0.00286739
R35203 DVSS.n11142 DVSS.n11141 0.00286739
R35204 DVSS.n16373 DVSS.n16372 0.00286739
R35205 DVSS.n16364 DVSS.n16363 0.00286739
R35206 DVSS.n4569 DVSS.n4568 0.00286111
R35207 DVSS.n4573 DVSS.n4572 0.00286111
R35208 DVSS.n4515 DVSS.n4514 0.00286111
R35209 DVSS.n4519 DVSS.n4518 0.00286111
R35210 DVSS.n4619 DVSS.n4618 0.00286111
R35211 DVSS.n4623 DVSS.n4622 0.00286111
R35212 DVSS.n5638 DVSS.n5637 0.00285947
R35213 DVSS.n5705 DVSS.n5704 0.00285947
R35214 DVSS.n5723 DVSS.n5722 0.00285947
R35215 DVSS.n4469 DVSS.n4468 0.00285947
R35216 DVSS.n4080 DVSS.n4079 0.00285947
R35217 DVSS.n6972 DVSS.n6971 0.00285947
R35218 DVSS.n7143 DVSS.n7142 0.00285947
R35219 DVSS.n7173 DVSS.n7172 0.00285947
R35220 DVSS.n865 DVSS.n864 0.00285947
R35221 DVSS.n5706 DVSS.n5705 0.00285947
R35222 DVSS.n4468 DVSS.n4467 0.00285947
R35223 DVSS.n10931 DVSS.n10930 0.00285947
R35224 DVSS.n10996 DVSS.n10995 0.00285947
R35225 DVSS.n11274 DVSS.n11273 0.00285947
R35226 DVSS.n11230 DVSS.n11229 0.00285947
R35227 DVSS.n11226 DVSS.n11225 0.00285947
R35228 DVSS.n9491 DVSS.n9490 0.00285947
R35229 DVSS.n9000 DVSS.n8999 0.00285947
R35230 DVSS.n12951 DVSS.n12950 0.00285947
R35231 DVSS.n12918 DVSS.n12917 0.00285947
R35232 DVSS.n12708 DVSS.n12707 0.00285947
R35233 DVSS.n12388 DVSS.n12387 0.00285947
R35234 DVSS.n12950 DVSS.n12949 0.00285947
R35235 DVSS.n9001 DVSS.n9000 0.00285947
R35236 DVSS.n9490 DVSS.n9489 0.00285947
R35237 DVSS.n10930 DVSS.n10929 0.00285947
R35238 DVSS.n10995 DVSS.n10994 0.00285947
R35239 DVSS.n5769 DVSS.n5768 0.00285947
R35240 DVSS.n11231 DVSS.n11230 0.00285947
R35241 DVSS.n11273 DVSS.n11272 0.00285947
R35242 DVSS.n11227 DVSS.n11226 0.00285947
R35243 DVSS.n5724 DVSS.n5723 0.00285947
R35244 DVSS.n17064 DVSS.n17063 0.00285947
R35245 DVSS.n16911 DVSS.n16910 0.00285947
R35246 DVSS.n17591 DVSS.n17590 0.00285947
R35247 DVSS.n17635 DVSS.n17634 0.00285947
R35248 DVSS.n17639 DVSS.n17638 0.00285947
R35249 DVSS.n15706 DVSS.n15705 0.00285947
R35250 DVSS.n14995 DVSS.n14994 0.00285947
R35251 DVSS.n13668 DVSS.n13667 0.00285947
R35252 DVSS.n13550 DVSS.n13549 0.00285947
R35253 DVSS.n13534 DVSS.n13533 0.00285947
R35254 DVSS.n20850 DVSS.n20849 0.00285947
R35255 DVSS.n15707 DVSS.n15706 0.00285947
R35256 DVSS.n14994 DVSS.n14993 0.00285947
R35257 DVSS.n17634 DVSS.n17633 0.00285947
R35258 DVSS.n17063 DVSS.n17062 0.00285947
R35259 DVSS.n16912 DVSS.n16911 0.00285947
R35260 DVSS.n17592 DVSS.n17591 0.00285947
R35261 DVSS.n17638 DVSS.n17637 0.00285947
R35262 DVSS.n13667 DVSS.n13666 0.00285947
R35263 DVSS.n7172 DVSS.n7171 0.00285947
R35264 DVSS.n13535 DVSS.n13534 0.00285947
R35265 DVSS.n10831 DVSS.n10830 0.00285947
R35266 DVSS.n11389 DVSS.n11388 0.00285947
R35267 DVSS.n11437 DVSS.n11436 0.00285947
R35268 DVSS.n11529 DVSS.n11528 0.00285947
R35269 DVSS.n11692 DVSS.n11691 0.00285947
R35270 DVSS.n13041 DVSS.n13040 0.00285947
R35271 DVSS.n12054 DVSS.n12053 0.00285947
R35272 DVSS.n66 DVSS.n65 0.00285947
R35273 DVSS.n21479 DVSS.n21478 0.00285947
R35274 DVSS.n13042 DVSS.n13041 0.00285947
R35275 DVSS.n11691 DVSS.n11690 0.00285947
R35276 DVSS.n11528 DVSS.n11527 0.00285947
R35277 DVSS.n11436 DVSS.n11435 0.00285947
R35278 DVSS.n10832 DVSS.n10831 0.00285947
R35279 DVSS.n11388 DVSS.n11387 0.00285947
R35280 DVSS.n4708 DVSS.n4707 0.00285947
R35281 DVSS.n4262 DVSS.n4261 0.00285947
R35282 DVSS.n3742 DVSS.n3741 0.00285947
R35283 DVSS.n3331 DVSS.n3330 0.00285947
R35284 DVSS.n3015 DVSS.n3014 0.00285947
R35285 DVSS.n3779 DVSS.n3778 0.00285947
R35286 DVSS.n3793 DVSS.n3792 0.00285947
R35287 DVSS.n4261 DVSS.n4260 0.00285947
R35288 DVSS.n9953 DVSS.n9952 0.00285947
R35289 DVSS.n9867 DVSS.n9866 0.00285947
R35290 DVSS.n11114 DVSS.n11113 0.00285947
R35291 DVSS.n11158 DVSS.n11157 0.00285947
R35292 DVSS.n11162 DVSS.n11161 0.00285947
R35293 DVSS.n9703 DVSS.n9702 0.00285947
R35294 DVSS.n9090 DVSS.n9089 0.00285947
R35295 DVSS.n13207 DVSS.n13206 0.00285947
R35296 DVSS.n13364 DVSS.n13363 0.00285947
R35297 DVSS.n13383 DVSS.n13382 0.00285947
R35298 DVSS.n21076 DVSS.n21075 0.00285947
R35299 DVSS.n13382 DVSS.n13381 0.00285947
R35300 DVSS.n9091 DVSS.n9090 0.00285947
R35301 DVSS.n9704 DVSS.n9703 0.00285947
R35302 DVSS.n11157 DVSS.n11156 0.00285947
R35303 DVSS.n9952 DVSS.n9951 0.00285947
R35304 DVSS.n9868 DVSS.n9867 0.00285947
R35305 DVSS.n11115 DVSS.n11114 0.00285947
R35306 DVSS.n11161 DVSS.n11160 0.00285947
R35307 DVSS.n13208 DVSS.n13207 0.00285947
R35308 DVSS.n17357 DVSS.n17356 0.00285947
R35309 DVSS.n17425 DVSS.n17424 0.00285947
R35310 DVSS.n16344 DVSS.n16343 0.00285947
R35311 DVSS.n16218 DVSS.n16217 0.00285947
R35312 DVSS.n7545 DVSS.n7544 0.00285947
R35313 DVSS.n18825 DVSS.n18824 0.00285947
R35314 DVSS.n18841 DVSS.n18840 0.00285947
R35315 DVSS.n1152 DVSS.n1151 0.00285947
R35316 DVSS.n16345 DVSS.n16344 0.00285947
R35317 DVSS.n18739 DVSS.n18738 0.00285947
R35318 DVSS.n18840 DVSS.n18839 0.00285947
R35319 DVSS.n16219 DVSS.n16218 0.00285947
R35320 DVSS.n17424 DVSS.n17423 0.00285947
R35321 DVSS.n16390 DVSS.n16389 0.00285947
R35322 DVSS.n5433 DVSS.n5432 0.00285947
R35323 DVSS.n6463 DVSS.n6462 0.00285947
R35324 DVSS.n6576 DVSS.n6575 0.00285947
R35325 DVSS.n3649 DVSS.n3648 0.00285947
R35326 DVSS.n18965 DVSS.n18964 0.00285947
R35327 DVSS.n543 DVSS.n542 0.00285947
R35328 DVSS.n6073 DVSS.n6072 0.00285947
R35329 DVSS.n6774 DVSS.n6773 0.00285947
R35330 DVSS.n3582 DVSS.n3581 0.00285947
R35331 DVSS.n6575 DVSS.n6574 0.00285947
R35332 DVSS.n6462 DVSS.n6461 0.00285947
R35333 DVSS.n12053 DVSS.n12052 0.00285947
R35334 DVSS.n12919 DVSS.n12918 0.00285947
R35335 DVSS.n13363 DVSS.n13362 0.00285947
R35336 DVSS.n13551 DVSS.n13550 0.00285947
R35337 DVSS.n18824 DVSS.n18823 0.00285947
R35338 DVSS.n7142 DVSS.n7141 0.00285947
R35339 DVSS.n3743 DVSS.n3742 0.00285947
R35340 DVSS.n3648 DVSS.n3647 0.00285947
R35341 DVSS.n12707 DVSS.n12706 0.00285947
R35342 DVSS.n3330 DVSS.n3329 0.00285947
R35343 DVSS.n65 DVSS.n64 0.00285947
R35344 DVSS.n18964 DVSS.n18963 0.00285947
R35345 DVSS.n21480 DVSS.n21479 0.00285947
R35346 DVSS.n12389 DVSS.n12388 0.00285947
R35347 DVSS.n21075 DVSS.n21074 0.00285947
R35348 DVSS.n20849 DVSS.n20848 0.00285947
R35349 DVSS.n1151 DVSS.n1150 0.00285947
R35350 DVSS.n864 DVSS.n863 0.00285947
R35351 DVSS.n542 DVSS.n541 0.00285947
R35352 DVSS.n17790 DVSS.n17789 0.0028295
R35353 DVSS.n17672 DVSS.n17671 0.0028295
R35354 DVSS.n15891 DVSS.n15890 0.0028295
R35355 DVSS.n17664 DVSS.n7655 0.0028295
R35356 DVSS.n12201 DVSS.n12200 0.00282847
R35357 DVSS.n16558 DVSS.n16557 0.00282394
R35358 DVSS.n16578 DVSS.n16577 0.00282394
R35359 DVSS.n16501 DVSS.n16500 0.00282394
R35360 DVSS.n16118 DVSS.n16117 0.00282394
R35361 DVSS.n17804 DVSS.n17803 0.00282394
R35362 DVSS.n17807 DVSS.n17806 0.00282394
R35363 DVSS.n17948 DVSS.n17947 0.00282394
R35364 DVSS.n18089 DVSS.n18088 0.00282394
R35365 DVSS.n18124 DVSS.n18123 0.00282394
R35366 DVSS.n18145 DVSS.n18144 0.00282394
R35367 DVSS.n18194 DVSS.n18193 0.00282394
R35368 DVSS.n7605 DVSS.n7604 0.00282394
R35369 DVSS.n18420 DVSS.n18419 0.00282394
R35370 DVSS.n18441 DVSS.n18440 0.00282394
R35371 DVSS.n18451 DVSS.n18450 0.00282394
R35372 DVSS.n18463 DVSS.n18462 0.00282394
R35373 DVSS.n18528 DVSS.n18527 0.00282394
R35374 DVSS.n14379 DVSS.n14378 0.00282394
R35375 DVSS.n19654 DVSS.n19653 0.00282394
R35376 DVSS.n16745 DVSS.n16744 0.00282394
R35377 DVSS.n16765 DVSS.n16764 0.00282394
R35378 DVSS.n16847 DVSS.n16846 0.00282394
R35379 DVSS.n15999 DVSS.n15998 0.00282394
R35380 DVSS.n15783 DVSS.n15782 0.00282394
R35381 DVSS.n15786 DVSS.n15785 0.00282394
R35382 DVSS.n15776 DVSS.n15775 0.00282394
R35383 DVSS.n15373 DVSS.n15372 0.00282394
R35384 DVSS.n15414 DVSS.n15413 0.00282394
R35385 DVSS.n15450 DVSS.n15449 0.00282394
R35386 DVSS.n15546 DVSS.n15545 0.00282394
R35387 DVSS.n15368 DVSS.n15367 0.00282394
R35388 DVSS.n15218 DVSS.n15217 0.00282394
R35389 DVSS.n15176 DVSS.n15175 0.00282394
R35390 DVSS.n15166 DVSS.n15165 0.00282394
R35391 DVSS.n15139 DVSS.n15138 0.00282394
R35392 DVSS.n13857 DVSS.n13856 0.00282394
R35393 DVSS.n14771 DVSS.n14770 0.00282394
R35394 DVSS.n19863 DVSS.n19862 0.00282394
R35395 DVSS.n10060 DVSS.n10059 0.0028235
R35396 DVSS.n2050 DVSS.n2049 0.00282169
R35397 DVSS.n1724 DVSS.n1723 0.00282169
R35398 DVSS.n6266 DVSS.n6265 0.00281429
R35399 DVSS.n1388 DVSS.n1387 0.00281
R35400 DVSS.n4146 DVSS.n4145 0.00281
R35401 DVSS.n4215 DVSS.n4214 0.00281
R35402 DVSS.n4169 DVSS.n4168 0.00281
R35403 DVSS.n9177 DVSS.n9176 0.00281
R35404 DVSS.n9217 DVSS.n9216 0.00281
R35405 DVSS.n9269 DVSS.n9268 0.00281
R35406 DVSS.n9322 DVSS.n9321 0.00281
R35407 DVSS.n9451 DVSS.n9450 0.00281
R35408 DVSS.n9442 DVSS.n9441 0.00281
R35409 DVSS.n21382 DVSS.n21381 0.00281
R35410 DVSS.n5732 DVSS.n5731 0.00280842
R35411 DVSS.n6518 DVSS.n6517 0.00280842
R35412 DVSS.n9144 DVSS.n9143 0.00280842
R35413 DVSS.n9584 DVSS.n9583 0.00280842
R35414 DVSS.n9756 DVSS.n9755 0.00280842
R35415 DVSS.n9776 DVSS.n9775 0.00280842
R35416 DVSS.n15716 DVSS.n15715 0.00280842
R35417 DVSS.n15859 DVSS.n15858 0.00280842
R35418 DVSS.n14986 DVSS.n14985 0.00280842
R35419 DVSS.n15613 DVSS.n15612 0.00280842
R35420 DVSS.n7133 DVSS.n7132 0.00280842
R35421 DVSS.n11429 DVSS.n11428 0.00280842
R35422 DVSS.n10756 DVSS.n10755 0.00280842
R35423 DVSS.n13145 DVSS.n13144 0.00280842
R35424 DVSS.n4038 DVSS.n4037 0.00280842
R35425 DVSS.n15040 DVSS.n15039 0.00280842
R35426 DVSS.n3997 DVSS.n3996 0.00280842
R35427 DVSS.n4122 DVSS.n4121 0.00280842
R35428 DVSS.n4348 DVSS.n4347 0.00280842
R35429 DVSS.n9802 DVSS.n9801 0.00280842
R35430 DVSS.n9713 DVSS.n9712 0.00280842
R35431 DVSS.n9610 DVSS.n9609 0.00280842
R35432 DVSS.n9101 DVSS.n9100 0.00280842
R35433 DVSS.n9045 DVSS.n9044 0.00280842
R35434 DVSS.n13354 DVSS.n13353 0.00280842
R35435 DVSS.n16291 DVSS.n16290 0.00280842
R35436 DVSS.n16252 DVSS.n16251 0.00280842
R35437 DVSS.n16131 DVSS.n16130 0.00280842
R35438 DVSS.n18385 DVSS.n18384 0.00280842
R35439 DVSS.n7503 DVSS.n7502 0.00280842
R35440 DVSS.n6440 DVSS.n6439 0.00280842
R35441 DVSS.n6351 DVSS.n6350 0.00280842
R35442 DVSS.n6662 DVSS.n6661 0.00280842
R35443 DVSS.n6723 DVSS.n6722 0.00280842
R35444 DVSS.n6844 DVSS.n6843 0.00280842
R35445 DVSS.n11024 DVSS.n11023 0.00280483
R35446 DVSS.n11195 DVSS.n11193 0.00280483
R35447 DVSS.n10035 DVSS.n10033 0.00280483
R35448 DVSS.n5566 DVSS.n5565 0.00280315
R35449 DVSS.n7153 DVSS.n7152 0.00280315
R35450 DVSS.n7177 DVSS.n7176 0.00280315
R35451 DVSS.n19245 DVSS.n19244 0.00280315
R35452 DVSS.n10207 DVSS.n10206 0.00280315
R35453 DVSS.n12732 DVSS.n12731 0.00280315
R35454 DVSS.n12723 DVSS.n12722 0.00280315
R35455 DVSS.n12722 DVSS.n12721 0.00280315
R35456 DVSS.n12486 DVSS.n12485 0.00280315
R35457 DVSS.n12455 DVSS.n12454 0.00280315
R35458 DVSS.n12454 DVSS.n12453 0.00280315
R35459 DVSS.n12397 DVSS.n12396 0.00280315
R35460 DVSS.n12203 DVSS.n12202 0.00280315
R35461 DVSS.n12199 DVSS.n12198 0.00280315
R35462 DVSS.n12179 DVSS.n12178 0.00280315
R35463 DVSS.n12178 DVSS.n12177 0.00280315
R35464 DVSS.n21248 DVSS.n21247 0.00280315
R35465 DVSS.n21292 DVSS.n21291 0.00280315
R35466 DVSS.n21212 DVSS.n21211 0.00280315
R35467 DVSS.n21221 DVSS.n21212 0.00280315
R35468 DVSS.n16952 DVSS.n16951 0.00280315
R35469 DVSS.n13540 DVSS.n13539 0.00280315
R35470 DVSS.n13530 DVSS.n13529 0.00280315
R35471 DVSS.n11407 DVSS.n11406 0.00280315
R35472 DVSS.n5219 DVSS.n5218 0.00280315
R35473 DVSS.n3354 DVSS.n3353 0.00280315
R35474 DVSS.n3346 DVSS.n3345 0.00280315
R35475 DVSS.n3345 DVSS.n3344 0.00280315
R35476 DVSS.n3111 DVSS.n3110 0.00280315
R35477 DVSS.n3081 DVSS.n3080 0.00280315
R35478 DVSS.n3080 DVSS.n3079 0.00280315
R35479 DVSS.n3023 DVSS.n3022 0.00280315
R35480 DVSS.n2833 DVSS.n2832 0.00280315
R35481 DVSS.n2828 DVSS.n2827 0.00280315
R35482 DVSS.n2807 DVSS.n2806 0.00280315
R35483 DVSS.n2806 DVSS.n2805 0.00280315
R35484 DVSS.n746 DVSS.n745 0.00280315
R35485 DVSS.n742 DVSS.n741 0.00280315
R35486 DVSS.n749 DVSS.n748 0.00280315
R35487 DVSS.n750 DVSS.n749 0.00280315
R35488 DVSS.n9908 DVSS.n9907 0.00280315
R35489 DVSS.n13374 DVSS.n13373 0.00280315
R35490 DVSS.n13387 DVSS.n13386 0.00280315
R35491 DVSS.n17261 DVSS.n17260 0.00280315
R35492 DVSS.n18835 DVSS.n18834 0.00280315
R35493 DVSS.n18845 DVSS.n18844 0.00280315
R35494 DVSS.n19516 DVSS.n19515 0.00280315
R35495 DVSS.n6330 DVSS.n6329 0.00280315
R35496 DVSS.n2350 DVSS.n2349 0.00279928
R35497 DVSS.n2388 DVSS.n2387 0.00279928
R35498 DVSS.n2349 DVSS.n2348 0.00279928
R35499 DVSS.n2387 DVSS.n2386 0.00279928
R35500 DVSS.n16647 DVSS.n16646 0.00279506
R35501 DVSS.n16119 DVSS.n16118 0.00279506
R35502 DVSS.n17749 DVSS.n17748 0.00279506
R35503 DVSS.n17803 DVSS.n17802 0.00279506
R35504 DVSS.n14378 DVSS.n14377 0.00279506
R35505 DVSS.n16120 DVSS.n16119 0.00279506
R35506 DVSS.n17802 DVSS.n17801 0.00279506
R35507 DVSS.n16646 DVSS.n16645 0.00279506
R35508 DVSS.n17748 DVSS.n17747 0.00279506
R35509 DVSS.n14377 DVSS.n14376 0.00279506
R35510 DVSS.n17176 DVSS.n17175 0.00279506
R35511 DVSS.n16000 DVSS.n15999 0.00279506
R35512 DVSS.n15914 DVSS.n15913 0.00279506
R35513 DVSS.n15782 DVSS.n15781 0.00279506
R35514 DVSS.n14772 DVSS.n14771 0.00279506
R35515 DVSS.n16001 DVSS.n16000 0.00279506
R35516 DVSS.n15781 DVSS.n15780 0.00279506
R35517 DVSS.n17177 DVSS.n17176 0.00279506
R35518 DVSS.n15915 DVSS.n15914 0.00279506
R35519 DVSS.n14773 DVSS.n14772 0.00279506
R35520 DVSS.n5564 DVSS.n5563 0.00277159
R35521 DVSS.n10205 DVSS.n10204 0.00277159
R35522 DVSS.n16950 DVSS.n16949 0.00277159
R35523 DVSS.n5217 DVSS.n5216 0.00277159
R35524 DVSS.n9906 DVSS.n9905 0.00277159
R35525 DVSS.n17259 DVSS.n17258 0.00277159
R35526 DVSS.n4442 DVSS.n4441 0.00277096
R35527 DVSS.n4394 DVSS.n4393 0.00277096
R35528 DVSS.n6958 DVSS.n6957 0.00277096
R35529 DVSS.n19119 DVSS.n19118 0.00277096
R35530 DVSS.n19200 DVSS.n19199 0.00277096
R35531 DVSS.n19286 DVSS.n19285 0.00277096
R35532 DVSS.n1041 DVSS.n1040 0.00277096
R35533 DVSS.n992 DVSS.n991 0.00277096
R35534 DVSS.n9518 DVSS.n9517 0.00277096
R35535 DVSS.n9571 DVSS.n9570 0.00277096
R35536 DVSS.n12947 DVSS.n12946 0.00277096
R35537 DVSS.n12890 DVSS.n12889 0.00277096
R35538 DVSS.n12838 DVSS.n12837 0.00277096
R35539 DVSS.n12407 DVSS.n12406 0.00277096
R35540 DVSS.n9570 DVSS.n9569 0.00277096
R35541 DVSS.n9519 DVSS.n9518 0.00277096
R35542 DVSS.n15679 DVSS.n15678 0.00277096
R35543 DVSS.n15626 DVSS.n15625 0.00277096
R35544 DVSS.n13845 DVSS.n13844 0.00277096
R35545 DVSS.n20119 DVSS.n20118 0.00277096
R35546 DVSS.n20211 DVSS.n20210 0.00277096
R35547 DVSS.n20300 DVSS.n20299 0.00277096
R35548 DVSS.n20842 DVSS.n20841 0.00277096
R35549 DVSS.n20806 DVSS.n20805 0.00277096
R35550 DVSS.n20754 DVSS.n20753 0.00277096
R35551 DVSS.n15678 DVSS.n15677 0.00277096
R35552 DVSS.n15627 DVSS.n15626 0.00277096
R35553 DVSS.n13846 DVSS.n13845 0.00277096
R35554 DVSS.n12946 DVSS.n12945 0.00277096
R35555 DVSS.n10814 DVSS.n10813 0.00277096
R35556 DVSS.n11556 DVSS.n11555 0.00277096
R35557 DVSS.n11609 DVSS.n11608 0.00277096
R35558 DVSS.n13046 DVSS.n13045 0.00277096
R35559 DVSS.n12075 DVSS.n12074 0.00277096
R35560 DVSS.n58 DVSS.n57 0.00277096
R35561 DVSS.n21539 DVSS.n21538 0.00277096
R35562 DVSS.n21487 DVSS.n21486 0.00277096
R35563 DVSS.n21451 DVSS.n21450 0.00277096
R35564 DVSS.n21399 DVSS.n21398 0.00277096
R35565 DVSS.n11608 DVSS.n11607 0.00277096
R35566 DVSS.n11557 DVSS.n11556 0.00277096
R35567 DVSS.n10815 DVSS.n10814 0.00277096
R35568 DVSS.n3782 DVSS.n3781 0.00277096
R35569 DVSS.n3499 DVSS.n3498 0.00277096
R35570 DVSS.n3450 DVSS.n3449 0.00277096
R35571 DVSS.n3033 DVSS.n3032 0.00277096
R35572 DVSS.n4336 DVSS.n4335 0.00277096
R35573 DVSS.n4288 DVSS.n4287 0.00277096
R35574 DVSS.n9676 DVSS.n9675 0.00277096
R35575 DVSS.n9623 DVSS.n9622 0.00277096
R35576 DVSS.n13187 DVSS.n13186 0.00277096
R35577 DVSS.n20402 DVSS.n20401 0.00277096
R35578 DVSS.n20482 DVSS.n20481 0.00277096
R35579 DVSS.n20574 DVSS.n20573 0.00277096
R35580 DVSS.n21068 DVSS.n21067 0.00277096
R35581 DVSS.n21032 DVSS.n21031 0.00277096
R35582 DVSS.n20980 DVSS.n20979 0.00277096
R35583 DVSS.n9675 DVSS.n9674 0.00277096
R35584 DVSS.n9624 DVSS.n9623 0.00277096
R35585 DVSS.n13186 DVSS.n13185 0.00277096
R35586 DVSS.n18579 DVSS.n18578 0.00277096
R35587 DVSS.n19393 DVSS.n19392 0.00277096
R35588 DVSS.n19471 DVSS.n19470 0.00277096
R35589 DVSS.n19557 DVSS.n19556 0.00277096
R35590 DVSS.n1256 DVSS.n1255 0.00277096
R35591 DVSS.n1208 DVSS.n1207 0.00277096
R35592 DVSS.n16192 DVSS.n16191 0.00277096
R35593 DVSS.n16143 DVSS.n16142 0.00277096
R35594 DVSS.n18578 DVSS.n18577 0.00277096
R35595 DVSS.n13045 DVSS.n13044 0.00277096
R35596 DVSS.n3783 DVSS.n3782 0.00277096
R35597 DVSS.n6957 DVSS.n6956 0.00277096
R35598 DVSS.n3579 DVSS.n3578 0.00277096
R35599 DVSS.n3561 DVSS.n3560 0.00277096
R35600 DVSS.n19005 DVSS.n19004 0.00277096
R35601 DVSS.n607 DVSS.n606 0.00277096
R35602 DVSS.n6602 DVSS.n6601 0.00277096
R35603 DVSS.n6651 DVSS.n6650 0.00277096
R35604 DVSS.n3578 DVSS.n3577 0.00277096
R35605 DVSS.n18958 DVSS.n18957 0.00277096
R35606 DVSS.n20210 DVSS.n20209 0.00277096
R35607 DVSS.n20481 DVSS.n20480 0.00277096
R35608 DVSS.n12839 DVSS.n12838 0.00277096
R35609 DVSS.n57 DVSS.n56 0.00277096
R35610 DVSS.n12076 DVSS.n12075 0.00277096
R35611 DVSS.n12891 DVSS.n12890 0.00277096
R35612 DVSS.n20401 DVSS.n20400 0.00277096
R35613 DVSS.n20118 DVSS.n20117 0.00277096
R35614 DVSS.n19470 DVSS.n19469 0.00277096
R35615 DVSS.n19199 DVSS.n19198 0.00277096
R35616 DVSS.n3451 DVSS.n3450 0.00277096
R35617 DVSS.n536 DVSS.n535 0.00277096
R35618 DVSS.n3034 DVSS.n3033 0.00277096
R35619 DVSS.n1145 DVSS.n1144 0.00277096
R35620 DVSS.n21488 DVSS.n21487 0.00277096
R35621 DVSS.n858 DVSS.n857 0.00277096
R35622 DVSS.n21540 DVSS.n21539 0.00277096
R35623 DVSS.n20575 DVSS.n20574 0.00277096
R35624 DVSS.n20301 DVSS.n20300 0.00277096
R35625 DVSS.n21067 DVSS.n21066 0.00277096
R35626 DVSS.n20841 DVSS.n20840 0.00277096
R35627 DVSS.n559 DVSS.n558 0.00277096
R35628 DVSS.n21452 DVSS.n21451 0.00277096
R35629 DVSS.n21033 DVSS.n21032 0.00277096
R35630 DVSS.n20807 DVSS.n20806 0.00277096
R35631 DVSS.n21400 DVSS.n21399 0.00277096
R35632 DVSS.n20755 DVSS.n20754 0.00277096
R35633 DVSS.n20981 DVSS.n20980 0.00277096
R35634 DVSS.n993 DVSS.n992 0.00277096
R35635 DVSS.n17457 DVSS.n17456 0.00275919
R35636 DVSS.n14257 DVSS.n14256 0.00275919
R35637 DVSS.n14282 DVSS.n14281 0.00275919
R35638 DVSS.n14311 DVSS.n14310 0.00275919
R35639 DVSS.n14397 DVSS.n14396 0.00275919
R35640 DVSS.n17538 DVSS.n17537 0.00275919
R35641 DVSS.n15882 DVSS.n15881 0.00275919
R35642 DVSS.n14692 DVSS.n14691 0.00275919
R35643 DVSS.n14753 DVSS.n14752 0.00275919
R35644 DVSS.n14858 DVSS.n14857 0.00275919
R35645 DVSS.n14841 DVSS.n14840 0.00275919
R35646 DVSS.n14824 DVSS.n14823 0.00275919
R35647 DVSS.n7718 DVSS.n7717 0.00275
R35648 DVSS.n15067 DVSS.n15066 0.00275
R35649 DVSS.n16049 DVSS.n16048 0.00275
R35650 DVSS.n17528 DVSS.n17527 0.00275
R35651 DVSS.n15264 DVSS.n15263 0.00275
R35652 DVSS.n18355 DVSS.n18354 0.00275
R35653 DVSS.n18076 DVSS.n18075 0.00275
R35654 DVSS.n17935 DVSS.n17934 0.00275
R35655 DVSS.n13972 DVSS.n13971 0.00275
R35656 DVSS DVSS.n21573 0.00275
R35657 DVSS.n6517 DVSS.n6516 0.00274945
R35658 DVSS.n4039 DVSS.n4038 0.00274945
R35659 DVSS.n7132 DVSS.n7131 0.00274945
R35660 DVSS.n6530 DVSS.n6529 0.00274945
R35661 DVSS.n4383 DVSS.n4382 0.00274945
R35662 DVSS.n4089 DVSS.n4088 0.00274945
R35663 DVSS.n5813 DVSS.n5812 0.00274945
R35664 DVSS.n11236 DVSS.n11235 0.00274945
R35665 DVSS.n9775 DVSS.n9774 0.00274945
R35666 DVSS.n9757 DVSS.n9756 0.00274945
R35667 DVSS.n9583 DVSS.n9582 0.00274945
R35668 DVSS.n9145 DVSS.n9144 0.00274945
R35669 DVSS.n13144 DVSS.n13143 0.00274945
R35670 DVSS.n11046 DVSS.n11045 0.00274945
R35671 DVSS.n17629 DVSS.n17628 0.00274945
R35672 DVSS.n15860 DVSS.n15859 0.00274945
R35673 DVSS.n15715 DVSS.n15714 0.00274945
R35674 DVSS.n15614 DVSS.n15613 0.00274945
R35675 DVSS.n14985 DVSS.n14984 0.00274945
R35676 DVSS.n15039 DVSS.n15038 0.00274945
R35677 DVSS.n16903 DVSS.n15872 0.00274945
R35678 DVSS.n10968 DVSS.n10967 0.00274945
R35679 DVSS.n17101 DVSS.n17100 0.00274945
R35680 DVSS.n5677 DVSS.n5676 0.00274945
R35681 DVSS.n4347 DVSS.n4346 0.00274945
R35682 DVSS.n4123 DVSS.n4122 0.00274945
R35683 DVSS.n3996 DVSS.n3995 0.00274945
R35684 DVSS.n11152 DVSS.n11151 0.00274945
R35685 DVSS.n9803 DVSS.n9802 0.00274945
R35686 DVSS.n9712 DVSS.n9711 0.00274945
R35687 DVSS.n9611 DVSS.n9610 0.00274945
R35688 DVSS.n9100 DVSS.n9099 0.00274945
R35689 DVSS.n9046 DVSS.n9045 0.00274945
R35690 DVSS.n13353 DVSS.n13352 0.00274945
R35691 DVSS.n11068 DVSS.n11067 0.00274945
R35692 DVSS.n9990 DVSS.n9989 0.00274945
R35693 DVSS.n17447 DVSS.n17446 0.00274945
R35694 DVSS.n16354 DVSS.n16353 0.00274945
R35695 DVSS.n16292 DVSS.n16291 0.00274945
R35696 DVSS.n16253 DVSS.n16252 0.00274945
R35697 DVSS.n16132 DVSS.n16131 0.00274945
R35698 DVSS.n18384 DVSS.n18383 0.00274945
R35699 DVSS.n7504 DVSS.n7503 0.00274945
R35700 DVSS.n18621 DVSS.n18620 0.00274945
R35701 DVSS.n18648 DVSS.n18647 0.00274945
R35702 DVSS.n18680 DVSS.n18679 0.00274945
R35703 DVSS.n17396 DVSS.n17395 0.00274945
R35704 DVSS.n5837 DVSS.n5836 0.00274945
R35705 DVSS.n6471 DVSS.n6470 0.00274945
R35706 DVSS.n6756 DVSS.n6755 0.00273544
R35707 DVSS.n6701 DVSS.n6700 0.00273544
R35708 DVSS.n2533 DVSS.n2532 0.00273544
R35709 DVSS.n6394 DVSS.n6393 0.00273544
R35710 DVSS.n6883 DVSS.n6882 0.00273544
R35711 DVSS.n4521 DVSS.n4520 0.00273544
R35712 DVSS.n6882 DVSS.n6881 0.00273544
R35713 DVSS.n6755 DVSS.n6754 0.00273544
R35714 DVSS.n6700 DVSS.n6699 0.00273544
R35715 DVSS.n2532 DVSS.n2531 0.00273544
R35716 DVSS.n6393 DVSS.n6392 0.00273544
R35717 DVSS.n4567 DVSS.n4566 0.00271192
R35718 DVSS.n6753 DVSS.n6752 0.00271192
R35719 DVSS.n6698 DVSS.n6697 0.00271192
R35720 DVSS.n2530 DVSS.n2529 0.00271192
R35721 DVSS.n4513 DVSS.n4512 0.00271192
R35722 DVSS.n6391 DVSS.n6390 0.00271192
R35723 DVSS.n6880 DVSS.n6879 0.00271192
R35724 DVSS.n4617 DVSS.n4616 0.00271192
R35725 DVSS.n8912 DVSS 0.0027
R35726 DVSS.n14424 DVSS.n14423 0.00268951
R35727 DVSS.n14425 DVSS.n14424 0.00268951
R35728 DVSS.n16064 DVSS.n16063 0.00268951
R35729 DVSS.n14392 DVSS.n14391 0.00268951
R35730 DVSS.n16065 DVSS.n16064 0.00268951
R35731 DVSS.n16541 DVSS.n16540 0.00268951
R35732 DVSS.n14391 DVSS.n14390 0.00268951
R35733 DVSS.n15956 DVSS.n15955 0.00268951
R35734 DVSS.n14758 DVSS.n14757 0.00268951
R35735 DVSS.n14703 DVSS.n14702 0.00268951
R35736 DVSS.n15957 DVSS.n15956 0.00268951
R35737 DVSS.n14704 DVSS.n14703 0.00268951
R35738 DVSS.n16728 DVSS.n16727 0.00268951
R35739 DVSS.n14759 DVSS.n14758 0.00268951
R35740 DVSS.n14256 DVSS.n14255 0.00268887
R35741 DVSS.n14281 DVSS.n14280 0.00268887
R35742 DVSS.n14310 DVSS.n14309 0.00268887
R35743 DVSS.n14859 DVSS.n14858 0.00268887
R35744 DVSS.n14842 DVSS.n14841 0.00268887
R35745 DVSS.n14825 DVSS.n14824 0.00268887
R35746 DVSS.n6267 DVSS.n6266 0.00268571
R35747 DVSS.n10955 DVSS.n10954 0.00268307
R35748 DVSS.n17088 DVSS.n17087 0.00268307
R35749 DVSS.n9977 DVSS.n9976 0.00268307
R35750 DVSS.n5693 DVSS.n5692 0.00268244
R35751 DVSS.n4420 DVSS.n4419 0.00268244
R35752 DVSS.n4415 DVSS.n4414 0.00268244
R35753 DVSS.n19178 DVSS.n19177 0.00268244
R35754 DVSS.n19259 DVSS.n19258 0.00268244
R35755 DVSS.n1014 DVSS.n1013 0.00268244
R35756 DVSS.n4421 DVSS.n4420 0.00268244
R35757 DVSS.n5692 DVSS.n5691 0.00268244
R35758 DVSS.n10983 DVSS.n10982 0.00268244
R35759 DVSS.n10986 DVSS.n10985 0.00268244
R35760 DVSS.n9541 DVSS.n9540 0.00268244
R35761 DVSS.n9549 DVSS.n9548 0.00268244
R35762 DVSS.n12868 DVSS.n12867 0.00268244
R35763 DVSS.n12861 DVSS.n12860 0.00268244
R35764 DVSS.n12489 DVSS.n12488 0.00268244
R35765 DVSS.n9540 DVSS.n9539 0.00268244
R35766 DVSS.n9548 DVSS.n9547 0.00268244
R35767 DVSS.n10987 DVSS.n10986 0.00268244
R35768 DVSS.n10982 DVSS.n10981 0.00268244
R35769 DVSS.n16924 DVSS.n16923 0.00268244
R35770 DVSS.n16921 DVSS.n16920 0.00268244
R35771 DVSS.n15656 DVSS.n15655 0.00268244
R35772 DVSS.n15648 DVSS.n15647 0.00268244
R35773 DVSS.n20181 DVSS.n20180 0.00268244
R35774 DVSS.n20188 DVSS.n20187 0.00268244
R35775 DVSS.n20278 DVSS.n20277 0.00268244
R35776 DVSS.n20270 DVSS.n20269 0.00268244
R35777 DVSS.n20784 DVSS.n20783 0.00268244
R35778 DVSS.n20776 DVSS.n20775 0.00268244
R35779 DVSS.n15657 DVSS.n15656 0.00268244
R35780 DVSS.n15649 DVSS.n15648 0.00268244
R35781 DVSS.n16920 DVSS.n16919 0.00268244
R35782 DVSS.n16925 DVSS.n16924 0.00268244
R35783 DVSS.n11579 DVSS.n11578 0.00268244
R35784 DVSS.n11587 DVSS.n11586 0.00268244
R35785 DVSS.n28 DVSS.n27 0.00268244
R35786 DVSS.n35 DVSS.n34 0.00268244
R35787 DVSS.n21517 DVSS.n21516 0.00268244
R35788 DVSS.n21509 DVSS.n21508 0.00268244
R35789 DVSS.n21429 DVSS.n21428 0.00268244
R35790 DVSS.n21421 DVSS.n21420 0.00268244
R35791 DVSS.n11578 DVSS.n11577 0.00268244
R35792 DVSS.n11586 DVSS.n11585 0.00268244
R35793 DVSS.n4656 DVSS.n4655 0.00268244
R35794 DVSS.n4657 DVSS.n4656 0.00268244
R35795 DVSS.n4315 DVSS.n4314 0.00268244
R35796 DVSS.n3477 DVSS.n3476 0.00268244
R35797 DVSS.n3472 DVSS.n3471 0.00268244
R35798 DVSS.n3114 DVSS.n3113 0.00268244
R35799 DVSS.n4309 DVSS.n4308 0.00268244
R35800 DVSS.n9880 DVSS.n9879 0.00268244
R35801 DVSS.n9877 DVSS.n9876 0.00268244
R35802 DVSS.n9653 DVSS.n9652 0.00268244
R35803 DVSS.n9645 DVSS.n9644 0.00268244
R35804 DVSS.n20452 DVSS.n20451 0.00268244
R35805 DVSS.n20459 DVSS.n20458 0.00268244
R35806 DVSS.n20552 DVSS.n20551 0.00268244
R35807 DVSS.n20544 DVSS.n20543 0.00268244
R35808 DVSS.n21010 DVSS.n21009 0.00268244
R35809 DVSS.n21002 DVSS.n21001 0.00268244
R35810 DVSS.n9654 DVSS.n9653 0.00268244
R35811 DVSS.n9646 DVSS.n9645 0.00268244
R35812 DVSS.n9876 DVSS.n9875 0.00268244
R35813 DVSS.n9881 DVSS.n9880 0.00268244
R35814 DVSS.n17412 DVSS.n17411 0.00268244
R35815 DVSS.n16164 DVSS.n16163 0.00268244
R35816 DVSS.n19530 DVSS.n19529 0.00268244
R35817 DVSS.n1229 DVSS.n1228 0.00268244
R35818 DVSS.n16171 DVSS.n16170 0.00268244
R35819 DVSS.n16165 DVSS.n16164 0.00268244
R35820 DVSS.n17411 DVSS.n17410 0.00268244
R35821 DVSS.n6630 DVSS.n6629 0.00268244
R35822 DVSS.n3539 DVSS.n3538 0.00268244
R35823 DVSS.n3534 DVSS.n3533 0.00268244
R35824 DVSS.n18978 DVSS.n18977 0.00268244
R35825 DVSS.n580 DVSS.n579 0.00268244
R35826 DVSS.n6623 DVSS.n6622 0.00268244
R35827 DVSS.n6629 DVSS.n6628 0.00268244
R35828 DVSS.n3540 DVSS.n3539 0.00268244
R35829 DVSS.n3478 DVSS.n3477 0.00268244
R35830 DVSS.n19172 DVSS.n19171 0.00268244
R35831 DVSS.n20460 DVSS.n20459 0.00268244
R35832 DVSS.n20451 DVSS.n20450 0.00268244
R35833 DVSS.n12869 DVSS.n12868 0.00268244
R35834 DVSS.n12860 DVSS.n12859 0.00268244
R35835 DVSS.n36 DVSS.n35 0.00268244
R35836 DVSS.n19449 DVSS.n19448 0.00268244
R35837 DVSS.n20189 DVSS.n20188 0.00268244
R35838 DVSS.n27 DVSS.n26 0.00268244
R35839 DVSS.n19443 DVSS.n19442 0.00268244
R35840 DVSS.n20180 DVSS.n20179 0.00268244
R35841 DVSS.n18984 DVSS.n18983 0.00268244
R35842 DVSS.n19536 DVSS.n19535 0.00268244
R35843 DVSS.n21518 DVSS.n21517 0.00268244
R35844 DVSS.n19265 DVSS.n19264 0.00268244
R35845 DVSS.n12490 DVSS.n12489 0.00268244
R35846 DVSS.n21510 DVSS.n21509 0.00268244
R35847 DVSS.n20545 DVSS.n20544 0.00268244
R35848 DVSS.n20271 DVSS.n20270 0.00268244
R35849 DVSS.n20553 DVSS.n20552 0.00268244
R35850 DVSS.n20279 DVSS.n20278 0.00268244
R35851 DVSS.n586 DVSS.n585 0.00268244
R35852 DVSS.n662 DVSS.n661 0.00268244
R35853 DVSS.n1235 DVSS.n1234 0.00268244
R35854 DVSS.n21285 DVSS.n21284 0.00268244
R35855 DVSS.n21430 DVSS.n21429 0.00268244
R35856 DVSS.n1020 DVSS.n1019 0.00268244
R35857 DVSS.n21422 DVSS.n21421 0.00268244
R35858 DVSS.n21304 DVSS.n21303 0.00268244
R35859 DVSS.n21003 DVSS.n21002 0.00268244
R35860 DVSS.n20777 DVSS.n20776 0.00268244
R35861 DVSS.n667 DVSS.n666 0.00268244
R35862 DVSS.n21011 DVSS.n21010 0.00268244
R35863 DVSS.n20785 DVSS.n20784 0.00268244
R35864 DVSS.n13297 DVSS.n13296 0.00267491
R35865 DVSS.n13296 DVSS.n13295 0.00267491
R35866 DVSS.n1395 DVSS.n1394 0.00263
R35867 DVSS.n4238 DVSS.n4237 0.00263
R35868 DVSS.n4207 DVSS.n4206 0.00263
R35869 DVSS.n4160 DVSS.n4159 0.00263
R35870 DVSS.n5772 DVSS.n5771 0.00262598
R35871 DVSS.n5741 DVSS.n5740 0.00262598
R35872 DVSS.n4046 DVSS.n4045 0.00262598
R35873 DVSS.n6986 DVSS.n6985 0.00262598
R35874 DVSS.n7111 DVSS.n7110 0.00262598
R35875 DVSS.n7148 DVSS.n7147 0.00262598
R35876 DVSS.n7198 DVSS.n7197 0.00262598
R35877 DVSS.n11277 DVSS.n11276 0.00262598
R35878 DVSS.n13137 DVSS.n13136 0.00262598
R35879 DVSS.n12921 DVSS.n12920 0.00262598
R35880 DVSS.n12835 DVSS.n12834 0.00262598
R35881 DVSS.n12774 DVSS.n12773 0.00262598
R35882 DVSS.n12756 DVSS.n12755 0.00262598
R35883 DVSS.n12751 DVSS.n12750 0.00262598
R35884 DVSS.n12495 DVSS.n12494 0.00262598
R35885 DVSS.n21245 DVSS.n21244 0.00262598
R35886 DVSS.n21208 DVSS.n21207 0.00262598
R35887 DVSS.n17588 DVSS.n17587 0.00262598
R35888 DVSS.n15032 DVSS.n15031 0.00262598
R35889 DVSS.n13652 DVSS.n13651 0.00262598
R35890 DVSS.n13570 DVSS.n13569 0.00262598
R35891 DVSS.n13545 DVSS.n13544 0.00262598
R35892 DVSS.n13522 DVSS.n13521 0.00262598
R35893 DVSS.n10774 DVSS.n10773 0.00262598
R35894 DVSS.n11385 DVSS.n11384 0.00262598
R35895 DVSS.n11452 DVSS.n11451 0.00262598
R35896 DVSS.n13064 DVSS.n13063 0.00262598
R35897 DVSS.n12051 DVSS.n12050 0.00262598
R35898 DVSS.n3989 DVSS.n3988 0.00262598
R35899 DVSS.n3745 DVSS.n3744 0.00262598
R35900 DVSS.n3447 DVSS.n3446 0.00262598
R35901 DVSS.n3386 DVSS.n3385 0.00262598
R35902 DVSS.n3369 DVSS.n3368 0.00262598
R35903 DVSS.n3364 DVSS.n3363 0.00262598
R35904 DVSS.n3119 DVSS.n3118 0.00262598
R35905 DVSS.n776 DVSS.n775 0.00262598
R35906 DVSS.n788 DVSS.n787 0.00262598
R35907 DVSS.n11111 DVSS.n11110 0.00262598
R35908 DVSS.n9053 DVSS.n9052 0.00262598
R35909 DVSS.n13223 DVSS.n13222 0.00262598
R35910 DVSS.n13262 DVSS.n13261 0.00262598
R35911 DVSS.n13369 DVSS.n13368 0.00262598
R35912 DVSS.n13402 DVSS.n13401 0.00262598
R35913 DVSS.n16393 DVSS.n16392 0.00262598
R35914 DVSS.n16362 DVSS.n16361 0.00262598
R35915 DVSS.n7511 DVSS.n7510 0.00262598
R35916 DVSS.n18753 DVSS.n18752 0.00262598
R35917 DVSS.n18790 DVSS.n18789 0.00262598
R35918 DVSS.n18830 DVSS.n18829 0.00262598
R35919 DVSS.n18858 DVSS.n18857 0.00262598
R35920 DVSS.n5500 DVSS.n5499 0.00262598
R35921 DVSS.n6070 DVSS.n6069 0.00262598
R35922 DVSS.n6447 DVSS.n6446 0.00262598
R35923 DVSS.n6837 DVSS.n6836 0.00262598
R35924 DVSS.n3646 DVSS.n3645 0.00262598
R35925 DVSS.n12539 DVSS.n12538 0.00261538
R35926 DVSS.n12663 DVSS.n12662 0.00261538
R35927 DVSS.n12571 DVSS.n12570 0.00261538
R35928 DVSS.n12375 DVSS.n12374 0.00261538
R35929 DVSS.n12283 DVSS.n12282 0.00261538
R35930 DVSS.n12258 DVSS.n12253 0.00261538
R35931 DVSS.n3163 DVSS.n3162 0.00261538
R35932 DVSS.n3287 DVSS.n3286 0.00261538
R35933 DVSS.n3195 DVSS.n3194 0.00261538
R35934 DVSS.n3002 DVSS.n3001 0.00261538
R35935 DVSS.n2910 DVSS.n2909 0.00261538
R35936 DVSS.n2885 DVSS.n2880 0.00261538
R35937 DVSS.n17478 DVSS.n17477 0.00261268
R35938 DVSS.n16070 DVSS.n16069 0.00261268
R35939 DVSS.n16069 DVSS.n16068 0.00261268
R35940 DVSS.n17885 DVSS.n17884 0.00261268
R35941 DVSS.n18026 DVSS.n18025 0.00261268
R35942 DVSS.n18107 DVSS.n18106 0.00261268
R35943 DVSS.n18111 DVSS.n18110 0.00261268
R35944 DVSS.n18127 DVSS.n18126 0.00261268
R35945 DVSS.n18263 DVSS.n18262 0.00261268
R35946 DVSS.n18243 DVSS.n18242 0.00261268
R35947 DVSS.n18181 DVSS.n18180 0.00261268
R35948 DVSS.n7577 DVSS.n7576 0.00261268
R35949 DVSS.n18471 DVSS.n18470 0.00261268
R35950 DVSS.n18511 DVSS.n18510 0.00261268
R35951 DVSS.n18556 DVSS.n18555 0.00261268
R35952 DVSS.n14387 DVSS.n14386 0.00261268
R35953 DVSS.n14401 DVSS.n14400 0.00261268
R35954 DVSS.n14465 DVSS.n14464 0.00261268
R35955 DVSS.n14515 DVSS.n14514 0.00261268
R35956 DVSS.n19670 DVSS.n19669 0.00261268
R35957 DVSS.n19805 DVSS.n19804 0.00261268
R35958 DVSS.n246 DVSS.n245 0.00261268
R35959 DVSS.n16819 DVSS.n16818 0.00261268
R35960 DVSS.n15962 DVSS.n15961 0.00261268
R35961 DVSS.n15961 DVSS.n15960 0.00261268
R35962 DVSS.n15814 DVSS.n15813 0.00261268
R35963 DVSS.n15748 DVSS.n15747 0.00261268
R35964 DVSS.n15385 DVSS.n15384 0.00261268
R35965 DVSS.n15389 DVSS.n15388 0.00261268
R35966 DVSS.n15417 DVSS.n15416 0.00261268
R35967 DVSS.n15477 DVSS.n15476 0.00261268
R35968 DVSS.n15497 DVSS.n15496 0.00261268
R35969 DVSS.n15559 DVSS.n15558 0.00261268
R35970 DVSS.n15232 DVSS.n15231 0.00261268
R35971 DVSS.n15131 DVSS.n15130 0.00261268
R35972 DVSS.n7752 DVSS.n7751 0.00261268
R35973 DVSS.n13920 DVSS.n13919 0.00261268
R35974 DVSS.n14763 DVSS.n14762 0.00261268
R35975 DVSS.n14727 DVSS.n14726 0.00261268
R35976 DVSS.n14657 DVSS.n14656 0.00261268
R35977 DVSS.n14612 DVSS.n14611 0.00261268
R35978 DVSS.n19885 DVSS.n19884 0.00261268
R35979 DVSS.n20030 DVSS.n20029 0.00261268
R35980 DVSS.n454 DVSS.n453 0.00261268
R35981 DVSS.n19312 DVSS.n19308 0.00260496
R35982 DVSS.n19574 DVSS.n19573 0.00260496
R35983 DVSS.n13915 DVSS.n13914 0.0026
R35984 DVSS.n16799 DVSS.n16798 0.0026
R35985 DVSS.n15114 DVSS.n15113 0.0026
R35986 DVSS.n7637 DVSS.n7636 0.0026
R35987 DVSS.n16007 DVSS.n16006 0.0026
R35988 DVSS.n15304 DVSS.n15303 0.0026
R35989 DVSS.n18297 DVSS.n18296 0.0026
R35990 DVSS.n18006 DVSS.n18005 0.0026
R35991 DVSS.n17865 DVSS.n17864 0.0026
R35992 DVSS.n9260 DVSS.n9259 0.0026
R35993 DVSS.n9313 DVSS.n9312 0.0026
R35994 DVSS.n9488 DVSS.n9487 0.0026
R35995 DVSS.n9431 DVSS.n8323 0.0026
R35996 DVSS.n21392 DVSS.n21391 0.0026
R35997 DVSS.n6989 DVSS.n6988 0.00259448
R35998 DVSS.n13649 DVSS.n13648 0.00259448
R35999 DVSS.n13226 DVSS.n13225 0.00259448
R36000 DVSS.n18756 DVSS.n18755 0.00259448
R36001 DVSS.n20133 DVSS.n20132 0.00259404
R36002 DVSS.n20416 DVSS.n20415 0.00259404
R36003 DVSS.n5665 DVSS.n5664 0.00259392
R36004 DVSS.n4448 DVSS.n4447 0.00259392
R36005 DVSS.n7206 DVSS.n7205 0.00259392
R36006 DVSS.n19292 DVSS.n19291 0.00259392
R36007 DVSS.n1047 DVSS.n1046 0.00259392
R36008 DVSS.n4449 DVSS.n4448 0.00259392
R36009 DVSS.n5664 DVSS.n5663 0.00259392
R36010 DVSS.n10957 DVSS.n10956 0.00259392
R36011 DVSS.n9511 DVSS.n9510 0.00259392
R36012 DVSS.n12898 DVSS.n12897 0.00259392
R36013 DVSS.n12703 DVSS.n12702 0.00259392
R36014 DVSS.n12431 DVSS.n12430 0.00259392
R36015 DVSS.n9510 DVSS.n9509 0.00259392
R36016 DVSS.n10956 DVSS.n10955 0.00259392
R36017 DVSS.n17090 DVSS.n17089 0.00259392
R36018 DVSS.n15686 DVSS.n15685 0.00259392
R36019 DVSS.n13509 DVSS.n13508 0.00259392
R36020 DVSS.n20308 DVSS.n20307 0.00259392
R36021 DVSS.n20814 DVSS.n20813 0.00259392
R36022 DVSS.n15687 DVSS.n15686 0.00259392
R36023 DVSS.n17089 DVSS.n17088 0.00259392
R36024 DVSS.n10802 DVSS.n10801 0.00259392
R36025 DVSS.n10778 DVSS.n10777 0.00259392
R36026 DVSS.n11441 DVSS.n11440 0.00259392
R36027 DVSS.n11549 DVSS.n11548 0.00259392
R36028 DVSS.n12083 DVSS.n12082 0.00259392
R36029 DVSS.n21547 DVSS.n21546 0.00259392
R36030 DVSS.n21459 DVSS.n21458 0.00259392
R36031 DVSS.n11548 DVSS.n11547 0.00259392
R36032 DVSS.n11440 DVSS.n11439 0.00259392
R36033 DVSS.n10779 DVSS.n10778 0.00259392
R36034 DVSS.n4684 DVSS.n4683 0.00259392
R36035 DVSS.n4685 DVSS.n4684 0.00259392
R36036 DVSS.n4282 DVSS.n4281 0.00259392
R36037 DVSS.n3505 DVSS.n3504 0.00259392
R36038 DVSS.n3326 DVSS.n3325 0.00259392
R36039 DVSS.n3057 DVSS.n3056 0.00259392
R36040 DVSS.n4281 DVSS.n4280 0.00259392
R36041 DVSS.n9979 DVSS.n9978 0.00259392
R36042 DVSS.n9683 DVSS.n9682 0.00259392
R36043 DVSS.n13411 DVSS.n13410 0.00259392
R36044 DVSS.n20582 DVSS.n20581 0.00259392
R36045 DVSS.n21040 DVSS.n21039 0.00259392
R36046 DVSS.n9684 DVSS.n9683 0.00259392
R36047 DVSS.n9978 DVSS.n9977 0.00259392
R36048 DVSS.n17384 DVSS.n17383 0.00259392
R36049 DVSS.n16198 DVSS.n16197 0.00259392
R36050 DVSS.n18866 DVSS.n18865 0.00259392
R36051 DVSS.n19563 DVSS.n19562 0.00259392
R36052 DVSS.n1262 DVSS.n1261 0.00259392
R36053 DVSS.n16199 DVSS.n16198 0.00259392
R36054 DVSS.n17383 DVSS.n17382 0.00259392
R36055 DVSS.n5462 DVSS.n5461 0.00259392
R36056 DVSS.n5504 DVSS.n5503 0.00259392
R36057 DVSS.n6458 DVSS.n6457 0.00259392
R36058 DVSS.n6596 DVSS.n6595 0.00259392
R36059 DVSS.n3567 DVSS.n3566 0.00259392
R36060 DVSS.n19011 DVSS.n19010 0.00259392
R36061 DVSS.n613 DVSS.n612 0.00259392
R36062 DVSS.n5461 DVSS.n5460 0.00259392
R36063 DVSS.n6595 DVSS.n6594 0.00259392
R36064 DVSS.n5504 DVSS.n5484 0.00259392
R36065 DVSS.n6459 DVSS.n6458 0.00259392
R36066 DVSS.n3568 DVSS.n3567 0.00259392
R36067 DVSS.n12084 DVSS.n12083 0.00259392
R36068 DVSS.n3506 DVSS.n3505 0.00259392
R36069 DVSS.n12899 DVSS.n12898 0.00259392
R36070 DVSS.n18867 DVSS.n18866 0.00259392
R36071 DVSS.n7207 DVSS.n7206 0.00259392
R36072 DVSS.n13412 DVSS.n13411 0.00259392
R36073 DVSS.n13510 DVSS.n13509 0.00259392
R36074 DVSS.n19012 DVSS.n19011 0.00259392
R36075 DVSS.n19564 DVSS.n19563 0.00259392
R36076 DVSS.n21548 DVSS.n21547 0.00259392
R36077 DVSS.n12704 DVSS.n12703 0.00259392
R36078 DVSS.n3327 DVSS.n3326 0.00259392
R36079 DVSS.n12432 DVSS.n12431 0.00259392
R36080 DVSS.n3058 DVSS.n3057 0.00259392
R36081 DVSS.n19293 DVSS.n19292 0.00259392
R36082 DVSS.n20309 DVSS.n20308 0.00259392
R36083 DVSS.n20583 DVSS.n20582 0.00259392
R36084 DVSS.n614 DVSS.n613 0.00259392
R36085 DVSS.n1263 DVSS.n1262 0.00259392
R36086 DVSS.n21460 DVSS.n21459 0.00259392
R36087 DVSS.n1048 DVSS.n1047 0.00259392
R36088 DVSS.n21041 DVSS.n21040 0.00259392
R36089 DVSS.n20815 DVSS.n20814 0.00259392
R36090 DVSS.n18273 DVSS.n18272 0.00258439
R36091 DVSS.n15467 DVSS.n15466 0.00258439
R36092 DVSS.n16667 DVSS.n16666 0.00258431
R36093 DVSS.n17156 DVSS.n17155 0.00258431
R36094 DVSS.n18150 DVSS.n18149 0.00258395
R36095 DVSS.n18469 DVSS.n18468 0.00258395
R36096 DVSS.n15455 DVSS.n15454 0.00258395
R36097 DVSS.n15133 DVSS.n15132 0.00258395
R36098 DVSS.n2375 DVSS.n2374 0.00257445
R36099 DVSS.n9259 DVSS.n9258 0.00257
R36100 DVSS.n9312 DVSS.n9311 0.00257
R36101 DVSS.n9488 DVSS.n9424 0.00257
R36102 DVSS.n9466 DVSS.n8323 0.00257
R36103 DVSS.n12103 DVSS.n12102 0.00257
R36104 DVSS.n21570 DVSS.n21569 0.00257
R36105 DVSS.n21392 DVSS.n21371 0.00257
R36106 DVSS.n3107 DVSS.n3106 0.00256281
R36107 DVSS.n6503 DVSS.n4478 0.00253439
R36108 DVSS.n5721 DVSS.n5720 0.00253439
R36109 DVSS.n5752 DVSS.n5751 0.00253439
R36110 DVSS.n5743 DVSS.n5742 0.00253439
R36111 DVSS.n11246 DVSS.n11245 0.00253439
R36112 DVSS.n11224 DVSS.n11223 0.00253439
R36113 DVSS.n11216 DVSS.n11215 0.00253439
R36114 DVSS.n11255 DVSS.n11254 0.00253439
R36115 DVSS.n17653 DVSS.n17652 0.00253439
R36116 DVSS.n17645 DVSS.n17640 0.00253439
R36117 DVSS.n9833 DVSS.n9832 0.00253439
R36118 DVSS.n11164 DVSS.n11163 0.00253439
R36119 DVSS.n16324 DVSS.n16323 0.00253439
R36120 DVSS.n16342 DVSS.n16341 0.00253439
R36121 DVSS.n16600 DVSS.n16599 0.002525
R36122 DVSS.n16603 DVSS.n16602 0.002525
R36123 DVSS.n18313 DVSS.n18312 0.002525
R36124 DVSS.n18316 DVSS.n18315 0.002525
R36125 DVSS.n5350 DVSS.n5349 0.00251117
R36126 DVSS.n17299 DVSS.n17298 0.00251117
R36127 DVSS.n17287 DVSS.n17285 0.00251117
R36128 DVSS.n16974 DVSS.n16971 0.00251117
R36129 DVSS.n16991 DVSS.n16990 0.00251117
R36130 DVSS.n10629 DVSS.n10628 0.00251117
R36131 DVSS.n1394 DVSS.n1393 0.00251
R36132 DVSS.n4237 DVSS.n4236 0.00251
R36133 DVSS.n4206 DVSS.n4205 0.00251
R36134 DVSS.n4159 DVSS.n4158 0.00251
R36135 DVSS.n3668 DVSS.n3667 0.00251
R36136 DVSS.n19021 DVSS.n19020 0.00251
R36137 DVSS.n630 DVSS.n629 0.00251
R36138 DVSS.n10985 DVSS.n10984 0.0025059
R36139 DVSS.n16922 DVSS.n16921 0.0025059
R36140 DVSS.n9878 DVSS.n9877 0.0025059
R36141 DVSS.n5632 DVSS.n5631 0.0025054
R36142 DVSS.n5801 DVSS.n5800 0.0025054
R36143 DVSS.n5762 DVSS.n5761 0.0025054
R36144 DVSS.n4074 DVSS.n4073 0.0025054
R36145 DVSS.n6978 DVSS.n6977 0.0025054
R36146 DVSS.n5802 DVSS.n5801 0.0025054
R36147 DVSS.n4073 DVSS.n4072 0.0025054
R36148 DVSS.n5631 DVSS.n5630 0.0025054
R36149 DVSS.n6979 DVSS.n6978 0.0025054
R36150 DVSS.n10923 DVSS.n10922 0.0025054
R36151 DVSS.n9849 DVSS.n9848 0.0025054
R36152 DVSS.n11265 DVSS.n11264 0.0025054
R36153 DVSS.n8992 DVSS.n8991 0.0025054
R36154 DVSS.n12959 DVSS.n12958 0.0025054
R36155 DVSS.n9850 DVSS.n9849 0.0025054
R36156 DVSS.n8993 DVSS.n8992 0.0025054
R36157 DVSS.n10922 DVSS.n10921 0.0025054
R36158 DVSS.n12958 DVSS.n12957 0.0025054
R36159 DVSS.n5763 DVSS.n5762 0.0025054
R36160 DVSS.n11266 DVSS.n11265 0.0025054
R36161 DVSS.n17056 DVSS.n17055 0.0025054
R36162 DVSS.n17557 DVSS.n17556 0.0025054
R36163 DVSS.n17600 DVSS.n17599 0.0025054
R36164 DVSS.n15003 DVSS.n15002 0.0025054
R36165 DVSS.n13659 DVSS.n13658 0.0025054
R36166 DVSS.n17556 DVSS.n17555 0.0025054
R36167 DVSS.n15002 DVSS.n15001 0.0025054
R36168 DVSS.n17055 DVSS.n17054 0.0025054
R36169 DVSS.n17599 DVSS.n17598 0.0025054
R36170 DVSS.n13660 DVSS.n13659 0.0025054
R36171 DVSS.n10839 DVSS.n10838 0.0025054
R36172 DVSS.n10783 DVSS.n10782 0.0025054
R36173 DVSS.n11397 DVSS.n11396 0.0025054
R36174 DVSS.n11700 DVSS.n11699 0.0025054
R36175 DVSS.n13033 DVSS.n13032 0.0025054
R36176 DVSS.n11699 DVSS.n11698 0.0025054
R36177 DVSS.n10784 DVSS.n10783 0.0025054
R36178 DVSS.n10840 DVSS.n10839 0.0025054
R36179 DVSS.n11396 DVSS.n11395 0.0025054
R36180 DVSS.n13034 DVSS.n13033 0.0025054
R36181 DVSS.n4702 DVSS.n4701 0.0025054
R36182 DVSS.n4701 DVSS.n4700 0.0025054
R36183 DVSS.n3800 DVSS.n3799 0.0025054
R36184 DVSS.n3772 DVSS.n3771 0.0025054
R36185 DVSS.n3799 DVSS.n3798 0.0025054
R36186 DVSS.n3773 DVSS.n3772 0.0025054
R36187 DVSS.n9945 DVSS.n9944 0.0025054
R36188 DVSS.n11080 DVSS.n11079 0.0025054
R36189 DVSS.n11123 DVSS.n11122 0.0025054
R36190 DVSS.n9082 DVSS.n9081 0.0025054
R36191 DVSS.n13216 DVSS.n13215 0.0025054
R36192 DVSS.n11079 DVSS.n11078 0.0025054
R36193 DVSS.n9083 DVSS.n9082 0.0025054
R36194 DVSS.n9944 DVSS.n9943 0.0025054
R36195 DVSS.n11122 DVSS.n11121 0.0025054
R36196 DVSS.n13215 DVSS.n13214 0.0025054
R36197 DVSS.n17351 DVSS.n17350 0.0025054
R36198 DVSS.n16422 DVSS.n16421 0.0025054
R36199 DVSS.n16383 DVSS.n16382 0.0025054
R36200 DVSS.n7538 DVSS.n7537 0.0025054
R36201 DVSS.n18746 DVSS.n18745 0.0025054
R36202 DVSS.n16423 DVSS.n16422 0.0025054
R36203 DVSS.n7539 DVSS.n7538 0.0025054
R36204 DVSS.n16384 DVSS.n16383 0.0025054
R36205 DVSS.n17350 DVSS.n17349 0.0025054
R36206 DVSS.n18745 DVSS.n18744 0.0025054
R36207 DVSS.n5427 DVSS.n5426 0.0025054
R36208 DVSS.n5481 DVSS.n5480 0.0025054
R36209 DVSS.n6080 DVSS.n6079 0.0025054
R36210 DVSS.n6781 DVSS.n6780 0.0025054
R36211 DVSS.n3589 DVSS.n3588 0.0025054
R36212 DVSS.n5426 DVSS.n5425 0.0025054
R36213 DVSS.n5480 DVSS.n5479 0.0025054
R36214 DVSS.n6780 DVSS.n6779 0.0025054
R36215 DVSS.n6079 DVSS.n6078 0.0025054
R36216 DVSS.n3588 DVSS.n3587 0.0025054
R36217 DVSS.n6881 DVSS.n6880 0.00248147
R36218 DVSS.n4568 DVSS.n4567 0.00248147
R36219 DVSS.n4618 DVSS.n4617 0.00248147
R36220 DVSS.n6754 DVSS.n6753 0.00248147
R36221 DVSS.n6699 DVSS.n6698 0.00248147
R36222 DVSS.n2531 DVSS.n2530 0.00248147
R36223 DVSS.n6392 DVSS.n6391 0.00248147
R36224 DVSS.n4514 DVSS.n4513 0.00248147
R36225 DVSS.n12133 DVSS.n12132 0.00248
R36226 DVSS.n20629 DVSS.n20628 0.00248
R36227 DVSS.n21264 DVSS.n21263 0.00248
R36228 DVSS.n16088 DVSS.n16087 0.00247852
R36229 DVSS.n15976 DVSS.n15975 0.00247852
R36230 DVSS.n16571 DVSS.n16570 0.00247839
R36231 DVSS.n19747 DVSS.n19746 0.00247839
R36232 DVSS.n18190 DVSS.n18189 0.00247839
R36233 DVSS.n18439 DVSS.n18438 0.00247839
R36234 DVSS.n16570 DVSS.n16569 0.00247839
R36235 DVSS.n16758 DVSS.n16757 0.00247839
R36236 DVSS.n15178 DVSS.n15177 0.00247839
R36237 DVSS.n19972 DVSS.n19971 0.00247839
R36238 DVSS.n15550 DVSS.n15549 0.00247839
R36239 DVSS.n16757 DVSS.n16756 0.00247839
R36240 DVSS.n19971 DVSS.n19970 0.00247839
R36241 DVSS.n19746 DVSS.n19745 0.00247839
R36242 DVSS.n6531 DVSS.n6530 0.00247541
R36243 DVSS.n4382 DVSS.n4381 0.00247541
R36244 DVSS.n4090 DVSS.n4089 0.00247541
R36245 DVSS.n5812 DVSS.n5811 0.00247541
R36246 DVSS.n11235 DVSS.n11234 0.00247541
R36247 DVSS.n11047 DVSS.n11046 0.00247541
R36248 DVSS.n17630 DVSS.n17629 0.00247541
R36249 DVSS.n13820 DVSS.n13819 0.00247541
R36250 DVSS.n13782 DVSS.n13781 0.00247541
R36251 DVSS.n13745 DVSS.n13744 0.00247541
R36252 DVSS.n13641 DVSS.n13640 0.00247541
R36253 DVSS.n17553 DVSS.n15872 0.00247541
R36254 DVSS.n7085 DVSS.n6996 0.00247541
R36255 DVSS.n11153 DVSS.n11152 0.00247541
R36256 DVSS.n11076 DVSS.n11068 0.00247541
R36257 DVSS.n17448 DVSS.n17447 0.00247541
R36258 DVSS.n18622 DVSS.n18621 0.00247541
R36259 DVSS.n18649 DVSS.n18648 0.00247541
R36260 DVSS.n18681 DVSS.n18680 0.00247541
R36261 DVSS.n18815 DVSS.n18814 0.00247541
R36262 DVSS.n16353 DVSS.n16352 0.00247541
R36263 DVSS.n10590 DVSS 0.00247183
R36264 DVSS.n10591 DVSS 0.00247183
R36265 DVSS.n5630 DVSS.n5629 0.00244882
R36266 DVSS.n5800 DVSS.n5799 0.00244882
R36267 DVSS.n5761 DVSS.n5760 0.00244882
R36268 DVSS.n6510 DVSS.n6509 0.00244882
R36269 DVSS.n4072 DVSS.n4071 0.00244882
R36270 DVSS.n6980 DVSS.n6979 0.00244882
R36271 DVSS.n19131 DVSS.n19130 0.00244882
R36272 DVSS.n10921 DVSS.n10920 0.00244882
R36273 DVSS.n9848 DVSS.n9847 0.00244882
R36274 DVSS.n11264 DVSS.n11263 0.00244882
R36275 DVSS.n9768 DVSS.n9767 0.00244882
R36276 DVSS.n8991 DVSS.n8990 0.00244882
R36277 DVSS.n12960 DVSS.n12959 0.00244882
R36278 DVSS.n12688 DVSS.n12687 0.00244882
R36279 DVSS.n12487 DVSS.n12486 0.00244882
R36280 DVSS.n12396 DVSS.n12395 0.00244882
R36281 DVSS.n12205 DVSS.n12204 0.00244882
R36282 DVSS.n21291 DVSS.n21290 0.00244882
R36283 DVSS.n21244 DVSS.n21243 0.00244882
R36284 DVSS.n17054 DVSS.n17053 0.00244882
R36285 DVSS.n17558 DVSS.n17557 0.00244882
R36286 DVSS.n17601 DVSS.n17600 0.00244882
R36287 DVSS.n15867 DVSS.n15866 0.00244882
R36288 DVSS.n15004 DVSS.n15003 0.00244882
R36289 DVSS.n13658 DVSS.n13657 0.00244882
R36290 DVSS.n20131 DVSS.n20130 0.00244882
R36291 DVSS.n10841 DVSS.n10840 0.00244882
R36292 DVSS.n10749 DVSS.n10748 0.00244882
R36293 DVSS.n11398 DVSS.n11397 0.00244882
R36294 DVSS.n11411 DVSS.n11410 0.00244882
R36295 DVSS.n11701 DVSS.n11700 0.00244882
R36296 DVSS.n13032 DVSS.n13031 0.00244882
R36297 DVSS.n4700 DVSS.n4699 0.00244882
R36298 DVSS.n3801 DVSS.n3800 0.00244882
R36299 DVSS.n3771 DVSS.n3770 0.00244882
R36300 DVSS.n3311 DVSS.n3310 0.00244882
R36301 DVSS.n3112 DVSS.n3111 0.00244882
R36302 DVSS.n3022 DVSS.n3021 0.00244882
R36303 DVSS.n2835 DVSS.n2834 0.00244882
R36304 DVSS.n741 DVSS.n740 0.00244882
R36305 DVSS.n775 DVSS.n774 0.00244882
R36306 DVSS.n9943 DVSS.n9942 0.00244882
R36307 DVSS.n11081 DVSS.n11080 0.00244882
R36308 DVSS.n11124 DVSS.n11123 0.00244882
R36309 DVSS.n9810 DVSS.n9809 0.00244882
R36310 DVSS.n9081 DVSS.n9080 0.00244882
R36311 DVSS.n13217 DVSS.n13216 0.00244882
R36312 DVSS.n20414 DVSS.n20413 0.00244882
R36313 DVSS.n17349 DVSS.n17348 0.00244882
R36314 DVSS.n16421 DVSS.n16420 0.00244882
R36315 DVSS.n16382 DVSS.n16381 0.00244882
R36316 DVSS.n16299 DVSS.n16298 0.00244882
R36317 DVSS.n7537 DVSS.n7536 0.00244882
R36318 DVSS.n18747 DVSS.n18746 0.00244882
R36319 DVSS.n19405 DVSS.n19404 0.00244882
R36320 DVSS.n5425 DVSS.n5424 0.00244882
R36321 DVSS.n5845 DVSS.n5844 0.00244882
R36322 DVSS.n6081 DVSS.n6080 0.00244882
R36323 DVSS.n6334 DVSS.n6333 0.00244882
R36324 DVSS.n6782 DVSS.n6781 0.00244882
R36325 DVSS.n3590 DVSS.n3589 0.00244882
R36326 DVSS.n14156 DVSS.n14155 0.00243571
R36327 DVSS.n13321 DVSS.n13320 0.00243571
R36328 DVSS.n13320 DVSS.n13319 0.00243571
R36329 DVSS.n14155 DVSS.n14154 0.00243571
R36330 DVSS.n7030 DVSS.n7029 0.00243571
R36331 DVSS.n7071 DVSS.n7070 0.00243571
R36332 DVSS.n7066 DVSS.n7065 0.00243571
R36333 DVSS.n13600 DVSS.n13599 0.00243571
R36334 DVSS.n13622 DVSS.n13621 0.00243571
R36335 DVSS.n13623 DVSS.n13622 0.00243571
R36336 DVSS.n13603 DVSS.n13600 0.00243571
R36337 DVSS.n7073 DVSS.n7071 0.00243571
R36338 DVSS.n7032 DVSS.n7030 0.00243571
R36339 DVSS.n7067 DVSS.n7066 0.00243571
R36340 DVSS.n4948 DVSS.n4947 0.00242857
R36341 DVSS.n4904 DVSS.n4903 0.00242857
R36342 DVSS.n4845 DVSS.n4843 0.00242857
R36343 DVSS.n6221 DVSS.n6220 0.00242857
R36344 DVSS.n6163 DVSS.n6162 0.00242857
R36345 DVSS.n14127 DVSS.n14126 0.00242
R36346 DVSS.n11999 DVSS.n11998 0.00242
R36347 DVSS.n19634 DVSS.n19633 0.00242
R36348 DVSS.n126 DVSS.n125 0.00242
R36349 DVSS.n21119 DVSS.n21118 0.00242
R36350 DVSS.n6992 DVSS.n6991 0.00241688
R36351 DVSS.n19133 DVSS.n19132 0.00241688
R36352 DVSS.n11278 DVSS.n11277 0.00241688
R36353 DVSS.n13136 DVSS.n13135 0.00241688
R36354 DVSS.n12752 DVSS.n12751 0.00241688
R36355 DVSS.n12686 DVSS.n12685 0.00241688
R36356 DVSS.n21210 DVSS.n21208 0.00241688
R36357 DVSS.n11279 DVSS.n11278 0.00241688
R36358 DVSS.n13135 DVSS.n13134 0.00241688
R36359 DVSS.n17587 DVSS.n17586 0.00241688
R36360 DVSS.n15031 DVSS.n15030 0.00241688
R36361 DVSS.n13646 DVSS.n13645 0.00241688
R36362 DVSS.n13571 DVSS.n13570 0.00241688
R36363 DVSS.n17586 DVSS.n17585 0.00241688
R36364 DVSS.n15030 DVSS.n15029 0.00241688
R36365 DVSS.n13572 DVSS.n13571 0.00241688
R36366 DVSS.n6991 DVSS.n6990 0.00241688
R36367 DVSS.n13647 DVSS.n13646 0.00241688
R36368 DVSS.n10752 DVSS.n10751 0.00241688
R36369 DVSS.n11384 DVSS.n11383 0.00241688
R36370 DVSS.n11451 DVSS.n11450 0.00241688
R36371 DVSS.n13065 DVSS.n13064 0.00241688
R36372 DVSS.n11450 DVSS.n11449 0.00241688
R36373 DVSS.n10753 DVSS.n10752 0.00241688
R36374 DVSS.n11383 DVSS.n11382 0.00241688
R36375 DVSS.n13066 DVSS.n13065 0.00241688
R36376 DVSS.n10615 DVSS.n10614 0.00241688
R36377 DVSS.n3746 DVSS.n3745 0.00241688
R36378 DVSS.n3365 DVSS.n3364 0.00241688
R36379 DVSS.n3309 DVSS.n3308 0.00241688
R36380 DVSS.n778 DVSS.n777 0.00241688
R36381 DVSS.n790 DVSS.n788 0.00241688
R36382 DVSS.n3747 DVSS.n3746 0.00241688
R36383 DVSS.n11110 DVSS.n11109 0.00241688
R36384 DVSS.n9054 DVSS.n9053 0.00241688
R36385 DVSS.n13229 DVSS.n13228 0.00241688
R36386 DVSS.n11109 DVSS.n11108 0.00241688
R36387 DVSS.n9055 DVSS.n9054 0.00241688
R36388 DVSS.n13228 DVSS.n13227 0.00241688
R36389 DVSS.n16394 DVSS.n16393 0.00241688
R36390 DVSS.n7512 DVSS.n7511 0.00241688
R36391 DVSS.n18759 DVSS.n18758 0.00241688
R36392 DVSS.n19407 DVSS.n19406 0.00241688
R36393 DVSS.n16395 DVSS.n16394 0.00241688
R36394 DVSS.n7513 DVSS.n7512 0.00241688
R36395 DVSS.n18758 DVSS.n18757 0.00241688
R36396 DVSS.n5328 DVSS.n5327 0.00241688
R36397 DVSS.n5842 DVSS.n5841 0.00241688
R36398 DVSS.n6069 DVSS.n6068 0.00241688
R36399 DVSS.n6448 DVSS.n6447 0.00241688
R36400 DVSS.n6836 DVSS.n6835 0.00241688
R36401 DVSS.n3645 DVSS.n3644 0.00241688
R36402 DVSS.n5841 DVSS.n5840 0.00241688
R36403 DVSS.n6068 DVSS.n6067 0.00241688
R36404 DVSS.n6835 DVSS.n6834 0.00241688
R36405 DVSS.n3644 DVSS.n3643 0.00241688
R36406 DVSS.n6449 DVSS.n6448 0.00241688
R36407 DVSS.n5327 DVSS.n5326 0.00241688
R36408 DVSS.n19132 DVSS.n19131 0.00241688
R36409 DVSS.n19406 DVSS.n19405 0.00241688
R36410 DVSS.n20415 DVSS.n20414 0.00241688
R36411 DVSS.n20132 DVSS.n20131 0.00241688
R36412 DVSS.n3366 DVSS.n3365 0.00241688
R36413 DVSS.n12753 DVSS.n12752 0.00241688
R36414 DVSS.n12685 DVSS.n12684 0.00241688
R36415 DVSS.n790 DVSS.n789 0.00241688
R36416 DVSS.n21210 DVSS.n21209 0.00241688
R36417 DVSS.n778 DVSS.n776 0.00241688
R36418 DVSS.n21246 DVSS.n21245 0.00241688
R36419 DVSS.n5773 DVSS.n5772 0.00241688
R36420 DVSS.n4048 DVSS.n4047 0.00241688
R36421 DVSS.n7109 DVSS.n7108 0.00241688
R36422 DVSS.n5774 DVSS.n5773 0.00241688
R36423 DVSS.n7110 DVSS.n7109 0.00241688
R36424 DVSS.n4047 DVSS.n4046 0.00241688
R36425 DVSS.n12922 DVSS.n12921 0.00241688
R36426 DVSS.n12923 DVSS.n12922 0.00241688
R36427 DVSS.n12050 DVSS.n12049 0.00241688
R36428 DVSS.n12049 DVSS.n12048 0.00241688
R36429 DVSS.n3987 DVSS.n3986 0.00241688
R36430 DVSS.n3988 DVSS.n3987 0.00241688
R36431 DVSS.n13260 DVSS.n13259 0.00241688
R36432 DVSS.n13261 DVSS.n13260 0.00241688
R36433 DVSS.n18789 DVSS.n18788 0.00241688
R36434 DVSS.n18788 DVSS.n18787 0.00241688
R36435 DVSS.n5733 DVSS.n5732 0.00241643
R36436 DVSS.n13821 DVSS.n13820 0.00241643
R36437 DVSS.n13783 DVSS.n13782 0.00241643
R36438 DVSS.n13746 DVSS.n13745 0.00241643
R36439 DVSS.n4672 DVSS.n4671 0.00241643
R36440 DVSS.n18814 DVSS.n18813 0.00241643
R36441 DVSS.n14490 DVSS.n14485 0.00241489
R36442 DVSS.n14472 DVSS.n14470 0.00241489
R36443 DVSS.n14081 DVSS.n14078 0.00241489
R36444 DVSS.n14650 DVSS.n14648 0.00241489
R36445 DVSS.n14172 DVSS.n14171 0.00241489
R36446 DVSS.n14734 DVSS.n14732 0.00241489
R36447 DVSS.n10896 DVSS.n10565 0.00240141
R36448 DVSS.n10879 DVSS.n10876 0.00240141
R36449 DVSS.n10412 DVSS.n10411 0.00240141
R36450 DVSS.n10471 DVSS.n10470 0.00240141
R36451 DVSS.n10897 DVSS.n10563 0.00240141
R36452 DVSS.n10880 DVSS.n10874 0.00240141
R36453 DVSS.n16569 DVSS.n16568 0.00240141
R36454 DVSS.n16574 DVSS.n16573 0.00240141
R36455 DVSS.n16579 DVSS.n16578 0.00240141
R36456 DVSS.n16669 DVSS.n16668 0.00240141
R36457 DVSS.n16703 DVSS.n16702 0.00240141
R36458 DVSS.n16509 DVSS.n16508 0.00240141
R36459 DVSS.n18238 DVSS.n18237 0.00240141
R36460 DVSS.n18236 DVSS.n18235 0.00240141
R36461 DVSS.n18235 DVSS.n18234 0.00240141
R36462 DVSS.n18222 DVSS.n18221 0.00240141
R36463 DVSS.n18455 DVSS.n18454 0.00240141
R36464 DVSS.n18466 DVSS.n18465 0.00240141
R36465 DVSS.n14402 DVSS.n14401 0.00240141
R36466 DVSS.n14409 DVSS.n14408 0.00240141
R36467 DVSS.n19659 DVSS.n19658 0.00240141
R36468 DVSS.n19685 DVSS.n19684 0.00240141
R36469 DVSS.n19696 DVSS.n19695 0.00240141
R36470 DVSS.n19775 DVSS.n19774 0.00240141
R36471 DVSS.n19764 DVSS.n19763 0.00240141
R36472 DVSS.n216 DVSS.n215 0.00240141
R36473 DVSS.n205 DVSS.n204 0.00240141
R36474 DVSS.n16756 DVSS.n16755 0.00240141
R36475 DVSS.n16761 DVSS.n16760 0.00240141
R36476 DVSS.n16766 DVSS.n16765 0.00240141
R36477 DVSS.n17154 DVSS.n17153 0.00240141
R36478 DVSS.n17120 DVSS.n17119 0.00240141
R36479 DVSS.n16855 DVSS.n16854 0.00240141
R36480 DVSS.n15502 DVSS.n15501 0.00240141
R36481 DVSS.n15504 DVSS.n15503 0.00240141
R36482 DVSS.n15505 DVSS.n15504 0.00240141
R36483 DVSS.n15518 DVSS.n15517 0.00240141
R36484 DVSS.n15162 DVSS.n15161 0.00240141
R36485 DVSS.n15136 DVSS.n15135 0.00240141
R36486 DVSS.n14726 DVSS.n14725 0.00240141
R36487 DVSS.n14719 DVSS.n14718 0.00240141
R36488 DVSS.n19868 DVSS.n19867 0.00240141
R36489 DVSS.n19904 DVSS.n19903 0.00240141
R36490 DVSS.n19915 DVSS.n19914 0.00240141
R36491 DVSS.n20000 DVSS.n19999 0.00240141
R36492 DVSS.n19989 DVSS.n19988 0.00240141
R36493 DVSS.n424 DVSS.n423 0.00240141
R36494 DVSS.n413 DVSS.n412 0.00240141
R36495 DVSS.n4242 DVSS.n4241 0.00239333
R36496 DVSS.n4243 DVSS.n4242 0.00239333
R36497 DVSS.n4244 DVSS.n4243 0.00239333
R36498 DVSS.n4245 DVSS.n4244 0.00239333
R36499 DVSS.n4246 DVSS.n4245 0.00239333
R36500 DVSS.n4247 DVSS.n4246 0.00239333
R36501 DVSS.n4248 DVSS.n4247 0.00239333
R36502 DVSS.n4249 DVSS.n4248 0.00239333
R36503 DVSS.n4255 DVSS.n4249 0.00239333
R36504 DVSS.n4255 DVSS.n4254 0.00239333
R36505 DVSS.n4254 DVSS.n4253 0.00239333
R36506 DVSS.n4253 DVSS.n4252 0.00239333
R36507 DVSS.n4252 DVSS.n4251 0.00239333
R36508 DVSS.n4251 DVSS.n4250 0.00239333
R36509 DVSS.n9346 DVSS.n9345 0.00239333
R36510 DVSS.n9347 DVSS.n9346 0.00239333
R36511 DVSS.n9348 DVSS.n9347 0.00239333
R36512 DVSS.n9349 DVSS.n9348 0.00239333
R36513 DVSS.n9350 DVSS.n9349 0.00239333
R36514 DVSS.n9351 DVSS.n9350 0.00239333
R36515 DVSS.n9352 DVSS.n9351 0.00239333
R36516 DVSS.n9353 DVSS.n9352 0.00239333
R36517 DVSS.n9354 DVSS.n9353 0.00239333
R36518 DVSS.n9355 DVSS.n9354 0.00239333
R36519 DVSS.n9356 DVSS.n9355 0.00239333
R36520 DVSS.n9357 DVSS.n9356 0.00239333
R36521 DVSS.n9358 DVSS.n9357 0.00239333
R36522 DVSS.n9359 DVSS.n9358 0.00239333
R36523 DVSS.n9360 DVSS.n9359 0.00239333
R36524 DVSS.n9361 DVSS.n9360 0.00239333
R36525 DVSS.n9362 DVSS.n9361 0.00239333
R36526 DVSS.n9363 DVSS.n9362 0.00239333
R36527 DVSS.n9364 DVSS.n9363 0.00239333
R36528 DVSS.n9365 DVSS.n9364 0.00239333
R36529 DVSS.n9366 DVSS.n9365 0.00239333
R36530 DVSS.n9367 DVSS.n9366 0.00239333
R36531 DVSS.n9368 DVSS.n9367 0.00239333
R36532 DVSS.n9369 DVSS.n9368 0.00239333
R36533 DVSS.n9370 DVSS.n9369 0.00239333
R36534 DVSS.n9371 DVSS.n9370 0.00239333
R36535 DVSS.n9372 DVSS.n9371 0.00239333
R36536 DVSS.n9373 DVSS.n9372 0.00239333
R36537 DVSS.n9374 DVSS.n9373 0.00239333
R36538 DVSS.n9375 DVSS.n9374 0.00239333
R36539 DVSS.n9376 DVSS.n9375 0.00239333
R36540 DVSS.n9377 DVSS.n9376 0.00239333
R36541 DVSS.n9378 DVSS.n9377 0.00239333
R36542 DVSS.n9379 DVSS.n9378 0.00239333
R36543 DVSS.n9380 DVSS.n9379 0.00239333
R36544 DVSS.n9381 DVSS.n9380 0.00239333
R36545 DVSS.n9382 DVSS.n9381 0.00239333
R36546 DVSS.n9383 DVSS.n9382 0.00239333
R36547 DVSS.n9384 DVSS.n9383 0.00239333
R36548 DVSS.n9385 DVSS.n9384 0.00239333
R36549 DVSS.n9386 DVSS.n9385 0.00239333
R36550 DVSS.n9387 DVSS.n9386 0.00239333
R36551 DVSS.n9388 DVSS.n9387 0.00239333
R36552 DVSS.n9389 DVSS.n9388 0.00239333
R36553 DVSS.n9390 DVSS.n9389 0.00239333
R36554 DVSS.n9391 DVSS.n9390 0.00239333
R36555 DVSS.n9392 DVSS.n9391 0.00239333
R36556 DVSS.n9393 DVSS.n9392 0.00239333
R36557 DVSS.n9394 DVSS.n9393 0.00239333
R36558 DVSS.n9395 DVSS.n9394 0.00239333
R36559 DVSS.n9396 DVSS.n9395 0.00239333
R36560 DVSS.n9397 DVSS.n9396 0.00239333
R36561 DVSS.n9398 DVSS.n9397 0.00239333
R36562 DVSS.n9399 DVSS.n9398 0.00239333
R36563 DVSS.n9400 DVSS.n9399 0.00239333
R36564 DVSS.n9401 DVSS.n9400 0.00239333
R36565 DVSS.n9402 DVSS.n9401 0.00239333
R36566 DVSS.n9403 DVSS.n9402 0.00239333
R36567 DVSS.n9404 DVSS.n9403 0.00239333
R36568 DVSS.n9405 DVSS.n9404 0.00239333
R36569 DVSS.n9406 DVSS.n9405 0.00239333
R36570 DVSS.n9407 DVSS.n9406 0.00239333
R36571 DVSS.n9408 DVSS.n9407 0.00239333
R36572 DVSS.n9409 DVSS.n9408 0.00239333
R36573 DVSS.n9410 DVSS.n9409 0.00239333
R36574 DVSS.n9411 DVSS.n9410 0.00239333
R36575 DVSS.n9412 DVSS.n9411 0.00239333
R36576 DVSS.n9413 DVSS.n9412 0.00239333
R36577 DVSS.n9414 DVSS.n9413 0.00239333
R36578 DVSS.n9415 DVSS.n9414 0.00239333
R36579 DVSS.n9416 DVSS.n9415 0.00239333
R36580 DVSS.n9417 DVSS.n9416 0.00239333
R36581 DVSS.n9418 DVSS.n9417 0.00239333
R36582 DVSS.n9419 DVSS.n9418 0.00239333
R36583 DVSS.n9420 DVSS.n9419 0.00239333
R36584 DVSS.n9421 DVSS.n9420 0.00239333
R36585 DVSS.n9484 DVSS.n9483 0.00239333
R36586 DVSS.n9483 DVSS.n9482 0.00239333
R36587 DVSS.n9482 DVSS.n9481 0.00239333
R36588 DVSS.n9481 DVSS.n9480 0.00239333
R36589 DVSS.n9480 DVSS.n9479 0.00239333
R36590 DVSS.n9479 DVSS.n9478 0.00239333
R36591 DVSS.n9478 DVSS.n9448 0.00239333
R36592 DVSS.n9447 DVSS.n9428 0.00239333
R36593 DVSS.n3666 DVSS.n3528 0.00239333
R36594 DVSS.n3670 DVSS.n3666 0.00239333
R36595 DVSS.n3674 DVSS.n3670 0.00239333
R36596 DVSS.n3677 DVSS.n3674 0.00239333
R36597 DVSS.n3680 DVSS.n3677 0.00239333
R36598 DVSS.n3683 DVSS.n3680 0.00239333
R36599 DVSS.n3686 DVSS.n3683 0.00239333
R36600 DVSS.n3696 DVSS.n3686 0.00239333
R36601 DVSS.n3724 DVSS.n3696 0.00239333
R36602 DVSS.n3724 DVSS.n3723 0.00239333
R36603 DVSS.n3723 DVSS.n3717 0.00239333
R36604 DVSS.n3717 DVSS.n3711 0.00239333
R36605 DVSS.n3711 DVSS.n3708 0.00239333
R36606 DVSS.n3708 DVSS.n3705 0.00239333
R36607 DVSS.n3701 DVSS.n1306 0.00239333
R36608 DVSS.n7232 DVSS.n1306 0.00239333
R36609 DVSS.n7234 DVSS.n7232 0.00239333
R36610 DVSS.n7248 DVSS.n7234 0.00239333
R36611 DVSS.n7251 DVSS.n7248 0.00239333
R36612 DVSS.n7254 DVSS.n7251 0.00239333
R36613 DVSS.n7257 DVSS.n7254 0.00239333
R36614 DVSS.n7260 DVSS.n7257 0.00239333
R36615 DVSS.n7263 DVSS.n7260 0.00239333
R36616 DVSS.n7266 DVSS.n7263 0.00239333
R36617 DVSS.n7269 DVSS.n7266 0.00239333
R36618 DVSS.n7272 DVSS.n7269 0.00239333
R36619 DVSS.n7275 DVSS.n7272 0.00239333
R36620 DVSS.n7278 DVSS.n7275 0.00239333
R36621 DVSS.n7281 DVSS.n7278 0.00239333
R36622 DVSS.n7284 DVSS.n7281 0.00239333
R36623 DVSS.n7288 DVSS.n7284 0.00239333
R36624 DVSS.n18891 DVSS.n7288 0.00239333
R36625 DVSS.n18893 DVSS.n18891 0.00239333
R36626 DVSS.n18907 DVSS.n18893 0.00239333
R36627 DVSS.n18910 DVSS.n18907 0.00239333
R36628 DVSS.n18913 DVSS.n18910 0.00239333
R36629 DVSS.n18918 DVSS.n18913 0.00239333
R36630 DVSS.n14090 DVSS.n14087 0.00239333
R36631 DVSS.n14093 DVSS.n14090 0.00239333
R36632 DVSS.n14096 DVSS.n14093 0.00239333
R36633 DVSS.n14099 DVSS.n14096 0.00239333
R36634 DVSS.n14102 DVSS.n14099 0.00239333
R36635 DVSS.n14105 DVSS.n14102 0.00239333
R36636 DVSS.n14108 DVSS.n14105 0.00239333
R36637 DVSS.n14111 DVSS.n14108 0.00239333
R36638 DVSS.n14115 DVSS.n14111 0.00239333
R36639 DVSS.n14134 DVSS.n14115 0.00239333
R36640 DVSS.n14535 DVSS.n14134 0.00239333
R36641 DVSS.n14593 DVSS.n14535 0.00239333
R36642 DVSS.n14593 DVSS.n14592 0.00239333
R36643 DVSS.n14592 DVSS.n14581 0.00239333
R36644 DVSS.n14581 DVSS.n14564 0.00239333
R36645 DVSS.n14564 DVSS.n14561 0.00239333
R36646 DVSS.n14561 DVSS.n14558 0.00239333
R36647 DVSS.n14558 DVSS.n14555 0.00239333
R36648 DVSS.n14555 DVSS.n14552 0.00239333
R36649 DVSS.n14552 DVSS.n14549 0.00239333
R36650 DVSS.n14549 DVSS.n14546 0.00239333
R36651 DVSS.n14546 DVSS.n14543 0.00239333
R36652 DVSS.n14543 DVSS.n14540 0.00239333
R36653 DVSS.n7902 DVSS.n7899 0.00239333
R36654 DVSS.n7905 DVSS.n7902 0.00239333
R36655 DVSS.n7908 DVSS.n7905 0.00239333
R36656 DVSS.n13498 DVSS.n7908 0.00239333
R36657 DVSS.n13498 DVSS.n13497 0.00239333
R36658 DVSS.n13497 DVSS.n13484 0.00239333
R36659 DVSS.n13484 DVSS.n13465 0.00239333
R36660 DVSS.n13465 DVSS.n13462 0.00239333
R36661 DVSS.n13462 DVSS.n13459 0.00239333
R36662 DVSS.n13459 DVSS.n13456 0.00239333
R36663 DVSS.n13456 DVSS.n13453 0.00239333
R36664 DVSS.n13453 DVSS.n13450 0.00239333
R36665 DVSS.n13450 DVSS.n13447 0.00239333
R36666 DVSS.n13447 DVSS.n13444 0.00239333
R36667 DVSS.n13444 DVSS.n13441 0.00239333
R36668 DVSS.n13441 DVSS.n13438 0.00239333
R36669 DVSS.n13438 DVSS.n13435 0.00239333
R36670 DVSS.n13435 DVSS.n13432 0.00239333
R36671 DVSS.n13432 DVSS.n13429 0.00239333
R36672 DVSS.n13429 DVSS.n13426 0.00239333
R36673 DVSS.n13426 DVSS.n7945 0.00239333
R36674 DVSS.n7945 DVSS.n7930 0.00239333
R36675 DVSS.n7930 DVSS.n7913 0.00239333
R36676 DVSS.n11992 DVSS.n11989 0.00239333
R36677 DVSS.n11995 DVSS.n11992 0.00239333
R36678 DVSS.n12001 DVSS.n11995 0.00239333
R36679 DVSS.n12012 DVSS.n12001 0.00239333
R36680 DVSS.n12123 DVSS.n12012 0.00239333
R36681 DVSS.n12123 DVSS.n12122 0.00239333
R36682 DVSS.n12122 DVSS.n12118 0.00239333
R36683 DVSS.n12118 DVSS.n12115 0.00239333
R36684 DVSS.n12016 DVSS.n12015 0.00239333
R36685 DVSS.n12108 DVSS.n12016 0.00239333
R36686 DVSS.n12108 DVSS.n12107 0.00239333
R36687 DVSS.n12107 DVSS.n12097 0.00239333
R36688 DVSS.n12097 DVSS.n12026 0.00239333
R36689 DVSS.n18938 DVSS.n18929 0.00239333
R36690 DVSS.n19023 DVSS.n18938 0.00239333
R36691 DVSS.n19027 DVSS.n19023 0.00239333
R36692 DVSS.n19030 DVSS.n19027 0.00239333
R36693 DVSS.n19033 DVSS.n19030 0.00239333
R36694 DVSS.n19036 DVSS.n19033 0.00239333
R36695 DVSS.n19039 DVSS.n19036 0.00239333
R36696 DVSS.n19049 DVSS.n19039 0.00239333
R36697 DVSS.n19060 DVSS.n19049 0.00239333
R36698 DVSS.n19066 DVSS.n19060 0.00239333
R36699 DVSS.n19072 DVSS.n19066 0.00239333
R36700 DVSS.n19075 DVSS.n19072 0.00239333
R36701 DVSS.n19078 DVSS.n19075 0.00239333
R36702 DVSS.n19081 DVSS.n19078 0.00239333
R36703 DVSS.n19091 DVSS.n19087 0.00239333
R36704 DVSS.n19307 DVSS.n19091 0.00239333
R36705 DVSS.n19314 DVSS.n19307 0.00239333
R36706 DVSS.n19317 DVSS.n19314 0.00239333
R36707 DVSS.n19320 DVSS.n19317 0.00239333
R36708 DVSS.n19323 DVSS.n19320 0.00239333
R36709 DVSS.n19326 DVSS.n19323 0.00239333
R36710 DVSS.n19329 DVSS.n19326 0.00239333
R36711 DVSS.n19332 DVSS.n19329 0.00239333
R36712 DVSS.n19335 DVSS.n19332 0.00239333
R36713 DVSS.n19338 DVSS.n19335 0.00239333
R36714 DVSS.n19341 DVSS.n19338 0.00239333
R36715 DVSS.n19344 DVSS.n19341 0.00239333
R36716 DVSS.n19347 DVSS.n19344 0.00239333
R36717 DVSS.n19350 DVSS.n19347 0.00239333
R36718 DVSS.n19353 DVSS.n19350 0.00239333
R36719 DVSS.n19357 DVSS.n19353 0.00239333
R36720 DVSS.n19376 DVSS.n19357 0.00239333
R36721 DVSS.n19576 DVSS.n19376 0.00239333
R36722 DVSS.n19582 DVSS.n19576 0.00239333
R36723 DVSS.n19585 DVSS.n19582 0.00239333
R36724 DVSS.n19588 DVSS.n19585 0.00239333
R36725 DVSS.n19593 DVSS.n19588 0.00239333
R36726 DVSS.n19600 DVSS.n19597 0.00239333
R36727 DVSS.n19603 DVSS.n19600 0.00239333
R36728 DVSS.n19606 DVSS.n19603 0.00239333
R36729 DVSS.n19609 DVSS.n19606 0.00239333
R36730 DVSS.n19612 DVSS.n19609 0.00239333
R36731 DVSS.n19615 DVSS.n19612 0.00239333
R36732 DVSS.n19618 DVSS.n19615 0.00239333
R36733 DVSS.n19621 DVSS.n19618 0.00239333
R36734 DVSS.n19631 DVSS.n19621 0.00239333
R36735 DVSS.n19818 DVSS.n19631 0.00239333
R36736 DVSS.n19831 DVSS.n19818 0.00239333
R36737 DVSS.n19839 DVSS.n19831 0.00239333
R36738 DVSS.n19850 DVSS.n19839 0.00239333
R36739 DVSS.n20049 DVSS.n19850 0.00239333
R36740 DVSS.n20052 DVSS.n20049 0.00239333
R36741 DVSS.n20055 DVSS.n20052 0.00239333
R36742 DVSS.n20058 DVSS.n20055 0.00239333
R36743 DVSS.n20061 DVSS.n20058 0.00239333
R36744 DVSS.n20064 DVSS.n20061 0.00239333
R36745 DVSS.n20067 DVSS.n20064 0.00239333
R36746 DVSS.n20070 DVSS.n20067 0.00239333
R36747 DVSS.n20073 DVSS.n20070 0.00239333
R36748 DVSS.n20078 DVSS.n20073 0.00239333
R36749 DVSS.n20085 DVSS.n20082 0.00239333
R36750 DVSS.n20088 DVSS.n20085 0.00239333
R36751 DVSS.n20091 DVSS.n20088 0.00239333
R36752 DVSS.n20102 DVSS.n20091 0.00239333
R36753 DVSS.n20112 DVSS.n20102 0.00239333
R36754 DVSS.n20329 DVSS.n20112 0.00239333
R36755 DVSS.n20332 DVSS.n20329 0.00239333
R36756 DVSS.n20335 DVSS.n20332 0.00239333
R36757 DVSS.n20338 DVSS.n20335 0.00239333
R36758 DVSS.n20341 DVSS.n20338 0.00239333
R36759 DVSS.n20344 DVSS.n20341 0.00239333
R36760 DVSS.n20347 DVSS.n20344 0.00239333
R36761 DVSS.n20350 DVSS.n20347 0.00239333
R36762 DVSS.n20353 DVSS.n20350 0.00239333
R36763 DVSS.n20356 DVSS.n20353 0.00239333
R36764 DVSS.n20359 DVSS.n20356 0.00239333
R36765 DVSS.n20362 DVSS.n20359 0.00239333
R36766 DVSS.n20365 DVSS.n20362 0.00239333
R36767 DVSS.n20367 DVSS.n20365 0.00239333
R36768 DVSS.n20379 DVSS.n20367 0.00239333
R36769 DVSS.n20598 DVSS.n20379 0.00239333
R36770 DVSS.n20614 DVSS.n20598 0.00239333
R36771 DVSS.n20619 DVSS.n20614 0.00239333
R36772 DVSS.n20672 DVSS.n20669 0.00239333
R36773 DVSS.n20669 DVSS.n20666 0.00239333
R36774 DVSS.n20666 DVSS.n20663 0.00239333
R36775 DVSS.n20663 DVSS.n20660 0.00239333
R36776 DVSS.n20660 DVSS.n20649 0.00239333
R36777 DVSS.n20649 DVSS.n20636 0.00239333
R36778 DVSS.n20636 DVSS.n20625 0.00239333
R36779 DVSS.n20625 DVSS.n20622 0.00239333
R36780 DVSS.n20622 DVSS.n2 0.00239333
R36781 DVSS.n21578 DVSS.n21575 0.00239333
R36782 DVSS.n21575 DVSS.n21563 0.00239333
R36783 DVSS.n21563 DVSS.n21562 0.00239333
R36784 DVSS.n21562 DVSS.n13 0.00239333
R36785 DVSS.n628 DVSS.n514 0.00239333
R36786 DVSS.n632 DVSS.n628 0.00239333
R36787 DVSS.n636 DVSS.n632 0.00239333
R36788 DVSS.n639 DVSS.n636 0.00239333
R36789 DVSS.n642 DVSS.n639 0.00239333
R36790 DVSS.n645 DVSS.n642 0.00239333
R36791 DVSS.n648 DVSS.n645 0.00239333
R36792 DVSS.n684 DVSS.n648 0.00239333
R36793 DVSS.n725 DVSS.n684 0.00239333
R36794 DVSS.n795 DVSS.n725 0.00239333
R36795 DVSS.n809 DVSS.n795 0.00239333
R36796 DVSS.n812 DVSS.n809 0.00239333
R36797 DVSS.n815 DVSS.n812 0.00239333
R36798 DVSS.n818 DVSS.n815 0.00239333
R36799 DVSS.n828 DVSS.n824 0.00239333
R36800 DVSS.n1063 DVSS.n828 0.00239333
R36801 DVSS.n1069 DVSS.n1063 0.00239333
R36802 DVSS.n1075 DVSS.n1069 0.00239333
R36803 DVSS.n1078 DVSS.n1075 0.00239333
R36804 DVSS.n1081 DVSS.n1078 0.00239333
R36805 DVSS.n1084 DVSS.n1081 0.00239333
R36806 DVSS.n1087 DVSS.n1084 0.00239333
R36807 DVSS.n1090 DVSS.n1087 0.00239333
R36808 DVSS.n1093 DVSS.n1090 0.00239333
R36809 DVSS.n1096 DVSS.n1093 0.00239333
R36810 DVSS.n1099 DVSS.n1096 0.00239333
R36811 DVSS.n1102 DVSS.n1099 0.00239333
R36812 DVSS.n1105 DVSS.n1102 0.00239333
R36813 DVSS.n1108 DVSS.n1105 0.00239333
R36814 DVSS.n1111 DVSS.n1108 0.00239333
R36815 DVSS.n1115 DVSS.n1111 0.00239333
R36816 DVSS.n1278 DVSS.n1115 0.00239333
R36817 DVSS.n1284 DVSS.n1278 0.00239333
R36818 DVSS.n1290 DVSS.n1284 0.00239333
R36819 DVSS.n1293 DVSS.n1290 0.00239333
R36820 DVSS.n1296 DVSS.n1293 0.00239333
R36821 DVSS.n1301 DVSS.n1296 0.00239333
R36822 DVSS.n87 DVSS.n84 0.00239333
R36823 DVSS.n90 DVSS.n87 0.00239333
R36824 DVSS.n93 DVSS.n90 0.00239333
R36825 DVSS.n96 DVSS.n93 0.00239333
R36826 DVSS.n99 DVSS.n96 0.00239333
R36827 DVSS.n102 DVSS.n99 0.00239333
R36828 DVSS.n105 DVSS.n102 0.00239333
R36829 DVSS.n108 DVSS.n105 0.00239333
R36830 DVSS.n118 DVSS.n108 0.00239333
R36831 DVSS.n122 DVSS.n118 0.00239333
R36832 DVSS.n267 DVSS.n122 0.00239333
R36833 DVSS.n275 DVSS.n267 0.00239333
R36834 DVSS.n286 DVSS.n275 0.00239333
R36835 DVSS.n474 DVSS.n286 0.00239333
R36836 DVSS.n477 DVSS.n474 0.00239333
R36837 DVSS.n480 DVSS.n477 0.00239333
R36838 DVSS.n483 DVSS.n480 0.00239333
R36839 DVSS.n486 DVSS.n483 0.00239333
R36840 DVSS.n489 DVSS.n486 0.00239333
R36841 DVSS.n492 DVSS.n489 0.00239333
R36842 DVSS.n495 DVSS.n492 0.00239333
R36843 DVSS.n498 DVSS.n495 0.00239333
R36844 DVSS.n503 DVSS.n498 0.00239333
R36845 DVSS.n20679 DVSS.n20676 0.00239333
R36846 DVSS.n20682 DVSS.n20679 0.00239333
R36847 DVSS.n20684 DVSS.n20682 0.00239333
R36848 DVSS.n20696 DVSS.n20684 0.00239333
R36849 DVSS.n20707 DVSS.n20696 0.00239333
R36850 DVSS.n20875 DVSS.n20707 0.00239333
R36851 DVSS.n20878 DVSS.n20875 0.00239333
R36852 DVSS.n20881 DVSS.n20878 0.00239333
R36853 DVSS.n20884 DVSS.n20881 0.00239333
R36854 DVSS.n20887 DVSS.n20884 0.00239333
R36855 DVSS.n20890 DVSS.n20887 0.00239333
R36856 DVSS.n20893 DVSS.n20890 0.00239333
R36857 DVSS.n20896 DVSS.n20893 0.00239333
R36858 DVSS.n20899 DVSS.n20896 0.00239333
R36859 DVSS.n20902 DVSS.n20899 0.00239333
R36860 DVSS.n20905 DVSS.n20902 0.00239333
R36861 DVSS.n20908 DVSS.n20905 0.00239333
R36862 DVSS.n20911 DVSS.n20908 0.00239333
R36863 DVSS.n20914 DVSS.n20911 0.00239333
R36864 DVSS.n20925 DVSS.n20914 0.00239333
R36865 DVSS.n20936 DVSS.n20925 0.00239333
R36866 DVSS.n21101 DVSS.n20936 0.00239333
R36867 DVSS.n21106 DVSS.n21101 0.00239333
R36868 DVSS.n21113 DVSS.n21110 0.00239333
R36869 DVSS.n21116 DVSS.n21113 0.00239333
R36870 DVSS.n21121 DVSS.n21116 0.00239333
R36871 DVSS.n21259 DVSS.n21121 0.00239333
R36872 DVSS.n21274 DVSS.n21259 0.00239333
R36873 DVSS.n21350 DVSS.n21274 0.00239333
R36874 DVSS.n21353 DVSS.n21350 0.00239333
R36875 DVSS.n21356 DVSS.n21353 0.00239333
R36876 DVSS.n21359 DVSS.n21356 0.00239333
R36877 DVSS.n21366 DVSS.n21359 0.00239333
R36878 DVSS.n21368 DVSS.n21367 0.00239333
R36879 DVSS.n21388 DVSS.n21387 0.00239333
R36880 DVSS.n3050 DVSS.n3049 0.00238571
R36881 DVSS.n16535 DVSS.n16534 0.00237282
R36882 DVSS.n16655 DVSS.n16654 0.00237282
R36883 DVSS.n14221 DVSS.n14220 0.00237282
R36884 DVSS.n14223 DVSS.n14222 0.00237282
R36885 DVSS.n14237 DVSS.n14236 0.00237282
R36886 DVSS.n14239 DVSS.n14238 0.00237282
R36887 DVSS.n14320 DVSS.n14319 0.00237282
R36888 DVSS.n14323 DVSS.n14322 0.00237282
R36889 DVSS.n14335 DVSS.n14334 0.00237282
R36890 DVSS.n14343 DVSS.n14342 0.00237282
R36891 DVSS.n14346 DVSS.n14345 0.00237282
R36892 DVSS.n14350 DVSS.n14349 0.00237282
R36893 DVSS.n14358 DVSS.n14357 0.00237282
R36894 DVSS.n14366 DVSS.n14365 0.00237282
R36895 DVSS.n14413 DVSS.n14412 0.00237282
R36896 DVSS.n19665 DVSS.n19664 0.00237282
R36897 DVSS.n14412 DVSS.n14411 0.00237282
R36898 DVSS.n14342 DVSS.n14335 0.00237282
R36899 DVSS.n14321 DVSS.n14320 0.00237282
R36900 DVSS.n14322 DVSS.n14321 0.00237282
R36901 DVSS.n14238 DVSS.n14237 0.00237282
R36902 DVSS.n14222 DVSS.n14221 0.00237282
R36903 DVSS.n18224 DVSS.n18223 0.00237282
R36904 DVSS.n14334 DVSS.n14325 0.00237282
R36905 DVSS.n14236 DVSS.n14227 0.00237282
R36906 DVSS.n14220 DVSS.n14219 0.00237282
R36907 DVSS.n16534 DVSS.n16533 0.00237282
R36908 DVSS.n19664 DVSS.n19659 0.00237282
R36909 DVSS.n14357 DVSS.n14356 0.00237282
R36910 DVSS.n14365 DVSS.n14358 0.00237282
R36911 DVSS.n14345 DVSS.n14344 0.00237282
R36912 DVSS.n14349 DVSS.n14346 0.00237282
R36913 DVSS.n16722 DVSS.n16721 0.00237282
R36914 DVSS.n14876 DVSS.n14875 0.00237282
R36915 DVSS.n14874 DVSS.n14873 0.00237282
R36916 DVSS.n14870 DVSS.n14869 0.00237282
R36917 DVSS.n14868 DVSS.n14867 0.00237282
R36918 DVSS.n14814 DVSS.n14813 0.00237282
R36919 DVSS.n14812 DVSS.n14811 0.00237282
R36920 DVSS.n14808 DVSS.n14807 0.00237282
R36921 DVSS.n14807 DVSS.n14806 0.00237282
R36922 DVSS.n14797 DVSS.n14796 0.00237282
R36923 DVSS.n14796 DVSS.n14795 0.00237282
R36924 DVSS.n14791 DVSS.n14785 0.00237282
R36925 DVSS.n14784 DVSS.n14783 0.00237282
R36926 DVSS.n14715 DVSS.n14714 0.00237282
R36927 DVSS.n19880 DVSS.n19879 0.00237282
R36928 DVSS.n19879 DVSS.n19868 0.00237282
R36929 DVSS.n14716 DVSS.n14715 0.00237282
R36930 DVSS.n14792 DVSS.n14791 0.00237282
R36931 DVSS.n14785 DVSS.n14784 0.00237282
R36932 DVSS.n14798 DVSS.n14797 0.00237282
R36933 DVSS.n15516 DVSS.n15515 0.00237282
R36934 DVSS.n14875 DVSS.n14874 0.00237282
R36935 DVSS.n14869 DVSS.n14868 0.00237282
R36936 DVSS.n14813 DVSS.n14812 0.00237282
R36937 DVSS.n14809 DVSS.n14808 0.00237282
R36938 DVSS.n14871 DVSS.n14870 0.00237282
R36939 DVSS.n14815 DVSS.n14814 0.00237282
R36940 DVSS.n14877 DVSS.n14876 0.00237282
R36941 DVSS.n14806 DVSS.n14799 0.00237282
R36942 DVSS.n14795 DVSS.n14794 0.00237282
R36943 DVSS.n16721 DVSS.n16720 0.00237282
R36944 DVSS.n17168 DVSS.n17167 0.00237282
R36945 DVSS.n14502 DVSS.n14501 0.00237282
R36946 DVSS.n14620 DVSS.n14619 0.00237282
R36947 DVSS DVSS.n9447 0.00236667
R36948 DVSS.n14570 DVSS.n14569 0.00236
R36949 DVSS.n12008 DVSS.n12007 0.00236
R36950 DVSS.n20040 DVSS.n20039 0.00236
R36951 DVSS.n20371 DVSS.n20370 0.00236
R36952 DVSS.n464 DVSS.n463 0.00236
R36953 DVSS.n20687 DVSS.n20686 0.00236
R36954 DVSS.n21255 DVSS.n21254 0.00236
R36955 DVSS DVSS.n8911 0.00235714
R36956 DVSS.n2364 DVSS.n2363 0.0023496
R36957 DVSS.n2402 DVSS.n2401 0.0023496
R36958 DVSS.n10402 DVSS.n10400 0.00233099
R36959 DVSS.n10461 DVSS.n10459 0.00233099
R36960 DVSS.n10559 DVSS.n10502 0.00233099
R36961 DVSS.n10887 DVSS.n10566 0.00233099
R36962 DVSS.n5267 DVSS.n5266 0.00233099
R36963 DVSS.n10403 DVSS.n10399 0.00233099
R36964 DVSS.n10462 DVSS.n10458 0.00233099
R36965 DVSS.n10560 DVSS.n10501 0.00233099
R36966 DVSS.n10886 DVSS.n10596 0.00233099
R36967 DVSS.n10883 DVSS.n10882 0.00233099
R36968 DVSS.n12472 DVSS.n12471 0.00232835
R36969 DVSS.n10770 DVSS.n10769 0.00232835
R36970 DVSS.n10771 DVSS.n10770 0.00232835
R36971 DVSS.n3098 DVSS.n3097 0.00232835
R36972 DVSS.n5496 DVSS.n5495 0.00232835
R36973 DVSS.n5497 DVSS.n5496 0.00232835
R36974 DVSS.n3097 DVSS.n3096 0.00232835
R36975 DVSS.n12471 DVSS.n12470 0.00232835
R36976 DVSS.n7715 DVSS.n7714 0.0023
R36977 DVSS.n1717 VSS 0.0023
R36978 DVSS.n2241 VSS 0.0023
R36979 DVSS.n2240 VSS 0.0023
R36980 DVSS.n1716 VSS 0.0023
R36981 DVSS.n16046 DVSS.n16045 0.0023
R36982 DVSS.n18305 DVSS 0.0023
R36983 DVSS.n10716 DVSS 0.0023
R36984 DVSS.n10717 DVSS 0.0023
R36985 DVSS.n8313 DVSS 0.0023
R36986 DVSS.n8314 DVSS 0.0023
R36987 DVSS DVSS.n12972 0.0023
R36988 DVSS.n12971 DVSS 0.0023
R36989 DVSS DVSS.n11306 0.0023
R36990 DVSS.n11305 DVSS 0.0023
R36991 DVSS.n8890 DVSS 0.0023
R36992 DVSS.n8889 DVSS 0.0023
R36993 DVSS.n3721 DVSS.n3720 0.0023
R36994 DVSS.n3715 DVSS.n3714 0.0023
R36995 DVSS.n19064 DVSS.n19063 0.0023
R36996 DVSS.n19070 DVSS.n19069 0.0023
R36997 DVSS.n793 DVSS.n792 0.0023
R36998 DVSS.n807 DVSS.n806 0.0023
R36999 DVSS.n5852 DVSS.n5851 0.00229713
R37000 DVSS DVSS.n21578 0.00227333
R37001 DVSS.n4450 DVSS.n4449 0.00227165
R37002 DVSS.n6988 DVSS.n6987 0.00227165
R37003 DVSS.n7089 DVSS.n7088 0.00227165
R37004 DVSS.n7152 DVSS.n7151 0.00227165
R37005 DVSS.n7208 DVSS.n7207 0.00227165
R37006 DVSS.n19148 DVSS.n19147 0.00227165
R37007 DVSS.n19294 DVSS.n19293 0.00227165
R37008 DVSS.n1049 DVSS.n1048 0.00227165
R37009 DVSS.n9509 DVSS.n9508 0.00227165
R37010 DVSS.n12900 DVSS.n12899 0.00227165
R37011 DVSS.n12720 DVSS.n12719 0.00227165
R37012 DVSS.n12682 DVSS.n12681 0.00227165
R37013 DVSS.n12679 DVSS.n12678 0.00227165
R37014 DVSS.n12433 DVSS.n12432 0.00227165
R37015 DVSS.n12176 DVSS.n12175 0.00227165
R37016 DVSS.n12175 DVSS.n12174 0.00227165
R37017 DVSS.n12157 DVSS.n12156 0.00227165
R37018 DVSS.n12155 DVSS.n12154 0.00227165
R37019 DVSS.n21196 DVSS.n21195 0.00227165
R37020 DVSS.n21296 DVSS.n21295 0.00227165
R37021 DVSS.n15688 DVSS.n15687 0.00227165
R37022 DVSS.n13650 DVSS.n13649 0.00227165
R37023 DVSS.n13594 DVSS.n13593 0.00227165
R37024 DVSS.n13541 DVSS.n13540 0.00227165
R37025 DVSS.n13511 DVSS.n13510 0.00227165
R37026 DVSS.n20159 DVSS.n20158 0.00227165
R37027 DVSS.n20310 DVSS.n20309 0.00227165
R37028 DVSS.n20816 DVSS.n20815 0.00227165
R37029 DVSS.n11547 DVSS.n11546 0.00227165
R37030 DVSS.n12085 DVSS.n12084 0.00227165
R37031 DVSS.n21549 DVSS.n21548 0.00227165
R37032 DVSS.n21461 DVSS.n21460 0.00227165
R37033 DVSS.n4280 DVSS.n4279 0.00227165
R37034 DVSS.n3507 DVSS.n3506 0.00227165
R37035 DVSS.n3343 DVSS.n3342 0.00227165
R37036 DVSS.n3306 DVSS.n3305 0.00227165
R37037 DVSS.n3303 DVSS.n3302 0.00227165
R37038 DVSS.n3059 DVSS.n3058 0.00227165
R37039 DVSS.n2804 DVSS.n2803 0.00227165
R37040 DVSS.n2803 DVSS.n2802 0.00227165
R37041 DVSS.n2785 DVSS.n2784 0.00227165
R37042 DVSS.n2783 DVSS.n2782 0.00227165
R37043 DVSS.n803 DVSS.n802 0.00227165
R37044 DVSS.n706 DVSS.n705 0.00227165
R37045 DVSS.n9685 DVSS.n9684 0.00227165
R37046 DVSS.n13225 DVSS.n13224 0.00227165
R37047 DVSS.n13238 DVSS.n13237 0.00227165
R37048 DVSS.n13373 DVSS.n13372 0.00227165
R37049 DVSS.n13413 DVSS.n13412 0.00227165
R37050 DVSS.n20430 DVSS.n20429 0.00227165
R37051 DVSS.n20584 DVSS.n20583 0.00227165
R37052 DVSS.n21042 DVSS.n21041 0.00227165
R37053 DVSS.n16200 DVSS.n16199 0.00227165
R37054 DVSS.n18755 DVSS.n18754 0.00227165
R37055 DVSS.n18768 DVSS.n18767 0.00227165
R37056 DVSS.n18834 DVSS.n18833 0.00227165
R37057 DVSS.n18868 DVSS.n18867 0.00227165
R37058 DVSS.n19422 DVSS.n19421 0.00227165
R37059 DVSS.n19565 DVSS.n19564 0.00227165
R37060 DVSS.n1264 DVSS.n1263 0.00227165
R37061 DVSS.n6594 DVSS.n6593 0.00227165
R37062 DVSS.n3569 DVSS.n3568 0.00227165
R37063 DVSS.n19013 DVSS.n19012 0.00227165
R37064 DVSS.n615 DVSS.n614 0.00227165
R37065 DVSS.n16087 DVSS.n16086 0.00226725
R37066 DVSS.n17777 DVSS.n17776 0.00226725
R37067 DVSS.n18109 DVSS.n18108 0.00226725
R37068 DVSS.n14492 DVSS.n14491 0.00226725
R37069 DVSS.n19683 DVSS.n19682 0.00226725
R37070 DVSS.n19756 DVSS.n19755 0.00226725
R37071 DVSS.n160 DVSS.n159 0.00226725
R37072 DVSS.n18108 DVSS.n18107 0.00226725
R37073 DVSS.n17776 DVSS.n17775 0.00226725
R37074 DVSS.n19682 DVSS.n19675 0.00226725
R37075 DVSS.n14491 DVSS.n14482 0.00226725
R37076 DVSS.n15975 DVSS.n15974 0.00226725
R37077 DVSS.n15886 DVSS.n15885 0.00226725
R37078 DVSS.n15387 DVSS.n15386 0.00226725
R37079 DVSS.n14632 DVSS.n14631 0.00226725
R37080 DVSS.n19901 DVSS.n19890 0.00226725
R37081 DVSS.n19981 DVSS.n19980 0.00226725
R37082 DVSS.n320 DVSS.n319 0.00226725
R37083 DVSS.n15386 DVSS.n15385 0.00226725
R37084 DVSS.n15887 DVSS.n15886 0.00226725
R37085 DVSS.n14633 DVSS.n14632 0.00226725
R37086 DVSS.n19902 DVSS.n19901 0.00226725
R37087 DVSS.n14460 DVSS.n14459 0.00226725
R37088 DVSS.n14662 DVSS.n14661 0.00226725
R37089 DVSS.n19980 DVSS.n19979 0.00226725
R37090 DVSS.n19755 DVSS.n19754 0.00226725
R37091 DVSS.n319 DVSS.n318 0.00226725
R37092 DVSS.n159 DVSS.n158 0.00226725
R37093 DVSS.n7246 DVSS.n7245 0.00224
R37094 DVSS.n18905 DVSS.n18904 0.00224
R37095 DVSS.n19580 DVSS.n19579 0.00224
R37096 DVSS.n1073 DVSS.n1072 0.00224
R37097 DVSS.n1288 DVSS.n1287 0.00224
R37098 DVSS.n5621 DVSS.n5620 0.00223982
R37099 DVSS.n19241 DVSS.n19240 0.00223982
R37100 DVSS.n5620 DVSS.n5619 0.00223982
R37101 DVSS.n10910 DVSS.n10909 0.00223982
R37102 DVSS.n12718 DVSS.n12717 0.00223982
R37103 DVSS.n12399 DVSS.n12398 0.00223982
R37104 DVSS.n21225 DVSS.n21224 0.00223982
R37105 DVSS.n10909 DVSS.n10908 0.00223982
R37106 DVSS.n17043 DVSS.n17042 0.00223982
R37107 DVSS.n20251 DVSS.n20250 0.00223982
R37108 DVSS.n17042 DVSS.n17041 0.00223982
R37109 DVSS.n10852 DVSS.n10851 0.00223982
R37110 DVSS.n10775 DVSS.n10774 0.00223982
R37111 DVSS.n10853 DVSS.n10852 0.00223982
R37112 DVSS.n10776 DVSS.n10775 0.00223982
R37113 DVSS.n5199 DVSS.n5198 0.00223982
R37114 DVSS.n5200 DVSS.n5199 0.00223982
R37115 DVSS.n3341 DVSS.n3340 0.00223982
R37116 DVSS.n3025 DVSS.n3024 0.00223982
R37117 DVSS.n747 DVSS.n744 0.00223982
R37118 DVSS.n754 DVSS.n753 0.00223982
R37119 DVSS.n19240 DVSS.n19239 0.00223982
R37120 DVSS.n20250 DVSS.n20249 0.00223982
R37121 DVSS.n9932 DVSS.n9931 0.00223982
R37122 DVSS.n20524 DVSS.n20523 0.00223982
R37123 DVSS.n20525 DVSS.n20524 0.00223982
R37124 DVSS.n9931 DVSS.n9930 0.00223982
R37125 DVSS.n17340 DVSS.n17339 0.00223982
R37126 DVSS.n19512 DVSS.n19511 0.00223982
R37127 DVSS.n19511 DVSS.n19510 0.00223982
R37128 DVSS.n17339 DVSS.n17338 0.00223982
R37129 DVSS.n5416 DVSS.n5415 0.00223982
R37130 DVSS.n5501 DVSS.n5500 0.00223982
R37131 DVSS.n5415 DVSS.n5414 0.00223982
R37132 DVSS.n5502 DVSS.n5501 0.00223982
R37133 DVSS.n3026 DVSS.n3025 0.00223982
R37134 DVSS.n12400 DVSS.n12399 0.00223982
R37135 DVSS.n3342 DVSS.n3341 0.00223982
R37136 DVSS.n12719 DVSS.n12718 0.00223982
R37137 DVSS.n747 DVSS.n746 0.00223982
R37138 DVSS.n21249 DVSS.n21248 0.00223982
R37139 DVSS.n21225 DVSS.n21223 0.00223982
R37140 DVSS.n754 DVSS.n752 0.00223982
R37141 DVSS.n2011 DVSS.n2010 0.00223571
R37142 DVSS.n2066 DVSS.n2063 0.00223571
R37143 DVSS.n2459 DVSS.n2458 0.00223571
R37144 DVSS.n1999 DVSS.n1998 0.00223571
R37145 DVSS.n1726 DVSS.n1725 0.00223571
R37146 DVSS.n10147 DVSS.n10146 0.00223571
R37147 DVSS.n10187 DVSS.n10186 0.00223571
R37148 DVSS.n10729 DVSS.n10660 0.00223571
R37149 DVSS.n10730 DVSS.n10658 0.00223571
R37150 DVSS.n13111 DVSS.n8291 0.00223571
R37151 DVSS.n13101 DVSS.n8294 0.00223571
R37152 DVSS.n8147 DVSS.n8146 0.00223571
R37153 DVSS.n8158 DVSS.n8157 0.00223571
R37154 DVSS.n8198 DVSS.n8197 0.00223571
R37155 DVSS.n8209 DVSS.n8208 0.00223571
R37156 DVSS.n8233 DVSS.n8232 0.00223571
R37157 DVSS.n13112 DVSS.n8289 0.00223571
R37158 DVSS.n8317 DVSS.n8316 0.00223571
R37159 DVSS.n13100 DVSS.n13099 0.00223571
R37160 DVSS.n12993 DVSS.n11737 0.00223571
R37161 DVSS.n13021 DVSS.n13018 0.00223571
R37162 DVSS.n11841 DVSS.n11840 0.00223571
R37163 DVSS.n11900 DVSS.n11899 0.00223571
R37164 DVSS.n11928 DVSS.n11927 0.00223571
R37165 DVSS.n12992 DVSS.n12991 0.00223571
R37166 DVSS.n12969 DVSS.n11733 0.00223571
R37167 DVSS.n13022 DVSS.n13016 0.00223571
R37168 DVSS.n11327 DVSS.n8342 0.00223571
R37169 DVSS.n11358 DVSS.n11355 0.00223571
R37170 DVSS.n8439 DVSS.n8438 0.00223571
R37171 DVSS.n8450 DVSS.n8449 0.00223571
R37172 DVSS.n8490 DVSS.n8489 0.00223571
R37173 DVSS.n8501 DVSS.n8500 0.00223571
R37174 DVSS.n8525 DVSS.n8524 0.00223571
R37175 DVSS.n11326 DVSS.n11325 0.00223571
R37176 DVSS.n11359 DVSS.n11353 0.00223571
R37177 DVSS.n6265 DVSS.n6264 0.00223571
R37178 DVSS.n8907 DVSS.n8906 0.00223571
R37179 DVSS.n8920 DVSS.n8919 0.00223571
R37180 DVSS.n8909 DVSS.n8908 0.00223571
R37181 DVSS.n12143 DVSS.n12138 0.00223077
R37182 DVSS.n12152 DVSS.n12151 0.00223077
R37183 DVSS.n12608 DVSS.n12603 0.00223077
R37184 DVSS.n12601 DVSS.n12600 0.00223077
R37185 DVSS.n12320 DVSS.n12315 0.00223077
R37186 DVSS.n12313 DVSS.n12312 0.00223077
R37187 DVSS.n12228 DVSS.n12223 0.00223077
R37188 DVSS.n21206 DVSS.n21205 0.00223077
R37189 DVSS.n2763 DVSS.n2758 0.00223077
R37190 DVSS.n2772 DVSS.n2771 0.00223077
R37191 DVSS.n3232 DVSS.n3227 0.00223077
R37192 DVSS.n3225 DVSS.n3224 0.00223077
R37193 DVSS.n2947 DVSS.n2942 0.00223077
R37194 DVSS.n2940 DVSS.n2939 0.00223077
R37195 DVSS.n2855 DVSS.n2852 0.00223077
R37196 DVSS.n882 DVSS.n877 0.00223077
R37197 DVSS.n1393 DVSS.n1391 0.00221
R37198 DVSS.n4236 DVSS.n4234 0.00221
R37199 DVSS.n4205 DVSS.n4203 0.00221
R37200 DVSS.n4158 DVSS.n4157 0.00221
R37201 DVSS.n3373 DVSS.n3372 0.0022086
R37202 DVSS.n711 DVSS.n709 0.00220857
R37203 DVSS.n11681 DVSS.n11680 0.00220306
R37204 DVSS.n11644 DVSS.n11643 0.00220306
R37205 DVSS.n11519 DVSS.n11518 0.00220306
R37206 DVSS.n11482 DVSS.n11481 0.00220306
R37207 DVSS.n11730 DVSS.n11729 0.00220306
R37208 DVSS.n5307 DVSS.n5269 0.00219014
R37209 DVSS.n5309 DVSS.n5308 0.00219014
R37210 DVSS.n5189 DVSS.n5188 0.00219014
R37211 DVSS.n5183 DVSS.n5182 0.00219014
R37212 DVSS.n5151 DVSS.n5150 0.00219014
R37213 DVSS.n5145 DVSS.n5144 0.00219014
R37214 DVSS.n5097 DVSS.n5096 0.00219014
R37215 DVSS.n5091 DVSS.n5090 0.00219014
R37216 DVSS.n10406 DVSS.n10405 0.00219014
R37217 DVSS.n10465 DVSS.n10464 0.00219014
R37218 DVSS.n10900 DVSS.n10562 0.00219014
R37219 DVSS.n16075 DVSS.n16074 0.00219014
R37220 DVSS.n18134 DVSS.n18133 0.00219014
R37221 DVSS.n18140 DVSS.n18139 0.00219014
R37222 DVSS.n18258 DVSS.n18257 0.00219014
R37223 DVSS.n18244 DVSS.n18243 0.00219014
R37224 DVSS.n18178 DVSS.n18177 0.00219014
R37225 DVSS.n18426 DVSS.n18425 0.00219014
R37226 DVSS.n18465 DVSS.n18464 0.00219014
R37227 DVSS.n14388 DVSS.n14387 0.00219014
R37228 DVSS.n14459 DVSS.n14458 0.00219014
R37229 DVSS.n14480 DVSS.n14479 0.00219014
R37230 DVSS.n14504 DVSS.n14503 0.00219014
R37231 DVSS.n19671 DVSS.n19670 0.00219014
R37232 DVSS.n19675 DVSS.n19674 0.00219014
R37233 DVSS.n19715 DVSS.n19714 0.00219014
R37234 DVSS.n19752 DVSS.n19751 0.00219014
R37235 DVSS.n19794 DVSS.n19793 0.00219014
R37236 DVSS.n146 DVSS.n145 0.00219014
R37237 DVSS.n235 DVSS.n234 0.00219014
R37238 DVSS.n186 DVSS.n185 0.00219014
R37239 DVSS.n15967 DVSS.n15966 0.00219014
R37240 DVSS.n15439 DVSS.n15438 0.00219014
R37241 DVSS.n15445 DVSS.n15444 0.00219014
R37242 DVSS.n15482 DVSS.n15481 0.00219014
R37243 DVSS.n15496 DVSS.n15495 0.00219014
R37244 DVSS.n15562 DVSS.n15561 0.00219014
R37245 DVSS.n15203 DVSS.n15202 0.00219014
R37246 DVSS.n15137 DVSS.n15136 0.00219014
R37247 DVSS.n14762 DVSS.n14761 0.00219014
R37248 DVSS.n14663 DVSS.n14662 0.00219014
R37249 DVSS.n14636 DVSS.n14635 0.00219014
R37250 DVSS.n14601 DVSS.n14600 0.00219014
R37251 DVSS.n19886 DVSS.n19885 0.00219014
R37252 DVSS.n19890 DVSS.n19889 0.00219014
R37253 DVSS.n19934 DVSS.n19933 0.00219014
R37254 DVSS.n19977 DVSS.n19976 0.00219014
R37255 DVSS.n20019 DVSS.n20018 0.00219014
R37256 DVSS.n306 DVSS.n305 0.00219014
R37257 DVSS.n443 DVSS.n442 0.00219014
R37258 DVSS.n394 DVSS.n393 0.00219014
R37259 DVSS.n9186 DVSS.n9185 0.00218
R37260 DVSS.n10063 DVSS.n10062 0.00217143
R37261 DVSS.n10127 DVSS.n10126 0.00217143
R37262 DVSS.n10175 DVSS.n10174 0.00217143
R37263 DVSS.n10725 DVSS.n10693 0.00217143
R37264 DVSS.n5058 DVSS.n4646 0.00217143
R37265 DVSS.n10056 DVSS.n10055 0.00217143
R37266 DVSS.n10064 DVSS.n10060 0.00217143
R37267 DVSS.n10076 DVSS.n10075 0.00217143
R37268 DVSS.n10078 DVSS.n10077 0.00217143
R37269 DVSS.n10121 DVSS.n10120 0.00217143
R37270 DVSS.n10128 DVSS.n10125 0.00217143
R37271 DVSS.n10137 DVSS.n10136 0.00217143
R37272 DVSS.n10169 DVSS.n10168 0.00217143
R37273 DVSS.n10176 DVSS.n10173 0.00217143
R37274 DVSS.n10189 DVSS.n10188 0.00217143
R37275 DVSS.n10724 DVSS.n10722 0.00217143
R37276 DVSS.n10733 DVSS.n10732 0.00217143
R37277 DVSS.n8149 DVSS.n8148 0.00217143
R37278 DVSS.n8200 DVSS.n8199 0.00217143
R37279 DVSS.n8286 DVSS.n8234 0.00217143
R37280 DVSS.n8320 DVSS.n8318 0.00217143
R37281 DVSS.n8150 DVSS.n8147 0.00217143
R37282 DVSS.n8159 DVSS.n8158 0.00217143
R37283 DVSS.n8201 DVSS.n8198 0.00217143
R37284 DVSS.n8210 DVSS.n8209 0.00217143
R37285 DVSS.n8287 DVSS.n8233 0.00217143
R37286 DVSS.n8295 DVSS.n8289 0.00217143
R37287 DVSS.n8321 DVSS.n8317 0.00217143
R37288 DVSS.n13099 DVSS.n13098 0.00217143
R37289 DVSS.n11831 DVSS.n11829 0.00217143
R37290 DVSS.n11890 DVSS.n11888 0.00217143
R37291 DVSS.n11981 DVSS.n11929 0.00217143
R37292 DVSS.n13002 DVSS.n11734 0.00217143
R37293 DVSS.n11832 DVSS.n11828 0.00217143
R37294 DVSS.n11891 DVSS.n11887 0.00217143
R37295 DVSS.n11982 DVSS.n11928 0.00217143
R37296 DVSS.n12991 DVSS.n12990 0.00217143
R37297 DVSS.n13003 DVSS.n11733 0.00217143
R37298 DVSS.n13016 DVSS.n13015 0.00217143
R37299 DVSS.n8441 DVSS.n8440 0.00217143
R37300 DVSS.n8492 DVSS.n8491 0.00217143
R37301 DVSS.n8583 DVSS.n8526 0.00217143
R37302 DVSS.n11336 DVSS.n8339 0.00217143
R37303 DVSS.n6044 DVSS.n6043 0.00217143
R37304 DVSS.n8442 DVSS.n8439 0.00217143
R37305 DVSS.n8451 DVSS.n8450 0.00217143
R37306 DVSS.n8493 DVSS.n8490 0.00217143
R37307 DVSS.n8502 DVSS.n8501 0.00217143
R37308 DVSS.n8584 DVSS.n8525 0.00217143
R37309 DVSS.n11325 DVSS.n11324 0.00217143
R37310 DVSS.n11337 DVSS.n8338 0.00217143
R37311 DVSS.n11362 DVSS.n11361 0.00217143
R37312 DVSS.n6326 DVSS.n6108 0.00217143
R37313 DVSS.n8692 DVSS.n8691 0.00217143
R37314 DVSS.n8696 DVSS.n8695 0.00217143
R37315 DVSS.n8710 DVSS.n8709 0.00217143
R37316 DVSS.n8712 DVSS.n8711 0.00217143
R37317 DVSS.n8753 DVSS.n8752 0.00217143
R37318 DVSS.n8759 DVSS.n8756 0.00217143
R37319 DVSS.n8771 DVSS.n8770 0.00217143
R37320 DVSS.n8773 DVSS.n8772 0.00217143
R37321 DVSS.n8798 DVSS.n8797 0.00217143
R37322 DVSS.n8860 DVSS.n8801 0.00217143
R37323 DVSS.n8921 DVSS.n8864 0.00217143
R37324 DVSS.n8868 DVSS.n8867 0.00217143
R37325 DVSS.n8899 DVSS.n8895 0.00217143
R37326 DVSS.n8903 DVSS.n8902 0.00217143
R37327 DVSS.n8705 DVSS.n8704 0.00217143
R37328 DVSS.n8758 DVSS.n8757 0.00217143
R37329 DVSS.n8859 DVSS.n8802 0.00217143
R37330 DVSS.n8898 DVSS.n8896 0.00217143
R37331 DVSS.n17801 DVSS.n17800 0.00216167
R37332 DVSS.n19646 DVSS.n19645 0.00216167
R37333 DVSS.n19713 DVSS.n19712 0.00216167
R37334 DVSS.n19791 DVSS.n19790 0.00216167
R37335 DVSS.n144 DVSS.n143 0.00216167
R37336 DVSS.n232 DVSS.n231 0.00216167
R37337 DVSS.n188 DVSS.n187 0.00216167
R37338 DVSS.n17800 DVSS.n17799 0.00216167
R37339 DVSS.n15780 DVSS.n15779 0.00216167
R37340 DVSS.n19855 DVSS.n19854 0.00216167
R37341 DVSS.n19931 DVSS.n19930 0.00216167
R37342 DVSS.n20016 DVSS.n20015 0.00216167
R37343 DVSS.n304 DVSS.n303 0.00216167
R37344 DVSS.n440 DVSS.n439 0.00216167
R37345 DVSS.n396 DVSS.n395 0.00216167
R37346 DVSS.n15779 DVSS.n7654 0.00216167
R37347 DVSS.n19712 DVSS.n19711 0.00216167
R37348 DVSS.n19854 DVSS.n19853 0.00216167
R37349 DVSS.n19645 DVSS.n19644 0.00216167
R37350 DVSS.n19932 DVSS.n19931 0.00216167
R37351 DVSS.n143 DVSS.n142 0.00216167
R37352 DVSS.n303 DVSS.n302 0.00216167
R37353 DVSS.n20017 DVSS.n20016 0.00216167
R37354 DVSS.n19792 DVSS.n19791 0.00216167
R37355 DVSS.n189 DVSS.n188 0.00216167
R37356 DVSS.n397 DVSS.n396 0.00216167
R37357 DVSS.n441 DVSS.n440 0.00216167
R37358 DVSS.n233 DVSS.n232 0.00216167
R37359 DVSS.n2047 DVSS.n2046 0.00215552
R37360 DVSS.n7092 DVSS.n7091 0.00215157
R37361 DVSS.n11229 DVSS.n11228 0.00215157
R37362 DVSS.n17636 DVSS.n17635 0.00215157
R37363 DVSS.n13591 DVSS.n13590 0.00215157
R37364 DVSS.n11159 DVSS.n11158 0.00215157
R37365 DVSS.n13241 DVSS.n13240 0.00215157
R37366 DVSS.n18771 DVSS.n18770 0.00215157
R37367 DVSS.n5562 DVSS.n5561 0.00215128
R37368 DVSS.n5784 DVSS.n5783 0.00215128
R37369 DVSS.n4057 DVSS.n4056 0.00215128
R37370 DVSS.n6961 DVSS.n6960 0.00215128
R37371 DVSS.n6963 DVSS.n6962 0.00215128
R37372 DVSS.n6967 DVSS.n6966 0.00215128
R37373 DVSS.n6969 DVSS.n6968 0.00215128
R37374 DVSS.n7100 DVSS.n7099 0.00215128
R37375 DVSS.n7201 DVSS.n7200 0.00215128
R37376 DVSS.n19143 DVSS.n19142 0.00215128
R37377 DVSS.n5783 DVSS.n5782 0.00215128
R37378 DVSS.n7099 DVSS.n7098 0.00215128
R37379 DVSS.n4058 DVSS.n4057 0.00215128
R37380 DVSS.n5563 DVSS.n5562 0.00215128
R37381 DVSS.n10204 DVSS.n10203 0.00215128
R37382 DVSS.n11290 DVSS.n11289 0.00215128
R37383 DVSS.n13124 DVSS.n13123 0.00215128
R37384 DVSS.n12934 DVSS.n12933 0.00215128
R37385 DVSS.n12725 DVSS.n12724 0.00215128
R37386 DVSS.n12401 DVSS.n12400 0.00215128
R37387 DVSS.n12935 DVSS.n12934 0.00215128
R37388 DVSS.n13123 DVSS.n13122 0.00215128
R37389 DVSS.n10203 DVSS.n10202 0.00215128
R37390 DVSS.n11291 DVSS.n11290 0.00215128
R37391 DVSS.n16949 DVSS.n16948 0.00215128
R37392 DVSS.n17575 DVSS.n17574 0.00215128
R37393 DVSS.n15019 DVSS.n15018 0.00215128
R37394 DVSS.n13842 DVSS.n13841 0.00215128
R37395 DVSS.n13841 DVSS.n13840 0.00215128
R37396 DVSS.n13832 DVSS.n13831 0.00215128
R37397 DVSS.n13830 DVSS.n13829 0.00215128
R37398 DVSS.n13704 DVSS.n13703 0.00215128
R37399 DVSS.n13702 DVSS.n13701 0.00215128
R37400 DVSS.n13698 DVSS.n13697 0.00215128
R37401 DVSS.n13697 DVSS.n13696 0.00215128
R37402 DVSS.n13687 DVSS.n13686 0.00215128
R37403 DVSS.n13686 DVSS.n13685 0.00215128
R37404 DVSS.n13678 DVSS.n13677 0.00215128
R37405 DVSS.n13671 DVSS.n13670 0.00215128
R37406 DVSS.n13583 DVSS.n13582 0.00215128
R37407 DVSS.n13519 DVSS.n13518 0.00215128
R37408 DVSS.n20154 DVSS.n20153 0.00215128
R37409 DVSS.n13584 DVSS.n13583 0.00215128
R37410 DVSS.n13699 DVSS.n13698 0.00215128
R37411 DVSS.n13703 DVSS.n13702 0.00215128
R37412 DVSS.n13831 DVSS.n13830 0.00215128
R37413 DVSS.n13833 DVSS.n13832 0.00215128
R37414 DVSS.n13705 DVSS.n13704 0.00215128
R37415 DVSS.n13843 DVSS.n13842 0.00215128
R37416 DVSS.n13840 DVSS.n13835 0.00215128
R37417 DVSS.n15018 DVSS.n15017 0.00215128
R37418 DVSS.n13696 DVSS.n13689 0.00215128
R37419 DVSS.n16948 DVSS.n16947 0.00215128
R37420 DVSS.n17574 DVSS.n17573 0.00215128
R37421 DVSS.n6968 DVSS.n6967 0.00215128
R37422 DVSS.n6962 DVSS.n6961 0.00215128
R37423 DVSS.n6966 DVSS.n6965 0.00215128
R37424 DVSS.n13677 DVSS.n13672 0.00215128
R37425 DVSS.n13672 DVSS.n13671 0.00215128
R37426 DVSS.n13688 DVSS.n13687 0.00215128
R37427 DVSS.n6960 DVSS.n6959 0.00215128
R37428 DVSS.n13685 DVSS.n13680 0.00215128
R37429 DVSS.n10607 DVSS.n10606 0.00215128
R37430 DVSS.n10613 DVSS.n10612 0.00215128
R37431 DVSS.n11372 DVSS.n11371 0.00215128
R37432 DVSS.n11415 DVSS.n11414 0.00215128
R37433 DVSS.n13077 DVSS.n13076 0.00215128
R37434 DVSS.n12038 DVSS.n12037 0.00215128
R37435 DVSS.n12037 DVSS.n12036 0.00215128
R37436 DVSS.n13078 DVSS.n13077 0.00215128
R37437 DVSS.n11371 DVSS.n11370 0.00215128
R37438 DVSS.n10612 DVSS.n10611 0.00215128
R37439 DVSS.n10608 DVSS.n10607 0.00215128
R37440 DVSS.n11414 DVSS.n11413 0.00215128
R37441 DVSS.n5216 DVSS.n5215 0.00215128
R37442 DVSS.n5215 DVSS.n5214 0.00215128
R37443 DVSS.n3978 DVSS.n3977 0.00215128
R37444 DVSS.n3756 DVSS.n3755 0.00215128
R37445 DVSS.n3348 DVSS.n3347 0.00215128
R37446 DVSS.n3027 DVSS.n3026 0.00215128
R37447 DVSS.n3757 DVSS.n3756 0.00215128
R37448 DVSS.n3977 DVSS.n3976 0.00215128
R37449 DVSS.n9905 DVSS.n9904 0.00215128
R37450 DVSS.n11098 DVSS.n11097 0.00215128
R37451 DVSS.n9066 DVSS.n9065 0.00215128
R37452 DVSS.n13190 DVSS.n13189 0.00215128
R37453 DVSS.n13192 DVSS.n13191 0.00215128
R37454 DVSS.n13201 DVSS.n13200 0.00215128
R37455 DVSS.n13204 DVSS.n13203 0.00215128
R37456 DVSS.n13249 DVSS.n13248 0.00215128
R37457 DVSS.n13405 DVSS.n13404 0.00215128
R37458 DVSS.n20425 DVSS.n20424 0.00215128
R37459 DVSS.n13248 DVSS.n13247 0.00215128
R37460 DVSS.n9067 DVSS.n9066 0.00215128
R37461 DVSS.n13191 DVSS.n13190 0.00215128
R37462 DVSS.n13189 DVSS.n13188 0.00215128
R37463 DVSS.n13202 DVSS.n13201 0.00215128
R37464 DVSS.n13203 DVSS.n13202 0.00215128
R37465 DVSS.n9904 DVSS.n9903 0.00215128
R37466 DVSS.n11097 DVSS.n11096 0.00215128
R37467 DVSS.n17258 DVSS.n17257 0.00215128
R37468 DVSS.n16404 DVSS.n16403 0.00215128
R37469 DVSS.n7522 DVSS.n7521 0.00215128
R37470 DVSS.n18582 DVSS.n18581 0.00215128
R37471 DVSS.n18584 DVSS.n18583 0.00215128
R37472 DVSS.n18600 DVSS.n18599 0.00215128
R37473 DVSS.n18602 DVSS.n18601 0.00215128
R37474 DVSS.n18691 DVSS.n18690 0.00215128
R37475 DVSS.n18693 DVSS.n18692 0.00215128
R37476 DVSS.n18703 DVSS.n18702 0.00215128
R37477 DVSS.n18705 DVSS.n18704 0.00215128
R37478 DVSS.n18708 DVSS.n18707 0.00215128
R37479 DVSS.n18710 DVSS.n18709 0.00215128
R37480 DVSS.n18726 DVSS.n18725 0.00215128
R37481 DVSS.n18736 DVSS.n18735 0.00215128
R37482 DVSS.n18779 DVSS.n18778 0.00215128
R37483 DVSS.n18861 DVSS.n18860 0.00215128
R37484 DVSS.n19417 DVSS.n19416 0.00215128
R37485 DVSS.n7523 DVSS.n7522 0.00215128
R37486 DVSS.n18583 DVSS.n18582 0.00215128
R37487 DVSS.n18601 DVSS.n18600 0.00215128
R37488 DVSS.n18692 DVSS.n18691 0.00215128
R37489 DVSS.n18704 DVSS.n18703 0.00215128
R37490 DVSS.n18709 DVSS.n18708 0.00215128
R37491 DVSS.n18735 DVSS.n18726 0.00215128
R37492 DVSS.n18778 DVSS.n18777 0.00215128
R37493 DVSS.n18725 DVSS.n18716 0.00215128
R37494 DVSS.n18702 DVSS.n18695 0.00215128
R37495 DVSS.n18599 DVSS.n18590 0.00215128
R37496 DVSS.n18690 DVSS.n18689 0.00215128
R37497 DVSS.n18581 DVSS.n18580 0.00215128
R37498 DVSS.n18707 DVSS.n18706 0.00215128
R37499 DVSS.n16405 DVSS.n16404 0.00215128
R37500 DVSS.n17257 DVSS.n17256 0.00215128
R37501 DVSS.n5321 DVSS.n5320 0.00215128
R37502 DVSS.n5325 DVSS.n5324 0.00215128
R37503 DVSS.n6059 DVSS.n6058 0.00215128
R37504 DVSS.n6337 DVSS.n6336 0.00215128
R37505 DVSS.n6826 DVSS.n6825 0.00215128
R37506 DVSS.n3635 DVSS.n3634 0.00215128
R37507 DVSS.n6058 DVSS.n6057 0.00215128
R37508 DVSS.n6825 DVSS.n6824 0.00215128
R37509 DVSS.n3634 DVSS.n3633 0.00215128
R37510 DVSS.n5320 DVSS.n5319 0.00215128
R37511 DVSS.n5324 DVSS.n5323 0.00215128
R37512 DVSS.n18860 DVSS.n18859 0.00215128
R37513 DVSS.n13520 DVSS.n13519 0.00215128
R37514 DVSS.n13404 DVSS.n13403 0.00215128
R37515 DVSS.n7200 DVSS.n7199 0.00215128
R37516 DVSS.n12402 DVSS.n12401 0.00215128
R37517 DVSS.n3028 DVSS.n3027 0.00215128
R37518 DVSS.n20529 DVSS.n20528 0.00215128
R37519 DVSS.n20255 DVSS.n20254 0.00215128
R37520 DVSS.n12726 DVSS.n12725 0.00215128
R37521 DVSS.n14523 DVSS.n14522 0.00215
R37522 DVSS.n19822 DVSS.n19821 0.00215
R37523 DVSS.n258 DVSS.n257 0.00215
R37524 DVSS.n10728 DVSS 0.00212857
R37525 DVSS.n19163 DVSS.n19162 0.00212162
R37526 DVSS.n19116 DVSS.n19114 0.00212162
R37527 DVSS.n19433 DVSS.n19432 0.00212162
R37528 DVSS.n19390 DVSS.n19389 0.00212162
R37529 DVSS.n20171 DVSS.n20170 0.00212162
R37530 DVSS.n20148 DVSS.n20146 0.00212162
R37531 DVSS.n20441 DVSS.n20440 0.00212162
R37532 DVSS.n20398 DVSS.n20397 0.00212162
R37533 DVSS.n10334 DVSS.n10333 0.00211972
R37534 DVSS.n10315 DVSS.n10314 0.00211972
R37535 DVSS.n10342 DVSS.n10341 0.00211972
R37536 DVSS.n4777 DVSS.n4776 0.00210714
R37537 DVSS.n4961 DVSS.n4960 0.00210714
R37538 DVSS.n4917 DVSS.n4916 0.00210714
R37539 DVSS.n4857 DVSS.n4856 0.00210714
R37540 DVSS.n10081 DVSS.n10080 0.00210714
R37541 DVSS.n10142 DVSS.n10141 0.00210714
R37542 DVSS.n10696 DVSS.n10695 0.00210714
R37543 DVSS.n6816 DVSS.n6815 0.00210714
R37544 DVSS.n3968 DVSS.n3967 0.00210714
R37545 DVSS.n3904 DVSS.n3903 0.00210714
R37546 DVSS.n3858 DVSS.n3857 0.00210714
R37547 DVSS.n3607 DVSS.n3606 0.00210714
R37548 DVSS.n2596 DVSS.n2595 0.00210714
R37549 DVSS.n11774 DVSS.n11773 0.00210714
R37550 DVSS.n5982 DVSS.n5981 0.00210714
R37551 DVSS.n5936 DVSS.n5935 0.00210714
R37552 DVSS.n6234 DVSS.n6233 0.00210714
R37553 DVSS.n6176 DVSS.n6175 0.00210714
R37554 DVSS.n8714 DVSS.n8713 0.00210714
R37555 DVSS.n8775 DVSS.n8774 0.00210714
R37556 DVSS.n8870 DVSS.n8869 0.00210714
R37557 DVSS.n5663 DVSS.n5662 0.00209449
R37558 DVSS.n5671 DVSS.n5670 0.00209449
R37559 DVSS.n4422 DVSS.n4421 0.00209449
R37560 DVSS.n4414 DVSS.n4413 0.00209449
R37561 DVSS.n7090 DVSS.n7089 0.00209449
R37562 DVSS.n7096 DVSS.n7095 0.00209449
R37563 DVSS.n19171 DVSS.n19170 0.00209449
R37564 DVSS.n19179 DVSS.n19178 0.00209449
R37565 DVSS.n19266 DVSS.n19265 0.00209449
R37566 DVSS.n19258 DVSS.n19257 0.00209449
R37567 DVSS.n1021 DVSS.n1020 0.00209449
R37568 DVSS.n1013 DVSS.n1012 0.00209449
R37569 DVSS.n10963 DVSS.n10962 0.00209449
R37570 DVSS.n9539 DVSS.n9538 0.00209449
R37571 DVSS.n9550 DVSS.n9549 0.00209449
R37572 DVSS.n12870 DVSS.n12869 0.00209449
R37573 DVSS.n12859 DVSS.n12858 0.00209449
R37574 DVSS.n12755 DVSS.n12754 0.00209449
R37575 DVSS.n12750 DVSS.n12749 0.00209449
R37576 DVSS.n12680 DVSS.n12679 0.00209449
R37577 DVSS.n12475 DVSS.n12474 0.00209449
R37578 DVSS.n12457 DVSS.n12456 0.00209449
R37579 DVSS.n12434 DVSS.n12433 0.00209449
R37580 DVSS.n12429 DVSS.n12428 0.00209449
R37581 DVSS.n12428 DVSS.n12427 0.00209449
R37582 DVSS.n12418 DVSS.n12417 0.00209449
R37583 DVSS.n12158 DVSS.n12157 0.00209449
R37584 DVSS.n21295 DVSS.n21294 0.00209449
R37585 DVSS.n21207 DVSS.n21201 0.00209449
R37586 DVSS.n17096 DVSS.n17095 0.00209449
R37587 DVSS.n15658 DVSS.n15657 0.00209449
R37588 DVSS.n15647 DVSS.n15646 0.00209449
R37589 DVSS.n13593 DVSS.n13592 0.00209449
R37590 DVSS.n13587 DVSS.n13586 0.00209449
R37591 DVSS.n20179 DVSS.n20178 0.00209449
R37592 DVSS.n20190 DVSS.n20189 0.00209449
R37593 DVSS.n20280 DVSS.n20279 0.00209449
R37594 DVSS.n20269 DVSS.n20268 0.00209449
R37595 DVSS.n20786 DVSS.n20785 0.00209449
R37596 DVSS.n20775 DVSS.n20774 0.00209449
R37597 DVSS.n10805 DVSS.n10804 0.00209449
R37598 DVSS.n10801 DVSS.n10800 0.00209449
R37599 DVSS.n11577 DVSS.n11576 0.00209449
R37600 DVSS.n11588 DVSS.n11587 0.00209449
R37601 DVSS.n26 DVSS.n25 0.00209449
R37602 DVSS.n37 DVSS.n36 0.00209449
R37603 DVSS.n21519 DVSS.n21518 0.00209449
R37604 DVSS.n21508 DVSS.n21507 0.00209449
R37605 DVSS.n21431 DVSS.n21430 0.00209449
R37606 DVSS.n21420 DVSS.n21419 0.00209449
R37607 DVSS.n4686 DVSS.n4685 0.00209449
R37608 DVSS.n4678 DVSS.n4677 0.00209449
R37609 DVSS.n4308 DVSS.n4307 0.00209449
R37610 DVSS.n4316 DVSS.n4315 0.00209449
R37611 DVSS.n3479 DVSS.n3478 0.00209449
R37612 DVSS.n3471 DVSS.n3470 0.00209449
R37613 DVSS.n3368 DVSS.n3367 0.00209449
R37614 DVSS.n3363 DVSS.n3362 0.00209449
R37615 DVSS.n3304 DVSS.n3303 0.00209449
R37616 DVSS.n3101 DVSS.n3100 0.00209449
R37617 DVSS.n3083 DVSS.n3082 0.00209449
R37618 DVSS.n3060 DVSS.n3059 0.00209449
R37619 DVSS.n3055 DVSS.n3054 0.00209449
R37620 DVSS.n3054 DVSS.n3053 0.00209449
R37621 DVSS.n3045 DVSS.n3044 0.00209449
R37622 DVSS.n2786 DVSS.n2785 0.00209449
R37623 DVSS.n669 DVSS.n668 0.00209449
R37624 DVSS.n705 DVSS.n704 0.00209449
R37625 DVSS.n787 DVSS.n786 0.00209449
R37626 DVSS.n9985 DVSS.n9984 0.00209449
R37627 DVSS.n9655 DVSS.n9654 0.00209449
R37628 DVSS.n9644 DVSS.n9643 0.00209449
R37629 DVSS.n13239 DVSS.n13238 0.00209449
R37630 DVSS.n13245 DVSS.n13244 0.00209449
R37631 DVSS.n20450 DVSS.n20449 0.00209449
R37632 DVSS.n20461 DVSS.n20460 0.00209449
R37633 DVSS.n20554 DVSS.n20553 0.00209449
R37634 DVSS.n20543 DVSS.n20542 0.00209449
R37635 DVSS.n21012 DVSS.n21011 0.00209449
R37636 DVSS.n21001 DVSS.n21000 0.00209449
R37637 DVSS.n17382 DVSS.n17381 0.00209449
R37638 DVSS.n17390 DVSS.n17389 0.00209449
R37639 DVSS.n16172 DVSS.n16171 0.00209449
R37640 DVSS.n16163 DVSS.n16162 0.00209449
R37641 DVSS.n18769 DVSS.n18768 0.00209449
R37642 DVSS.n18775 DVSS.n18774 0.00209449
R37643 DVSS.n19442 DVSS.n19441 0.00209449
R37644 DVSS.n19450 DVSS.n19449 0.00209449
R37645 DVSS.n19537 DVSS.n19536 0.00209449
R37646 DVSS.n19529 DVSS.n19528 0.00209449
R37647 DVSS.n1236 DVSS.n1235 0.00209449
R37648 DVSS.n1228 DVSS.n1227 0.00209449
R37649 DVSS.n5458 DVSS.n5457 0.00209449
R37650 DVSS.n5463 DVSS.n5462 0.00209449
R37651 DVSS.n6622 DVSS.n6621 0.00209449
R37652 DVSS.n6631 DVSS.n6630 0.00209449
R37653 DVSS.n3541 DVSS.n3540 0.00209449
R37654 DVSS.n3533 DVSS.n3532 0.00209449
R37655 DVSS.n18985 DVSS.n18984 0.00209449
R37656 DVSS.n18977 DVSS.n18976 0.00209449
R37657 DVSS.n587 DVSS.n586 0.00209449
R37658 DVSS.n579 DVSS.n578 0.00209449
R37659 DVSS.n9208 DVSS.n9207 0.00209
R37660 DVSS.n7221 DVSS.n7220 0.00209
R37661 DVSS.n18881 DVSS.n18880 0.00209
R37662 DVSS.n14586 DVSS.n14585 0.00209
R37663 DVSS.n19100 DVSS.n19099 0.00209
R37664 DVSS.n19366 DVSS.n19365 0.00209
R37665 DVSS.n19844 DVSS.n19843 0.00209
R37666 DVSS.n837 DVSS.n836 0.00209
R37667 DVSS.n1124 DVSS.n1123 0.00209
R37668 DVSS.n281 DVSS.n280 0.00209
R37669 DVSS.n16092 DVSS.n16091 0.002075
R37670 DVSS.n16094 DVSS.n16093 0.002075
R37671 DVSS.n15433 DVSS.n15432 0.002075
R37672 DVSS.n18279 DVSS.n18278 0.002075
R37673 DVSS.n18328 DVSS.n18327 0.002075
R37674 DVSS.n18347 DVSS.n18346 0.002075
R37675 DVSS.n11989 DVSS.n80 0.00207333
R37676 DVSS.n20673 DVSS.n20672 0.00207333
R37677 DVSS.n21110 DVSS.n21107 0.00207333
R37678 DVSS.n5642 DVSS.n5641 0.00206274
R37679 DVSS.n5736 DVSS.n5735 0.00206274
R37680 DVSS.n4465 DVSS.n4464 0.00206274
R37681 DVSS.n7188 DVSS.n7187 0.00206274
R37682 DVSS.n19168 DVSS.n19153 0.00206274
R37683 DVSS.n869 DVSS.n868 0.00206274
R37684 DVSS.n4464 DVSS.n4463 0.00206274
R37685 DVSS.n5641 DVSS.n5640 0.00206274
R37686 DVSS.n10935 DVSS.n10934 0.00206274
R37687 DVSS.n11243 DVSS.n11242 0.00206274
R37688 DVSS.n11239 DVSS.n11238 0.00206274
R37689 DVSS.n9495 DVSS.n9494 0.00206274
R37690 DVSS.n12914 DVSS.n12913 0.00206274
R37691 DVSS.n12776 DVSS.n12775 0.00206274
R37692 DVSS.n12458 DVSS.n12457 0.00206274
R37693 DVSS.n12200 DVSS.n12199 0.00206274
R37694 DVSS.n21131 DVSS.n21130 0.00206274
R37695 DVSS.n9494 DVSS.n9493 0.00206274
R37696 DVSS.n10934 DVSS.n10933 0.00206274
R37697 DVSS.n11244 DVSS.n11243 0.00206274
R37698 DVSS.n11240 DVSS.n11239 0.00206274
R37699 DVSS.n5737 DVSS.n5736 0.00206274
R37700 DVSS.n19169 DVSS.n19168 0.00206274
R37701 DVSS.n17068 DVSS.n17067 0.00206274
R37702 DVSS.n17621 DVSS.n17620 0.00206274
R37703 DVSS.n17626 DVSS.n17625 0.00206274
R37704 DVSS.n15702 DVSS.n15701 0.00206274
R37705 DVSS.n13525 DVSS.n13524 0.00206274
R37706 DVSS.n20177 DVSS.n20176 0.00206274
R37707 DVSS.n20261 DVSS.n20260 0.00206274
R37708 DVSS.n20854 DVSS.n20853 0.00206274
R37709 DVSS.n15703 DVSS.n15702 0.00206274
R37710 DVSS.n17067 DVSS.n17066 0.00206274
R37711 DVSS.n17625 DVSS.n17624 0.00206274
R37712 DVSS.n17622 DVSS.n17621 0.00206274
R37713 DVSS.n20176 DVSS.n20164 0.00206274
R37714 DVSS.n7187 DVSS.n7180 0.00206274
R37715 DVSS.n13526 DVSS.n13525 0.00206274
R37716 DVSS.n10827 DVSS.n10826 0.00206274
R37717 DVSS.n11533 DVSS.n11532 0.00206274
R37718 DVSS.n12058 DVSS.n12057 0.00206274
R37719 DVSS.n70 DVSS.n69 0.00206274
R37720 DVSS.n21475 DVSS.n21474 0.00206274
R37721 DVSS.n11532 DVSS.n11531 0.00206274
R37722 DVSS.n10828 DVSS.n10827 0.00206274
R37723 DVSS.n4712 DVSS.n4711 0.00206274
R37724 DVSS.n4711 DVSS.n4710 0.00206274
R37725 DVSS.n4266 DVSS.n4265 0.00206274
R37726 DVSS.n3738 DVSS.n3737 0.00206274
R37727 DVSS.n3388 DVSS.n3387 0.00206274
R37728 DVSS.n3084 DVSS.n3083 0.00206274
R37729 DVSS.n2829 DVSS.n2828 0.00206274
R37730 DVSS.n2811 DVSS.n2810 0.00206274
R37731 DVSS.n4265 DVSS.n4264 0.00206274
R37732 DVSS.n9957 DVSS.n9956 0.00206274
R37733 DVSS.n11145 DVSS.n11144 0.00206274
R37734 DVSS.n11149 DVSS.n11148 0.00206274
R37735 DVSS.n9699 DVSS.n9698 0.00206274
R37736 DVSS.n13392 DVSS.n13391 0.00206274
R37737 DVSS.n20448 DVSS.n20447 0.00206274
R37738 DVSS.n20534 DVSS.n20533 0.00206274
R37739 DVSS.n21080 DVSS.n21079 0.00206274
R37740 DVSS.n13391 DVSS.n13390 0.00206274
R37741 DVSS.n9700 DVSS.n9699 0.00206274
R37742 DVSS.n11144 DVSS.n11143 0.00206274
R37743 DVSS.n9956 DVSS.n9955 0.00206274
R37744 DVSS.n11148 DVSS.n11147 0.00206274
R37745 DVSS.n20447 DVSS.n20435 0.00206274
R37746 DVSS.n17361 DVSS.n17360 0.00206274
R37747 DVSS.n16357 DVSS.n16356 0.00206274
R37748 DVSS.n16214 DVSS.n16213 0.00206274
R37749 DVSS.n18850 DVSS.n18849 0.00206274
R37750 DVSS.n19440 DVSS.n19439 0.00206274
R37751 DVSS.n19521 DVSS.n19520 0.00206274
R37752 DVSS.n1156 DVSS.n1155 0.00206274
R37753 DVSS.n16358 DVSS.n16357 0.00206274
R37754 DVSS.n18849 DVSS.n18848 0.00206274
R37755 DVSS.n16215 DVSS.n16214 0.00206274
R37756 DVSS.n17360 DVSS.n17359 0.00206274
R37757 DVSS.n19439 DVSS.n19427 0.00206274
R37758 DVSS.n5437 DVSS.n5436 0.00206274
R37759 DVSS.n6580 DVSS.n6579 0.00206274
R37760 DVSS.n3653 DVSS.n3652 0.00206274
R37761 DVSS.n18969 DVSS.n18968 0.00206274
R37762 DVSS.n547 DVSS.n546 0.00206274
R37763 DVSS.n6579 DVSS.n6578 0.00206274
R37764 DVSS.n5436 DVSS.n5435 0.00206274
R37765 DVSS.n12915 DVSS.n12914 0.00206274
R37766 DVSS.n12057 DVSS.n12056 0.00206274
R37767 DVSS.n3739 DVSS.n3738 0.00206274
R37768 DVSS.n3652 DVSS.n3651 0.00206274
R37769 DVSS.n3085 DVSS.n3084 0.00206274
R37770 DVSS.n12459 DVSS.n12458 0.00206274
R37771 DVSS.n19250 DVSS.n19249 0.00206274
R37772 DVSS.n12777 DVSS.n12776 0.00206274
R37773 DVSS.n69 DVSS.n68 0.00206274
R37774 DVSS.n20260 DVSS.n20259 0.00206274
R37775 DVSS.n20535 DVSS.n20534 0.00206274
R37776 DVSS.n3389 DVSS.n3388 0.00206274
R37777 DVSS.n18968 DVSS.n18967 0.00206274
R37778 DVSS.n2812 DVSS.n2811 0.00206274
R37779 DVSS.n12183 DVSS.n12182 0.00206274
R37780 DVSS.n21476 DVSS.n21475 0.00206274
R37781 DVSS.n21079 DVSS.n21078 0.00206274
R37782 DVSS.n20853 DVSS.n20852 0.00206274
R37783 DVSS.n1155 DVSS.n1154 0.00206274
R37784 DVSS.n868 DVSS.n867 0.00206274
R37785 DVSS.n546 DVSS.n545 0.00206274
R37786 DVSS.n2830 DVSS.n2829 0.00206274
R37787 DVSS.n715 DVSS.n714 0.00206274
R37788 DVSS.n21131 DVSS.n21129 0.00206274
R37789 DVSS.n13474 DVSS.n13473 0.00206
R37790 DVSS.n7920 DVSS.n7919 0.00206
R37791 DVSS.n20320 DVSS.n20319 0.00206
R37792 DVSS.n20605 DVSS.n20604 0.00206
R37793 DVSS.n20865 DVSS.n20864 0.00206
R37794 DVSS.n21091 DVSS.n21090 0.00206
R37795 DVSS.n16695 DVSS.n16694 0.00205609
R37796 DVSS.n16073 DVSS.n16072 0.00205609
R37797 DVSS.n18241 DVSS.n18240 0.00205609
R37798 DVSS.n18215 DVSS.n18214 0.00205609
R37799 DVSS.n19699 DVSS.n19698 0.00205609
R37800 DVSS.n19777 DVSS.n19776 0.00205609
R37801 DVSS.n130 DVSS.n129 0.00205609
R37802 DVSS.n218 DVSS.n217 0.00205609
R37803 DVSS.n202 DVSS.n201 0.00205609
R37804 DVSS.n18242 DVSS.n18241 0.00205609
R37805 DVSS.n18216 DVSS.n18215 0.00205609
R37806 DVSS.n18267 DVSS.n18266 0.00205609
R37807 DVSS.n18121 DVSS.n18120 0.00205609
R37808 DVSS.n16694 DVSS.n16693 0.00205609
R37809 DVSS.n17128 DVSS.n17127 0.00205609
R37810 DVSS.n15965 DVSS.n15964 0.00205609
R37811 DVSS.n15499 DVSS.n15498 0.00205609
R37812 DVSS.n15525 DVSS.n15524 0.00205609
R37813 DVSS.n19918 DVSS.n19917 0.00205609
R37814 DVSS.n20002 DVSS.n20001 0.00205609
R37815 DVSS.n290 DVSS.n289 0.00205609
R37816 DVSS.n426 DVSS.n425 0.00205609
R37817 DVSS.n410 DVSS.n409 0.00205609
R37818 DVSS.n15524 DVSS.n15523 0.00205609
R37819 DVSS.n15473 DVSS.n15472 0.00205609
R37820 DVSS.n15411 DVSS.n15410 0.00205609
R37821 DVSS.n15498 DVSS.n15497 0.00205609
R37822 DVSS.n17129 DVSS.n17128 0.00205609
R37823 DVSS.n19917 DVSS.n19916 0.00205609
R37824 DVSS.n19698 DVSS.n19697 0.00205609
R37825 DVSS.n19778 DVSS.n19777 0.00205609
R37826 DVSS.n20003 DVSS.n20002 0.00205609
R37827 DVSS.n289 DVSS.n288 0.00205609
R37828 DVSS.n129 DVSS.n128 0.00205609
R37829 DVSS.n219 DVSS.n218 0.00205609
R37830 DVSS.n427 DVSS.n426 0.00205609
R37831 DVSS.n411 DVSS.n410 0.00205609
R37832 DVSS.n203 DVSS.n202 0.00205609
R37833 DVSS.n10413 DVSS.n10412 0.0020493
R37834 DVSS.n10416 DVSS.n10415 0.0020493
R37835 DVSS.n10472 DVSS.n10471 0.0020493
R37836 DVSS.n10475 DVSS.n10474 0.0020493
R37837 DVSS.n10568 DVSS.n10563 0.0020493
R37838 DVSS.n10571 DVSS.n10570 0.0020493
R37839 DVSS.n4643 DVSS.n4639 0.00204286
R37840 DVSS.n4644 DVSS.n4638 0.00204286
R37841 DVSS.n4964 DVSS.n4963 0.00204286
R37842 DVSS.n4920 DVSS.n4919 0.00204286
R37843 DVSS.n4860 DVSS.n4859 0.00204286
R37844 DVSS.n4771 DVSS.n4770 0.00204286
R37845 DVSS.n4767 DVSS.n4766 0.00204286
R37846 DVSS.n6813 DVSS.n6808 0.00204286
R37847 DVSS.n3965 DVSS.n3930 0.00204286
R37848 DVSS.n6815 DVSS.n6814 0.00204286
R37849 DVSS.n3967 DVSS.n3966 0.00204286
R37850 DVSS.n3903 DVSS.n3902 0.00204286
R37851 DVSS.n3857 DVSS.n3856 0.00204286
R37852 DVSS.n8098 DVSS.n8097 0.00204286
R37853 DVSS.n8101 DVSS.n8100 0.00204286
R37854 DVSS.n3612 DVSS.n3608 0.00204286
R37855 DVSS.n2604 DVSS.n2597 0.00204286
R37856 DVSS.n3613 DVSS.n3607 0.00204286
R37857 DVSS.n2605 DVSS.n2596 0.00204286
R37858 DVSS.n2695 DVSS.n2694 0.00204286
R37859 DVSS.n2689 DVSS.n2688 0.00204286
R37860 DVSS.n2641 DVSS.n2640 0.00204286
R37861 DVSS.n2635 DVSS.n2634 0.00204286
R37862 DVSS.n11835 DVSS.n11834 0.00204286
R37863 DVSS.n11894 DVSS.n11893 0.00204286
R37864 DVSS.n5910 DVSS.n5872 0.00204286
R37865 DVSS.n6047 DVSS.n6046 0.00204286
R37866 DVSS.n5981 DVSS.n5980 0.00204286
R37867 DVSS.n5935 DVSS.n5934 0.00204286
R37868 DVSS.n8390 DVSS.n8389 0.00204286
R37869 DVSS.n8393 DVSS.n8392 0.00204286
R37870 DVSS.n6106 DVSS.n6101 0.00204286
R37871 DVSS.n6236 DVSS.n6235 0.00204286
R37872 DVSS.n6178 DVSS.n6177 0.00204286
R37873 DVSS.n8640 DVSS.n8639 0.00204286
R37874 DVSS.n8643 DVSS.n8642 0.00204286
R37875 DVSS.n6105 DVSS.n6102 0.00204286
R37876 DVSS.n3412 DVSS.n3394 0.00203846
R37877 DVSS.n12800 DVSS.n12799 0.00203846
R37878 DVSS.n934 DVSS.n933 0.00203846
R37879 DVSS.n21182 DVSS.n21181 0.00203846
R37880 DVSS.n5388 DVSS.n5387 0.00200838
R37881 DVSS.n10264 DVSS.n10263 0.00200838
R37882 DVSS.n10362 DVSS.n10360 0.00197887
R37883 DVSS.n5238 DVSS.n5237 0.00197887
R37884 DVSS.n5190 DVSS.n5189 0.00197887
R37885 DVSS.n5155 DVSS.n5154 0.00197887
R37886 DVSS.n5152 DVSS.n5151 0.00197887
R37887 DVSS.n5101 DVSS.n5100 0.00197887
R37888 DVSS.n5098 DVSS.n5097 0.00197887
R37889 DVSS.n10363 DVSS.n10358 0.00197887
R37890 DVSS.n16536 DVSS.n16535 0.00197887
R37891 DVSS.n16549 DVSS.n16548 0.00197887
R37892 DVSS.n16645 DVSS.n16644 0.00197887
R37893 DVSS.n17474 DVSS.n17473 0.00197887
R37894 DVSS.n16107 DVSS.n16106 0.00197887
R37895 DVSS.n17750 DVSS.n17749 0.00197887
R37896 DVSS.n17757 DVSS.n17756 0.00197887
R37897 DVSS.n17786 DVSS.n17785 0.00197887
R37898 DVSS.n18100 DVSS.n18099 0.00197887
R37899 DVSS.n18102 DVSS.n18101 0.00197887
R37900 DVSS.n18103 DVSS.n18102 0.00197887
R37901 DVSS.n18128 DVSS.n18127 0.00197887
R37902 DVSS.n18131 DVSS.n18130 0.00197887
R37903 DVSS.n18271 DVSS.n18270 0.00197887
R37904 DVSS.n18219 DVSS.n18218 0.00197887
R37905 DVSS.n18212 DVSS.n18211 0.00197887
R37906 DVSS.n18188 DVSS.n18187 0.00197887
R37907 DVSS.n18427 DVSS.n18426 0.00197887
R37908 DVSS.n18464 DVSS.n18463 0.00197887
R37909 DVSS.n14368 DVSS.n14367 0.00197887
R37910 DVSS.n14408 DVSS.n14407 0.00197887
R37911 DVSS.n14456 DVSS.n14455 0.00197887
R37912 DVSS.n19657 DVSS.n19656 0.00197887
R37913 DVSS.n157 DVSS.n156 0.00197887
R37914 DVSS.n16723 DVSS.n16722 0.00197887
R37915 DVSS.n16736 DVSS.n16735 0.00197887
R37916 DVSS.n17178 DVSS.n17177 0.00197887
R37917 DVSS.n16815 DVSS.n16814 0.00197887
R37918 DVSS.n15988 DVSS.n15987 0.00197887
R37919 DVSS.n15913 DVSS.n15912 0.00197887
R37920 DVSS.n15906 DVSS.n15905 0.00197887
R37921 DVSS.n15877 DVSS.n15876 0.00197887
R37922 DVSS.n15378 DVSS.n15377 0.00197887
R37923 DVSS.n15380 DVSS.n15379 0.00197887
R37924 DVSS.n15381 DVSS.n15380 0.00197887
R37925 DVSS.n15418 DVSS.n15417 0.00197887
R37926 DVSS.n15421 DVSS.n15420 0.00197887
R37927 DVSS.n15469 DVSS.n15468 0.00197887
R37928 DVSS.n15521 DVSS.n15520 0.00197887
R37929 DVSS.n15528 DVSS.n15527 0.00197887
R37930 DVSS.n15552 DVSS.n15551 0.00197887
R37931 DVSS.n15202 DVSS.n15201 0.00197887
R37932 DVSS.n15138 DVSS.n15137 0.00197887
R37933 DVSS.n14782 DVSS.n14781 0.00197887
R37934 DVSS.n14720 DVSS.n14719 0.00197887
R37935 DVSS.n14666 DVSS.n14665 0.00197887
R37936 DVSS.n19866 DVSS.n19865 0.00197887
R37937 DVSS.n317 DVSS.n316 0.00197887
R37938 DVSS.n4806 DVSS.n4805 0.00197857
R37939 DVSS.n4811 DVSS.n4810 0.00197857
R37940 DVSS.n4773 DVSS.n4772 0.00197857
R37941 DVSS.n8088 DVSS.n8087 0.00197857
R37942 DVSS.n8066 DVSS.n8065 0.00197857
R37943 DVSS.n8071 DVSS.n8070 0.00197857
R37944 DVSS.n8096 DVSS.n8095 0.00197857
R37945 DVSS.n11766 DVSS.n11765 0.00197857
R37946 DVSS.n11750 DVSS.n11749 0.00197857
R37947 DVSS.n11767 DVSS.n11764 0.00197857
R37948 DVSS.n8380 DVSS.n8379 0.00197857
R37949 DVSS.n8358 DVSS.n8357 0.00197857
R37950 DVSS.n8363 DVSS.n8362 0.00197857
R37951 DVSS.n8388 DVSS.n8387 0.00197857
R37952 DVSS.n8603 DVSS.n8602 0.00197857
R37953 DVSS.n8638 DVSS.n8637 0.00197857
R37954 DVSS.n8630 DVSS.n8629 0.00197857
R37955 DVSS.n6506 DVSS.n6505 0.0019742
R37956 DVSS.n4439 DVSS.n4438 0.0019742
R37957 DVSS.n4397 DVSS.n4396 0.0019742
R37958 DVSS.n19123 DVSS.n19122 0.0019742
R37959 DVSS.n19196 DVSS.n19195 0.0019742
R37960 DVSS.n19282 DVSS.n19281 0.0019742
R37961 DVSS.n855 DVSS.n854 0.0019742
R37962 DVSS.n1037 DVSS.n1036 0.0019742
R37963 DVSS.n996 DVSS.n995 0.0019742
R37964 DVSS.n4398 DVSS.n4397 0.0019742
R37965 DVSS.n4438 DVSS.n4437 0.0019742
R37966 DVSS.n9765 DVSS.n9764 0.0019742
R37967 DVSS.n9523 DVSS.n9522 0.0019742
R37968 DVSS.n9567 DVSS.n9566 0.0019742
R37969 DVSS.n12886 DVSS.n12885 0.0019742
R37970 DVSS.n12842 DVSS.n12841 0.0019742
R37971 DVSS.n21125 DVSS.n21124 0.0019742
R37972 DVSS.n9566 DVSS.n9565 0.0019742
R37973 DVSS.n9522 DVSS.n9521 0.0019742
R37974 DVSS.n9764 DVSS.n8926 0.0019742
R37975 DVSS.n6505 DVSS.n6504 0.0019742
R37976 DVSS.n15870 DVSS.n15869 0.0019742
R37977 DVSS.n15674 DVSS.n15673 0.0019742
R37978 DVSS.n15630 DVSS.n15629 0.0019742
R37979 DVSS.n20123 DVSS.n20122 0.0019742
R37980 DVSS.n20207 DVSS.n20206 0.0019742
R37981 DVSS.n20296 DVSS.n20295 0.0019742
R37982 DVSS.n20838 DVSS.n20837 0.0019742
R37983 DVSS.n20802 DVSS.n20801 0.0019742
R37984 DVSS.n20758 DVSS.n20757 0.0019742
R37985 DVSS.n15631 DVSS.n15630 0.0019742
R37986 DVSS.n15675 DVSS.n15674 0.0019742
R37987 DVSS.n15871 DVSS.n15870 0.0019742
R37988 DVSS.n11561 DVSS.n11560 0.0019742
R37989 DVSS.n11605 DVSS.n11604 0.0019742
R37990 DVSS.n12071 DVSS.n12070 0.0019742
R37991 DVSS.n54 DVSS.n53 0.0019742
R37992 DVSS.n21535 DVSS.n21534 0.0019742
R37993 DVSS.n21491 DVSS.n21490 0.0019742
R37994 DVSS.n21447 DVSS.n21446 0.0019742
R37995 DVSS.n21403 DVSS.n21402 0.0019742
R37996 DVSS.n11604 DVSS.n11603 0.0019742
R37997 DVSS.n11560 DVSS.n11559 0.0019742
R37998 DVSS.n4292 DVSS.n4291 0.0019742
R37999 DVSS.n4333 DVSS.n4332 0.0019742
R38000 DVSS.n3495 DVSS.n3494 0.0019742
R38001 DVSS.n3454 DVSS.n3453 0.0019742
R38002 DVSS.n717 DVSS.n716 0.0019742
R38003 DVSS.n4332 DVSS.n4331 0.0019742
R38004 DVSS.n4291 DVSS.n4290 0.0019742
R38005 DVSS.n9813 DVSS.n9812 0.0019742
R38006 DVSS.n9671 DVSS.n9670 0.0019742
R38007 DVSS.n9627 DVSS.n9626 0.0019742
R38008 DVSS.n20406 DVSS.n20405 0.0019742
R38009 DVSS.n20478 DVSS.n20477 0.0019742
R38010 DVSS.n20570 DVSS.n20569 0.0019742
R38011 DVSS.n21064 DVSS.n21063 0.0019742
R38012 DVSS.n21028 DVSS.n21027 0.0019742
R38013 DVSS.n20984 DVSS.n20983 0.0019742
R38014 DVSS.n9814 DVSS.n9813 0.0019742
R38015 DVSS.n9628 DVSS.n9627 0.0019742
R38016 DVSS.n9672 DVSS.n9671 0.0019742
R38017 DVSS.n16303 DVSS.n16302 0.0019742
R38018 DVSS.n16188 DVSS.n16187 0.0019742
R38019 DVSS.n16146 DVSS.n16145 0.0019742
R38020 DVSS.n19397 DVSS.n19396 0.0019742
R38021 DVSS.n19467 DVSS.n19466 0.0019742
R38022 DVSS.n19553 DVSS.n19552 0.0019742
R38023 DVSS.n1142 DVSS.n1141 0.0019742
R38024 DVSS.n1252 DVSS.n1251 0.0019742
R38025 DVSS.n1211 DVSS.n1210 0.0019742
R38026 DVSS.n16304 DVSS.n16303 0.0019742
R38027 DVSS.n16147 DVSS.n16146 0.0019742
R38028 DVSS.n16189 DVSS.n16188 0.0019742
R38029 DVSS.n6606 DVSS.n6605 0.0019742
R38030 DVSS.n6648 DVSS.n6647 0.0019742
R38031 DVSS.n3557 DVSS.n3556 0.0019742
R38032 DVSS.n18955 DVSS.n18954 0.0019742
R38033 DVSS.n19001 DVSS.n19000 0.0019742
R38034 DVSS.n533 DVSS.n532 0.0019742
R38035 DVSS.n603 DVSS.n602 0.0019742
R38036 DVSS.n562 DVSS.n561 0.0019742
R38037 DVSS.n6647 DVSS.n6646 0.0019742
R38038 DVSS.n6605 DVSS.n6604 0.0019742
R38039 DVSS.n18954 DVSS.n18953 0.0019742
R38040 DVSS.n3455 DVSS.n3454 0.0019742
R38041 DVSS.n19195 DVSS.n19194 0.0019742
R38042 DVSS.n19466 DVSS.n19465 0.0019742
R38043 DVSS.n20206 DVSS.n20205 0.0019742
R38044 DVSS.n20477 DVSS.n20476 0.0019742
R38045 DVSS.n12843 DVSS.n12842 0.0019742
R38046 DVSS.n53 DVSS.n52 0.0019742
R38047 DVSS.n12072 DVSS.n12071 0.0019742
R38048 DVSS.n12887 DVSS.n12886 0.0019742
R38049 DVSS.n20405 DVSS.n20404 0.0019742
R38050 DVSS.n20122 DVSS.n20121 0.0019742
R38051 DVSS.n19396 DVSS.n19395 0.0019742
R38052 DVSS.n19122 DVSS.n19121 0.0019742
R38053 DVSS.n3496 DVSS.n3495 0.0019742
R38054 DVSS.n3558 DVSS.n3557 0.0019742
R38055 DVSS.n532 DVSS.n531 0.0019742
R38056 DVSS.n1141 DVSS.n1140 0.0019742
R38057 DVSS.n21492 DVSS.n21491 0.0019742
R38058 DVSS.n854 DVSS.n853 0.0019742
R38059 DVSS.n21536 DVSS.n21535 0.0019742
R38060 DVSS.n20571 DVSS.n20570 0.0019742
R38061 DVSS.n20297 DVSS.n20296 0.0019742
R38062 DVSS.n19554 DVSS.n19553 0.0019742
R38063 DVSS.n19283 DVSS.n19282 0.0019742
R38064 DVSS.n19002 DVSS.n19001 0.0019742
R38065 DVSS.n21063 DVSS.n21062 0.0019742
R38066 DVSS.n20837 DVSS.n20836 0.0019742
R38067 DVSS.n563 DVSS.n562 0.0019742
R38068 DVSS.n678 DVSS.n677 0.0019742
R38069 DVSS.n1212 DVSS.n1211 0.0019742
R38070 DVSS.n21328 DVSS.n21327 0.0019742
R38071 DVSS.n21125 DVSS.n21123 0.0019742
R38072 DVSS.n21448 DVSS.n21447 0.0019742
R38073 DVSS.n21308 DVSS.n21307 0.0019742
R38074 DVSS.n21029 DVSS.n21028 0.0019742
R38075 DVSS.n20803 DVSS.n20802 0.0019742
R38076 DVSS.n1253 DVSS.n1252 0.0019742
R38077 DVSS.n1038 DVSS.n1037 0.0019742
R38078 DVSS.n672 DVSS.n671 0.0019742
R38079 DVSS.n604 DVSS.n603 0.0019742
R38080 DVSS.n21404 DVSS.n21403 0.0019742
R38081 DVSS.n20985 DVSS.n20984 0.0019742
R38082 DVSS.n20759 DVSS.n20758 0.0019742
R38083 DVSS.n997 DVSS.n996 0.0019742
R38084 DVSS.n20641 DVSS.n20640 0.00197
R38085 DVSS.n20082 DVSS.n20079 0.00196667
R38086 DVSS.n14162 DVSS.n14160 0.00195724
R38087 DVSS.n14741 DVSS.n14740 0.00195724
R38088 DVSS.n14160 DVSS.n14159 0.00195724
R38089 DVSS.n14742 DVSS.n14741 0.00195724
R38090 DVSS.n17755 DVSS.n17754 0.00195058
R38091 DVSS.n15908 DVSS.n15907 0.00195058
R38092 DVSS.n16666 DVSS.n16665 0.0019505
R38093 DVSS.n16706 DVSS.n16705 0.0019505
R38094 DVSS.n14517 DVSS.n14516 0.0019505
R38095 DVSS.n19807 DVSS.n19806 0.0019505
R38096 DVSS.n248 DVSS.n247 0.0019505
R38097 DVSS.n18233 DVSS.n18232 0.0019505
R38098 DVSS.n17117 DVSS.n17116 0.0019505
R38099 DVSS.n15507 DVSS.n15506 0.0019505
R38100 DVSS.n14614 DVSS.n14613 0.0019505
R38101 DVSS.n20032 DVSS.n20031 0.0019505
R38102 DVSS.n456 DVSS.n455 0.0019505
R38103 DVSS.n17157 DVSS.n17156 0.0019505
R38104 DVSS.n17116 DVSS.n17115 0.0019505
R38105 DVSS.n16707 DVSS.n16706 0.0019505
R38106 DVSS.n14518 DVSS.n14517 0.0019505
R38107 DVSS.n14615 DVSS.n14614 0.0019505
R38108 DVSS.n19808 DVSS.n19807 0.0019505
R38109 DVSS.n20033 DVSS.n20032 0.0019505
R38110 DVSS.n249 DVSS.n248 0.0019505
R38111 DVSS.n457 DVSS.n456 0.0019505
R38112 DVSS.n5696 DVSS.n5695 0.00191732
R38113 DVSS.n4441 DVSS.n4440 0.00191732
R38114 DVSS.n4395 DVSS.n4394 0.00191732
R38115 DVSS.n7093 DVSS.n7092 0.00191732
R38116 DVSS.n7147 DVSS.n7146 0.00191732
R38117 DVSS.n7178 DVSS.n7177 0.00191732
R38118 DVSS.n19120 DVSS.n19119 0.00191732
R38119 DVSS.n19149 DVSS.n19148 0.00191732
R38120 DVSS.n19153 DVSS.n19152 0.00191732
R38121 DVSS.n19198 DVSS.n19197 0.00191732
R38122 DVSS.n19247 DVSS.n19246 0.00191732
R38123 DVSS.n19285 DVSS.n19284 0.00191732
R38124 DVSS.n857 DVSS.n856 0.00191732
R38125 DVSS.n1040 DVSS.n1039 0.00191732
R38126 DVSS.n994 DVSS.n993 0.00191732
R38127 DVSS.n9520 DVSS.n9519 0.00191732
R38128 DVSS.n9569 DVSS.n9568 0.00191732
R38129 DVSS.n12889 DVSS.n12888 0.00191732
R38130 DVSS.n12840 DVSS.n12839 0.00191732
R38131 DVSS.n12833 DVSS.n12832 0.00191732
R38132 DVSS.n12731 DVSS.n12730 0.00191732
R38133 DVSS.n12700 DVSS.n12699 0.00191732
R38134 DVSS.n12493 DVSS.n12492 0.00191732
R38135 DVSS.n12448 DVSS.n12447 0.00191732
R38136 DVSS.n12427 DVSS.n12426 0.00191732
R38137 DVSS.n12209 DVSS.n12208 0.00191732
R38138 DVSS.n12174 DVSS.n12173 0.00191732
R38139 DVSS.n12156 DVSS.n12155 0.00191732
R38140 DVSS.n21223 DVSS.n21222 0.00191732
R38141 DVSS.n15677 DVSS.n15676 0.00191732
R38142 DVSS.n15628 DVSS.n15627 0.00191732
R38143 DVSS.n13590 DVSS.n13589 0.00191732
R38144 DVSS.n13546 DVSS.n13545 0.00191732
R38145 DVSS.n13529 DVSS.n13528 0.00191732
R38146 DVSS.n20120 DVSS.n20119 0.00191732
R38147 DVSS.n20160 DVSS.n20159 0.00191732
R38148 DVSS.n20164 DVSS.n20163 0.00191732
R38149 DVSS.n20209 DVSS.n20208 0.00191732
R38150 DVSS.n20257 DVSS.n20256 0.00191732
R38151 DVSS.n20299 DVSS.n20298 0.00191732
R38152 DVSS.n20840 DVSS.n20839 0.00191732
R38153 DVSS.n20805 DVSS.n20804 0.00191732
R38154 DVSS.n20756 DVSS.n20755 0.00191732
R38155 DVSS.n10794 DVSS.n10793 0.00191732
R38156 DVSS.n10791 DVSS.n10790 0.00191732
R38157 DVSS.n10790 DVSS.n10789 0.00191732
R38158 DVSS.n10782 DVSS.n10781 0.00191732
R38159 DVSS.n10780 DVSS.n10779 0.00191732
R38160 DVSS.n11558 DVSS.n11557 0.00191732
R38161 DVSS.n11607 DVSS.n11606 0.00191732
R38162 DVSS.n12074 DVSS.n12073 0.00191732
R38163 DVSS.n56 DVSS.n55 0.00191732
R38164 DVSS.n21538 DVSS.n21537 0.00191732
R38165 DVSS.n21489 DVSS.n21488 0.00191732
R38166 DVSS.n21450 DVSS.n21449 0.00191732
R38167 DVSS.n21401 DVSS.n21400 0.00191732
R38168 DVSS.n4653 DVSS.n4652 0.00191732
R38169 DVSS.n4289 DVSS.n4288 0.00191732
R38170 DVSS.n4335 DVSS.n4334 0.00191732
R38171 DVSS.n3498 DVSS.n3497 0.00191732
R38172 DVSS.n3452 DVSS.n3451 0.00191732
R38173 DVSS.n3445 DVSS.n3444 0.00191732
R38174 DVSS.n3353 DVSS.n3352 0.00191732
R38175 DVSS.n3323 DVSS.n3322 0.00191732
R38176 DVSS.n3117 DVSS.n3116 0.00191732
R38177 DVSS.n3075 DVSS.n3074 0.00191732
R38178 DVSS.n3053 DVSS.n3052 0.00191732
R38179 DVSS.n2839 DVSS.n2838 0.00191732
R38180 DVSS.n2802 DVSS.n2801 0.00191732
R38181 DVSS.n2784 DVSS.n2783 0.00191732
R38182 DVSS.n752 DVSS.n751 0.00191732
R38183 DVSS.n9674 DVSS.n9673 0.00191732
R38184 DVSS.n9625 DVSS.n9624 0.00191732
R38185 DVSS.n13242 DVSS.n13241 0.00191732
R38186 DVSS.n13368 DVSS.n13367 0.00191732
R38187 DVSS.n13388 DVSS.n13387 0.00191732
R38188 DVSS.n20403 DVSS.n20402 0.00191732
R38189 DVSS.n20431 DVSS.n20430 0.00191732
R38190 DVSS.n20435 DVSS.n20434 0.00191732
R38191 DVSS.n20480 DVSS.n20479 0.00191732
R38192 DVSS.n20531 DVSS.n20530 0.00191732
R38193 DVSS.n20573 DVSS.n20572 0.00191732
R38194 DVSS.n21066 DVSS.n21065 0.00191732
R38195 DVSS.n21031 DVSS.n21030 0.00191732
R38196 DVSS.n20982 DVSS.n20981 0.00191732
R38197 DVSS.n17415 DVSS.n17414 0.00191732
R38198 DVSS.n16191 DVSS.n16190 0.00191732
R38199 DVSS.n16144 DVSS.n16143 0.00191732
R38200 DVSS.n18772 DVSS.n18771 0.00191732
R38201 DVSS.n18829 DVSS.n18828 0.00191732
R38202 DVSS.n18846 DVSS.n18845 0.00191732
R38203 DVSS.n19394 DVSS.n19393 0.00191732
R38204 DVSS.n19423 DVSS.n19422 0.00191732
R38205 DVSS.n19427 DVSS.n19426 0.00191732
R38206 DVSS.n19469 DVSS.n19468 0.00191732
R38207 DVSS.n19518 DVSS.n19517 0.00191732
R38208 DVSS.n19556 DVSS.n19555 0.00191732
R38209 DVSS.n1144 DVSS.n1143 0.00191732
R38210 DVSS.n1255 DVSS.n1254 0.00191732
R38211 DVSS.n1209 DVSS.n1208 0.00191732
R38212 DVSS.n5470 DVSS.n5469 0.00191732
R38213 DVSS.n5473 DVSS.n5472 0.00191732
R38214 DVSS.n5474 DVSS.n5473 0.00191732
R38215 DVSS.n5482 DVSS.n5481 0.00191732
R38216 DVSS.n5484 DVSS.n5483 0.00191732
R38217 DVSS.n6603 DVSS.n6602 0.00191732
R38218 DVSS.n6650 DVSS.n6649 0.00191732
R38219 DVSS.n3560 DVSS.n3559 0.00191732
R38220 DVSS.n18957 DVSS.n18956 0.00191732
R38221 DVSS.n19004 DVSS.n19003 0.00191732
R38222 DVSS.n535 DVSS.n534 0.00191732
R38223 DVSS.n606 DVSS.n605 0.00191732
R38224 DVSS.n560 DVSS.n559 0.00191732
R38225 DVSS.n4959 DVSS.n4958 0.00191429
R38226 DVSS.n4915 DVSS.n4914 0.00191429
R38227 DVSS.n4855 DVSS.n4854 0.00191429
R38228 DVSS.n4785 DVSS.n4784 0.00191429
R38229 DVSS.n8085 DVSS.n8084 0.00191429
R38230 DVSS.n11842 DVSS.n11841 0.00191429
R38231 DVSS.n11845 DVSS.n11844 0.00191429
R38232 DVSS.n11901 DVSS.n11900 0.00191429
R38233 DVSS.n11904 DVSS.n11903 0.00191429
R38234 DVSS.n8377 DVSS.n8376 0.00191429
R38235 DVSS.n6232 DVSS.n6231 0.00191429
R38236 DVSS.n6174 DVSS.n6173 0.00191429
R38237 DVSS.n8626 DVSS.n8625 0.00191429
R38238 DVSS.n2049 DVSS.n2048 0.00191342
R38239 DVSS.n1726 DVSS.n1724 0.00191342
R38240 DVSS.n10059 DVSS.n10058 0.0019116
R38241 DVSS.n21566 DVSS 0.00191
R38242 DVSS.n5261 DVSS.n5260 0.00190845
R38243 DVSS.n10309 DVSS.n10308 0.00190845
R38244 DVSS.n10367 DVSS.n10366 0.00190845
R38245 DVSS.n2358 DVSS.n2357 0.00189982
R38246 DVSS.n2408 DVSS.n2407 0.00189982
R38247 DVSS.n2063 DVSS.n2062 0.00189982
R38248 DVSS.n2062 DVSS.n2061 0.00189982
R38249 DVSS.n2001 DVSS.n2000 0.00189982
R38250 DVSS.n2409 DVSS.n2408 0.00189982
R38251 DVSS.n2000 DVSS.n1999 0.00189982
R38252 DVSS.n4424 DVSS.n4423 0.00188565
R38253 DVSS.n4412 DVSS.n4411 0.00188565
R38254 DVSS.n19182 DVSS.n19181 0.00188565
R38255 DVSS.n19268 DVSS.n19267 0.00188565
R38256 DVSS.n841 DVSS.n840 0.00188565
R38257 DVSS.n1023 DVSS.n1022 0.00188565
R38258 DVSS.n1010 DVSS.n1009 0.00188565
R38259 DVSS.n4411 DVSS.n4410 0.00188565
R38260 DVSS.n4425 DVSS.n4424 0.00188565
R38261 DVSS.n9537 DVSS.n9536 0.00188565
R38262 DVSS.n9553 DVSS.n9552 0.00188565
R38263 DVSS.n12873 DVSS.n12872 0.00188565
R38264 DVSS.n12856 DVSS.n12855 0.00188565
R38265 DVSS.n12692 DVSS.n12691 0.00188565
R38266 DVSS.n12482 DVSS.n12481 0.00188565
R38267 DVSS.n12452 DVSS.n12451 0.00188565
R38268 DVSS.n12449 DVSS.n12448 0.00188565
R38269 DVSS.n21241 DVSS.n21240 0.00188565
R38270 DVSS.n9536 DVSS.n9535 0.00188565
R38271 DVSS.n9552 DVSS.n9551 0.00188565
R38272 DVSS.n15660 DVSS.n15659 0.00188565
R38273 DVSS.n15644 DVSS.n15643 0.00188565
R38274 DVSS.n20193 DVSS.n20192 0.00188565
R38275 DVSS.n20282 DVSS.n20281 0.00188565
R38276 DVSS.n20824 DVSS.n20823 0.00188565
R38277 DVSS.n20788 DVSS.n20787 0.00188565
R38278 DVSS.n20772 DVSS.n20771 0.00188565
R38279 DVSS.n15661 DVSS.n15660 0.00188565
R38280 DVSS.n15645 DVSS.n15644 0.00188565
R38281 DVSS.n10788 DVSS.n10787 0.00188565
R38282 DVSS.n10736 DVSS.n10735 0.00188565
R38283 DVSS.n11410 DVSS.n11409 0.00188565
R38284 DVSS.n11575 DVSS.n11574 0.00188565
R38285 DVSS.n11591 DVSS.n11590 0.00188565
R38286 DVSS.n23 DVSS.n22 0.00188565
R38287 DVSS.n40 DVSS.n39 0.00188565
R38288 DVSS.n21521 DVSS.n21520 0.00188565
R38289 DVSS.n21505 DVSS.n21504 0.00188565
R38290 DVSS.n21433 DVSS.n21432 0.00188565
R38291 DVSS.n21417 DVSS.n21416 0.00188565
R38292 DVSS.n11574 DVSS.n11573 0.00188565
R38293 DVSS.n11590 DVSS.n11589 0.00188565
R38294 DVSS.n10735 DVSS.n10734 0.00188565
R38295 DVSS.n11409 DVSS.n11408 0.00188565
R38296 DVSS.n10789 DVSS.n10788 0.00188565
R38297 DVSS.n4306 DVSS.n4305 0.00188565
R38298 DVSS.n4319 DVSS.n4318 0.00188565
R38299 DVSS.n3482 DVSS.n3481 0.00188565
R38300 DVSS.n3468 DVSS.n3467 0.00188565
R38301 DVSS.n3315 DVSS.n3314 0.00188565
R38302 DVSS.n3078 DVSS.n3077 0.00188565
R38303 DVSS.n3076 DVSS.n3075 0.00188565
R38304 DVSS.n772 DVSS.n771 0.00188565
R38305 DVSS.n804 DVSS.n799 0.00188565
R38306 DVSS.n4305 DVSS.n4304 0.00188565
R38307 DVSS.n4318 DVSS.n4317 0.00188565
R38308 DVSS.n9657 DVSS.n9656 0.00188565
R38309 DVSS.n9641 DVSS.n9640 0.00188565
R38310 DVSS.n20464 DVSS.n20463 0.00188565
R38311 DVSS.n20556 DVSS.n20555 0.00188565
R38312 DVSS.n21050 DVSS.n21049 0.00188565
R38313 DVSS.n21014 DVSS.n21013 0.00188565
R38314 DVSS.n20998 DVSS.n20997 0.00188565
R38315 DVSS.n9658 DVSS.n9657 0.00188565
R38316 DVSS.n9642 DVSS.n9641 0.00188565
R38317 DVSS.n16174 DVSS.n16173 0.00188565
R38318 DVSS.n16160 DVSS.n16159 0.00188565
R38319 DVSS.n19453 DVSS.n19452 0.00188565
R38320 DVSS.n19539 DVSS.n19538 0.00188565
R38321 DVSS.n1128 DVSS.n1127 0.00188565
R38322 DVSS.n1238 DVSS.n1237 0.00188565
R38323 DVSS.n1225 DVSS.n1224 0.00188565
R38324 DVSS.n16175 DVSS.n16174 0.00188565
R38325 DVSS.n16161 DVSS.n16160 0.00188565
R38326 DVSS.n5476 DVSS.n5475 0.00188565
R38327 DVSS.n5858 DVSS.n5857 0.00188565
R38328 DVSS.n6333 DVSS.n6332 0.00188565
R38329 DVSS.n6620 DVSS.n6619 0.00188565
R38330 DVSS.n6634 DVSS.n6633 0.00188565
R38331 DVSS.n3543 DVSS.n3542 0.00188565
R38332 DVSS.n18941 DVSS.n18940 0.00188565
R38333 DVSS.n18987 DVSS.n18986 0.00188565
R38334 DVSS.n519 DVSS.n518 0.00188565
R38335 DVSS.n589 DVSS.n588 0.00188565
R38336 DVSS.n576 DVSS.n575 0.00188565
R38337 DVSS.n6619 DVSS.n6618 0.00188565
R38338 DVSS.n6332 DVSS.n6331 0.00188565
R38339 DVSS.n6633 DVSS.n6632 0.00188565
R38340 DVSS.n5857 DVSS.n5856 0.00188565
R38341 DVSS.n5475 DVSS.n5474 0.00188565
R38342 DVSS.n3544 DVSS.n3543 0.00188565
R38343 DVSS.n39 DVSS.n38 0.00188565
R38344 DVSS.n12857 DVSS.n12856 0.00188565
R38345 DVSS.n20463 DVSS.n20462 0.00188565
R38346 DVSS.n20192 DVSS.n20191 0.00188565
R38347 DVSS.n19452 DVSS.n19451 0.00188565
R38348 DVSS.n19181 DVSS.n19180 0.00188565
R38349 DVSS.n3469 DVSS.n3468 0.00188565
R38350 DVSS.n18940 DVSS.n18939 0.00188565
R38351 DVSS.n24 DVSS.n23 0.00188565
R38352 DVSS.n12872 DVSS.n12871 0.00188565
R38353 DVSS.n3481 DVSS.n3480 0.00188565
R38354 DVSS.n18988 DVSS.n18987 0.00188565
R38355 DVSS.n3316 DVSS.n3315 0.00188565
R38356 DVSS.n3108 DVSS.n3107 0.00188565
R38357 DVSS.n19540 DVSS.n19539 0.00188565
R38358 DVSS.n12693 DVSS.n12692 0.00188565
R38359 DVSS.n12483 DVSS.n12482 0.00188565
R38360 DVSS.n21522 DVSS.n21521 0.00188565
R38361 DVSS.n19269 DVSS.n19268 0.00188565
R38362 DVSS.n21506 DVSS.n21505 0.00188565
R38363 DVSS.n12450 DVSS.n12449 0.00188565
R38364 DVSS.n12451 DVSS.n12450 0.00188565
R38365 DVSS.n21049 DVSS.n21048 0.00188565
R38366 DVSS.n20823 DVSS.n20822 0.00188565
R38367 DVSS.n1127 DVSS.n1126 0.00188565
R38368 DVSS.n840 DVSS.n839 0.00188565
R38369 DVSS.n518 DVSS.n517 0.00188565
R38370 DVSS.n20557 DVSS.n20556 0.00188565
R38371 DVSS.n20283 DVSS.n20282 0.00188565
R38372 DVSS.n590 DVSS.n589 0.00188565
R38373 DVSS.n1239 DVSS.n1238 0.00188565
R38374 DVSS.n21434 DVSS.n21433 0.00188565
R38375 DVSS.n1024 DVSS.n1023 0.00188565
R38376 DVSS.n772 DVSS.n769 0.00188565
R38377 DVSS.n21418 DVSS.n21417 0.00188565
R38378 DVSS.n21128 DVSS.n21127 0.00188565
R38379 DVSS.n20999 DVSS.n20998 0.00188565
R38380 DVSS.n20773 DVSS.n20772 0.00188565
R38381 DVSS.n1226 DVSS.n1225 0.00188565
R38382 DVSS.n1011 DVSS.n1010 0.00188565
R38383 DVSS.n799 DVSS.n798 0.00188565
R38384 DVSS.n577 DVSS.n576 0.00188565
R38385 DVSS.n21015 DVSS.n21014 0.00188565
R38386 DVSS.n20789 DVSS.n20788 0.00188565
R38387 DVSS.n2010 DVSS.n2009 0.00187029
R38388 DVSS.n2459 DVSS.n1903 0.00187029
R38389 DVSS.n4952 DVSS.n4951 0.00186769
R38390 DVSS.n4951 DVSS.n4950 0.00186769
R38391 DVSS.n4947 DVSS.n4946 0.00186769
R38392 DVSS.n4944 DVSS.n4943 0.00186769
R38393 DVSS.n4849 DVSS.n4848 0.00186769
R38394 DVSS.n4847 DVSS.n4846 0.00186769
R38395 DVSS.n4843 DVSS.n4842 0.00186769
R38396 DVSS.n4841 DVSS.n4840 0.00186769
R38397 DVSS.n10125 DVSS.n10124 0.00186769
R38398 DVSS.n10131 DVSS.n10130 0.00186769
R38399 DVSS.n10134 DVSS.n10133 0.00186769
R38400 DVSS.n6272 DVSS.n6271 0.00186769
R38401 DVSS.n6225 DVSS.n6224 0.00186769
R38402 DVSS.n6224 DVSS.n6223 0.00186769
R38403 DVSS.n6219 DVSS.n6218 0.00186769
R38404 DVSS.n6218 DVSS.n6217 0.00186769
R38405 DVSS.n6168 DVSS.n6167 0.00186769
R38406 DVSS.n6165 DVSS.n6164 0.00186769
R38407 DVSS.n6161 DVSS.n6160 0.00186769
R38408 DVSS.n6159 DVSS.n6158 0.00186769
R38409 DVSS.n8695 DVSS.n8694 0.00186769
R38410 DVSS.n8701 DVSS.n8700 0.00186769
R38411 DVSS.n8756 DVSS.n8755 0.00186769
R38412 DVSS.n8763 DVSS.n8762 0.00186769
R38413 DVSS.n6220 DVSS.n6219 0.00186769
R38414 DVSS.n6223 DVSS.n6222 0.00186769
R38415 DVSS.n6217 DVSS.n6216 0.00186769
R38416 DVSS.n6226 DVSS.n6225 0.00186769
R38417 DVSS.n8702 DVSS.n8701 0.00186769
R38418 DVSS.n8694 DVSS.n8693 0.00186769
R38419 DVSS.n4946 DVSS.n4945 0.00186769
R38420 DVSS.n4953 DVSS.n4952 0.00186769
R38421 DVSS.n4945 DVSS.n4944 0.00186769
R38422 DVSS.n4950 DVSS.n4949 0.00186769
R38423 DVSS.n6273 DVSS.n6272 0.00186769
R38424 DVSS.n8755 DVSS.n8754 0.00186769
R38425 DVSS.n8762 DVSS.n8761 0.00186769
R38426 DVSS.n10133 DVSS.n10132 0.00186769
R38427 DVSS.n10124 DVSS.n10123 0.00186769
R38428 DVSS.n10132 DVSS.n10131 0.00186769
R38429 DVSS.n6166 DVSS.n6165 0.00186769
R38430 DVSS.n6162 DVSS.n6161 0.00186769
R38431 DVSS.n4842 DVSS.n4841 0.00186769
R38432 DVSS.n4850 DVSS.n4849 0.00186769
R38433 DVSS.n4848 DVSS.n4847 0.00186769
R38434 DVSS.n4840 DVSS.n4839 0.00186769
R38435 DVSS.n6167 DVSS.n6166 0.00186769
R38436 DVSS.n6160 DVSS.n6159 0.00186769
R38437 DVSS.n4908 DVSS.n4907 0.00186769
R38438 DVSS.n4906 DVSS.n4905 0.00186769
R38439 DVSS.n4902 DVSS.n4901 0.00186769
R38440 DVSS.n4900 DVSS.n4899 0.00186769
R38441 DVSS.n10068 DVSS.n10067 0.00186769
R38442 DVSS.n10070 DVSS.n10069 0.00186769
R38443 DVSS.n10173 DVSS.n10172 0.00186769
R38444 DVSS.n10180 DVSS.n10179 0.00186769
R38445 DVSS.n10182 DVSS.n10181 0.00186769
R38446 DVSS.n4909 DVSS.n4908 0.00186769
R38447 DVSS.n4903 DVSS.n4902 0.00186769
R38448 DVSS.n10179 DVSS.n10178 0.00186769
R38449 DVSS.n6268 DVSS.n6267 0.00186769
R38450 DVSS.n6263 DVSS.n6262 0.00186769
R38451 DVSS.n8700 DVSS.n8699 0.00186769
R38452 DVSS.n8765 DVSS.n8764 0.00186769
R38453 DVSS.n8800 DVSS.n8799 0.00186769
R38454 DVSS.n8925 DVSS.n8863 0.00186769
R38455 DVSS.n8924 DVSS.n8923 0.00186769
R38456 DVSS.n8801 DVSS.n8800 0.00186769
R38457 DVSS.n8925 DVSS.n8924 0.00186769
R38458 DVSS.n8863 DVSS.n8862 0.00186769
R38459 DVSS.n8699 DVSS.n8698 0.00186769
R38460 DVSS.n10067 DVSS.n10066 0.00186769
R38461 DVSS.n10069 DVSS.n10068 0.00186769
R38462 DVSS.n10181 DVSS.n10180 0.00186769
R38463 DVSS.n10172 DVSS.n10171 0.00186769
R38464 DVSS.n4901 DVSS.n4900 0.00186769
R38465 DVSS.n4907 DVSS.n4906 0.00186769
R38466 DVSS.n6271 DVSS.n6268 0.00186769
R38467 DVSS.n6264 DVSS.n6263 0.00186769
R38468 DVSS.n8764 DVSS.n8763 0.00186769
R38469 DVSS.n2009 DVSS.n2008 0.00186509
R38470 DVSS.n1903 DVSS.n1902 0.00186509
R38471 DVSS.n19597 DVSS.n19594 0.00186
R38472 DVSS.n21237 DVSS.n21233 0.00185432
R38473 DVSS.n17211 DVSS.n17210 0.00185
R38474 DVSS.n15152 DVSS.n15151 0.00185
R38475 DVSS.n15110 DVSS.n15109 0.00185
R38476 DVSS.n2369 DVSS.n2368 0.00185
R38477 DVSS.n2396 DVSS.n2395 0.00185
R38478 DVSS.n17689 DVSS.n17688 0.00185
R38479 DVSS.n4751 DVSS.n4749 0.00185
R38480 DVSS.n4789 DVSS.n4788 0.00185
R38481 DVSS.n4746 DVSS.n4745 0.00185
R38482 DVSS.n8114 DVSS.n8112 0.00185
R38483 DVSS.n8082 DVSS.n8081 0.00185
R38484 DVSS.n8115 DVSS.n8110 0.00185
R38485 DVSS.n8118 DVSS.n8117 0.00185
R38486 DVSS.n11791 DVSS.n11789 0.00185
R38487 DVSS.n2699 DVSS.n2698 0.00185
R38488 DVSS.n2696 DVSS.n2695 0.00185
R38489 DVSS.n2645 DVSS.n2644 0.00185
R38490 DVSS.n2642 DVSS.n2641 0.00185
R38491 DVSS.n11792 DVSS.n11787 0.00185
R38492 DVSS.n8406 DVSS.n8404 0.00185
R38493 DVSS.n8374 DVSS.n8373 0.00185
R38494 DVSS.n8407 DVSS.n8402 0.00185
R38495 DVSS.n8410 DVSS.n8409 0.00185
R38496 DVSS.n8623 DVSS.n8622 0.00185
R38497 DVSS.n8663 DVSS.n8662 0.00185
R38498 DVSS.n8659 DVSS.n8657 0.00185
R38499 DVSS.n14912 DVSS.n14911 0.00185
R38500 DVSS DVSS.n21366 0.00184667
R38501 DVSS.n12546 DVSS.n12541 0.00184615
R38502 DVSS.n12670 DVSS.n12665 0.00184615
R38503 DVSS.n12578 DVSS.n12573 0.00184615
R38504 DVSS.n12382 DVSS.n12377 0.00184615
R38505 DVSS.n12290 DVSS.n12285 0.00184615
R38506 DVSS.n12251 DVSS.n12250 0.00184615
R38507 DVSS.n3170 DVSS.n3165 0.00184615
R38508 DVSS.n3294 DVSS.n3289 0.00184615
R38509 DVSS.n3202 DVSS.n3197 0.00184615
R38510 DVSS.n3009 DVSS.n3004 0.00184615
R38511 DVSS.n2917 DVSS.n2912 0.00184615
R38512 DVSS.n2878 DVSS.n2877 0.00184615
R38513 DVSS.n16673 DVSS.n16672 0.00184491
R38514 DVSS.n16114 DVSS.n16113 0.00184491
R38515 DVSS.n18448 DVSS.n18447 0.00184491
R38516 DVSS.n14382 DVSS.n14381 0.00184491
R38517 DVSS.n16115 DVSS.n16114 0.00184491
R38518 DVSS.n18240 DVSS.n18239 0.00184491
R38519 DVSS.n18429 DVSS.n18428 0.00184491
R38520 DVSS.n18447 DVSS.n18446 0.00184491
R38521 DVSS.n14381 DVSS.n14380 0.00184491
R38522 DVSS.n15995 DVSS.n15994 0.00184491
R38523 DVSS.n15500 DVSS.n15499 0.00184491
R38524 DVSS.n15200 DVSS.n15199 0.00184491
R38525 DVSS.n15169 DVSS.n15168 0.00184491
R38526 DVSS.n14768 DVSS.n14767 0.00184491
R38527 DVSS.n15996 DVSS.n15995 0.00184491
R38528 DVSS.n15170 DVSS.n15169 0.00184491
R38529 DVSS.n17150 DVSS.n17149 0.00184491
R38530 DVSS.n14769 DVSS.n14768 0.00184491
R38531 DVSS.n19749 DVSS.n19748 0.00184491
R38532 DVSS.n19975 DVSS.n19974 0.00184491
R38533 DVSS.n19750 DVSS.n19749 0.00184491
R38534 DVSS.n19974 DVSS.n19973 0.00184491
R38535 DVSS.n10330 DVSS.n10329 0.00183803
R38536 DVSS.n10345 DVSS.n10344 0.00183803
R38537 DVSS.n10349 DVSS.n10348 0.00183803
R38538 DVSS.n10593 DVSS.n10592 0.00183803
R38539 DVSS.n10596 DVSS.n10595 0.00183803
R38540 DVSS.n10139 DVSS.n10138 0.00183556
R38541 DVSS.n10191 DVSS.n10190 0.00183556
R38542 DVSS.n10192 DVSS.n10191 0.00183556
R38543 DVSS.n10140 DVSS.n10139 0.00183556
R38544 DVSS.n19303 DVSS.n19302 0.00182
R38545 DVSS.n19372 DVSS.n19371 0.00182
R38546 DVSS.n12015 DVSS 0.00180667
R38547 DVSS.n5676 DVSS.n5675 0.0017971
R38548 DVSS.n4452 DVSS.n4451 0.0017971
R38549 DVSS.n7210 DVSS.n7209 0.0017971
R38550 DVSS.n19297 DVSS.n19296 0.0017971
R38551 DVSS.n1051 DVSS.n1050 0.0017971
R38552 DVSS.n4453 DVSS.n4452 0.0017971
R38553 DVSS.n5675 DVSS.n5674 0.0017971
R38554 DVSS.n10967 DVSS.n10966 0.0017971
R38555 DVSS.n9507 DVSS.n9506 0.0017971
R38556 DVSS.n12902 DVSS.n12901 0.0017971
R38557 DVSS.n12727 DVSS.n12726 0.0017971
R38558 DVSS.n12414 DVSS.n12413 0.0017971
R38559 DVSS.n12181 DVSS.n12180 0.0017971
R38560 DVSS.n9506 DVSS.n9505 0.0017971
R38561 DVSS.n10966 DVSS.n10965 0.0017971
R38562 DVSS.n17100 DVSS.n17099 0.0017971
R38563 DVSS.n15690 DVSS.n15689 0.0017971
R38564 DVSS.n13513 DVSS.n13512 0.0017971
R38565 DVSS.n20312 DVSS.n20311 0.0017971
R38566 DVSS.n20818 DVSS.n20817 0.0017971
R38567 DVSS.n15691 DVSS.n15690 0.0017971
R38568 DVSS.n17099 DVSS.n17098 0.0017971
R38569 DVSS.n11423 DVSS.n11422 0.0017971
R38570 DVSS.n11545 DVSS.n11544 0.0017971
R38571 DVSS.n12087 DVSS.n12086 0.0017971
R38572 DVSS.n21551 DVSS.n21550 0.0017971
R38573 DVSS.n21463 DVSS.n21462 0.0017971
R38574 DVSS.n11544 DVSS.n11543 0.0017971
R38575 DVSS.n11422 DVSS.n11421 0.0017971
R38576 DVSS.n4673 DVSS.n4672 0.0017971
R38577 DVSS.n4674 DVSS.n4673 0.0017971
R38578 DVSS.n4278 DVSS.n4277 0.0017971
R38579 DVSS.n3509 DVSS.n3508 0.0017971
R38580 DVSS.n3041 DVSS.n3040 0.0017971
R38581 DVSS.n2809 DVSS.n2808 0.0017971
R38582 DVSS.n4277 DVSS.n4276 0.0017971
R38583 DVSS.n9989 DVSS.n9988 0.0017971
R38584 DVSS.n9687 DVSS.n9686 0.0017971
R38585 DVSS.n13415 DVSS.n13414 0.0017971
R38586 DVSS.n20586 DVSS.n20585 0.0017971
R38587 DVSS.n21044 DVSS.n21043 0.0017971
R38588 DVSS.n9688 DVSS.n9687 0.0017971
R38589 DVSS.n9988 DVSS.n9987 0.0017971
R38590 DVSS.n17395 DVSS.n17394 0.0017971
R38591 DVSS.n16202 DVSS.n16201 0.0017971
R38592 DVSS.n18870 DVSS.n18869 0.0017971
R38593 DVSS.n19568 DVSS.n19567 0.0017971
R38594 DVSS.n1266 DVSS.n1265 0.0017971
R38595 DVSS.n16203 DVSS.n16202 0.0017971
R38596 DVSS.n17394 DVSS.n17393 0.0017971
R38597 DVSS.n6345 DVSS.n6344 0.0017971
R38598 DVSS.n6592 DVSS.n6591 0.0017971
R38599 DVSS.n3571 DVSS.n3570 0.0017971
R38600 DVSS.n19015 DVSS.n19014 0.0017971
R38601 DVSS.n617 DVSS.n616 0.0017971
R38602 DVSS.n6591 DVSS.n6590 0.0017971
R38603 DVSS.n6344 DVSS.n6343 0.0017971
R38604 DVSS.n3572 DVSS.n3571 0.0017971
R38605 DVSS.n12088 DVSS.n12087 0.0017971
R38606 DVSS.n3510 DVSS.n3509 0.0017971
R38607 DVSS.n12903 DVSS.n12902 0.0017971
R38608 DVSS.n18871 DVSS.n18870 0.0017971
R38609 DVSS.n7211 DVSS.n7210 0.0017971
R38610 DVSS.n13416 DVSS.n13415 0.0017971
R38611 DVSS.n13514 DVSS.n13513 0.0017971
R38612 DVSS.n19016 DVSS.n19015 0.0017971
R38613 DVSS.n3350 DVSS.n3349 0.0017971
R38614 DVSS.n12728 DVSS.n12727 0.0017971
R38615 DVSS.n3040 DVSS.n3039 0.0017971
R38616 DVSS.n12413 DVSS.n12412 0.0017971
R38617 DVSS.n21552 DVSS.n21551 0.0017971
R38618 DVSS.n19296 DVSS.n19295 0.0017971
R38619 DVSS.n19567 DVSS.n19566 0.0017971
R38620 DVSS.n20313 DVSS.n20312 0.0017971
R38621 DVSS.n20587 DVSS.n20586 0.0017971
R38622 DVSS.n618 DVSS.n617 0.0017971
R38623 DVSS.n2810 DVSS.n2809 0.0017971
R38624 DVSS.n1267 DVSS.n1266 0.0017971
R38625 DVSS.n21464 DVSS.n21463 0.0017971
R38626 DVSS.n1052 DVSS.n1051 0.0017971
R38627 DVSS.n21045 DVSS.n21044 0.0017971
R38628 DVSS.n20819 DVSS.n20818 0.0017971
R38629 DVSS.n13491 DVSS.n13490 0.00179
R38630 DVSS.n7937 DVSS.n7936 0.00179
R38631 DVSS.n20107 DVSS.n20106 0.00179
R38632 DVSS.n20593 DVSS.n20592 0.00179
R38633 DVSS.n20702 DVSS.n20701 0.00179
R38634 DVSS.n20931 DVSS.n20930 0.00179
R38635 DVSS.n4988 DVSS.n4987 0.00178571
R38636 DVSS.n11744 DVSS.n11743 0.00178571
R38637 DVSS.n11763 DVSS.n11762 0.00178571
R38638 DVSS.n11776 DVSS.n11775 0.00178571
R38639 DVSS.n11796 DVSS.n11795 0.00178571
R38640 DVSS.n6038 DVSS.n6037 0.00178571
R38641 DVSS.n6286 DVSS.n6285 0.00178571
R38642 DVSS.n10575 DVSS.n10574 0.00176761
R38643 DVSS.n10867 DVSS.n10866 0.00176761
R38644 DVSS.n10326 DVSS.n10325 0.00176761
R38645 DVSS.n10335 DVSS.n10332 0.00176761
R38646 DVSS.n10422 DVSS.n10421 0.00176761
R38647 DVSS.n10481 DVSS.n10480 0.00176761
R38648 DVSS.n10577 DVSS.n10576 0.00176761
R38649 DVSS.n10868 DVSS.n10864 0.00176761
R38650 DVSS.n16525 DVSS.n16524 0.00176761
R38651 DVSS.n16079 DVSS.n16078 0.00176761
R38652 DVSS.n17745 DVSS.n17744 0.00176761
R38653 DVSS.n18099 DVSS.n18098 0.00176761
R38654 DVSS.n18110 DVSS.n18109 0.00176761
R38655 DVSS.n18206 DVSS.n18205 0.00176761
R38656 DVSS.n18456 DVSS.n18455 0.00176761
R38657 DVSS.n18481 DVSS.n18480 0.00176761
R38658 DVSS.n18491 DVSS.n18490 0.00176761
R38659 DVSS.n14386 DVSS.n14385 0.00176761
R38660 DVSS.n14405 DVSS.n14404 0.00176761
R38661 DVSS.n14415 DVSS.n14414 0.00176761
R38662 DVSS.n19669 DVSS.n19668 0.00176761
R38663 DVSS.n16712 DVSS.n16711 0.00176761
R38664 DVSS.n15971 DVSS.n15970 0.00176761
R38665 DVSS.n15918 DVSS.n15917 0.00176761
R38666 DVSS.n15377 DVSS.n15376 0.00176761
R38667 DVSS.n15388 DVSS.n15387 0.00176761
R38668 DVSS.n15534 DVSS.n15533 0.00176761
R38669 DVSS.n15161 DVSS.n15160 0.00176761
R38670 DVSS.n15121 DVSS.n15120 0.00176761
R38671 DVSS.n7732 DVSS.n7731 0.00176761
R38672 DVSS.n14764 DVSS.n14763 0.00176761
R38673 DVSS.n14723 DVSS.n14722 0.00176761
R38674 DVSS.n14713 DVSS.n14712 0.00176761
R38675 DVSS.n19884 DVSS.n19883 0.00176761
R38676 DVSS.n3702 DVSS.n3701 0.00175333
R38677 DVSS.n19087 DVSS.n19082 0.00175333
R38678 DVSS.n824 DVSS.n819 0.00175333
R38679 DVSS.n5591 DVSS.n5590 0.00174016
R38680 DVSS.n5639 DVSS.n5638 0.00174016
R38681 DVSS.n5704 DVSS.n5703 0.00174016
R38682 DVSS.n5770 DVSS.n5769 0.00174016
R38683 DVSS.n4467 DVSS.n4466 0.00174016
R38684 DVSS.n4081 DVSS.n4080 0.00174016
R38685 DVSS.n6971 DVSS.n6970 0.00174016
R38686 DVSS.n7095 DVSS.n7094 0.00174016
R38687 DVSS.n7144 DVSS.n7143 0.00174016
R38688 DVSS.n19135 DVSS.n19134 0.00174016
R38689 DVSS.n19246 DVSS.n19245 0.00174016
R38690 DVSS.n866 DVSS.n865 0.00174016
R38691 DVSS.n10275 DVSS.n10274 0.00174016
R38692 DVSS.n10932 DVSS.n10931 0.00174016
R38693 DVSS.n10994 DVSS.n10993 0.00174016
R38694 DVSS.n11275 DVSS.n11274 0.00174016
R38695 DVSS.n9492 DVSS.n9491 0.00174016
R38696 DVSS.n9002 DVSS.n9001 0.00174016
R38697 DVSS.n12949 DVSS.n12948 0.00174016
R38698 DVSS.n12917 DVSS.n12916 0.00174016
R38699 DVSS.n12836 DVSS.n12835 0.00174016
R38700 DVSS.n12834 DVSS.n12833 0.00174016
R38701 DVSS.n12820 DVSS.n12819 0.00174016
R38702 DVSS.n12681 DVSS.n12680 0.00174016
R38703 DVSS.n12496 DVSS.n12495 0.00174016
R38704 DVSS.n12494 DVSS.n12493 0.00174016
R38705 DVSS.n12456 DVSS.n12455 0.00174016
R38706 DVSS.n12404 DVSS.n12403 0.00174016
R38707 DVSS.n12184 DVSS.n12183 0.00174016
R38708 DVSS.n12180 DVSS.n12179 0.00174016
R38709 DVSS.n21307 DVSS.n21306 0.00174016
R38710 DVSS.n21240 DVSS.n21239 0.00174016
R38711 DVSS.n21310 DVSS.n21309 0.00174016
R38712 DVSS.n21301 DVSS.n21300 0.00174016
R38713 DVSS.n21297 DVSS.n21296 0.00174016
R38714 DVSS.n17014 DVSS.n17013 0.00174016
R38715 DVSS.n17065 DVSS.n17064 0.00174016
R38716 DVSS.n16913 DVSS.n16912 0.00174016
R38717 DVSS.n17590 DVSS.n17589 0.00174016
R38718 DVSS.n15705 DVSS.n15704 0.00174016
R38719 DVSS.n14993 DVSS.n14992 0.00174016
R38720 DVSS.n13669 DVSS.n13668 0.00174016
R38721 DVSS.n13588 DVSS.n13587 0.00174016
R38722 DVSS.n13549 DVSS.n13548 0.00174016
R38723 DVSS.n20134 DVSS.n20133 0.00174016
R38724 DVSS.n20851 DVSS.n20850 0.00174016
R38725 DVSS.n10635 DVSS.n10634 0.00174016
R38726 DVSS.n10830 DVSS.n10829 0.00174016
R38727 DVSS.n10772 DVSS.n10771 0.00174016
R38728 DVSS.n11387 DVSS.n11386 0.00174016
R38729 DVSS.n11530 DVSS.n11529 0.00174016
R38730 DVSS.n11690 DVSS.n11689 0.00174016
R38731 DVSS.n13043 DVSS.n13042 0.00174016
R38732 DVSS.n12055 DVSS.n12054 0.00174016
R38733 DVSS.n67 DVSS.n66 0.00174016
R38734 DVSS.n21478 DVSS.n21477 0.00174016
R38735 DVSS.n5230 DVSS.n5229 0.00174016
R38736 DVSS.n4709 DVSS.n4708 0.00174016
R38737 DVSS.n4263 DVSS.n4262 0.00174016
R38738 DVSS.n3792 DVSS.n3791 0.00174016
R38739 DVSS.n3780 DVSS.n3779 0.00174016
R38740 DVSS.n3741 DVSS.n3740 0.00174016
R38741 DVSS.n3448 DVSS.n3447 0.00174016
R38742 DVSS.n3446 DVSS.n3445 0.00174016
R38743 DVSS.n3432 DVSS.n3431 0.00174016
R38744 DVSS.n3305 DVSS.n3304 0.00174016
R38745 DVSS.n3120 DVSS.n3119 0.00174016
R38746 DVSS.n3118 DVSS.n3117 0.00174016
R38747 DVSS.n3082 DVSS.n3081 0.00174016
R38748 DVSS.n3030 DVSS.n3029 0.00174016
R38749 DVSS.n2813 DVSS.n2812 0.00174016
R38750 DVSS.n2808 DVSS.n2807 0.00174016
R38751 DVSS.n671 DVSS.n670 0.00174016
R38752 DVSS.n771 DVSS.n770 0.00174016
R38753 DVSS.n780 DVSS.n779 0.00174016
R38754 DVSS.n664 DVSS.n663 0.00174016
R38755 DVSS.n707 DVSS.n706 0.00174016
R38756 DVSS.n9918 DVSS.n9917 0.00174016
R38757 DVSS.n9954 DVSS.n9953 0.00174016
R38758 DVSS.n9869 DVSS.n9868 0.00174016
R38759 DVSS.n11113 DVSS.n11112 0.00174016
R38760 DVSS.n9702 DVSS.n9701 0.00174016
R38761 DVSS.n9092 DVSS.n9091 0.00174016
R38762 DVSS.n13206 DVSS.n13205 0.00174016
R38763 DVSS.n13244 DVSS.n13243 0.00174016
R38764 DVSS.n13365 DVSS.n13364 0.00174016
R38765 DVSS.n20417 DVSS.n20416 0.00174016
R38766 DVSS.n21077 DVSS.n21076 0.00174016
R38767 DVSS.n17309 DVSS.n17308 0.00174016
R38768 DVSS.n17358 DVSS.n17357 0.00174016
R38769 DVSS.n17423 DVSS.n17422 0.00174016
R38770 DVSS.n16391 DVSS.n16390 0.00174016
R38771 DVSS.n16217 DVSS.n16216 0.00174016
R38772 DVSS.n7546 DVSS.n7545 0.00174016
R38773 DVSS.n18738 DVSS.n18737 0.00174016
R38774 DVSS.n18774 DVSS.n18773 0.00174016
R38775 DVSS.n18826 DVSS.n18825 0.00174016
R38776 DVSS.n19409 DVSS.n19408 0.00174016
R38777 DVSS.n19517 DVSS.n19516 0.00174016
R38778 DVSS.n1153 DVSS.n1152 0.00174016
R38779 DVSS.n5322 DVSS.n5321 0.00174016
R38780 DVSS.n5394 DVSS.n5393 0.00174016
R38781 DVSS.n5434 DVSS.n5433 0.00174016
R38782 DVSS.n5498 DVSS.n5497 0.00174016
R38783 DVSS.n6072 DVSS.n6071 0.00174016
R38784 DVSS.n6577 DVSS.n6576 0.00174016
R38785 DVSS.n6773 DVSS.n6772 0.00174016
R38786 DVSS.n3581 DVSS.n3580 0.00174016
R38787 DVSS.n3650 DVSS.n3649 0.00174016
R38788 DVSS.n18966 DVSS.n18965 0.00174016
R38789 DVSS.n544 DVSS.n543 0.00174016
R38790 DVSS.n16547 DVSS.n16546 0.00173932
R38791 DVSS.n16066 DVSS.n16065 0.00173932
R38792 DVSS.n17754 DVSS.n17753 0.00173932
R38793 DVSS.n18274 DVSS.n18273 0.00173932
R38794 DVSS.n16546 DVSS.n16545 0.00173932
R38795 DVSS.n16734 DVSS.n16733 0.00173932
R38796 DVSS.n15958 DVSS.n15957 0.00173932
R38797 DVSS.n15466 DVSS.n15465 0.00173932
R38798 DVSS.n15909 DVSS.n15908 0.00173932
R38799 DVSS.n16733 DVSS.n16732 0.00173932
R38800 DVSS DVSS.n21564 0.00173
R38801 DVSS.n21574 DVSS 0.00173
R38802 DVSS.n2336 DVSS.n2335 0.00172143
R38803 DVSS.n2413 DVSS.n2007 0.00172143
R38804 DVSS.n10719 DVSS.n10718 0.00172143
R38805 DVSS.n10722 DVSS.n10721 0.00172143
R38806 DVSS.n11304 DVSS.n11303 0.00172143
R38807 DVSS.n11301 DVSS.n8338 0.00172143
R38808 DVSS.n8892 DVSS.n8891 0.00172143
R38809 DVSS.n8895 DVSS.n8894 0.00172143
R38810 DVSS.n5796 DVSS.n5795 0.00170855
R38811 DVSS.n4070 DVSS.n4069 0.00170855
R38812 DVSS.n6983 DVSS.n6982 0.00170855
R38813 DVSS.n5797 DVSS.n5796 0.00170855
R38814 DVSS.n4069 DVSS.n4068 0.00170855
R38815 DVSS.n6982 DVSS.n6981 0.00170855
R38816 DVSS.n5570 DVSS.n5569 0.00170855
R38817 DVSS.n5758 DVSS.n5757 0.00170855
R38818 DVSS.n19244 DVSS.n19243 0.00170855
R38819 DVSS.n5569 DVSS.n5568 0.00170855
R38820 DVSS.n9844 DVSS.n9843 0.00170855
R38821 DVSS.n11261 DVSS.n11260 0.00170855
R38822 DVSS.n8988 DVSS.n8987 0.00170855
R38823 DVSS.n12963 DVSS.n12962 0.00170855
R38824 DVSS.n12422 DVSS.n12421 0.00170855
R38825 DVSS.n21228 DVSS.n21227 0.00170855
R38826 DVSS.n9845 DVSS.n9844 0.00170855
R38827 DVSS.n8989 DVSS.n8988 0.00170855
R38828 DVSS.n10210 DVSS.n10209 0.00170855
R38829 DVSS.n12962 DVSS.n12961 0.00170855
R38830 DVSS.n11262 DVSS.n11261 0.00170855
R38831 DVSS.n5759 DVSS.n5758 0.00170855
R38832 DVSS.n17562 DVSS.n17561 0.00170855
R38833 DVSS.n17604 DVSS.n17603 0.00170855
R38834 DVSS.n15007 DVSS.n15006 0.00170855
R38835 DVSS.n13655 DVSS.n13654 0.00170855
R38836 DVSS.n20254 DVSS.n20253 0.00170855
R38837 DVSS.n17561 DVSS.n17560 0.00170855
R38838 DVSS.n15006 DVSS.n15005 0.00170855
R38839 DVSS.n17603 DVSS.n17602 0.00170855
R38840 DVSS.n16955 DVSS.n16954 0.00170855
R38841 DVSS.n13656 DVSS.n13655 0.00170855
R38842 DVSS.n10617 DVSS.n10616 0.00170855
R38843 DVSS.n10741 DVSS.n10740 0.00170855
R38844 DVSS.n11401 DVSS.n11400 0.00170855
R38845 DVSS.n11418 DVSS.n11417 0.00170855
R38846 DVSS.n11448 DVSS.n11447 0.00170855
R38847 DVSS.n11704 DVSS.n11703 0.00170855
R38848 DVSS.n13029 DVSS.n13028 0.00170855
R38849 DVSS.n11703 DVSS.n11702 0.00170855
R38850 DVSS.n11400 DVSS.n11399 0.00170855
R38851 DVSS.n10740 DVSS.n10739 0.00170855
R38852 DVSS.n11417 DVSS.n11416 0.00170855
R38853 DVSS.n11447 DVSS.n11446 0.00170855
R38854 DVSS.n13030 DVSS.n13029 0.00170855
R38855 DVSS.n5223 DVSS.n5222 0.00170855
R38856 DVSS.n5222 DVSS.n5221 0.00170855
R38857 DVSS.n3804 DVSS.n3803 0.00170855
R38858 DVSS.n3768 DVSS.n3767 0.00170855
R38859 DVSS.n3049 DVSS.n3048 0.00170855
R38860 DVSS.n758 DVSS.n757 0.00170855
R38861 DVSS.n3803 DVSS.n3802 0.00170855
R38862 DVSS.n3769 DVSS.n3768 0.00170855
R38863 DVSS.n11085 DVSS.n11084 0.00170855
R38864 DVSS.n11127 DVSS.n11126 0.00170855
R38865 DVSS.n9078 DVSS.n9077 0.00170855
R38866 DVSS.n13220 DVSS.n13219 0.00170855
R38867 DVSS.n20528 DVSS.n20527 0.00170855
R38868 DVSS.n11084 DVSS.n11083 0.00170855
R38869 DVSS.n9079 DVSS.n9078 0.00170855
R38870 DVSS.n11126 DVSS.n11125 0.00170855
R38871 DVSS.n9911 DVSS.n9910 0.00170855
R38872 DVSS.n13219 DVSS.n13218 0.00170855
R38873 DVSS.n17265 DVSS.n17264 0.00170855
R38874 DVSS.n16417 DVSS.n16416 0.00170855
R38875 DVSS.n16379 DVSS.n16378 0.00170855
R38876 DVSS.n7534 DVSS.n7533 0.00170855
R38877 DVSS.n18750 DVSS.n18749 0.00170855
R38878 DVSS.n19515 DVSS.n19514 0.00170855
R38879 DVSS.n16418 DVSS.n16417 0.00170855
R38880 DVSS.n7535 DVSS.n7534 0.00170855
R38881 DVSS.n16380 DVSS.n16379 0.00170855
R38882 DVSS.n17264 DVSS.n17263 0.00170855
R38883 DVSS.n18749 DVSS.n18748 0.00170855
R38884 DVSS.n5330 DVSS.n5329 0.00170855
R38885 DVSS.n5853 DVSS.n5852 0.00170855
R38886 DVSS.n6084 DVSS.n6083 0.00170855
R38887 DVSS.n6340 DVSS.n6339 0.00170855
R38888 DVSS.n6451 DVSS.n6450 0.00170855
R38889 DVSS.n6785 DVSS.n6784 0.00170855
R38890 DVSS.n3593 DVSS.n3592 0.00170855
R38891 DVSS.n6339 DVSS.n6338 0.00170855
R38892 DVSS.n6784 DVSS.n6783 0.00170855
R38893 DVSS.n5329 DVSS.n5328 0.00170855
R38894 DVSS.n6083 DVSS.n6082 0.00170855
R38895 DVSS.n3592 DVSS.n3591 0.00170855
R38896 DVSS.n6452 DVSS.n6451 0.00170855
R38897 DVSS.n19243 DVSS.n19242 0.00170855
R38898 DVSS.n19514 DVSS.n19513 0.00170855
R38899 DVSS.n12423 DVSS.n12422 0.00170855
R38900 DVSS.n20527 DVSS.n20526 0.00170855
R38901 DVSS.n20253 DVSS.n20252 0.00170855
R38902 DVSS.n758 DVSS.n755 0.00170855
R38903 DVSS.n7240 DVSS.n7239 0.0017
R38904 DVSS.n18899 DVSS.n18898 0.0017
R38905 DVSS.n18915 DVSS.n18914 0.0017
R38906 DVSS.n19591 DVSS.n19590 0.0017
R38907 DVSS.n1067 DVSS.n1066 0.0017
R38908 DVSS.n1282 DVSS.n1281 0.0017
R38909 DVSS.n1299 DVSS.n1298 0.0017
R38910 DVSS.n1300 DVSS.n1297 0.0017
R38911 DVSS.n19592 DVSS.n19589 0.0017
R38912 DVSS.n18917 DVSS.n18916 0.0017
R38913 DVSS.n10864 DVSS.n10863 0.00169718
R38914 DVSS.n2333 DVSS.n2045 0.00165714
R38915 DVSS.n2335 DVSS.n2334 0.00165714
R38916 DVSS.n2007 DVSS.n2006 0.00165714
R38917 DVSS.n10105 DVSS.n10104 0.00165714
R38918 DVSS.n10700 DVSS.n10699 0.00165714
R38919 DVSS.n10651 DVSS.n10650 0.00165714
R38920 DVSS.n4782 DVSS.n4781 0.00165714
R38921 DVSS.n10652 DVSS.n10647 0.00165714
R38922 DVSS.n8300 DVSS.n8299 0.00165714
R38923 DVSS.n13094 DVSS.n13093 0.00165714
R38924 DVSS.n8089 DVSS.n8086 0.00165714
R38925 DVSS.n8166 DVSS.n8165 0.00165714
R38926 DVSS.n8217 DVSS.n8216 0.00165714
R38927 DVSS.n8302 DVSS.n8301 0.00165714
R38928 DVSS.n13095 DVSS.n13091 0.00165714
R38929 DVSS.n12986 DVSS.n12985 0.00165714
R38930 DVSS.n13011 DVSS.n13010 0.00165714
R38931 DVSS.n11851 DVSS.n11850 0.00165714
R38932 DVSS.n11910 DVSS.n11909 0.00165714
R38933 DVSS.n12987 DVSS.n12983 0.00165714
R38934 DVSS.n13012 DVSS.n13008 0.00165714
R38935 DVSS.n11320 DVSS.n11319 0.00165714
R38936 DVSS.n11346 DVSS.n11345 0.00165714
R38937 DVSS.n8381 DVSS.n8378 0.00165714
R38938 DVSS.n8458 DVSS.n8457 0.00165714
R38939 DVSS.n8509 DVSS.n8508 0.00165714
R38940 DVSS.n11321 DVSS.n11317 0.00165714
R38941 DVSS.n11347 DVSS.n11343 0.00165714
R38942 DVSS.n8631 DVSS.n8628 0.00165714
R38943 DVSS.n8332 DVSS.n8326 0.00165714
R38944 DVSS.n8874 DVSS.n8873 0.00165714
R38945 DVSS.n8331 DVSS.n8329 0.00165714
R38946 DVSS.n16538 DVSS.n16537 0.00163371
R38947 DVSS.n14215 DVSS.n14214 0.00163371
R38948 DVSS.n14216 DVSS.n14215 0.00163371
R38949 DVSS.n16537 DVSS.n16536 0.00163371
R38950 DVSS.n16725 DVSS.n16724 0.00163371
R38951 DVSS.n14882 DVSS.n14881 0.00163371
R38952 DVSS.n16724 DVSS.n16723 0.00163371
R38953 DVSS.n14881 DVSS.n14880 0.00163371
R38954 DVSS.n5062 DVSS.n5061 0.00162676
R38955 DVSS.n5178 DVSS.n5177 0.00162676
R38956 DVSS.n5140 DVSS.n5139 0.00162676
R38957 DVSS.n5086 DVSS.n5085 0.00162676
R38958 DVSS.n10355 DVSS.n10354 0.00162676
R38959 DVSS.n10356 DVSS.n10355 0.00162676
R38960 DVSS.n10874 DVSS.n10873 0.00162676
R38961 DVSS.n10871 DVSS.n10870 0.00162676
R38962 DVSS.n15397 DVSS.n15396 0.001625
R38963 DVSS.n18294 DVSS.n18293 0.001625
R38964 DVSS.n18304 DVSS.n18303 0.001625
R38965 DVSS.n5589 DVSS.n5588 0.00161999
R38966 DVSS.n5588 DVSS.n5587 0.00161999
R38967 DVSS.n10273 DVSS.n10272 0.00161999
R38968 DVSS.n12825 DVSS.n12824 0.00161999
R38969 DVSS.n12460 DVSS.n12459 0.00161999
R38970 DVSS.n21268 DVSS.n21267 0.00161999
R38971 DVSS.n10272 DVSS.n10271 0.00161999
R38972 DVSS.n17012 DVSS.n17011 0.00161999
R38973 DVSS.n17011 DVSS.n17010 0.00161999
R38974 DVSS.n10610 DVSS.n10609 0.00161999
R38975 DVSS.n10633 DVSS.n10632 0.00161999
R38976 DVSS.n10810 DVSS.n10809 0.00161999
R38977 DVSS.n11443 DVSS.n11442 0.00161999
R38978 DVSS.n11442 DVSS.n11441 0.00161999
R38979 DVSS.n10632 DVSS.n10631 0.00161999
R38980 DVSS.n10811 DVSS.n10810 0.00161999
R38981 DVSS.n10609 DVSS.n10608 0.00161999
R38982 DVSS.n5228 DVSS.n5227 0.00161999
R38983 DVSS.n5227 DVSS.n5226 0.00161999
R38984 DVSS.n3437 DVSS.n3436 0.00161999
R38985 DVSS.n3086 DVSS.n3085 0.00161999
R38986 DVSS.n711 DVSS.n710 0.00161999
R38987 DVSS.n12824 DVSS.n12823 0.00161999
R38988 DVSS.n3436 DVSS.n3435 0.00161999
R38989 DVSS.n9916 DVSS.n9915 0.00161999
R38990 DVSS.n9915 DVSS.n9914 0.00161999
R38991 DVSS.n17307 DVSS.n17306 0.00161999
R38992 DVSS.n17306 DVSS.n17305 0.00161999
R38993 DVSS.n5392 DVSS.n5391 0.00161999
R38994 DVSS.n5453 DVSS.n5452 0.00161999
R38995 DVSS.n6456 DVSS.n6455 0.00161999
R38996 DVSS.n6457 DVSS.n6456 0.00161999
R38997 DVSS.n5391 DVSS.n5390 0.00161999
R38998 DVSS.n5452 DVSS.n5451 0.00161999
R38999 DVSS.n12461 DVSS.n12460 0.00161999
R39000 DVSS.n3087 DVSS.n3086 0.00161999
R39001 DVSS.n21268 DVSS.n21266 0.00161999
R39002 DVSS.n4570 DVSS.n4569 0.00161111
R39003 DVSS.n11021 DVSS.n11020 0.00161111
R39004 DVSS.n4516 DVSS.n4515 0.00161111
R39005 DVSS.n11191 DVSS.n11190 0.00161111
R39006 DVSS.n4620 DVSS.n4619 0.00161111
R39007 DVSS.n10031 DVSS.n10030 0.00161111
R39008 DVSS.n4807 DVSS.n4803 0.00159286
R39009 DVSS.n10153 DVSS.n10152 0.00159286
R39010 DVSS.n10647 DVSS.n10646 0.00159286
R39011 DVSS.n8167 DVSS.n8166 0.00159286
R39012 DVSS.n8218 DVSS.n8217 0.00159286
R39013 DVSS.n8303 DVSS.n8302 0.00159286
R39014 DVSS.n13091 DVSS.n13090 0.00159286
R39015 DVSS.n12983 DVSS.n12982 0.00159286
R39016 DVSS.n13008 DVSS.n13007 0.00159286
R39017 DVSS.n8459 DVSS.n8458 0.00159286
R39018 DVSS.n8510 DVSS.n8509 0.00159286
R39019 DVSS.n11317 DVSS.n11316 0.00159286
R39020 DVSS.n11343 DVSS.n11342 0.00159286
R39021 DVSS.n8608 DVSS.n8607 0.00159286
R39022 DVSS.n8722 DVSS.n8721 0.00159286
R39023 DVSS.n8783 DVSS.n8782 0.00159286
R39024 DVSS.n8878 DVSS.n8877 0.00159286
R39025 DVSS.n8326 DVSS.n8325 0.00159286
R39026 DVSS.n2048 DVSS.n2047 0.00157975
R39027 DVSS.n5555 DVSS.n5554 0.00156299
R39028 DVSS.n5781 DVSS.n5780 0.00156299
R39029 DVSS.n5727 DVSS.n5726 0.00156299
R39030 DVSS.n4055 DVSS.n4054 0.00156299
R39031 DVSS.n6987 DVSS.n6986 0.00156299
R39032 DVSS.n7102 DVSS.n7101 0.00156299
R39033 DVSS.n19147 DVSS.n19146 0.00156299
R39034 DVSS.n10194 DVSS.n10193 0.00156299
R39035 DVSS.n11288 DVSS.n11287 0.00156299
R39036 DVSS.n13126 DVSS.n13125 0.00156299
R39037 DVSS.n12932 DVSS.n12931 0.00156299
R39038 DVSS.n12729 DVSS.n12728 0.00156299
R39039 DVSS.n12386 DVSS.n12214 0.00156299
R39040 DVSS.n21317 DVSS.n21316 0.00156299
R39041 DVSS.n21327 DVSS.n21326 0.00156299
R39042 DVSS.n21222 DVSS.n21221 0.00156299
R39043 DVSS.n16939 DVSS.n16938 0.00156299
R39044 DVSS.n17577 DVSS.n17576 0.00156299
R39045 DVSS.n15021 DVSS.n15020 0.00156299
R39046 DVSS.n13651 DVSS.n13650 0.00156299
R39047 DVSS.n13581 DVSS.n13580 0.00156299
R39048 DVSS.n20158 DVSS.n20157 0.00156299
R39049 DVSS.n10598 DVSS.n10597 0.00156299
R39050 DVSS.n10611 DVSS.n10610 0.00156299
R39051 DVSS.n10773 DVSS.n10772 0.00156299
R39052 DVSS.n11374 DVSS.n11373 0.00156299
R39053 DVSS.n11433 DVSS.n11432 0.00156299
R39054 DVSS.n13075 DVSS.n13074 0.00156299
R39055 DVSS.n12040 DVSS.n12039 0.00156299
R39056 DVSS.n5208 DVSS.n5207 0.00156299
R39057 DVSS.n3980 DVSS.n3979 0.00156299
R39058 DVSS.n3754 DVSS.n3753 0.00156299
R39059 DVSS.n3351 DVSS.n3350 0.00156299
R39060 DVSS.n3013 DVSS.n2844 0.00156299
R39061 DVSS.n675 DVSS.n674 0.00156299
R39062 DVSS.n677 DVSS.n676 0.00156299
R39063 DVSS.n751 DVSS.n750 0.00156299
R39064 DVSS.n9895 DVSS.n9894 0.00156299
R39065 DVSS.n11100 DVSS.n11099 0.00156299
R39066 DVSS.n9064 DVSS.n9063 0.00156299
R39067 DVSS.n13224 DVSS.n13223 0.00156299
R39068 DVSS.n13251 DVSS.n13250 0.00156299
R39069 DVSS.n20429 DVSS.n20428 0.00156299
R39070 DVSS.n17250 DVSS.n17249 0.00156299
R39071 DVSS.n16402 DVSS.n16401 0.00156299
R39072 DVSS.n16348 DVSS.n16347 0.00156299
R39073 DVSS.n7520 DVSS.n7519 0.00156299
R39074 DVSS.n18754 DVSS.n18753 0.00156299
R39075 DVSS.n18781 DVSS.n18780 0.00156299
R39076 DVSS.n19421 DVSS.n19420 0.00156299
R39077 DVSS.n5313 DVSS.n5312 0.00156299
R39078 DVSS.n5323 DVSS.n5322 0.00156299
R39079 DVSS.n5499 DVSS.n5498 0.00156299
R39080 DVSS.n6061 DVSS.n6060 0.00156299
R39081 DVSS.n6466 DVSS.n6465 0.00156299
R39082 DVSS.n6828 DVSS.n6827 0.00156299
R39083 DVSS.n3637 DVSS.n3636 0.00156299
R39084 DVSS.n5066 DVSS.n5063 0.00155634
R39085 DVSS.n5067 DVSS.n5062 0.00155634
R39086 DVSS.n5070 DVSS.n5069 0.00155634
R39087 DVSS.n5310 DVSS.n5309 0.00155634
R39088 DVSS.n5244 DVSS.n5243 0.00155634
R39089 DVSS.n5161 DVSS.n5160 0.00155634
R39090 DVSS.n5107 DVSS.n5106 0.00155634
R39091 DVSS.n10396 DVSS.n10395 0.00155634
R39092 DVSS.n10399 DVSS.n10398 0.00155634
R39093 DVSS.n10455 DVSS.n10454 0.00155634
R39094 DVSS.n10458 DVSS.n10457 0.00155634
R39095 DVSS.n10498 DVSS.n10497 0.00155634
R39096 DVSS.n10501 DVSS.n10500 0.00155634
R39097 DVSS.n16568 DVSS.n16567 0.00155634
R39098 DVSS.n16572 DVSS.n16571 0.00155634
R39099 DVSS.n16577 DVSS.n16576 0.00155634
R39100 DVSS.n16662 DVSS.n16661 0.00155634
R39101 DVSS.n16104 DVSS.n16103 0.00155634
R39102 DVSS.n16063 DVSS.n16062 0.00155634
R39103 DVSS.n16061 DVSS.n16060 0.00155634
R39104 DVSS.n17733 DVSS.n17732 0.00155634
R39105 DVSS.n18105 DVSS.n18104 0.00155634
R39106 DVSS.n18138 DVSS.n18137 0.00155634
R39107 DVSS.n18269 DVSS.n18268 0.00155634
R39108 DVSS.n18257 DVSS.n18256 0.00155634
R39109 DVSS.n18203 DVSS.n18202 0.00155634
R39110 DVSS.n14458 DVSS.n14457 0.00155634
R39111 DVSS.n14476 DVSS.n14475 0.00155634
R39112 DVSS.n19674 DVSS.n19673 0.00155634
R39113 DVSS.n16755 DVSS.n16754 0.00155634
R39114 DVSS.n16759 DVSS.n16758 0.00155634
R39115 DVSS.n16764 DVSS.n16763 0.00155634
R39116 DVSS.n17161 DVSS.n17160 0.00155634
R39117 DVSS.n15985 DVSS.n15984 0.00155634
R39118 DVSS.n15955 DVSS.n15954 0.00155634
R39119 DVSS.n15953 DVSS.n15952 0.00155634
R39120 DVSS.n15930 DVSS.n15929 0.00155634
R39121 DVSS.n15383 DVSS.n15382 0.00155634
R39122 DVSS.n15443 DVSS.n15442 0.00155634
R39123 DVSS.n15471 DVSS.n15470 0.00155634
R39124 DVSS.n15483 DVSS.n15482 0.00155634
R39125 DVSS.n15537 DVSS.n15536 0.00155634
R39126 DVSS.n14664 DVSS.n14663 0.00155634
R39127 DVSS.n14644 DVSS.n14639 0.00155634
R39128 DVSS.n19889 DVSS.n19888 0.00155634
R39129 DVSS.n10086 DVSS.n10085 0.00154636
R39130 DVSS.n10704 DVSS.n10703 0.00154636
R39131 DVSS.n10705 DVSS.n10704 0.00154636
R39132 DVSS.n10087 DVSS.n10086 0.00154636
R39133 DVSS DVSS.n10888 0.00153286
R39134 DVSS.n6955 DVSS.n6954 0.00153143
R39135 DVSS.n5565 DVSS.n5564 0.00153143
R39136 DVSS.n12945 DVSS.n12944 0.00153143
R39137 DVSS.n12709 DVSS.n12708 0.00153143
R39138 DVSS.n10206 DVSS.n10205 0.00153143
R39139 DVSS.n13847 DVSS.n13846 0.00153143
R39140 DVSS.n16951 DVSS.n16950 0.00153143
R39141 DVSS.n13848 DVSS.n13847 0.00153143
R39142 DVSS.n12944 DVSS.n12943 0.00153143
R39143 DVSS.n10816 DVSS.n10815 0.00153143
R39144 DVSS.n10768 DVSS.n10767 0.00153143
R39145 DVSS.n10765 DVSS.n10764 0.00153143
R39146 DVSS.n13047 DVSS.n13046 0.00153143
R39147 DVSS.n13048 DVSS.n13047 0.00153143
R39148 DVSS.n10769 DVSS.n10768 0.00153143
R39149 DVSS.n10766 DVSS.n10765 0.00153143
R39150 DVSS.n10817 DVSS.n10816 0.00153143
R39151 DVSS.n5218 DVSS.n5217 0.00153143
R39152 DVSS.n3785 DVSS.n3784 0.00153143
R39153 DVSS.n3332 DVSS.n3331 0.00153143
R39154 DVSS.n3035 DVSS.n3034 0.00153143
R39155 DVSS.n784 DVSS.n782 0.00153143
R39156 DVSS.n13185 DVSS.n13184 0.00153143
R39157 DVSS.n13184 DVSS.n13183 0.00153143
R39158 DVSS.n9907 DVSS.n9906 0.00153143
R39159 DVSS.n18577 DVSS.n18576 0.00153143
R39160 DVSS.n18576 DVSS.n18575 0.00153143
R39161 DVSS.n17260 DVSS.n17259 0.00153143
R39162 DVSS.n3784 DVSS.n3783 0.00153143
R39163 DVSS.n6956 DVSS.n6955 0.00153143
R39164 DVSS.n5448 DVSS.n5447 0.00153143
R39165 DVSS.n5495 DVSS.n5494 0.00153143
R39166 DVSS.n5491 DVSS.n5490 0.00153143
R39167 DVSS.n3577 DVSS.n3576 0.00153143
R39168 DVSS.n5447 DVSS.n5446 0.00153143
R39169 DVSS.n5492 DVSS.n5491 0.00153143
R39170 DVSS.n5494 DVSS.n5493 0.00153143
R39171 DVSS.n3576 DVSS.n3575 0.00153143
R39172 DVSS.n3036 DVSS.n3035 0.00153143
R39173 DVSS.n12409 DVSS.n12408 0.00153143
R39174 DVSS.n12710 DVSS.n12709 0.00153143
R39175 DVSS.n3333 DVSS.n3332 0.00153143
R39176 DVSS.n784 DVSS.n783 0.00153143
R39177 DVSS.n21199 DVSS.n21198 0.00153143
R39178 DVSS.n21189 DVSS.n21188 0.00153143
R39179 DVSS.n703 DVSS.n702 0.00153143
R39180 DVSS.n4763 DVSS.n4762 0.00152857
R39181 DVSS.n4628 DVSS.n4627 0.00152857
R39182 DVSS.n4869 DVSS.n4868 0.00152857
R39183 DVSS.n4759 DVSS.n4758 0.00152857
R39184 DVSS.n10089 DVSS.n10088 0.00152857
R39185 DVSS.n10156 DVSS.n10155 0.00152857
R39186 DVSS.n10707 DVSS.n10706 0.00152857
R39187 DVSS.n10658 DVSS.n10657 0.00152857
R39188 DVSS.n10655 DVSS.n10654 0.00152857
R39189 DVSS.n6791 DVSS.n6790 0.00152857
R39190 DVSS.n3815 DVSS.n3814 0.00152857
R39191 DVSS.n3913 DVSS.n3912 0.00152857
R39192 DVSS.n3867 DVSS.n3866 0.00152857
R39193 DVSS.n8107 DVSS.n8106 0.00152857
R39194 DVSS.n8108 DVSS.n8107 0.00152857
R39195 DVSS.n3599 DVSS.n3598 0.00152857
R39196 DVSS.n2588 DVSS.n2587 0.00152857
R39197 DVSS.n2684 DVSS.n2683 0.00152857
R39198 DVSS.n2630 DVSS.n2629 0.00152857
R39199 DVSS.n11784 DVSS.n11783 0.00152857
R39200 DVSS.n11785 DVSS.n11784 0.00152857
R39201 DVSS.n5863 DVSS.n5862 0.00152857
R39202 DVSS.n5991 DVSS.n5990 0.00152857
R39203 DVSS.n5945 DVSS.n5944 0.00152857
R39204 DVSS.n8399 DVSS.n8398 0.00152857
R39205 DVSS.n8400 DVSS.n8399 0.00152857
R39206 DVSS.n11353 DVSS.n11352 0.00152857
R39207 DVSS.n11350 DVSS.n11349 0.00152857
R39208 DVSS.n6090 DVSS.n6089 0.00152857
R39209 DVSS.n6245 DVSS.n6244 0.00152857
R39210 DVSS.n6187 DVSS.n6186 0.00152857
R39211 DVSS.n8652 DVSS.n8651 0.00152857
R39212 DVSS.n8724 DVSS.n8723 0.00152857
R39213 DVSS.n8785 DVSS.n8784 0.00152857
R39214 DVSS.n8880 DVSS.n8879 0.00152857
R39215 DVSS.n8906 DVSS.n8905 0.00152857
R39216 DVSS.n8335 DVSS.n8334 0.00152857
R39217 DVSS.n8648 DVSS.n8647 0.00152857
R39218 DVSS.n18115 DVSS.n18114 0.00152817
R39219 DVSS.n15405 DVSS.n15404 0.00152817
R39220 DVSS.n16563 DVSS.n16562 0.00152811
R39221 DVSS.n16100 DVSS.n16099 0.00152811
R39222 DVSS.n16562 DVSS.n16561 0.00152811
R39223 DVSS.n16750 DVSS.n16749 0.00152811
R39224 DVSS.n15981 DVSS.n15980 0.00152811
R39225 DVSS.n16749 DVSS.n16748 0.00152811
R39226 DVSS.n4973 DVSS.n4972 0.00151423
R39227 DVSS.n4929 DVSS.n4928 0.00151423
R39228 DVSS.n4930 DVSS.n4929 0.00151423
R39229 DVSS.n4974 DVSS.n4973 0.00151423
R39230 DVSS.n5379 DVSS.n5378 0.00150559
R39231 DVSS.n5370 DVSS.n5369 0.00150559
R39232 DVSS.n5585 DVSS.n5582 0.00150559
R39233 DVSS.n5581 DVSS.n5579 0.00150559
R39234 DVSS.n17270 DVSS.n17267 0.00150559
R39235 DVSS.n17274 DVSS.n17273 0.00150559
R39236 DVSS.n17004 DVSS.n17001 0.00150559
R39237 DVSS.n17030 DVSS.n17029 0.00150559
R39238 DVSS.n10224 DVSS.n10221 0.00150559
R39239 DVSS.n10237 DVSS.n10236 0.00150559
R39240 DVSS.n10256 DVSS.n10253 0.00150559
R39241 DVSS.n10291 DVSS.n10290 0.00150559
R39242 DVSS.n10322 DVSS.n10320 0.00148592
R39243 DVSS.n10322 DVSS.n10321 0.00148592
R39244 DVSS.n10317 DVSS.n10316 0.00148592
R39245 DVSS.n10318 DVSS.n10317 0.00148592
R39246 DVSS.n10323 DVSS.n10318 0.00148592
R39247 DVSS.n10324 DVSS.n10323 0.00148592
R39248 DVSS.n7039 DVSS.n7037 0.00147867
R39249 DVSS.n7078 DVSS.n7077 0.00147867
R39250 DVSS.n13609 DVSS.n13608 0.00147867
R39251 DVSS.n13629 DVSS.n13628 0.00147867
R39252 DVSS.n13632 DVSS.n13629 0.00147867
R39253 DVSS.n13612 DVSS.n13609 0.00147867
R39254 DVSS.n7079 DVSS.n7078 0.00147867
R39255 DVSS.n7037 DVSS.n7036 0.00147867
R39256 DVSS.n4631 DVSS.n4629 0.00146429
R39257 DVSS.n4969 DVSS.n4966 0.00146429
R39258 DVSS.n4925 DVSS.n4922 0.00146429
R39259 DVSS.n4865 DVSS.n4862 0.00146429
R39260 DVSS.n4632 DVSS.n4628 0.00146429
R39261 DVSS.n4635 DVSS.n4634 0.00146429
R39262 DVSS.n4638 DVSS.n4637 0.00146429
R39263 DVSS.n4976 DVSS.n4975 0.00146429
R39264 DVSS.n4932 DVSS.n4931 0.00146429
R39265 DVSS.n4872 DVSS.n4871 0.00146429
R39266 DVSS.n4756 DVSS.n4755 0.00146429
R39267 DVSS.n6795 DVSS.n6792 0.00146429
R39268 DVSS.n3823 DVSS.n3816 0.00146429
R39269 DVSS.n3910 DVSS.n3907 0.00146429
R39270 DVSS.n3864 DVSS.n3861 0.00146429
R39271 DVSS.n6796 DVSS.n6791 0.00146429
R39272 DVSS.n3824 DVSS.n3815 0.00146429
R39273 DVSS.n3912 DVSS.n3911 0.00146429
R39274 DVSS.n3866 DVSS.n3865 0.00146429
R39275 DVSS.n3602 DVSS.n3600 0.00146429
R39276 DVSS.n2591 DVSS.n2589 0.00146429
R39277 DVSS.n2704 DVSS.n2701 0.00146429
R39278 DVSS.n2650 DVSS.n2647 0.00146429
R39279 DVSS.n3603 DVSS.n3599 0.00146429
R39280 DVSS.n2592 DVSS.n2588 0.00146429
R39281 DVSS.n2706 DVSS.n2705 0.00146429
R39282 DVSS.n2652 DVSS.n2651 0.00146429
R39283 DVSS.n11825 DVSS.n11824 0.00146429
R39284 DVSS.n11828 DVSS.n11827 0.00146429
R39285 DVSS.n11884 DVSS.n11883 0.00146429
R39286 DVSS.n11887 DVSS.n11886 0.00146429
R39287 DVSS.n5867 DVSS.n5864 0.00146429
R39288 DVSS.n5988 DVSS.n5985 0.00146429
R39289 DVSS.n5942 DVSS.n5939 0.00146429
R39290 DVSS.n5868 DVSS.n5863 0.00146429
R39291 DVSS.n5871 DVSS.n5870 0.00146429
R39292 DVSS.n6048 DVSS.n6047 0.00146429
R39293 DVSS.n5990 DVSS.n5989 0.00146429
R39294 DVSS.n5944 DVSS.n5943 0.00146429
R39295 DVSS.n6095 DVSS.n6090 0.00146429
R39296 DVSS.n6098 DVSS.n6097 0.00146429
R39297 DVSS.n6101 DVSS.n6100 0.00146429
R39298 DVSS.n6247 DVSS.n6246 0.00146429
R39299 DVSS.n6189 DVSS.n6188 0.00146429
R39300 DVSS.n8654 DVSS.n8653 0.00146429
R39301 DVSS.n6094 DVSS.n6091 0.00146429
R39302 DVSS.n6241 DVSS.n6238 0.00146429
R39303 DVSS.n6183 DVSS.n6180 0.00146429
R39304 DVSS.n12501 DVSS.n12500 0.00146154
R39305 DVSS.n12516 DVSS.n12511 0.00146154
R39306 DVSS.n12640 DVSS.n12635 0.00146154
R39307 DVSS.n12625 DVSS.n12624 0.00146154
R39308 DVSS.n12352 DVSS.n12347 0.00146154
R39309 DVSS.n12337 DVSS.n12336 0.00146154
R39310 DVSS.n21325 DVSS.n21323 0.00146154
R39311 DVSS.n21161 DVSS.n21145 0.00146154
R39312 DVSS.n3125 DVSS.n3124 0.00146154
R39313 DVSS.n3140 DVSS.n3135 0.00146154
R39314 DVSS.n3264 DVSS.n3259 0.00146154
R39315 DVSS.n3249 DVSS.n3248 0.00146154
R39316 DVSS.n2979 DVSS.n2974 0.00146154
R39317 DVSS.n2964 DVSS.n2963 0.00146154
R39318 DVSS.n899 DVSS.n898 0.00146154
R39319 DVSS.n926 DVSS.n909 0.00146154
R39320 DVSS.n3411 DVSS.n3410 0.00146154
R39321 DVSS.n12792 DVSS.n12791 0.00146154
R39322 DVSS.n14538 DVSS.n14537 0.00146
R39323 DVSS.n20075 DVSS.n20074 0.00146
R39324 DVSS.n501 DVSS.n500 0.00146
R39325 DVSS.n502 DVSS.n499 0.00146
R39326 DVSS.n20077 DVSS.n20076 0.00146
R39327 DVSS.n14539 DVSS.n14536 0.00146
R39328 DVSS.n7169 DVSS.n7167 0.00145745
R39329 DVSS.n7186 DVSS.n7184 0.00145745
R39330 DVSS.n7307 DVSS.n7302 0.00145745
R39331 DVSS.n7316 DVSS.n7314 0.00145745
R39332 DVSS.n7873 DVSS.n7871 0.00145745
R39333 DVSS.n7883 DVSS.n7881 0.00145745
R39334 DVSS.n7962 DVSS.n7959 0.00145745
R39335 DVSS.n13377 DVSS.n13376 0.00145745
R39336 DVSS.n7061 DVSS.n7060 0.00145745
R39337 DVSS.n7051 DVSS.n7050 0.00145745
R39338 DVSS.n13302 DVSS.n13300 0.00145745
R39339 DVSS.n13314 DVSS.n13313 0.00145745
R39340 DVSS.n2343 DVSS.n2342 0.00144995
R39341 DVSS.n5617 DVSS.n5616 0.00144287
R39342 DVSS.n5616 DVSS.n5615 0.00144287
R39343 DVSS.n10906 DVSS.n10905 0.00144287
R39344 DVSS.n12762 DVSS.n12761 0.00144287
R39345 DVSS.n12391 DVSS.n12390 0.00144287
R39346 DVSS.n21134 DVSS.n21133 0.00144287
R39347 DVSS.n10905 DVSS.n10904 0.00144287
R39348 DVSS.n17039 DVSS.n17038 0.00144287
R39349 DVSS.n17038 DVSS.n17037 0.00144287
R39350 DVSS.n10856 DVSS.n10855 0.00144287
R39351 DVSS.n10857 DVSS.n10856 0.00144287
R39352 DVSS.n5203 DVSS.n5202 0.00144287
R39353 DVSS.n5204 DVSS.n5203 0.00144287
R39354 DVSS.n3374 DVSS.n3373 0.00144287
R39355 DVSS.n3017 DVSS.n3016 0.00144287
R39356 DVSS.n713 DVSS.n712 0.00144287
R39357 DVSS.n9928 DVSS.n9927 0.00144287
R39358 DVSS.n9927 DVSS.n9926 0.00144287
R39359 DVSS.n17336 DVSS.n17335 0.00144287
R39360 DVSS.n17335 DVSS.n17334 0.00144287
R39361 DVSS.n5412 DVSS.n5411 0.00144287
R39362 DVSS.n5411 DVSS.n5410 0.00144287
R39363 DVSS.n12761 DVSS.n12760 0.00144287
R39364 DVSS.n12390 DVSS.n12389 0.00144287
R39365 DVSS.n21134 DVSS.n21132 0.00144287
R39366 DVSS.n14721 DVSS.n14720 0.0014225
R39367 DVSS.n16101 DVSS.n16100 0.0014225
R39368 DVSS.n18468 DVSS.n18467 0.0014225
R39369 DVSS.n19667 DVSS.n19666 0.0014225
R39370 DVSS.n18217 DVSS.n18216 0.0014225
R39371 DVSS.n18467 DVSS.n18466 0.0014225
R39372 DVSS.n16648 DVSS.n16647 0.0014225
R39373 DVSS.n16102 DVSS.n16101 0.0014225
R39374 DVSS.n14407 DVSS.n14406 0.0014225
R39375 DVSS.n19666 DVSS.n19665 0.0014225
R39376 DVSS.n15982 DVSS.n15981 0.0014225
R39377 DVSS.n15523 DVSS.n15522 0.0014225
R39378 DVSS.n15134 DVSS.n15133 0.0014225
R39379 DVSS.n19882 DVSS.n19881 0.0014225
R39380 DVSS.n19881 DVSS.n19880 0.0014225
R39381 DVSS.n15135 DVSS.n15134 0.0014225
R39382 DVSS.n17175 DVSS.n17174 0.0014225
R39383 DVSS.n15983 DVSS.n15982 0.0014225
R39384 DVSS.n5514 DVSS.n5513 0.00141663
R39385 DVSS.n10041 DVSS.n10040 0.00141663
R39386 DVSS.n10040 DVSS.n10039 0.00141663
R39387 DVSS.n5513 DVSS.n5512 0.00141663
R39388 DVSS.n5066 DVSS.n5065 0.00141549
R39389 DVSS.n5242 DVSS.n5241 0.00141549
R39390 DVSS.n5159 DVSS.n5158 0.00141549
R39391 DVSS.n5105 DVSS.n5104 0.00141549
R39392 DVSS.n5068 DVSS.n5067 0.00141549
R39393 DVSS.n5243 DVSS.n5239 0.00141549
R39394 DVSS.n5160 DVSS.n5156 0.00141549
R39395 DVSS.n5106 DVSS.n5102 0.00141549
R39396 DVSS DVSS.n12999 0.00141429
R39397 DVSS.n9307 DVSS.n9306 0.00140496
R39398 DVSS.n9306 DVSS.n9305 0.00140496
R39399 DVSS.n20098 DVSS.n20097 0.00140496
R39400 DVSS.n20375 DVSS.n20374 0.00140496
R39401 DVSS.n19578 DVSS.n19577 0.00140496
R39402 DVSS.n19310 DVSS.n19309 0.00140496
R39403 DVSS.n19573 DVSS.n19572 0.00140496
R39404 DVSS.n20097 DVSS.n20096 0.00140496
R39405 DVSS.n20374 DVSS.n20373 0.00140496
R39406 DVSS.n20690 DVSS.n20689 0.00140496
R39407 DVSS.n20919 DVSS.n20918 0.00140496
R39408 DVSS.n20920 DVSS.n20919 0.00140496
R39409 DVSS.n20691 DVSS.n20690 0.00140496
R39410 DVSS.n1280 DVSS.n1279 0.00140496
R39411 DVSS.n1065 DVSS.n1064 0.00140496
R39412 DVSS.n1071 DVSS.n1070 0.00140496
R39413 DVSS.n1286 DVSS.n1285 0.00140496
R39414 DVSS.n20700 DVSS.n20699 0.00140496
R39415 DVSS.n20929 DVSS.n20928 0.00140496
R39416 DVSS.n17218 DVSS.n17217 0.0014
R39417 DVSS.n17226 DVSS.n17225 0.0014
R39418 DVSS.n17229 DVSS.n17228 0.0014
R39419 DVSS.n17231 DVSS.n17230 0.0014
R39420 DVSS.n15186 DVSS.n15185 0.0014
R39421 DVSS.n15145 DVSS.n15144 0.0014
R39422 DVSS.n2381 DVSS.n2380 0.0014
R39423 DVSS.n17696 DVSS.n17695 0.0014
R39424 DVSS.n4795 DVSS.n4792 0.0014
R39425 DVSS.n4795 DVSS.n4794 0.0014
R39426 DVSS.n4800 DVSS.n4799 0.0014
R39427 DVSS.n4799 DVSS.n4798 0.0014
R39428 DVSS.n4796 DVSS.n4791 0.0014
R39429 DVSS.n8078 DVSS.n8076 0.0014
R39430 DVSS.n8078 DVSS.n8077 0.0014
R39431 DVSS.n8073 DVSS.n8072 0.0014
R39432 DVSS.n8074 DVSS.n8073 0.0014
R39433 DVSS.n8079 DVSS.n8074 0.0014
R39434 DVSS.n8080 DVSS.n8079 0.0014
R39435 DVSS.n11757 DVSS.n11755 0.0014
R39436 DVSS.n11757 DVSS.n11756 0.0014
R39437 DVSS.n11752 DVSS.n11751 0.0014
R39438 DVSS.n11753 DVSS.n11752 0.0014
R39439 DVSS.n11758 DVSS.n11753 0.0014
R39440 DVSS.n11759 DVSS.n11758 0.0014
R39441 DVSS.n8370 DVSS.n8368 0.0014
R39442 DVSS.n8370 DVSS.n8369 0.0014
R39443 DVSS.n8365 DVSS.n8364 0.0014
R39444 DVSS.n8366 DVSS.n8365 0.0014
R39445 DVSS.n8371 DVSS.n8366 0.0014
R39446 DVSS.n8372 DVSS.n8371 0.0014
R39447 DVSS.n8612 DVSS.n8611 0.0014
R39448 DVSS.n8613 DVSS.n8612 0.0014
R39449 DVSS.n8620 DVSS.n8619 0.0014
R39450 DVSS.n8618 DVSS.n8616 0.0014
R39451 DVSS.n8618 DVSS.n8617 0.0014
R39452 DVSS.n7241 DVSS.n7240 0.0014
R39453 DVSS.n18900 DVSS.n18899 0.0014
R39454 DVSS.n19312 DVSS.n19311 0.0014
R39455 DVSS.n12093 DVSS.n12092 0.00138997
R39456 DVSS.n12094 DVSS.n12093 0.00138997
R39457 DVSS.n5623 DVSS.n5622 0.00138583
R39458 DVSS.n7146 DVSS.n7145 0.00138583
R39459 DVSS.n7174 DVSS.n7173 0.00138583
R39460 DVSS.n19152 DVSS.n19151 0.00138583
R39461 DVSS.n10912 DVSS.n10911 0.00138583
R39462 DVSS.n12757 DVSS.n12756 0.00138583
R39463 DVSS.n12730 DVSS.n12729 0.00138583
R39464 DVSS.n12714 DVSS.n12713 0.00138583
R39465 DVSS.n12463 DVSS.n12462 0.00138583
R39466 DVSS.n12447 DVSS.n12446 0.00138583
R39467 DVSS.n12446 DVSS.n12445 0.00138583
R39468 DVSS.n12186 DVSS.n12185 0.00138583
R39469 DVSS.n12173 DVSS.n12172 0.00138583
R39470 DVSS.n12172 DVSS.n12171 0.00138583
R39471 DVSS.n21326 DVSS.n21317 0.00138583
R39472 DVSS.n21187 DVSS.n21186 0.00138583
R39473 DVSS.n21185 DVSS.n21184 0.00138583
R39474 DVSS.n21143 DVSS.n21142 0.00138583
R39475 DVSS.n17045 DVSS.n17044 0.00138583
R39476 DVSS.n13547 DVSS.n13546 0.00138583
R39477 DVSS.n13533 DVSS.n13532 0.00138583
R39478 DVSS.n20163 DVSS.n20162 0.00138583
R39479 DVSS.n10850 DVSS.n10849 0.00138583
R39480 DVSS.n10763 DVSS.n10762 0.00138583
R39481 DVSS.n10760 DVSS.n10759 0.00138583
R39482 DVSS.n5197 DVSS.n5196 0.00138583
R39483 DVSS.n3370 DVSS.n3369 0.00138583
R39484 DVSS.n3352 DVSS.n3351 0.00138583
R39485 DVSS.n3337 DVSS.n3336 0.00138583
R39486 DVSS.n3089 DVSS.n3088 0.00138583
R39487 DVSS.n3074 DVSS.n3073 0.00138583
R39488 DVSS.n3073 DVSS.n3072 0.00138583
R39489 DVSS.n2815 DVSS.n2814 0.00138583
R39490 DVSS.n2801 DVSS.n2800 0.00138583
R39491 DVSS.n2800 DVSS.n2799 0.00138583
R39492 DVSS.n676 DVSS.n675 0.00138583
R39493 DVSS.n701 DVSS.n700 0.00138583
R39494 DVSS.n699 DVSS.n698 0.00138583
R39495 DVSS.n696 DVSS.n695 0.00138583
R39496 DVSS.n9934 DVSS.n9933 0.00138583
R39497 DVSS.n13367 DVSS.n13366 0.00138583
R39498 DVSS.n13384 DVSS.n13383 0.00138583
R39499 DVSS.n20434 DVSS.n20433 0.00138583
R39500 DVSS.n17342 DVSS.n17341 0.00138583
R39501 DVSS.n18828 DVSS.n18827 0.00138583
R39502 DVSS.n18842 DVSS.n18841 0.00138583
R39503 DVSS.n19426 DVSS.n19425 0.00138583
R39504 DVSS.n5418 DVSS.n5417 0.00138583
R39505 DVSS.n5489 DVSS.n5488 0.00138583
R39506 DVSS.n5486 DVSS.n5485 0.00138583
R39507 DVSS.n4870 DVSS.n4869 0.00138568
R39508 DVSS.n4757 DVSS.n4756 0.00138568
R39509 DVSS.n4758 DVSS.n4757 0.00138568
R39510 DVSS.n4871 DVSS.n4870 0.00138568
R39511 DVSS.n7150 DVSS.n7149 0.00135432
R39512 DVSS.n13543 DVSS.n13542 0.00135432
R39513 DVSS.n13371 DVSS.n13370 0.00135432
R39514 DVSS.n18832 DVSS.n18831 0.00135432
R39515 DVSS.n5788 DVSS.n5787 0.0013543
R39516 DVSS.n4061 DVSS.n4060 0.0013543
R39517 DVSS.n19145 DVSS.n19144 0.0013543
R39518 DVSS.n5787 DVSS.n5786 0.0013543
R39519 DVSS.n4062 DVSS.n4061 0.0013543
R39520 DVSS.n11294 DVSS.n11293 0.0013543
R39521 DVSS.n13120 DVSS.n13119 0.0013543
R39522 DVSS.n12938 DVSS.n12937 0.0013543
R39523 DVSS.n12717 DVSS.n12716 0.0013543
R39524 DVSS.n12473 DVSS.n12472 0.0013543
R39525 DVSS.n12467 DVSS.n12466 0.0013543
R39526 DVSS.n12193 DVSS.n12192 0.0013543
R39527 DVSS.n12189 DVSS.n12188 0.0013543
R39528 DVSS.n12939 DVSS.n12938 0.0013543
R39529 DVSS.n13119 DVSS.n13118 0.0013543
R39530 DVSS.n11295 DVSS.n11294 0.0013543
R39531 DVSS.n19144 DVSS.n19143 0.0013543
R39532 DVSS.n17571 DVSS.n17570 0.0013543
R39533 DVSS.n15015 DVSS.n15014 0.0013543
R39534 DVSS.n20156 DVSS.n20155 0.0013543
R39535 DVSS.n20155 DVSS.n20154 0.0013543
R39536 DVSS.n15014 DVSS.n15013 0.0013543
R39537 DVSS.n17570 DVSS.n17569 0.0013543
R39538 DVSS.n11368 DVSS.n11367 0.0013543
R39539 DVSS.n11413 DVSS.n11412 0.0013543
R39540 DVSS.n11425 DVSS.n11424 0.0013543
R39541 DVSS.n13081 DVSS.n13080 0.0013543
R39542 DVSS.n12034 DVSS.n12033 0.0013543
R39543 DVSS.n12033 DVSS.n12032 0.0013543
R39544 DVSS.n13082 DVSS.n13081 0.0013543
R39545 DVSS.n11412 DVSS.n11411 0.0013543
R39546 DVSS.n11367 DVSS.n11366 0.0013543
R39547 DVSS.n11424 DVSS.n11423 0.0013543
R39548 DVSS.n3974 DVSS.n3973 0.0013543
R39549 DVSS.n3761 DVSS.n3760 0.0013543
R39550 DVSS.n3340 DVSS.n3339 0.0013543
R39551 DVSS.n3099 DVSS.n3098 0.0013543
R39552 DVSS.n3093 DVSS.n3092 0.0013543
R39553 DVSS.n2822 DVSS.n2821 0.0013543
R39554 DVSS.n2818 DVSS.n2817 0.0013543
R39555 DVSS.n3973 DVSS.n3972 0.0013543
R39556 DVSS.n3760 DVSS.n3759 0.0013543
R39557 DVSS.n11094 DVSS.n11093 0.0013543
R39558 DVSS.n9070 DVSS.n9069 0.0013543
R39559 DVSS.n20427 DVSS.n20426 0.0013543
R39560 DVSS.n20426 DVSS.n20425 0.0013543
R39561 DVSS.n9071 DVSS.n9070 0.0013543
R39562 DVSS.n11093 DVSS.n11092 0.0013543
R39563 DVSS.n16408 DVSS.n16407 0.0013543
R39564 DVSS.n7526 DVSS.n7525 0.0013543
R39565 DVSS.n19419 DVSS.n19418 0.0013543
R39566 DVSS.n19418 DVSS.n19417 0.0013543
R39567 DVSS.n7527 DVSS.n7526 0.0013543
R39568 DVSS.n16409 DVSS.n16408 0.0013543
R39569 DVSS.n6055 DVSS.n6054 0.0013543
R39570 DVSS.n6346 DVSS.n6345 0.0013543
R39571 DVSS.n6822 DVSS.n6821 0.0013543
R39572 DVSS.n3630 DVSS.n3629 0.0013543
R39573 DVSS.n6054 DVSS.n6053 0.0013543
R39574 DVSS.n6335 DVSS.n6334 0.0013543
R39575 DVSS.n6821 DVSS.n6820 0.0013543
R39576 DVSS.n3631 DVSS.n3630 0.0013543
R39577 DVSS.n6347 DVSS.n6346 0.0013543
R39578 DVSS.n3094 DVSS.n3093 0.0013543
R39579 DVSS.n12468 DVSS.n12467 0.0013543
R39580 DVSS.n3100 DVSS.n3099 0.0013543
R39581 DVSS.n12474 DVSS.n12473 0.0013543
R39582 DVSS.n3339 DVSS.n3338 0.0013543
R39583 DVSS.n12716 DVSS.n12715 0.0013543
R39584 DVSS.n2819 DVSS.n2818 0.0013543
R39585 DVSS.n12190 DVSS.n12189 0.0013543
R39586 DVSS.n12194 DVSS.n12193 0.0013543
R39587 DVSS.n2823 DVSS.n2822 0.0013543
R39588 DVSS.n10155 DVSS.n10154 0.00135354
R39589 DVSS.n10154 DVSS.n10153 0.00135354
R39590 DVSS.n10353 DVSS.n10352 0.00134507
R39591 DVSS.n5061 DVSS.n5060 0.00134507
R39592 DVSS.n5247 DVSS.n5246 0.00134507
R39593 DVSS.n5246 DVSS.n5245 0.00134507
R39594 DVSS.n5179 DVSS.n5178 0.00134507
R39595 DVSS.n5164 DVSS.n5163 0.00134507
R39596 DVSS.n5163 DVSS.n5162 0.00134507
R39597 DVSS.n5141 DVSS.n5140 0.00134507
R39598 DVSS.n5110 DVSS.n5109 0.00134507
R39599 DVSS.n5109 DVSS.n5108 0.00134507
R39600 DVSS.n5087 DVSS.n5086 0.00134507
R39601 DVSS.n10354 DVSS.n10350 0.00134507
R39602 DVSS.n10357 DVSS.n10356 0.00134507
R39603 DVSS.n10398 DVSS.n10397 0.00134507
R39604 DVSS.n10424 DVSS.n10423 0.00134507
R39605 DVSS.n10457 DVSS.n10456 0.00134507
R39606 DVSS.n10483 DVSS.n10482 0.00134507
R39607 DVSS.n10500 DVSS.n10499 0.00134507
R39608 DVSS.n10579 DVSS.n10578 0.00134507
R39609 DVSS.n16540 DVSS.n16539 0.00134507
R39610 DVSS.n16543 DVSS.n16542 0.00134507
R39611 DVSS.n16644 DVSS.n16643 0.00134507
R39612 DVSS.n16657 DVSS.n16656 0.00134507
R39613 DVSS.n16671 DVSS.n16670 0.00134507
R39614 DVSS.n16677 DVSS.n16676 0.00134507
R39615 DVSS.n16678 DVSS.n16677 0.00134507
R39616 DVSS.n16680 DVSS.n16679 0.00134507
R39617 DVSS.n17747 DVSS.n17746 0.00134507
R39618 DVSS.n17751 DVSS.n17750 0.00134507
R39619 DVSS.n18154 DVSS.n18153 0.00134507
R39620 DVSS.n18157 DVSS.n18156 0.00134507
R39621 DVSS.n18158 DVSS.n18157 0.00134507
R39622 DVSS.n18213 DVSS.n18212 0.00134507
R39623 DVSS.n18199 DVSS.n18198 0.00134507
R39624 DVSS.n18431 DVSS.n18430 0.00134507
R39625 DVSS.n18444 DVSS.n18443 0.00134507
R39626 DVSS.n14394 DVSS.n14393 0.00134507
R39627 DVSS.n14477 DVSS.n14476 0.00134507
R39628 DVSS.n14481 DVSS.n14480 0.00134507
R39629 DVSS.n19658 DVSS.n19657 0.00134507
R39630 DVSS.n19672 DVSS.n19671 0.00134507
R39631 DVSS.n19748 DVSS.n19747 0.00134507
R39632 DVSS.n16727 DVSS.n16726 0.00134507
R39633 DVSS.n16730 DVSS.n16729 0.00134507
R39634 DVSS.n17179 DVSS.n17178 0.00134507
R39635 DVSS.n17166 DVSS.n17165 0.00134507
R39636 DVSS.n17152 DVSS.n17151 0.00134507
R39637 DVSS.n17146 DVSS.n17145 0.00134507
R39638 DVSS.n17145 DVSS.n17144 0.00134507
R39639 DVSS.n17143 DVSS.n17142 0.00134507
R39640 DVSS.n15916 DVSS.n15915 0.00134507
R39641 DVSS.n15912 DVSS.n15911 0.00134507
R39642 DVSS.n15459 DVSS.n15458 0.00134507
R39643 DVSS.n15462 DVSS.n15461 0.00134507
R39644 DVSS.n15463 DVSS.n15462 0.00134507
R39645 DVSS.n15527 DVSS.n15526 0.00134507
R39646 DVSS.n15541 DVSS.n15540 0.00134507
R39647 DVSS.n15198 DVSS.n15197 0.00134507
R39648 DVSS.n15173 DVSS.n15172 0.00134507
R39649 DVSS.n14756 DVSS.n14755 0.00134507
R39650 DVSS.n14639 DVSS.n14638 0.00134507
R39651 DVSS.n14635 DVSS.n14634 0.00134507
R39652 DVSS.n19867 DVSS.n19866 0.00134507
R39653 DVSS.n19887 DVSS.n19886 0.00134507
R39654 DVSS.n19973 DVSS.n19972 0.00134507
R39655 DVSS.n9169 DVSS.n9168 0.00134497
R39656 DVSS.n9170 DVSS.n9169 0.00134497
R39657 DVSS.n9477 DVSS 0.00134
R39658 DVSS DVSS.n9474 0.00134
R39659 DVSS DVSS.n12110 0.00134
R39660 DVSS.n12109 DVSS 0.00134
R39661 DVSS.n4631 DVSS.n4630 0.00133571
R39662 DVSS.n4969 DVSS.n4968 0.00133571
R39663 DVSS.n4925 DVSS.n4924 0.00133571
R39664 DVSS.n4865 DVSS.n4864 0.00133571
R39665 DVSS.n4633 DVSS.n4632 0.00133571
R39666 DVSS.n4970 DVSS.n4965 0.00133571
R39667 DVSS.n4926 DVSS.n4921 0.00133571
R39668 DVSS.n4866 DVSS.n4861 0.00133571
R39669 DVSS.n4801 DVSS.n4800 0.00133571
R39670 DVSS.n4798 DVSS.n4797 0.00133571
R39671 DVSS.n4753 DVSS.n4752 0.00133571
R39672 DVSS.n6795 DVSS.n6794 0.00133571
R39673 DVSS.n3823 DVSS.n3822 0.00133571
R39674 DVSS.n3910 DVSS.n3909 0.00133571
R39675 DVSS.n3864 DVSS.n3863 0.00133571
R39676 DVSS.n6797 DVSS.n6796 0.00133571
R39677 DVSS.n3825 DVSS.n3824 0.00133571
R39678 DVSS.n3911 DVSS.n3906 0.00133571
R39679 DVSS.n3865 DVSS.n3860 0.00133571
R39680 DVSS.n3602 DVSS.n3601 0.00133571
R39681 DVSS.n2591 DVSS.n2590 0.00133571
R39682 DVSS.n2704 DVSS.n2703 0.00133571
R39683 DVSS.n2650 DVSS.n2649 0.00133571
R39684 DVSS.n3604 DVSS.n3603 0.00133571
R39685 DVSS.n2593 DVSS.n2592 0.00133571
R39686 DVSS.n2705 DVSS.n2700 0.00133571
R39687 DVSS.n2651 DVSS.n2646 0.00133571
R39688 DVSS.n5867 DVSS.n5865 0.00133571
R39689 DVSS.n5988 DVSS.n5987 0.00133571
R39690 DVSS.n5942 DVSS.n5941 0.00133571
R39691 DVSS.n5869 DVSS.n5868 0.00133571
R39692 DVSS.n5989 DVSS.n5984 0.00133571
R39693 DVSS.n5943 DVSS.n5938 0.00133571
R39694 DVSS.n6096 DVSS.n6095 0.00133571
R39695 DVSS.n6242 DVSS.n6237 0.00133571
R39696 DVSS.n6184 DVSS.n6179 0.00133571
R39697 DVSS.n8611 DVSS.n8610 0.00133571
R39698 DVSS.n8614 DVSS.n8613 0.00133571
R39699 DVSS.n8660 DVSS.n8656 0.00133571
R39700 DVSS.n6094 DVSS.n6093 0.00133571
R39701 DVSS.n6241 DVSS.n6240 0.00133571
R39702 DVSS.n6183 DVSS.n6182 0.00133571
R39703 DVSS.n5835 DVSS.n5834 0.00133333
R39704 DVSS.n11029 DVSS.n11028 0.00133333
R39705 DVSS.n6473 DVSS.n6472 0.00133333
R39706 DVSS.n11202 DVSS.n11201 0.00133333
R39707 DVSS.n16675 DVSS.n16674 0.00131688
R39708 DVSS.n17770 DVSS.n17769 0.00131688
R39709 DVSS.n18493 DVSS.n18492 0.00131688
R39710 DVSS.n19760 DVSS.n19759 0.00131688
R39711 DVSS.n164 DVSS.n163 0.00131688
R39712 DVSS.n18183 DVSS.n18182 0.00131688
R39713 DVSS.n18446 DVSS.n18445 0.00131688
R39714 DVSS.n16674 DVSS.n16673 0.00131688
R39715 DVSS.n17769 DVSS.n17768 0.00131688
R39716 DVSS.n14473 DVSS.n14468 0.00131688
R39717 DVSS.n17148 DVSS.n17147 0.00131688
R39718 DVSS.n15893 DVSS.n15892 0.00131688
R39719 DVSS.n15557 DVSS.n15556 0.00131688
R39720 DVSS.n15171 DVSS.n15170 0.00131688
R39721 DVSS.n7734 DVSS.n7733 0.00131688
R39722 DVSS.n19985 DVSS.n19984 0.00131688
R39723 DVSS.n324 DVSS.n323 0.00131688
R39724 DVSS.n14653 DVSS.n14652 0.00131688
R39725 DVSS.n15894 DVSS.n15893 0.00131688
R39726 DVSS.n17149 DVSS.n17148 0.00131688
R39727 DVSS.n14638 DVSS.n14637 0.00131688
R39728 DVSS.n14478 DVSS.n14477 0.00131688
R39729 DVSS.n19759 DVSS.n19758 0.00131688
R39730 DVSS.n19984 DVSS.n19983 0.00131688
R39731 DVSS.n323 DVSS.n322 0.00131688
R39732 DVSS.n163 DVSS.n162 0.00131688
R39733 DVSS.n9225 DVSS.n9224 0.00131498
R39734 DVSS.n9224 DVSS.n9223 0.00131498
R39735 DVSS.n20044 DVSS.n20043 0.00131498
R39736 DVSS.n20045 DVSS.n20044 0.00131498
R39737 DVSS.n468 DVSS.n467 0.00131498
R39738 DVSS.n469 DVSS.n468 0.00131498
R39739 DVSS.n9264 DVSS.n9263 0.00131
R39740 DVSS.n9317 DVSS.n9316 0.00131
R39741 DVSS.n9485 DVSS.n9427 0.00131
R39742 DVSS.n9446 DVSS.n9430 0.00131
R39743 DVSS.n9254 DVSS.n9253 0.00131
R39744 DVSS.n9266 DVSS.n9265 0.00131
R39745 DVSS.n9319 DVSS.n9318 0.00131
R39746 DVSS.n9342 DVSS.n9341 0.00131
R39747 DVSS.n9486 DVSS.n9425 0.00131
R39748 DVSS.n9472 DVSS.n9471 0.00131
R39749 DVSS.n9445 DVSS.n9444 0.00131
R39750 DVSS.n12126 DVSS.n12125 0.00131
R39751 DVSS.n12101 DVSS.n12100 0.00131
R39752 DVSS.n12095 DVSS.n12094 0.00131
R39753 DVSS.n19302 DVSS.n19301 0.00131
R39754 DVSS.n19311 DVSS.n19310 0.00131
R39755 DVSS.n19579 DVSS.n19578 0.00131
R39756 DVSS.n20105 DVSS.n20104 0.00131
R39757 DVSS.n20106 DVSS.n20105 0.00131
R39758 DVSS.n20591 DVSS.n20381 0.00131
R39759 DVSS.n20592 DVSS.n20591 0.00131
R39760 DVSS.n20646 DVSS.n20645 0.00131
R39761 DVSS.n21568 DVSS.n21567 0.00131
R39762 DVSS.n21559 DVSS.n21558 0.00131
R39763 DVSS.n1066 DVSS.n1065 0.00131
R39764 DVSS.n1072 DVSS.n1071 0.00131
R39765 DVSS.n1281 DVSS.n1280 0.00131
R39766 DVSS.n1287 DVSS.n1286 0.00131
R39767 DVSS.n20701 DVSS.n20700 0.00131
R39768 DVSS.n20930 DVSS.n20929 0.00131
R39769 DVSS.n21272 DVSS.n21271 0.00131
R39770 DVSS.n21361 DVSS.n77 0.00131
R39771 DVSS.n21390 DVSS.n21384 0.00131
R39772 DVSS.n20706 DVSS.n20698 0.00131
R39773 DVSS.n20935 DVSS.n20927 0.00131
R39774 DVSS.n21273 DVSS.n21261 0.00131
R39775 DVSS.n21389 DVSS.n21386 0.00131
R39776 DVSS.n20111 DVSS.n20110 0.00131
R39777 DVSS.n20597 DVSS.n20596 0.00131
R39778 DVSS.n20648 DVSS.n20647 0.00131
R39779 DVSS.n21561 DVSS.n21560 0.00131
R39780 DVSS.n13496 DVSS.n13495 0.00131
R39781 DVSS.n7944 DVSS.n7943 0.00131
R39782 DVSS.n12124 DVSS.n11986 0.00131
R39783 DVSS.n12096 DVSS.n12028 0.00131
R39784 DVSS.n9256 DVSS.n9255 0.00128
R39785 DVSS.n9309 DVSS.n9308 0.00128
R39786 DVSS.n9422 DVSS.n9343 0.00128
R39787 DVSS.n9469 DVSS.n9467 0.00128
R39788 DVSS.n9257 DVSS.n9254 0.00128
R39789 DVSS.n9267 DVSS.n9266 0.00128
R39790 DVSS.n9310 DVSS.n9307 0.00128
R39791 DVSS.n9320 DVSS.n9319 0.00128
R39792 DVSS.n9423 DVSS.n9342 0.00128
R39793 DVSS.n9449 DVSS.n9425 0.00128
R39794 DVSS.n9471 DVSS.n9470 0.00128
R39795 DVSS.n9444 DVSS.n9443 0.00128
R39796 DVSS.n13501 DVSS.n13500 0.00128
R39797 DVSS.n13494 DVSS.n13493 0.00128
R39798 DVSS.n13424 DVSS.n13422 0.00128
R39799 DVSS.n7942 DVSS.n7941 0.00128
R39800 DVSS.n12009 DVSS.n12004 0.00128
R39801 DVSS.n12104 DVSS.n12101 0.00128
R39802 DVSS.n20095 DVSS.n20094 0.00128
R39803 DVSS.n20100 DVSS.n20098 0.00128
R39804 DVSS.n20109 DVSS.n20108 0.00128
R39805 DVSS.n20317 DVSS.n20115 0.00128
R39806 DVSS.n20372 DVSS.n20371 0.00128
R39807 DVSS.n20377 DVSS.n20375 0.00128
R39808 DVSS.n20595 DVSS.n20594 0.00128
R39809 DVSS.n20602 DVSS.n20601 0.00128
R39810 DVSS.n20658 DVSS.n20656 0.00128
R39811 DVSS.n21571 DVSS.n21568 0.00128
R39812 DVSS.n21558 DVSS.n21557 0.00128
R39813 DVSS.n20688 DVSS.n20687 0.00128
R39814 DVSS.n20693 DVSS.n20691 0.00128
R39815 DVSS.n20705 DVSS.n20704 0.00128
R39816 DVSS.n20917 DVSS.n20916 0.00128
R39817 DVSS.n20922 DVSS.n20920 0.00128
R39818 DVSS.n20934 DVSS.n20933 0.00128
R39819 DVSS.n21256 DVSS.n21192 0.00128
R39820 DVSS.n21370 DVSS.n77 0.00128
R39821 DVSS.n21384 DVSS.n21383 0.00128
R39822 DVSS.n20695 DVSS.n20685 0.00128
R39823 DVSS.n20924 DVSS.n20915 0.00128
R39824 DVSS.n21258 DVSS.n21122 0.00128
R39825 DVSS.n21369 DVSS.n78 0.00128
R39826 DVSS.n20101 DVSS.n20092 0.00128
R39827 DVSS.n20378 DVSS.n20368 0.00128
R39828 DVSS.n20659 DVSS.n20650 0.00128
R39829 DVSS.n21573 DVSS.n21572 0.00128
R39830 DVSS.n13499 DVSS.n7895 0.00128
R39831 DVSS.n13425 DVSS.n7946 0.00128
R39832 DVSS.n12011 DVSS.n12002 0.00128
R39833 DVSS.n12106 DVSS.n12098 0.00128
R39834 DVSS.n10425 DVSS.n10424 0.00127465
R39835 DVSS.n10484 DVSS.n10483 0.00127465
R39836 DVSS.n10580 DVSS.n10579 0.00127465
R39837 DVSS.n10863 DVSS.n10862 0.00127465
R39838 DVSS.n4763 DVSS.n4761 0.00127143
R39839 DVSS.n4627 DVSS.n4626 0.00127143
R39840 DVSS.n4975 DVSS.n4974 0.00127143
R39841 DVSS.n4931 DVSS.n4930 0.00127143
R39842 DVSS.n4765 DVSS.n4764 0.00127143
R39843 DVSS.n8105 DVSS.n8104 0.00127143
R39844 DVSS.n6790 DVSS.n6789 0.00127143
R39845 DVSS.n3814 DVSS.n3813 0.00127143
R39846 DVSS.n3914 DVSS.n3913 0.00127143
R39847 DVSS.n3868 DVSS.n3867 0.00127143
R39848 DVSS.n8106 DVSS.n8102 0.00127143
R39849 DVSS.n8109 DVSS.n8108 0.00127143
R39850 DVSS.n11782 DVSS.n11781 0.00127143
R39851 DVSS.n3598 DVSS.n3597 0.00127143
R39852 DVSS.n2587 DVSS.n2586 0.00127143
R39853 DVSS.n2709 DVSS.n2708 0.00127143
R39854 DVSS.n2708 DVSS.n2707 0.00127143
R39855 DVSS.n2685 DVSS.n2684 0.00127143
R39856 DVSS.n2655 DVSS.n2654 0.00127143
R39857 DVSS.n2654 DVSS.n2653 0.00127143
R39858 DVSS.n2631 DVSS.n2630 0.00127143
R39859 DVSS.n11783 DVSS.n11779 0.00127143
R39860 DVSS.n11786 DVSS.n11785 0.00127143
R39861 DVSS.n11827 DVSS.n11826 0.00127143
R39862 DVSS.n11853 DVSS.n11852 0.00127143
R39863 DVSS.n11886 DVSS.n11885 0.00127143
R39864 DVSS.n11912 DVSS.n11911 0.00127143
R39865 DVSS.n8397 DVSS.n8396 0.00127143
R39866 DVSS.n5862 DVSS.n5861 0.00127143
R39867 DVSS.n5992 DVSS.n5991 0.00127143
R39868 DVSS.n5946 DVSS.n5945 0.00127143
R39869 DVSS.n8398 DVSS.n8394 0.00127143
R39870 DVSS.n8401 DVSS.n8400 0.00127143
R39871 DVSS.n6089 DVSS.n6088 0.00127143
R39872 DVSS.n6246 DVSS.n6245 0.00127143
R39873 DVSS.n6188 DVSS.n6187 0.00127143
R39874 DVSS.n8649 DVSS.n8644 0.00127143
R39875 DVSS.n8653 DVSS.n8652 0.00127143
R39876 DVSS.n8648 DVSS.n8646 0.00127143
R39877 DVSS.n20748 DVSS.n20747 0.00126575
R39878 DVSS.n20974 DVSS.n20973 0.00126575
R39879 DVSS.n5646 DVSS.n5645 0.00126573
R39880 DVSS.n5745 DVSS.n5744 0.00126573
R39881 DVSS.n4461 DVSS.n4460 0.00126573
R39882 DVSS.n7171 DVSS.n7170 0.00126573
R39883 DVSS.n19254 DVSS.n19253 0.00126573
R39884 DVSS.n873 DVSS.n872 0.00126573
R39885 DVSS.n4460 DVSS.n4459 0.00126573
R39886 DVSS.n5645 DVSS.n5644 0.00126573
R39887 DVSS.n10939 DVSS.n10938 0.00126573
R39888 DVSS.n11253 DVSS.n11252 0.00126573
R39889 DVSS.n11248 DVSS.n11247 0.00126573
R39890 DVSS.n9499 DVSS.n9498 0.00126573
R39891 DVSS.n12910 DVSS.n12909 0.00126573
R39892 DVSS.n12759 DVSS.n12758 0.00126573
R39893 DVSS.n9498 DVSS.n9497 0.00126573
R39894 DVSS.n10938 DVSS.n10937 0.00126573
R39895 DVSS.n11249 DVSS.n11248 0.00126573
R39896 DVSS.n5746 DVSS.n5745 0.00126573
R39897 DVSS.n11252 DVSS.n11251 0.00126573
R39898 DVSS.n17072 DVSS.n17071 0.00126573
R39899 DVSS.n17612 DVSS.n17611 0.00126573
R39900 DVSS.n17617 DVSS.n17616 0.00126573
R39901 DVSS.n15698 DVSS.n15697 0.00126573
R39902 DVSS.n13536 DVSS.n13535 0.00126573
R39903 DVSS.n20265 DVSS.n20264 0.00126573
R39904 DVSS.n20858 DVSS.n20857 0.00126573
R39905 DVSS.n15699 DVSS.n15698 0.00126573
R39906 DVSS.n17613 DVSS.n17612 0.00126573
R39907 DVSS.n17071 DVSS.n17070 0.00126573
R39908 DVSS.n17616 DVSS.n17615 0.00126573
R39909 DVSS.n7170 DVSS.n7155 0.00126573
R39910 DVSS.n13537 DVSS.n13536 0.00126573
R39911 DVSS.n10823 DVSS.n10822 0.00126573
R39912 DVSS.n10785 DVSS.n10784 0.00126573
R39913 DVSS.n11537 DVSS.n11536 0.00126573
R39914 DVSS.n12062 DVSS.n12061 0.00126573
R39915 DVSS.n74 DVSS.n73 0.00126573
R39916 DVSS.n21471 DVSS.n21470 0.00126573
R39917 DVSS.n11536 DVSS.n11535 0.00126573
R39918 DVSS.n10786 DVSS.n10785 0.00126573
R39919 DVSS.n10824 DVSS.n10823 0.00126573
R39920 DVSS.n4716 DVSS.n4715 0.00126573
R39921 DVSS.n4715 DVSS.n4714 0.00126573
R39922 DVSS.n4270 DVSS.n4269 0.00126573
R39923 DVSS.n3734 DVSS.n3733 0.00126573
R39924 DVSS.n2831 DVSS.n2830 0.00126573
R39925 DVSS.n4269 DVSS.n4268 0.00126573
R39926 DVSS.n9961 DVSS.n9960 0.00126573
R39927 DVSS.n11135 DVSS.n11134 0.00126573
R39928 DVSS.n11140 DVSS.n11139 0.00126573
R39929 DVSS.n9695 DVSS.n9694 0.00126573
R39930 DVSS.n13381 DVSS.n13380 0.00126573
R39931 DVSS.n20539 DVSS.n20538 0.00126573
R39932 DVSS.n21084 DVSS.n21083 0.00126573
R39933 DVSS.n13380 DVSS.n13379 0.00126573
R39934 DVSS.n9696 DVSS.n9695 0.00126573
R39935 DVSS.n11136 DVSS.n11135 0.00126573
R39936 DVSS.n9960 DVSS.n9959 0.00126573
R39937 DVSS.n11139 DVSS.n11138 0.00126573
R39938 DVSS.n17365 DVSS.n17364 0.00126573
R39939 DVSS.n16366 DVSS.n16365 0.00126573
R39940 DVSS.n16210 DVSS.n16209 0.00126573
R39941 DVSS.n18839 DVSS.n18838 0.00126573
R39942 DVSS.n19525 DVSS.n19524 0.00126573
R39943 DVSS.n1160 DVSS.n1159 0.00126573
R39944 DVSS.n16367 DVSS.n16366 0.00126573
R39945 DVSS.n18838 DVSS.n18837 0.00126573
R39946 DVSS.n16211 DVSS.n16210 0.00126573
R39947 DVSS.n17364 DVSS.n17363 0.00126573
R39948 DVSS.n5441 DVSS.n5440 0.00126573
R39949 DVSS.n5479 DVSS.n5478 0.00126573
R39950 DVSS.n6584 DVSS.n6583 0.00126573
R39951 DVSS.n3657 DVSS.n3656 0.00126573
R39952 DVSS.n18973 DVSS.n18972 0.00126573
R39953 DVSS.n551 DVSS.n550 0.00126573
R39954 DVSS.n6583 DVSS.n6582 0.00126573
R39955 DVSS.n5440 DVSS.n5439 0.00126573
R39956 DVSS.n5478 DVSS.n5477 0.00126573
R39957 DVSS.n12061 DVSS.n12060 0.00126573
R39958 DVSS.n12911 DVSS.n12910 0.00126573
R39959 DVSS.n3735 DVSS.n3734 0.00126573
R39960 DVSS.n3656 DVSS.n3655 0.00126573
R39961 DVSS.n3372 DVSS.n3371 0.00126573
R39962 DVSS.n73 DVSS.n72 0.00126573
R39963 DVSS.n20538 DVSS.n20537 0.00126573
R39964 DVSS.n20264 DVSS.n20263 0.00126573
R39965 DVSS.n19524 DVSS.n19523 0.00126573
R39966 DVSS.n19253 DVSS.n19252 0.00126573
R39967 DVSS.n18972 DVSS.n18971 0.00126573
R39968 DVSS.n12760 DVSS.n12759 0.00126573
R39969 DVSS.n21472 DVSS.n21471 0.00126573
R39970 DVSS.n12202 DVSS.n12201 0.00126573
R39971 DVSS.n21083 DVSS.n21082 0.00126573
R39972 DVSS.n20857 DVSS.n20856 0.00126573
R39973 DVSS.n1159 DVSS.n1158 0.00126573
R39974 DVSS.n872 DVSS.n871 0.00126573
R39975 DVSS.n2832 DVSS.n2831 0.00126573
R39976 DVSS.n550 DVSS.n549 0.00126573
R39977 DVSS.n9200 DVSS.n9199 0.00125
R39978 DVSS.n1401 DVSS.n1400 0.00125
R39979 DVSS.n4259 DVSS.n4258 0.00125
R39980 DVSS.n4213 DVSS.n4212 0.00125
R39981 DVSS.n4167 DVSS.n4166 0.00125
R39982 DVSS.n3662 DVSS.n3661 0.00125
R39983 DVSS.n3714 DVSS.n3713 0.00125
R39984 DVSS.n18933 DVSS.n18932 0.00125
R39985 DVSS.n19069 DVSS.n19068 0.00125
R39986 DVSS.n19103 DVSS.n19102 0.00125
R39987 DVSS.n19369 DVSS.n19368 0.00125
R39988 DVSS.n20319 DVSS.n20318 0.00125
R39989 DVSS.n20604 DVSS.n20603 0.00125
R39990 DVSS.n623 DVSS.n622 0.00125
R39991 DVSS.n806 DVSS.n805 0.00125
R39992 DVSS.n1057 DVSS.n1056 0.00125
R39993 DVSS.n1272 DVSS.n1271 0.00125
R39994 DVSS.n20864 DVSS.n20863 0.00125
R39995 DVSS.n21090 DVSS.n21089 0.00125
R39996 DVSS.n274 DVSS.n273 0.00125
R39997 DVSS.n19838 DVSS.n19837 0.00125
R39998 DVSS.n14594 DVSS.n14084 0.00125
R39999 DVSS.n4747 DVSS.n4746 0.00122499
R40000 DVSS.n4748 DVSS.n4747 0.00122499
R40001 DVSS.n6136 DVSS.n6135 0.00122499
R40002 DVSS.n6130 DVSS.n6129 0.00122499
R40003 DVSS.n6122 DVSS.n6121 0.00122499
R40004 DVSS.n6116 DVSS.n6115 0.00122499
R40005 DVSS.n6110 DVSS.n6109 0.00122499
R40006 DVSS.n6125 DVSS.n6124 0.00122499
R40007 DVSS.n1398 DVSS.n1396 0.00122
R40008 DVSS.n4256 DVSS.n4239 0.00122
R40009 DVSS.n4210 DVSS.n4208 0.00122
R40010 DVSS.n4164 DVSS.n4161 0.00122
R40011 DVSS.n1400 DVSS.n1399 0.00122
R40012 DVSS.n4258 DVSS.n4257 0.00122
R40013 DVSS.n4212 DVSS.n4211 0.00122
R40014 DVSS.n4166 DVSS.n4165 0.00122
R40015 DVSS.n9204 DVSS.n9203 0.00122
R40016 DVSS.n9207 DVSS.n9206 0.00122
R40017 DVSS.n3664 DVSS.n3662 0.00122
R40018 DVSS.n3727 DVSS.n3726 0.00122
R40019 DVSS.n7238 DVSS.n7237 0.00122
R40020 DVSS.n18897 DVSS.n18896 0.00122
R40021 DVSS.n13488 DVSS.n13487 0.00122
R40022 DVSS.n7934 DVSS.n7933 0.00122
R40023 DVSS.n7911 DVSS.n7910 0.00122
R40024 DVSS.n11998 DVSS.n11997 0.00122
R40025 DVSS.n12004 DVSS.n12003 0.00122
R40026 DVSS.n18935 DVSS.n18933 0.00122
R40027 DVSS.n19057 DVSS.n19055 0.00122
R40028 DVSS.n19101 DVSS.n19100 0.00122
R40029 DVSS.n19367 DVSS.n19366 0.00122
R40030 DVSS.n19843 DVSS.n19842 0.00122
R40031 DVSS.n20616 DVSS.n20615 0.00122
R40032 DVSS.n20653 DVSS.n20652 0.00122
R40033 DVSS.n20656 DVSS.n20655 0.00122
R40034 DVSS.n625 DVSS.n623 0.00122
R40035 DVSS.n722 DVSS.n720 0.00122
R40036 DVSS.n838 DVSS.n837 0.00122
R40037 DVSS.n1125 DVSS.n1124 0.00122
R40038 DVSS.n280 DVSS.n279 0.00122
R40039 DVSS.n21104 DVSS.n21103 0.00122
R40040 DVSS.n21118 DVSS.n21117 0.00122
R40041 DVSS.n21192 DVSS.n21191 0.00122
R40042 DVSS.n627 DVSS.n515 0.00122
R40043 DVSS.n724 DVSS.n685 0.00122
R40044 DVSS.n1062 DVSS.n829 0.00122
R40045 DVSS.n1277 DVSS.n1116 0.00122
R40046 DVSS.n21105 DVSS.n21102 0.00122
R40047 DVSS.n18937 DVSS.n18930 0.00122
R40048 DVSS.n19059 DVSS.n19050 0.00122
R40049 DVSS.n19306 DVSS.n19092 0.00122
R40050 DVSS.n19375 DVSS.n19358 0.00122
R40051 DVSS.n20618 DVSS.n20617 0.00122
R40052 DVSS.n3665 DVSS.n3529 0.00122
R40053 DVSS.n3725 DVSS.n3516 0.00122
R40054 DVSS.n7231 DVSS.n1307 0.00122
R40055 DVSS.n18890 DVSS.n7289 0.00122
R40056 DVSS.n7912 DVSS.n7909 0.00122
R40057 DVSS.n16690 DVSS.n16689 0.00121126
R40058 DVSS.n16701 DVSS.n16700 0.00121126
R40059 DVSS.n16523 DVSS.n16522 0.00121126
R40060 DVSS.n16514 DVSS.n16513 0.00121126
R40061 DVSS.n16505 DVSS.n16504 0.00121126
R40062 DVSS.n17792 DVSS.n17791 0.00121126
R40063 DVSS.n18265 DVSS.n18264 0.00121126
R40064 DVSS.n18191 DVSS.n18190 0.00121126
R40065 DVSS.n14244 DVSS.n14243 0.00121126
R40066 DVSS.n14269 DVSS.n14268 0.00121126
R40067 DVSS.n14294 DVSS.n14293 0.00121126
R40068 DVSS.n14390 DVSS.n14389 0.00121126
R40069 DVSS.n14431 DVSS.n14430 0.00121126
R40070 DVSS.n14464 DVSS.n14463 0.00121126
R40071 DVSS.n19650 DVSS.n19649 0.00121126
R40072 DVSS.n19709 DVSS.n19708 0.00121126
R40073 DVSS.n19720 DVSS.n19719 0.00121126
R40074 DVSS.n19723 DVSS.n19722 0.00121126
R40075 DVSS.n19787 DVSS.n19786 0.00121126
R40076 DVSS.n140 DVSS.n139 0.00121126
R40077 DVSS.n228 DVSS.n227 0.00121126
R40078 DVSS.n192 DVSS.n191 0.00121126
R40079 DVSS.n174 DVSS.n173 0.00121126
R40080 DVSS.n14293 DVSS.n14292 0.00121126
R40081 DVSS.n14268 DVSS.n14267 0.00121126
R40082 DVSS.n14243 DVSS.n14242 0.00121126
R40083 DVSS.n18192 DVSS.n18191 0.00121126
R40084 DVSS.n18266 DVSS.n18265 0.00121126
R40085 DVSS.n18143 DVSS.n18142 0.00121126
R40086 DVSS.n18476 DVSS.n18475 0.00121126
R40087 DVSS.n17736 DVSS.n17735 0.00121126
R40088 DVSS.n17793 DVSS.n17792 0.00121126
R40089 DVSS.n14430 DVSS.n14429 0.00121126
R40090 DVSS.n14463 DVSS.n14462 0.00121126
R40091 DVSS.n14389 DVSS.n14388 0.00121126
R40092 DVSS.n17133 DVSS.n17132 0.00121126
R40093 DVSS.n17122 DVSS.n17121 0.00121126
R40094 DVSS.n16868 DVSS.n16867 0.00121126
R40095 DVSS.n16859 DVSS.n16858 0.00121126
R40096 DVSS.n16851 DVSS.n16850 0.00121126
R40097 DVSS.n17666 DVSS.n17665 0.00121126
R40098 DVSS.n15448 DVSS.n15447 0.00121126
R40099 DVSS.n15475 DVSS.n15474 0.00121126
R40100 DVSS.n15549 DVSS.n15548 0.00121126
R40101 DVSS.n15126 DVSS.n15125 0.00121126
R40102 DVSS.n14863 DVSS.n14862 0.00121126
R40103 DVSS.n14846 DVSS.n14845 0.00121126
R40104 DVSS.n14829 DVSS.n14828 0.00121126
R40105 DVSS.n14761 DVSS.n14760 0.00121126
R40106 DVSS.n14697 DVSS.n14696 0.00121126
R40107 DVSS.n14658 DVSS.n14657 0.00121126
R40108 DVSS.n19859 DVSS.n19858 0.00121126
R40109 DVSS.n19928 DVSS.n19927 0.00121126
R40110 DVSS.n19939 DVSS.n19938 0.00121126
R40111 DVSS.n19942 DVSS.n19941 0.00121126
R40112 DVSS.n20012 DVSS.n20011 0.00121126
R40113 DVSS.n300 DVSS.n299 0.00121126
R40114 DVSS.n436 DVSS.n435 0.00121126
R40115 DVSS.n400 DVSS.n399 0.00121126
R40116 DVSS.n382 DVSS.n381 0.00121126
R40117 DVSS.n15548 DVSS.n15547 0.00121126
R40118 DVSS.n15474 DVSS.n15473 0.00121126
R40119 DVSS.n14864 DVSS.n14863 0.00121126
R40120 DVSS.n14847 DVSS.n14846 0.00121126
R40121 DVSS.n14830 DVSS.n14829 0.00121126
R40122 DVSS.n15927 DVSS.n15926 0.00121126
R40123 DVSS.n17667 DVSS.n17666 0.00121126
R40124 DVSS.n14760 DVSS.n14759 0.00121126
R40125 DVSS.n14698 DVSS.n14697 0.00121126
R40126 DVSS.n14659 DVSS.n14658 0.00121126
R40127 DVSS.n16504 DVSS.n16503 0.00121126
R40128 DVSS.n16850 DVSS.n16849 0.00121126
R40129 DVSS.n16513 DVSS.n16512 0.00121126
R40130 DVSS.n16522 DVSS.n16521 0.00121126
R40131 DVSS.n16691 DVSS.n16690 0.00121126
R40132 DVSS.n17132 DVSS.n17131 0.00121126
R40133 DVSS.n16700 DVSS.n16699 0.00121126
R40134 DVSS.n17123 DVSS.n17122 0.00121126
R40135 DVSS.n16867 DVSS.n16866 0.00121126
R40136 DVSS.n16860 DVSS.n16859 0.00121126
R40137 DVSS.n19938 DVSS.n19937 0.00121126
R40138 DVSS.n19719 DVSS.n19718 0.00121126
R40139 DVSS.n383 DVSS.n382 0.00121126
R40140 DVSS.n175 DVSS.n174 0.00121126
R40141 DVSS.n19941 DVSS.n19940 0.00121126
R40142 DVSS.n19722 DVSS.n19721 0.00121126
R40143 DVSS.n19708 DVSS.n19707 0.00121126
R40144 DVSS.n19927 DVSS.n19926 0.00121126
R40145 DVSS.n19858 DVSS.n19857 0.00121126
R40146 DVSS.n19649 DVSS.n19648 0.00121126
R40147 DVSS.n139 DVSS.n138 0.00121126
R40148 DVSS.n299 DVSS.n298 0.00121126
R40149 DVSS.n20013 DVSS.n20012 0.00121126
R40150 DVSS.n19788 DVSS.n19787 0.00121126
R40151 DVSS.n193 DVSS.n192 0.00121126
R40152 DVSS.n401 DVSS.n400 0.00121126
R40153 DVSS.n437 DVSS.n436 0.00121126
R40154 DVSS.n229 DVSS.n228 0.00121126
R40155 DVSS.n9178 DVSS.n9177 0.00120999
R40156 DVSS.n9179 DVSS.n9178 0.00120999
R40157 DVSS.n5567 DVSS.n5566 0.00120866
R40158 DVSS.n5571 DVSS.n5570 0.00120866
R40159 DVSS.n5628 DVSS.n5627 0.00120866
R40160 DVSS.n6994 DVSS.n6993 0.00120866
R40161 DVSS.n7094 DVSS.n7093 0.00120866
R40162 DVSS.n7175 DVSS.n7174 0.00120866
R40163 DVSS.n7179 DVSS.n7178 0.00120866
R40164 DVSS.n19136 DVSS.n19135 0.00120866
R40165 DVSS.n19150 DVSS.n19149 0.00120866
R40166 DVSS.n19242 DVSS.n19241 0.00120866
R40167 DVSS.n10208 DVSS.n10207 0.00120866
R40168 DVSS.n10211 DVSS.n10210 0.00120866
R40169 DVSS.n10919 DVSS.n10918 0.00120866
R40170 DVSS.n12745 DVSS.n12744 0.00120866
R40171 DVSS.n12721 DVSS.n12720 0.00120866
R40172 DVSS.n12465 DVSS.n12464 0.00120866
R40173 DVSS.n12210 DVSS.n12209 0.00120866
R40174 DVSS.n12207 DVSS.n12206 0.00120866
R40175 DVSS.n21288 DVSS.n21287 0.00120866
R40176 DVSS.n21284 DVSS.n21283 0.00120866
R40177 DVSS.n16953 DVSS.n16952 0.00120866
R40178 DVSS.n16956 DVSS.n16955 0.00120866
R40179 DVSS.n17052 DVSS.n17051 0.00120866
R40180 DVSS.n13644 DVSS.n13643 0.00120866
R40181 DVSS.n13589 DVSS.n13588 0.00120866
R40182 DVSS.n13532 DVSS.n13531 0.00120866
R40183 DVSS.n13528 DVSS.n13527 0.00120866
R40184 DVSS.n20135 DVSS.n20134 0.00120866
R40185 DVSS.n20161 DVSS.n20160 0.00120866
R40186 DVSS.n20252 DVSS.n20251 0.00120866
R40187 DVSS.n10614 DVSS.n10613 0.00120866
R40188 DVSS.n10618 DVSS.n10617 0.00120866
R40189 DVSS.n10843 DVSS.n10842 0.00120866
R40190 DVSS.n11420 DVSS.n11419 0.00120866
R40191 DVSS.n5220 DVSS.n5219 0.00120866
R40192 DVSS.n5224 DVSS.n5223 0.00120866
R40193 DVSS.n5192 DVSS.n5191 0.00120866
R40194 DVSS.n3358 DVSS.n3357 0.00120866
R40195 DVSS.n3344 DVSS.n3343 0.00120866
R40196 DVSS.n3091 DVSS.n3090 0.00120866
R40197 DVSS.n2840 DVSS.n2839 0.00120866
R40198 DVSS.n2837 DVSS.n2836 0.00120866
R40199 DVSS.n738 DVSS.n737 0.00120866
R40200 DVSS.n661 DVSS.n660 0.00120866
R40201 DVSS.n9909 DVSS.n9908 0.00120866
R40202 DVSS.n9912 DVSS.n9911 0.00120866
R40203 DVSS.n9941 DVSS.n9940 0.00120866
R40204 DVSS.n13231 DVSS.n13230 0.00120866
R40205 DVSS.n13243 DVSS.n13242 0.00120866
R40206 DVSS.n13385 DVSS.n13384 0.00120866
R40207 DVSS.n13389 DVSS.n13388 0.00120866
R40208 DVSS.n20418 DVSS.n20417 0.00120866
R40209 DVSS.n20432 DVSS.n20431 0.00120866
R40210 DVSS.n20526 DVSS.n20525 0.00120866
R40211 DVSS.n17262 DVSS.n17261 0.00120866
R40212 DVSS.n17266 DVSS.n17265 0.00120866
R40213 DVSS.n17347 DVSS.n17346 0.00120866
R40214 DVSS.n18761 DVSS.n18760 0.00120866
R40215 DVSS.n18773 DVSS.n18772 0.00120866
R40216 DVSS.n18843 DVSS.n18842 0.00120866
R40217 DVSS.n18847 DVSS.n18846 0.00120866
R40218 DVSS.n19410 DVSS.n19409 0.00120866
R40219 DVSS.n19424 DVSS.n19423 0.00120866
R40220 DVSS.n19513 DVSS.n19512 0.00120866
R40221 DVSS.n5326 DVSS.n5325 0.00120866
R40222 DVSS.n5331 DVSS.n5330 0.00120866
R40223 DVSS.n5423 DVSS.n5422 0.00120866
R40224 DVSS.n6342 DVSS.n6341 0.00120866
R40225 DVSS.n4972 DVSS.n4971 0.00120714
R40226 DVSS.n4928 DVSS.n4927 0.00120714
R40227 DVSS.n4868 DVSS.n4867 0.00120714
R40228 DVSS.n4760 DVSS.n4759 0.00120714
R40229 DVSS.n10088 DVSS.n10087 0.00120714
R40230 DVSS.n10706 DVSS.n10705 0.00120714
R40231 DVSS.n10646 DVSS.n10645 0.00120714
R40232 DVSS.n8168 DVSS.n8167 0.00120714
R40233 DVSS.n8219 DVSS.n8218 0.00120714
R40234 DVSS.n8304 DVSS.n8303 0.00120714
R40235 DVSS.n13090 DVSS.n13089 0.00120714
R40236 DVSS.n11854 DVSS.n11853 0.00120714
R40237 DVSS.n11913 DVSS.n11912 0.00120714
R40238 DVSS.n12982 DVSS.n12981 0.00120714
R40239 DVSS.n13007 DVSS.n13006 0.00120714
R40240 DVSS.n8460 DVSS.n8459 0.00120714
R40241 DVSS.n8511 DVSS.n8510 0.00120714
R40242 DVSS.n11316 DVSS.n11315 0.00120714
R40243 DVSS.n11342 DVSS.n11341 0.00120714
R40244 DVSS.n6244 DVSS.n6243 0.00120714
R40245 DVSS.n6186 DVSS.n6185 0.00120714
R40246 DVSS.n8651 DVSS.n8650 0.00120714
R40247 DVSS.n8723 DVSS.n8722 0.00120714
R40248 DVSS.n8784 DVSS.n8783 0.00120714
R40249 DVSS.n8879 DVSS.n8878 0.00120714
R40250 DVSS.n8325 DVSS.n8324 0.00120714
R40251 DVSS.n10420 DVSS.n10419 0.00120422
R40252 DVSS.n10479 DVSS.n10478 0.00120422
R40253 DVSS.n10575 DVSS.n10573 0.00120422
R40254 DVSS.n10867 DVSS.n10865 0.00120422
R40255 DVSS.n5311 DVSS.n5310 0.00120422
R40256 DVSS.n10421 DVSS.n10417 0.00120422
R40257 DVSS.n10480 DVSS.n10476 0.00120422
R40258 DVSS.n10576 DVSS.n10572 0.00120422
R40259 DVSS.n10873 DVSS.n10872 0.00120422
R40260 DVSS.n10869 DVSS.n10868 0.00120422
R40261 DVSS.n9174 DVSS.n9173 0.00119
R40262 DVSS.n9193 DVSS.n9192 0.00119
R40263 DVSS.n9176 DVSS.n9175 0.00119
R40264 DVSS.n9202 DVSS.n9201 0.00119
R40265 DVSS.n7236 DVSS.n7235 0.00119
R40266 DVSS.n18895 DVSS.n18894 0.00119
R40267 DVSS.n14596 DVSS.n14595 0.00119
R40268 DVSS.n13490 DVSS.n13489 0.00119
R40269 DVSS.n7936 DVSS.n7935 0.00119
R40270 DVSS.n19626 DVSS.n19625 0.00119
R40271 DVSS.n19826 DVSS.n19825 0.00119
R40272 DVSS.n19836 DVSS.n19835 0.00119
R40273 DVSS.n113 DVSS.n112 0.00119
R40274 DVSS.n262 DVSS.n261 0.00119
R40275 DVSS.n272 DVSS.n271 0.00119
R40276 DVSS.n117 DVSS.n110 0.00119
R40277 DVSS.n266 DVSS.n123 0.00119
R40278 DVSS.n19630 DVSS.n19623 0.00119
R40279 DVSS.n19830 DVSS.n19819 0.00119
R40280 DVSS.n14114 DVSS.n14113 0.00119
R40281 DVSS.n14534 DVSS.n14135 0.00119
R40282 DVSS.n4222 DVSS.n4221 0.00117999
R40283 DVSS.n9216 DVSS.n9215 0.00117999
R40284 DVSS.n4223 DVSS.n4222 0.00117999
R40285 DVSS.n9215 DVSS.n9214 0.00117999
R40286 DVSS.n3522 DVSS.n3521 0.00117999
R40287 DVSS.n3690 DVSS.n3689 0.00117999
R40288 DVSS.n3689 DVSS.n3688 0.00117999
R40289 DVSS.n3521 DVSS.n3520 0.00117999
R40290 DVSS.n19044 DVSS.n19043 0.00117999
R40291 DVSS.n19043 DVSS.n19042 0.00117999
R40292 DVSS.n679 DVSS.n652 0.00117999
R40293 DVSS.n652 DVSS.n651 0.00117999
R40294 DVSS.n5658 DVSS.n5657 0.00117716
R40295 DVSS.n5669 DVSS.n5668 0.00117716
R40296 DVSS.n5680 DVSS.n5679 0.00117716
R40297 DVSS.n5690 DVSS.n5689 0.00117716
R40298 DVSS.n5701 DVSS.n5700 0.00117716
R40299 DVSS.n5718 DVSS.n5717 0.00117716
R40300 DVSS.n4435 DVSS.n4434 0.00117716
R40301 DVSS.n4401 DVSS.n4400 0.00117716
R40302 DVSS.n7115 DVSS.n7114 0.00117716
R40303 DVSS.n19127 DVSS.n19126 0.00117716
R40304 DVSS.n19192 DVSS.n19191 0.00117716
R40305 DVSS.n19203 DVSS.n19202 0.00117716
R40306 DVSS.n19206 DVSS.n19205 0.00117716
R40307 DVSS.n19278 DVSS.n19277 0.00117716
R40308 DVSS.n851 DVSS.n850 0.00117716
R40309 DVSS.n1033 DVSS.n1032 0.00117716
R40310 DVSS.n1000 DVSS.n999 0.00117716
R40311 DVSS.n981 DVSS.n980 0.00117716
R40312 DVSS.n4402 DVSS.n4401 0.00117716
R40313 DVSS.n4434 DVSS.n4433 0.00117716
R40314 DVSS.n10951 DVSS.n10950 0.00117716
R40315 DVSS.n10961 DVSS.n10960 0.00117716
R40316 DVSS.n10971 DVSS.n10970 0.00117716
R40317 DVSS.n10980 DVSS.n10979 0.00117716
R40318 DVSS.n10991 DVSS.n10990 0.00117716
R40319 DVSS.n11221 DVSS.n11220 0.00117716
R40320 DVSS.n9527 DVSS.n9526 0.00117716
R40321 DVSS.n9563 DVSS.n9562 0.00117716
R40322 DVSS.n12882 DVSS.n12881 0.00117716
R40323 DVSS.n12846 DVSS.n12845 0.00117716
R40324 DVSS.n12701 DVSS.n12700 0.00117716
R40325 DVSS.n12683 DVSS.n12682 0.00117716
R40326 DVSS.n12480 DVSS.n12479 0.00117716
R40327 DVSS.n12424 DVSS.n12423 0.00117716
R40328 DVSS.n12415 DVSS.n12414 0.00117716
R40329 DVSS.n21237 DVSS.n21236 0.00117716
R40330 DVSS.n21344 DVSS.n21343 0.00117716
R40331 DVSS.n9562 DVSS.n9561 0.00117716
R40332 DVSS.n9526 DVSS.n9525 0.00117716
R40333 DVSS.n11222 DVSS.n11221 0.00117716
R40334 DVSS.n5719 DVSS.n5718 0.00117716
R40335 DVSS.n17084 DVSS.n17083 0.00117716
R40336 DVSS.n17094 DVSS.n17093 0.00117716
R40337 DVSS.n16936 DVSS.n16935 0.00117716
R40338 DVSS.n16927 DVSS.n16926 0.00117716
R40339 DVSS.n16916 DVSS.n16915 0.00117716
R40340 DVSS.n17647 DVSS.n17646 0.00117716
R40341 DVSS.n15670 DVSS.n15669 0.00117716
R40342 DVSS.n15634 DVSS.n15633 0.00117716
R40343 DVSS.n13825 DVSS.n13824 0.00117716
R40344 DVSS.n13787 DVSS.n13786 0.00117716
R40345 DVSS.n13750 DVSS.n13749 0.00117716
R40346 DVSS.n13565 DVSS.n13564 0.00117716
R40347 DVSS.n20127 DVSS.n20126 0.00117716
R40348 DVSS.n20203 DVSS.n20202 0.00117716
R40349 DVSS.n20214 DVSS.n20213 0.00117716
R40350 DVSS.n20217 DVSS.n20216 0.00117716
R40351 DVSS.n20292 DVSS.n20291 0.00117716
R40352 DVSS.n20834 DVSS.n20833 0.00117716
R40353 DVSS.n20798 DVSS.n20797 0.00117716
R40354 DVSS.n20762 DVSS.n20761 0.00117716
R40355 DVSS.n20743 DVSS.n20742 0.00117716
R40356 DVSS.n15635 DVSS.n15634 0.00117716
R40357 DVSS.n15671 DVSS.n15670 0.00117716
R40358 DVSS.n13751 DVSS.n13750 0.00117716
R40359 DVSS.n13788 DVSS.n13787 0.00117716
R40360 DVSS.n13826 DVSS.n13825 0.00117716
R40361 DVSS.n17648 DVSS.n17647 0.00117716
R40362 DVSS.n13566 DVSS.n13565 0.00117716
R40363 DVSS.n7116 DVSS.n7115 0.00117716
R40364 DVSS.n7151 DVSS.n7150 0.00117716
R40365 DVSS.n13542 DVSS.n13541 0.00117716
R40366 DVSS.n6990 DVSS.n6989 0.00117716
R40367 DVSS.n13648 DVSS.n13647 0.00117716
R40368 DVSS.n10809 DVSS.n10808 0.00117716
R40369 DVSS.n10798 DVSS.n10797 0.00117716
R40370 DVSS.n10745 DVSS.n10744 0.00117716
R40371 DVSS.n11565 DVSS.n11564 0.00117716
R40372 DVSS.n11601 DVSS.n11600 0.00117716
R40373 DVSS.n12067 DVSS.n12066 0.00117716
R40374 DVSS.n50 DVSS.n49 0.00117716
R40375 DVSS.n21531 DVSS.n21530 0.00117716
R40376 DVSS.n21495 DVSS.n21494 0.00117716
R40377 DVSS.n21443 DVSS.n21442 0.00117716
R40378 DVSS.n21407 DVSS.n21406 0.00117716
R40379 DVSS.n11600 DVSS.n11599 0.00117716
R40380 DVSS.n11564 DVSS.n11563 0.00117716
R40381 DVSS.n10808 DVSS.n10807 0.00117716
R40382 DVSS.n10746 DVSS.n10745 0.00117716
R40383 DVSS.n5700 DVSS.n5699 0.00117716
R40384 DVSS.n16917 DVSS.n16916 0.00117716
R40385 DVSS.n10990 DVSS.n10989 0.00117716
R40386 DVSS.n5679 DVSS.n5678 0.00117716
R40387 DVSS.n10970 DVSS.n10969 0.00117716
R40388 DVSS.n16937 DVSS.n16936 0.00117716
R40389 DVSS.n5657 DVSS.n5656 0.00117716
R40390 DVSS.n17083 DVSS.n17082 0.00117716
R40391 DVSS.n10950 DVSS.n10949 0.00117716
R40392 DVSS.n10960 DVSS.n10959 0.00117716
R40393 DVSS.n16928 DVSS.n16927 0.00117716
R40394 DVSS.n10979 DVSS.n10978 0.00117716
R40395 DVSS.n10799 DVSS.n10798 0.00117716
R40396 DVSS.n17093 DVSS.n17092 0.00117716
R40397 DVSS.n5668 DVSS.n5667 0.00117716
R40398 DVSS.n5689 DVSS.n5688 0.00117716
R40399 DVSS.n4691 DVSS.n4690 0.00117716
R40400 DVSS.n4681 DVSS.n4680 0.00117716
R40401 DVSS.n4669 DVSS.n4668 0.00117716
R40402 DVSS.n4660 DVSS.n4659 0.00117716
R40403 DVSS.n4648 DVSS.n4647 0.00117716
R40404 DVSS.n4649 DVSS.n4648 0.00117716
R40405 DVSS.n4670 DVSS.n4669 0.00117716
R40406 DVSS.n4692 DVSS.n4691 0.00117716
R40407 DVSS.n4680 DVSS.n4679 0.00117716
R40408 DVSS.n4659 DVSS.n4658 0.00117716
R40409 DVSS.n4296 DVSS.n4295 0.00117716
R40410 DVSS.n4329 DVSS.n4328 0.00117716
R40411 DVSS.n3491 DVSS.n3490 0.00117716
R40412 DVSS.n3458 DVSS.n3457 0.00117716
R40413 DVSS.n3324 DVSS.n3323 0.00117716
R40414 DVSS.n3307 DVSS.n3306 0.00117716
R40415 DVSS.n3106 DVSS.n3105 0.00117716
R40416 DVSS.n3042 DVSS.n3041 0.00117716
R40417 DVSS.n764 DVSS.n763 0.00117716
R40418 DVSS.n768 DVSS.n767 0.00117716
R40419 DVSS.n732 DVSS.n731 0.00117716
R40420 DVSS.n4328 DVSS.n4327 0.00117716
R40421 DVSS.n4295 DVSS.n4294 0.00117716
R40422 DVSS.n19202 DVSS.n19201 0.00117716
R40423 DVSS.n20213 DVSS.n20212 0.00117716
R40424 DVSS.n9973 DVSS.n9972 0.00117716
R40425 DVSS.n9983 DVSS.n9982 0.00117716
R40426 DVSS.n9892 DVSS.n9891 0.00117716
R40427 DVSS.n9883 DVSS.n9882 0.00117716
R40428 DVSS.n9872 DVSS.n9871 0.00117716
R40429 DVSS.n9839 DVSS.n9838 0.00117716
R40430 DVSS.n9667 DVSS.n9666 0.00117716
R40431 DVSS.n9631 DVSS.n9630 0.00117716
R40432 DVSS.n13266 DVSS.n13265 0.00117716
R40433 DVSS.n20410 DVSS.n20409 0.00117716
R40434 DVSS.n20474 DVSS.n20473 0.00117716
R40435 DVSS.n20485 DVSS.n20484 0.00117716
R40436 DVSS.n20488 DVSS.n20487 0.00117716
R40437 DVSS.n20566 DVSS.n20565 0.00117716
R40438 DVSS.n21060 DVSS.n21059 0.00117716
R40439 DVSS.n21024 DVSS.n21023 0.00117716
R40440 DVSS.n20988 DVSS.n20987 0.00117716
R40441 DVSS.n20969 DVSS.n20968 0.00117716
R40442 DVSS.n20484 DVSS.n20483 0.00117716
R40443 DVSS.n9873 DVSS.n9872 0.00117716
R40444 DVSS.n9632 DVSS.n9631 0.00117716
R40445 DVSS.n9668 DVSS.n9667 0.00117716
R40446 DVSS.n9893 DVSS.n9892 0.00117716
R40447 DVSS.n9972 DVSS.n9971 0.00117716
R40448 DVSS.n9884 DVSS.n9883 0.00117716
R40449 DVSS.n9982 DVSS.n9981 0.00117716
R40450 DVSS.n9838 DVSS.n9837 0.00117716
R40451 DVSS.n13227 DVSS.n13226 0.00117716
R40452 DVSS.n13267 DVSS.n13266 0.00117716
R40453 DVSS.n13372 DVSS.n13371 0.00117716
R40454 DVSS.n982 DVSS.n981 0.00117716
R40455 DVSS.n20744 DVSS.n20743 0.00117716
R40456 DVSS.n20970 DVSS.n20969 0.00117716
R40457 DVSS.n17377 DVSS.n17376 0.00117716
R40458 DVSS.n17388 DVSS.n17387 0.00117716
R40459 DVSS.n17399 DVSS.n17398 0.00117716
R40460 DVSS.n17409 DVSS.n17408 0.00117716
R40461 DVSS.n17420 DVSS.n17419 0.00117716
R40462 DVSS.n16331 DVSS.n16330 0.00117716
R40463 DVSS.n16184 DVSS.n16183 0.00117716
R40464 DVSS.n16150 DVSS.n16149 0.00117716
R40465 DVSS.n18607 DVSS.n18606 0.00117716
R40466 DVSS.n18634 DVSS.n18633 0.00117716
R40467 DVSS.n18661 DVSS.n18660 0.00117716
R40468 DVSS.n18795 DVSS.n18794 0.00117716
R40469 DVSS.n19401 DVSS.n19400 0.00117716
R40470 DVSS.n19463 DVSS.n19462 0.00117716
R40471 DVSS.n19474 DVSS.n19473 0.00117716
R40472 DVSS.n19477 DVSS.n19476 0.00117716
R40473 DVSS.n19549 DVSS.n19548 0.00117716
R40474 DVSS.n1138 DVSS.n1137 0.00117716
R40475 DVSS.n1248 DVSS.n1247 0.00117716
R40476 DVSS.n1215 DVSS.n1214 0.00117716
R40477 DVSS.n1197 DVSS.n1196 0.00117716
R40478 DVSS.n19473 DVSS.n19472 0.00117716
R40479 DVSS.n17419 DVSS.n17418 0.00117716
R40480 DVSS.n16151 DVSS.n16150 0.00117716
R40481 DVSS.n18606 DVSS.n18605 0.00117716
R40482 DVSS.n18633 DVSS.n18632 0.00117716
R40483 DVSS.n18660 DVSS.n18659 0.00117716
R40484 DVSS.n18794 DVSS.n18793 0.00117716
R40485 DVSS.n16185 DVSS.n16184 0.00117716
R40486 DVSS.n17398 DVSS.n17397 0.00117716
R40487 DVSS.n17376 DVSS.n17375 0.00117716
R40488 DVSS.n17387 DVSS.n17386 0.00117716
R40489 DVSS.n17408 DVSS.n17407 0.00117716
R40490 DVSS.n16330 DVSS.n16329 0.00117716
R40491 DVSS.n18757 DVSS.n18756 0.00117716
R40492 DVSS.n18833 DVSS.n18832 0.00117716
R40493 DVSS.n1198 DVSS.n1197 0.00117716
R40494 DVSS.n5454 DVSS.n5453 0.00117716
R40495 DVSS.n5466 DVSS.n5465 0.00117716
R40496 DVSS.n5849 DVSS.n5848 0.00117716
R40497 DVSS.n6610 DVSS.n6609 0.00117716
R40498 DVSS.n6644 DVSS.n6643 0.00117716
R40499 DVSS.n3553 DVSS.n3552 0.00117716
R40500 DVSS.n18951 DVSS.n18950 0.00117716
R40501 DVSS.n18997 DVSS.n18996 0.00117716
R40502 DVSS.n529 DVSS.n528 0.00117716
R40503 DVSS.n599 DVSS.n598 0.00117716
R40504 DVSS.n566 DVSS.n565 0.00117716
R40505 DVSS.n6643 DVSS.n6642 0.00117716
R40506 DVSS.n6609 DVSS.n6608 0.00117716
R40507 DVSS.n5465 DVSS.n5464 0.00117716
R40508 DVSS.n5455 DVSS.n5454 0.00117716
R40509 DVSS.n5848 DVSS.n5847 0.00117716
R40510 DVSS.n18950 DVSS.n18949 0.00117716
R40511 DVSS.n20487 DVSS.n20486 0.00117716
R40512 DVSS.n20216 DVSS.n20215 0.00117716
R40513 DVSS.n19476 DVSS.n19475 0.00117716
R40514 DVSS.n19205 DVSS.n19204 0.00117716
R40515 DVSS.n3459 DVSS.n3458 0.00117716
R40516 DVSS.n19191 DVSS.n19190 0.00117716
R40517 DVSS.n19462 DVSS.n19461 0.00117716
R40518 DVSS.n20473 DVSS.n20472 0.00117716
R40519 DVSS.n12847 DVSS.n12846 0.00117716
R40520 DVSS.n49 DVSS.n48 0.00117716
R40521 DVSS.n20202 DVSS.n20201 0.00117716
R40522 DVSS.n19400 DVSS.n19399 0.00117716
R40523 DVSS.n12068 DVSS.n12067 0.00117716
R40524 DVSS.n12883 DVSS.n12882 0.00117716
R40525 DVSS.n20409 DVSS.n20408 0.00117716
R40526 DVSS.n20126 DVSS.n20125 0.00117716
R40527 DVSS.n19126 DVSS.n19125 0.00117716
R40528 DVSS.n3492 DVSS.n3491 0.00117716
R40529 DVSS.n3554 DVSS.n3553 0.00117716
R40530 DVSS.n528 DVSS.n527 0.00117716
R40531 DVSS.n3325 DVSS.n3324 0.00117716
R40532 DVSS.n3051 DVSS.n3050 0.00117716
R40533 DVSS.n1137 DVSS.n1136 0.00117716
R40534 DVSS.n12702 DVSS.n12701 0.00117716
R40535 DVSS.n12425 DVSS.n12424 0.00117716
R40536 DVSS.n21496 DVSS.n21495 0.00117716
R40537 DVSS.n850 DVSS.n849 0.00117716
R40538 DVSS.n21532 DVSS.n21531 0.00117716
R40539 DVSS.n12684 DVSS.n12683 0.00117716
R40540 DVSS.n20567 DVSS.n20566 0.00117716
R40541 DVSS.n20293 DVSS.n20292 0.00117716
R40542 DVSS.n19550 DVSS.n19549 0.00117716
R40543 DVSS.n19279 DVSS.n19278 0.00117716
R40544 DVSS.n18998 DVSS.n18997 0.00117716
R40545 DVSS.n12481 DVSS.n12480 0.00117716
R40546 DVSS.n3043 DVSS.n3042 0.00117716
R40547 DVSS.n12416 DVSS.n12415 0.00117716
R40548 DVSS.n21059 DVSS.n21058 0.00117716
R40549 DVSS.n20833 DVSS.n20832 0.00117716
R40550 DVSS.n567 DVSS.n566 0.00117716
R40551 DVSS.n1216 DVSS.n1215 0.00117716
R40552 DVSS.n21444 DVSS.n21443 0.00117716
R40553 DVSS.n21233 DVSS.n21232 0.00117716
R40554 DVSS.n21025 DVSS.n21024 0.00117716
R40555 DVSS.n20799 DVSS.n20798 0.00117716
R40556 DVSS.n1249 DVSS.n1248 0.00117716
R40557 DVSS.n1034 DVSS.n1033 0.00117716
R40558 DVSS.n768 DVSS.n764 0.00117716
R40559 DVSS.n763 DVSS.n762 0.00117716
R40560 DVSS.n600 DVSS.n599 0.00117716
R40561 DVSS.n21408 DVSS.n21407 0.00117716
R40562 DVSS.n20989 DVSS.n20988 0.00117716
R40563 DVSS.n20763 DVSS.n20762 0.00117716
R40564 DVSS.n1001 DVSS.n1000 0.00117716
R40565 DVSS.n731 DVSS.n730 0.00117716
R40566 DVSS.n15426 DVSS.n15425 0.001175
R40567 DVSS.n18286 DVSS.n18285 0.001175
R40568 DVSS.n18335 DVSS.n18334 0.001175
R40569 DVSS.n18340 DVSS.n18339 0.001175
R40570 DVSS.n9277 DVSS.n9276 0.00116499
R40571 DVSS.n9459 DVSS.n9458 0.00116499
R40572 DVSS.n9433 DVSS.n9432 0.00116499
R40573 DVSS.n9458 DVSS.n9457 0.00116499
R40574 DVSS.n9276 DVSS.n9275 0.00116499
R40575 DVSS.n9434 DVSS.n9433 0.00116499
R40576 DVSS.n20323 DVSS.n20322 0.00116499
R40577 DVSS.n20608 DVSS.n20607 0.00116499
R40578 DVSS.n20631 DVSS.n20630 0.00116499
R40579 DVSS.n8 DVSS.n7 0.00116499
R40580 DVSS.n20632 DVSS.n20631 0.00116499
R40581 DVSS.n9 DVSS.n8 0.00116499
R40582 DVSS.n20609 DVSS.n20608 0.00116499
R40583 DVSS.n20324 DVSS.n20323 0.00116499
R40584 DVSS.n20868 DVSS.n20867 0.00116499
R40585 DVSS.n21094 DVSS.n21093 0.00116499
R40586 DVSS.n21314 DVSS.n21313 0.00116499
R40587 DVSS.n21374 DVSS.n21373 0.00116499
R40588 DVSS.n21345 DVSS.n21314 0.00116499
R40589 DVSS.n21375 DVSS.n21374 0.00116499
R40590 DVSS.n21095 DVSS.n21094 0.00116499
R40591 DVSS.n20869 DVSS.n20868 0.00116499
R40592 DVSS.n4809 DVSS.n4808 0.00116071
R40593 DVSS.n4787 DVSS.n4786 0.00116071
R40594 DVSS.n4810 DVSS.n4809 0.00116071
R40595 DVSS.n4788 DVSS.n4787 0.00116071
R40596 DVSS.n9190 DVSS.n9189 0.00116
R40597 DVSS.n7229 DVSS.n7227 0.00116
R40598 DVSS.n18889 DVSS.n18887 0.00116
R40599 DVSS.n13472 DVSS.n13471 0.00116
R40600 DVSS.n7940 DVSS.n7939 0.00116
R40601 DVSS.n7918 DVSS.n7917 0.00116
R40602 DVSS.n19304 DVSS.n19104 0.00116
R40603 DVSS.n19373 DVSS.n19370 0.00116
R40604 DVSS.n19823 DVSS.n19822 0.00116
R40605 DVSS.n1060 DVSS.n1058 0.00116
R40606 DVSS.n1275 DVSS.n1273 0.00116
R40607 DVSS.n259 DVSS.n258 0.00116
R40608 DVSS.n2005 DVSS.n2004 0.00114286
R40609 DVSS.n2333 DVSS.n2332 0.00114286
R40610 DVSS.n2334 DVSS.n2044 0.00114286
R40611 DVSS.n2006 DVSS.n2002 0.00114286
R40612 DVSS.n10104 DVSS.n10103 0.00114286
R40613 DVSS.n10149 DVSS.n10148 0.00114286
R40614 DVSS.n10700 DVSS.n10698 0.00114286
R40615 DVSS.n10651 DVSS.n10648 0.00114286
R40616 DVSS.n4637 DVSS.n4636 0.00114286
R40617 DVSS.n10083 DVSS.n10082 0.00114286
R40618 DVSS.n10085 DVSS.n10084 0.00114286
R40619 DVSS.n10150 DVSS.n10143 0.00114286
R40620 DVSS.n10152 DVSS.n10151 0.00114286
R40621 DVSS.n10701 DVSS.n10697 0.00114286
R40622 DVSS.n10703 DVSS.n10702 0.00114286
R40623 DVSS.n10657 DVSS.n10656 0.00114286
R40624 DVSS.n10653 DVSS.n10652 0.00114286
R40625 DVSS.n8164 DVSS.n8163 0.00114286
R40626 DVSS.n8215 DVSS.n8214 0.00114286
R40627 DVSS.n8300 DVSS.n8298 0.00114286
R40628 DVSS.n13094 DVSS.n13092 0.00114286
R40629 DVSS.n8165 DVSS.n8161 0.00114286
R40630 DVSS.n8216 DVSS.n8212 0.00114286
R40631 DVSS.n8301 DVSS.n8297 0.00114286
R40632 DVSS.n13096 DVSS.n13095 0.00114286
R40633 DVSS.n11849 DVSS.n11848 0.00114286
R40634 DVSS.n11908 DVSS.n11907 0.00114286
R40635 DVSS.n12986 DVSS.n12984 0.00114286
R40636 DVSS.n13011 DVSS.n13009 0.00114286
R40637 DVSS.n11850 DVSS.n11846 0.00114286
R40638 DVSS.n11909 DVSS.n11905 0.00114286
R40639 DVSS.n12988 DVSS.n12987 0.00114286
R40640 DVSS.n13013 DVSS.n13012 0.00114286
R40641 DVSS.n8456 DVSS.n8455 0.00114286
R40642 DVSS.n8507 DVSS.n8506 0.00114286
R40643 DVSS.n11320 DVSS.n11318 0.00114286
R40644 DVSS.n11346 DVSS.n11344 0.00114286
R40645 DVSS.n6049 DVSS.n6048 0.00114286
R40646 DVSS.n8457 DVSS.n8453 0.00114286
R40647 DVSS.n8508 DVSS.n8504 0.00114286
R40648 DVSS.n11322 DVSS.n11321 0.00114286
R40649 DVSS.n11352 DVSS.n11351 0.00114286
R40650 DVSS.n11348 DVSS.n11347 0.00114286
R40651 DVSS.n6100 DVSS.n6099 0.00114286
R40652 DVSS.n8719 DVSS.n8715 0.00114286
R40653 DVSS.n8721 DVSS.n8720 0.00114286
R40654 DVSS.n8780 DVSS.n8776 0.00114286
R40655 DVSS.n8782 DVSS.n8781 0.00114286
R40656 DVSS.n8875 DVSS.n8871 0.00114286
R40657 DVSS.n8877 DVSS.n8876 0.00114286
R40658 DVSS.n8905 DVSS.n8336 0.00114286
R40659 DVSS.n8333 DVSS.n8332 0.00114286
R40660 DVSS.n8718 DVSS.n8717 0.00114286
R40661 DVSS.n8779 DVSS.n8778 0.00114286
R40662 DVSS.n8874 DVSS.n8872 0.00114286
R40663 DVSS.n8331 DVSS.n8327 0.00114286
R40664 DVSS.n3705 DVSS.n3702 0.00114
R40665 DVSS.n19082 DVSS.n19081 0.00114
R40666 DVSS.n819 DVSS.n818 0.00114
R40667 DVSS.n16532 DVSS.n16531 0.0011338
R40668 DVSS.n16580 DVSS.n16579 0.0011338
R40669 DVSS.n16586 DVSS.n16585 0.0011338
R40670 DVSS.n16071 DVSS.n16070 0.0011338
R40671 DVSS.n17767 DVSS.n17766 0.0011338
R40672 DVSS.n18119 DVSS.n18118 0.0011338
R40673 DVSS.n18152 DVSS.n18151 0.0011338
R40674 DVSS.n18262 DVSS.n18261 0.0011338
R40675 DVSS.n18205 DVSS.n18204 0.0011338
R40676 DVSS.n18200 DVSS.n18199 0.0011338
R40677 DVSS.n18195 DVSS.n18194 0.0011338
R40678 DVSS.n18186 DVSS.n18185 0.0011338
R40679 DVSS.n18433 DVSS.n18432 0.0011338
R40680 DVSS.n18436 DVSS.n18435 0.0011338
R40681 DVSS.n18450 DVSS.n18449 0.0011338
R40682 DVSS.n18488 DVSS.n18487 0.0011338
R40683 DVSS.n18496 DVSS.n18495 0.0011338
R40684 DVSS.n14422 DVSS.n14421 0.0011338
R40685 DVSS.n14501 DVSS.n14500 0.0011338
R40686 DVSS.n16719 DVSS.n16718 0.0011338
R40687 DVSS.n16767 DVSS.n16766 0.0011338
R40688 DVSS.n16773 DVSS.n16772 0.0011338
R40689 DVSS.n15963 DVSS.n15962 0.0011338
R40690 DVSS.n15896 DVSS.n15895 0.0011338
R40691 DVSS.n15409 DVSS.n15408 0.0011338
R40692 DVSS.n15457 DVSS.n15456 0.0011338
R40693 DVSS.n15478 DVSS.n15477 0.0011338
R40694 DVSS.n15535 DVSS.n15534 0.0011338
R40695 DVSS.n15540 DVSS.n15539 0.0011338
R40696 DVSS.n15545 DVSS.n15544 0.0011338
R40697 DVSS.n15554 DVSS.n15553 0.0011338
R40698 DVSS.n15196 DVSS.n15195 0.0011338
R40699 DVSS.n15193 DVSS.n15192 0.0011338
R40700 DVSS.n15167 DVSS.n15166 0.0011338
R40701 DVSS.n7729 DVSS.n7728 0.0011338
R40702 DVSS.n7737 DVSS.n7736 0.0011338
R40703 DVSS.n14706 DVSS.n14705 0.0011338
R40704 DVSS.n14621 DVSS.n14620 0.0011338
R40705 DVSS.n9220 DVSS.n9218 0.00113
R40706 DVSS.n9187 DVSS.n9186 0.00113
R40707 DVSS.n9221 DVSS.n9217 0.00113
R40708 DVSS.n3719 DVSS.n3718 0.00113
R40709 DVSS.n7223 DVSS.n7222 0.00113
R40710 DVSS.n7226 DVSS.n7225 0.00113
R40711 DVSS.n18883 DVSS.n18882 0.00113
R40712 DVSS.n18886 DVSS.n18885 0.00113
R40713 DVSS.n12006 DVSS.n12005 0.00113
R40714 DVSS.n19062 DVSS.n19061 0.00113
R40715 DVSS.n20640 DVSS.n20639 0.00113
R40716 DVSS.n791 DVSS.n726 0.00113
R40717 DVSS.n21253 DVSS.n21238 0.00113
R40718 DVSS.n473 DVSS.n287 0.00113
R40719 DVSS.n20048 DVSS.n19851 0.00113
R40720 DVSS.n14580 DVSS.n14565 0.00113
R40721 DVSS.n5351 DVSS.n5332 0.00112569
R40722 DVSS.n1370 DVSS.n1369 0.00112569
R40723 DVSS.n5351 DVSS.n5350 0.00112569
R40724 DVSS.n1369 DVSS.n1368 0.00112569
R40725 DVSS.n16551 DVSS.n16550 0.00110563
R40726 DVSS.n16583 DVSS.n16582 0.00110563
R40727 DVSS.n16685 DVSS.n16684 0.00110563
R40728 DVSS.n17784 DVSS.n17783 0.00110563
R40729 DVSS.n18249 DVSS.n18248 0.00110563
R40730 DVSS.n18207 DVSS.n18206 0.00110563
R40731 DVSS.n14262 DVSS.n14261 0.00110563
R40732 DVSS.n14287 DVSS.n14286 0.00110563
R40733 DVSS.n14316 DVSS.n14315 0.00110563
R40734 DVSS.n14403 DVSS.n14402 0.00110563
R40735 DVSS.n14450 DVSS.n14449 0.00110563
R40736 DVSS.n14498 DVSS.n14497 0.00110563
R40737 DVSS.n19703 DVSS.n19702 0.00110563
R40738 DVSS.n19781 DVSS.n19780 0.00110563
R40739 DVSS.n134 DVSS.n133 0.00110563
R40740 DVSS.n222 DVSS.n221 0.00110563
R40741 DVSS.n198 DVSS.n197 0.00110563
R40742 DVSS.n18250 DVSS.n18249 0.00110563
R40743 DVSS.n18114 DVSS.n18113 0.00110563
R40744 DVSS.n18208 DVSS.n18207 0.00110563
R40745 DVSS.n14261 DVSS.n14260 0.00110563
R40746 DVSS.n14286 DVSS.n14285 0.00110563
R40747 DVSS.n14315 DVSS.n14314 0.00110563
R40748 DVSS.n16684 DVSS.n16683 0.00110563
R40749 DVSS.n16552 DVSS.n16551 0.00110563
R40750 DVSS.n17783 DVSS.n17782 0.00110563
R40751 DVSS.n14449 DVSS.n14448 0.00110563
R40752 DVSS.n14497 DVSS.n14492 0.00110563
R40753 DVSS.n14404 DVSS.n14403 0.00110563
R40754 DVSS.n16739 DVSS.n16738 0.00110563
R40755 DVSS.n17139 DVSS.n17138 0.00110563
R40756 DVSS.n15879 DVSS.n15878 0.00110563
R40757 DVSS.n15491 DVSS.n15490 0.00110563
R40758 DVSS.n15533 DVSS.n15532 0.00110563
R40759 DVSS.n14853 DVSS.n14852 0.00110563
R40760 DVSS.n14836 DVSS.n14835 0.00110563
R40761 DVSS.n14819 DVSS.n14818 0.00110563
R40762 DVSS.n14724 DVSS.n14723 0.00110563
R40763 DVSS.n14672 DVSS.n14671 0.00110563
R40764 DVSS.n14631 DVSS.n14630 0.00110563
R40765 DVSS.n19922 DVSS.n19921 0.00110563
R40766 DVSS.n20006 DVSS.n20005 0.00110563
R40767 DVSS.n294 DVSS.n293 0.00110563
R40768 DVSS.n430 DVSS.n429 0.00110563
R40769 DVSS.n406 DVSS.n405 0.00110563
R40770 DVSS.n14725 DVSS.n14724 0.00110563
R40771 DVSS.n15532 DVSS.n15531 0.00110563
R40772 DVSS.n15490 DVSS.n15489 0.00110563
R40773 DVSS.n15404 DVSS.n15403 0.00110563
R40774 DVSS.n14854 DVSS.n14853 0.00110563
R40775 DVSS.n14837 DVSS.n14836 0.00110563
R40776 DVSS.n14820 DVSS.n14819 0.00110563
R40777 DVSS.n16770 DVSS.n16769 0.00110563
R40778 DVSS.n16738 DVSS.n16737 0.00110563
R40779 DVSS.n17138 DVSS.n17137 0.00110563
R40780 DVSS.n15880 DVSS.n15879 0.00110563
R40781 DVSS.n14673 DVSS.n14672 0.00110563
R40782 DVSS.n14630 DVSS.n14623 0.00110563
R40783 DVSS.n19921 DVSS.n19920 0.00110563
R40784 DVSS.n19702 DVSS.n19701 0.00110563
R40785 DVSS.n19865 DVSS.n19864 0.00110563
R40786 DVSS.n19656 DVSS.n19655 0.00110563
R40787 DVSS.n19782 DVSS.n19781 0.00110563
R40788 DVSS.n20007 DVSS.n20006 0.00110563
R40789 DVSS.n293 DVSS.n292 0.00110563
R40790 DVSS.n133 DVSS.n132 0.00110563
R40791 DVSS.n223 DVSS.n222 0.00110563
R40792 DVSS.n431 DVSS.n430 0.00110563
R40793 DVSS.n407 DVSS.n406 0.00110563
R40794 DVSS.n199 DVSS.n198 0.00110563
R40795 DVSS.n14576 DVSS.n14575 0.001105
R40796 DVSS.n14577 DVSS.n14576 0.001105
R40797 DVSS.n14121 DVSS.n14120 0.0011
R40798 DVSS.n14528 DVSS.n14527 0.0011
R40799 DVSS.n14599 DVSS.n14598 0.0011
R40800 DVSS.n14575 DVSS.n14574 0.0011
R40801 DVSS.n4962 DVSS.n4961 0.00109643
R40802 DVSS.n4919 DVSS.n4918 0.00109643
R40803 DVSS.n4858 DVSS.n4857 0.00109643
R40804 DVSS.n4768 DVSS.n4767 0.00109643
R40805 DVSS.n4918 DVSS.n4917 0.00109643
R40806 DVSS.n4769 DVSS.n4768 0.00109643
R40807 DVSS.n4963 DVSS.n4962 0.00109643
R40808 DVSS.n4859 DVSS.n4858 0.00109643
R40809 DVSS.n5609 DVSS.n5601 0.00108858
R40810 DVSS.n5662 DVSS.n5661 0.00108858
R40811 DVSS.n5672 DVSS.n5671 0.00108858
R40812 DVSS.n5684 DVSS.n5683 0.00108858
R40813 DVSS.n5694 DVSS.n5693 0.00108858
R40814 DVSS.n5729 DVSS.n5728 0.00108858
R40815 DVSS.n4428 DVSS.n4427 0.00108858
R40816 DVSS.n4408 DVSS.n4407 0.00108858
R40817 DVSS.n4407 DVSS.n4406 0.00108858
R40818 DVSS.n4429 DVSS.n4428 0.00108858
R40819 DVSS.n5695 DVSS.n5694 0.00108858
R40820 DVSS.n5673 DVSS.n5672 0.00108858
R40821 DVSS.n5661 DVSS.n5660 0.00108858
R40822 DVSS.n5610 DVSS.n5609 0.00108858
R40823 DVSS.n5730 DVSS.n5729 0.00108858
R40824 DVSS.n10293 DVSS.n10292 0.00108858
R40825 DVSS.n12876 DVSS.n12875 0.00108858
R40826 DVSS.n10292 DVSS.n10284 0.00108858
R40827 DVSS.n17032 DVSS.n17031 0.00108858
R40828 DVSS.n20749 DVSS.n20748 0.00108858
R40829 DVSS.n17031 DVSS.n17023 0.00108858
R40830 DVSS.n5233 DVSS.n5232 0.00108858
R40831 DVSS.n4665 DVSS.n4664 0.00108858
R40832 DVSS.n4654 DVSS.n4653 0.00108858
R40833 DVSS.n4655 DVSS.n4654 0.00108858
R40834 DVSS.n5232 DVSS.n5231 0.00108858
R40835 DVSS.n9921 DVSS.n9920 0.00108858
R40836 DVSS.n20975 DVSS.n20974 0.00108858
R40837 DVSS.n9920 DVSS.n9919 0.00108858
R40838 DVSS.n17329 DVSS.n17328 0.00108858
R40839 DVSS.n17380 DVSS.n17379 0.00108858
R40840 DVSS.n17403 DVSS.n17402 0.00108858
R40841 DVSS.n17414 DVSS.n17413 0.00108858
R40842 DVSS.n1204 DVSS.n1203 0.00108858
R40843 DVSS.n17413 DVSS.n17412 0.00108858
R40844 DVSS.n17328 DVSS.n17319 0.00108858
R40845 DVSS.n17381 DVSS.n17380 0.00108858
R40846 DVSS.n12877 DVSS.n12876 0.00108858
R40847 DVSS.n1203 DVSS.n1202 0.00108858
R40848 DVSS.n5652 DVSS.n5651 0.00108858
R40849 DVSS.n5747 DVSS.n5746 0.00108858
R40850 DVSS.n5738 DVSS.n5737 0.00108858
R40851 DVSS.n5725 DVSS.n5724 0.00108858
R40852 DVSS.n5715 DVSS.n5714 0.00108858
R40853 DVSS.n6509 DVSS.n6508 0.00108858
R40854 DVSS.n7138 DVSS.n7137 0.00108858
R40855 DVSS.n19186 DVSS.n19185 0.00108858
R40856 DVSS.n19272 DVSS.n19271 0.00108858
R40857 DVSS.n845 DVSS.n844 0.00108858
R40858 DVSS.n1027 DVSS.n1026 0.00108858
R40859 DVSS.n1006 DVSS.n1005 0.00108858
R40860 DVSS.n987 DVSS.n986 0.00108858
R40861 DVSS.n5651 DVSS.n5650 0.00108858
R40862 DVSS.n10945 DVSS.n10944 0.00108858
R40863 DVSS.n10975 DVSS.n10974 0.00108858
R40864 DVSS.n11232 DVSS.n11231 0.00108858
R40865 DVSS.n11219 DVSS.n11218 0.00108858
R40866 DVSS.n9767 DVSS.n9766 0.00108858
R40867 DVSS.n9533 DVSS.n9532 0.00108858
R40868 DVSS.n9557 DVSS.n9556 0.00108858
R40869 DVSS.n12852 DVSS.n12851 0.00108858
R40870 DVSS.n12694 DVSS.n12693 0.00108858
R40871 DVSS.n12491 DVSS.n12490 0.00108858
R40872 DVSS.n12163 DVSS.n12162 0.00108858
R40873 DVSS.n21293 DVSS.n21292 0.00108858
R40874 DVSS.n21299 DVSS.n21298 0.00108858
R40875 DVSS.n9532 DVSS.n9531 0.00108858
R40876 DVSS.n9556 DVSS.n9555 0.00108858
R40877 DVSS.n10954 DVSS.n10953 0.00108858
R40878 DVSS.n10964 DVSS.n10963 0.00108858
R40879 DVSS.n10944 DVSS.n10943 0.00108858
R40880 DVSS.n10984 DVSS.n10983 0.00108858
R40881 DVSS.n11233 DVSS.n11232 0.00108858
R40882 DVSS.n6508 DVSS.n6507 0.00108858
R40883 DVSS.n11241 DVSS.n11240 0.00108858
R40884 DVSS.n5748 DVSS.n5747 0.00108858
R40885 DVSS.n11250 DVSS.n11249 0.00108858
R40886 DVSS.n5739 DVSS.n5738 0.00108858
R40887 DVSS.n5726 DVSS.n5725 0.00108858
R40888 DVSS.n11228 DVSS.n11227 0.00108858
R40889 DVSS.n5716 DVSS.n5715 0.00108858
R40890 DVSS.n17078 DVSS.n17077 0.00108858
R40891 DVSS.n17633 DVSS.n17632 0.00108858
R40892 DVSS.n17650 DVSS.n17649 0.00108858
R40893 DVSS.n15664 DVSS.n15663 0.00108858
R40894 DVSS.n15640 DVSS.n15639 0.00108858
R40895 DVSS.n13794 DVSS.n13793 0.00108858
R40896 DVSS.n13757 DVSS.n13756 0.00108858
R40897 DVSS.n13709 DVSS.n13708 0.00108858
R40898 DVSS.n13555 DVSS.n13554 0.00108858
R40899 DVSS.n20197 DVSS.n20196 0.00108858
R40900 DVSS.n20286 DVSS.n20285 0.00108858
R40901 DVSS.n20828 DVSS.n20827 0.00108858
R40902 DVSS.n20792 DVSS.n20791 0.00108858
R40903 DVSS.n20768 DVSS.n20767 0.00108858
R40904 DVSS.n15665 DVSS.n15664 0.00108858
R40905 DVSS.n15641 DVSS.n15640 0.00108858
R40906 DVSS.n15868 DVSS.n15867 0.00108858
R40907 DVSS.n13795 DVSS.n13794 0.00108858
R40908 DVSS.n13758 DVSS.n13757 0.00108858
R40909 DVSS.n13710 DVSS.n13709 0.00108858
R40910 DVSS.n17632 DVSS.n17631 0.00108858
R40911 DVSS.n17077 DVSS.n17076 0.00108858
R40912 DVSS.n17087 DVSS.n17086 0.00108858
R40913 DVSS.n17097 DVSS.n17096 0.00108858
R40914 DVSS.n16923 DVSS.n16922 0.00108858
R40915 DVSS.n17615 DVSS.n17614 0.00108858
R40916 DVSS.n17624 DVSS.n17623 0.00108858
R40917 DVSS.n17637 DVSS.n17636 0.00108858
R40918 DVSS.n7137 DVSS.n7136 0.00108858
R40919 DVSS.n13556 DVSS.n13555 0.00108858
R40920 DVSS.n7196 DVSS.n7188 0.00108858
R40921 DVSS.n13524 DVSS.n13523 0.00108858
R40922 DVSS.n7091 DVSS.n7090 0.00108858
R40923 DVSS.n13592 DVSS.n13591 0.00108858
R40924 DVSS.n10642 DVSS.n10641 0.00108858
R40925 DVSS.n10750 DVSS.n10749 0.00108858
R40926 DVSS.n10742 DVSS.n10741 0.00108858
R40927 DVSS.n11431 DVSS.n11430 0.00108858
R40928 DVSS.n11434 DVSS.n11433 0.00108858
R40929 DVSS.n11571 DVSS.n11570 0.00108858
R40930 DVSS.n11595 DVSS.n11594 0.00108858
R40931 DVSS.n20 DVSS.n19 0.00108858
R40932 DVSS.n44 DVSS.n43 0.00108858
R40933 DVSS.n21525 DVSS.n21524 0.00108858
R40934 DVSS.n21501 DVSS.n21500 0.00108858
R40935 DVSS.n21437 DVSS.n21436 0.00108858
R40936 DVSS.n21413 DVSS.n21412 0.00108858
R40937 DVSS.n11570 DVSS.n11569 0.00108858
R40938 DVSS.n11594 DVSS.n11593 0.00108858
R40939 DVSS.n11435 DVSS.n11434 0.00108858
R40940 DVSS.n10751 DVSS.n10750 0.00108858
R40941 DVSS.n10641 DVSS.n10636 0.00108858
R40942 DVSS.n10804 DVSS.n10803 0.00108858
R40943 DVSS.n10743 DVSS.n10742 0.00108858
R40944 DVSS.n4697 DVSS.n4696 0.00108858
R40945 DVSS.n4687 DVSS.n4686 0.00108858
R40946 DVSS.n4676 DVSS.n4675 0.00108858
R40947 DVSS.n4677 DVSS.n4676 0.00108858
R40948 DVSS.n4698 DVSS.n4697 0.00108858
R40949 DVSS.n4688 DVSS.n4687 0.00108858
R40950 DVSS.n4302 DVSS.n4301 0.00108858
R40951 DVSS.n4323 DVSS.n4322 0.00108858
R40952 DVSS.n3485 DVSS.n3484 0.00108858
R40953 DVSS.n3464 DVSS.n3463 0.00108858
R40954 DVSS.n3317 DVSS.n3316 0.00108858
R40955 DVSS.n3066 DVSS.n3065 0.00108858
R40956 DVSS.n2791 DVSS.n2790 0.00108858
R40957 DVSS.n743 DVSS.n742 0.00108858
R40958 DVSS.n709 DVSS.n708 0.00108858
R40959 DVSS.n4301 DVSS.n4300 0.00108858
R40960 DVSS.n4322 DVSS.n4321 0.00108858
R40961 DVSS.n9967 DVSS.n9966 0.00108858
R40962 DVSS.n11156 DVSS.n11155 0.00108858
R40963 DVSS.n9836 DVSS.n9835 0.00108858
R40964 DVSS.n9661 DVSS.n9660 0.00108858
R40965 DVSS.n9637 DVSS.n9636 0.00108858
R40966 DVSS.n13240 DVSS.n13239 0.00108858
R40967 DVSS.n13359 DVSS.n13358 0.00108858
R40968 DVSS.n20468 DVSS.n20467 0.00108858
R40969 DVSS.n20560 DVSS.n20559 0.00108858
R40970 DVSS.n21054 DVSS.n21053 0.00108858
R40971 DVSS.n21018 DVSS.n21017 0.00108858
R40972 DVSS.n20994 DVSS.n20993 0.00108858
R40973 DVSS.n13400 DVSS.n13392 0.00108858
R40974 DVSS.n9811 DVSS.n9810 0.00108858
R40975 DVSS.n9662 DVSS.n9661 0.00108858
R40976 DVSS.n9638 DVSS.n9637 0.00108858
R40977 DVSS.n11155 DVSS.n11154 0.00108858
R40978 DVSS.n11147 DVSS.n11146 0.00108858
R40979 DVSS.n9986 DVSS.n9985 0.00108858
R40980 DVSS.n9966 DVSS.n9965 0.00108858
R40981 DVSS.n9879 DVSS.n9878 0.00108858
R40982 DVSS.n9976 DVSS.n9975 0.00108858
R40983 DVSS.n11138 DVSS.n11137 0.00108858
R40984 DVSS.n11160 DVSS.n11159 0.00108858
R40985 DVSS.n13358 DVSS.n13357 0.00108858
R40986 DVSS.n17371 DVSS.n17370 0.00108858
R40987 DVSS.n17392 DVSS.n17391 0.00108858
R40988 DVSS.n16368 DVSS.n16367 0.00108858
R40989 DVSS.n16359 DVSS.n16358 0.00108858
R40990 DVSS.n16350 DVSS.n16349 0.00108858
R40991 DVSS.n16346 DVSS.n16345 0.00108858
R40992 DVSS.n16327 DVSS.n16326 0.00108858
R40993 DVSS.n16300 DVSS.n16299 0.00108858
R40994 DVSS.n16178 DVSS.n16177 0.00108858
R40995 DVSS.n16156 DVSS.n16155 0.00108858
R40996 DVSS.n18627 DVSS.n18626 0.00108858
R40997 DVSS.n18654 DVSS.n18653 0.00108858
R40998 DVSS.n18686 DVSS.n18685 0.00108858
R40999 DVSS.n18820 DVSS.n18819 0.00108858
R41000 DVSS.n19457 DVSS.n19456 0.00108858
R41001 DVSS.n19543 DVSS.n19542 0.00108858
R41002 DVSS.n1132 DVSS.n1131 0.00108858
R41003 DVSS.n1242 DVSS.n1241 0.00108858
R41004 DVSS.n1221 DVSS.n1220 0.00108858
R41005 DVSS.n16301 DVSS.n16300 0.00108858
R41006 DVSS.n16179 DVSS.n16178 0.00108858
R41007 DVSS.n18856 DVSS.n18850 0.00108858
R41008 DVSS.n18770 DVSS.n18769 0.00108858
R41009 DVSS.n16157 DVSS.n16156 0.00108858
R41010 DVSS.n18626 DVSS.n18625 0.00108858
R41011 DVSS.n18653 DVSS.n18652 0.00108858
R41012 DVSS.n18685 DVSS.n18684 0.00108858
R41013 DVSS.n17391 DVSS.n17390 0.00108858
R41014 DVSS.n17370 DVSS.n17369 0.00108858
R41015 DVSS.n16369 DVSS.n16368 0.00108858
R41016 DVSS.n16360 DVSS.n16359 0.00108858
R41017 DVSS.n16351 DVSS.n16350 0.00108858
R41018 DVSS.n16347 DVSS.n16346 0.00108858
R41019 DVSS.n16328 DVSS.n16327 0.00108858
R41020 DVSS.n18819 DVSS.n18818 0.00108858
R41021 DVSS.n5405 DVSS.n5404 0.00108858
R41022 DVSS.n5460 DVSS.n5459 0.00108858
R41023 DVSS.n5844 DVSS.n5843 0.00108858
R41024 DVSS.n5851 DVSS.n5850 0.00108858
R41025 DVSS.n6469 DVSS.n6468 0.00108858
R41026 DVSS.n6464 DVSS.n6463 0.00108858
R41027 DVSS.n6616 DVSS.n6615 0.00108858
R41028 DVSS.n6638 DVSS.n6637 0.00108858
R41029 DVSS.n3547 DVSS.n3546 0.00108858
R41030 DVSS.n18945 DVSS.n18944 0.00108858
R41031 DVSS.n18991 DVSS.n18990 0.00108858
R41032 DVSS.n523 DVSS.n522 0.00108858
R41033 DVSS.n593 DVSS.n592 0.00108858
R41034 DVSS.n572 DVSS.n571 0.00108858
R41035 DVSS.n5459 DVSS.n5458 0.00108858
R41036 DVSS.n5843 DVSS.n5842 0.00108858
R41037 DVSS.n6615 DVSS.n6614 0.00108858
R41038 DVSS.n6637 DVSS.n6636 0.00108858
R41039 DVSS.n5404 DVSS.n5395 0.00108858
R41040 DVSS.n6468 DVSS.n6467 0.00108858
R41041 DVSS.n6465 DVSS.n6464 0.00108858
R41042 DVSS.n3548 DVSS.n3547 0.00108858
R41043 DVSS.n43 DVSS.n42 0.00108858
R41044 DVSS.n12853 DVSS.n12852 0.00108858
R41045 DVSS.n20467 DVSS.n20466 0.00108858
R41046 DVSS.n20196 DVSS.n20195 0.00108858
R41047 DVSS.n19456 DVSS.n19455 0.00108858
R41048 DVSS.n19185 DVSS.n19184 0.00108858
R41049 DVSS.n3465 DVSS.n3464 0.00108858
R41050 DVSS.n18944 DVSS.n18943 0.00108858
R41051 DVSS.n19 DVSS.n18 0.00108858
R41052 DVSS.n3486 DVSS.n3485 0.00108858
R41053 DVSS.n18992 DVSS.n18991 0.00108858
R41054 DVSS.n3116 DVSS.n3115 0.00108858
R41055 DVSS.n19544 DVSS.n19543 0.00108858
R41056 DVSS.n12492 DVSS.n12491 0.00108858
R41057 DVSS.n21526 DVSS.n21525 0.00108858
R41058 DVSS.n19273 DVSS.n19272 0.00108858
R41059 DVSS.n12695 DVSS.n12694 0.00108858
R41060 DVSS.n3318 DVSS.n3317 0.00108858
R41061 DVSS.n21502 DVSS.n21501 0.00108858
R41062 DVSS.n12440 DVSS.n12439 0.00108858
R41063 DVSS.n21053 DVSS.n21052 0.00108858
R41064 DVSS.n20827 DVSS.n20826 0.00108858
R41065 DVSS.n1131 DVSS.n1130 0.00108858
R41066 DVSS.n844 DVSS.n843 0.00108858
R41067 DVSS.n3067 DVSS.n3066 0.00108858
R41068 DVSS.n522 DVSS.n521 0.00108858
R41069 DVSS.n20561 DVSS.n20560 0.00108858
R41070 DVSS.n20287 DVSS.n20286 0.00108858
R41071 DVSS.n594 DVSS.n593 0.00108858
R41072 DVSS.n744 DVSS.n743 0.00108858
R41073 DVSS.n988 DVSS.n987 0.00108858
R41074 DVSS.n1243 DVSS.n1242 0.00108858
R41075 DVSS.n21438 DVSS.n21437 0.00108858
R41076 DVSS.n1028 DVSS.n1027 0.00108858
R41077 DVSS.n2790 DVSS.n2789 0.00108858
R41078 DVSS.n12162 DVSS.n12161 0.00108858
R41079 DVSS.n21414 DVSS.n21413 0.00108858
R41080 DVSS.n20995 DVSS.n20994 0.00108858
R41081 DVSS.n21019 DVSS.n21018 0.00108858
R41082 DVSS.n20769 DVSS.n20768 0.00108858
R41083 DVSS.n20793 DVSS.n20792 0.00108858
R41084 DVSS.n1222 DVSS.n1221 0.00108858
R41085 DVSS.n1007 DVSS.n1006 0.00108858
R41086 DVSS.n573 DVSS.n572 0.00108858
R41087 DVSS.n12115 DVSS 0.00108667
R41088 DVSS.n2336 DVSS.n2043 0.00107857
R41089 DVSS.n2414 DVSS.n2413 0.00107857
R41090 DVSS.n12531 DVSS.n12530 0.00107692
R41091 DVSS.n12655 DVSS.n12654 0.00107692
R41092 DVSS.n12367 DVSS.n12366 0.00107692
R41093 DVSS.n12275 DVSS.n12274 0.00107692
R41094 DVSS.n12266 DVSS.n12261 0.00107692
R41095 DVSS.n3155 DVSS.n3154 0.00107692
R41096 DVSS.n3279 DVSS.n3278 0.00107692
R41097 DVSS.n2994 DVSS.n2993 0.00107692
R41098 DVSS.n2902 DVSS.n2901 0.00107692
R41099 DVSS.n2893 DVSS.n2888 0.00107692
R41100 DVSS.n14526 DVSS.n14525 0.001075
R41101 DVSS.n14527 DVSS.n14526 0.001075
R41102 DVSS.n19825 DVSS.n19824 0.001075
R41103 DVSS.n19824 DVSS.n19823 0.001075
R41104 DVSS.n260 DVSS.n259 0.001075
R41105 DVSS.n261 DVSS.n260 0.001075
R41106 DVSS.n14524 DVSS.n14523 0.00107
R41107 DVSS.n14532 DVSS.n14530 0.00107
R41108 DVSS.n14585 DVSS.n14584 0.00107
R41109 DVSS.n19829 DVSS.n19827 0.00107
R41110 DVSS.n265 DVSS.n263 0.00107
R41111 DVSS.n4571 DVSS.n4570 0.00106944
R41112 DVSS.n6758 DVSS.n6757 0.00106944
R41113 DVSS.n6703 DVSS.n6702 0.00106944
R41114 DVSS.n2535 DVSS.n2534 0.00106944
R41115 DVSS.n4518 DVSS.n4517 0.00106944
R41116 DVSS.n6396 DVSS.n6395 0.00106944
R41117 DVSS.n6885 DVSS.n6884 0.00106944
R41118 DVSS.n4622 DVSS.n4621 0.00106944
R41119 DVSS.n4621 DVSS.n4620 0.00106944
R41120 DVSS.n4517 DVSS.n4516 0.00106944
R41121 DVSS.n6395 DVSS.n6394 0.00106944
R41122 DVSS.n2534 DVSS.n2533 0.00106944
R41123 DVSS.n6702 DVSS.n6701 0.00106944
R41124 DVSS.n6757 DVSS.n6756 0.00106944
R41125 DVSS.n6884 DVSS.n6883 0.00106944
R41126 DVSS.n4572 DVSS.n4571 0.00106944
R41127 DVSS.n10080 DVSS.n10079 0.00106429
R41128 DVSS.n10079 DVSS.n10078 0.00106429
R41129 DVSS.n5262 DVSS.n5261 0.00106338
R41130 DVSS.n10595 DVSS.n10594 0.00106338
R41131 DVSS.n21367 DVSS 0.00104667
R41132 DVSS.n9272 DVSS.n9271 0.00104
R41133 DVSS.n9325 DVSS.n9324 0.00104
R41134 DVSS.n9454 DVSS.n9453 0.00104
R41135 DVSS.n9439 DVSS.n9438 0.00104
R41136 DVSS.n9194 DVSS.n9191 0.00104
R41137 DVSS.n9274 DVSS.n9273 0.00104
R41138 DVSS.n9327 DVSS.n9326 0.00104
R41139 DVSS.n9456 DVSS.n9455 0.00104
R41140 DVSS.n9440 DVSS.n9435 0.00104
R41141 DVSS.n12131 DVSS.n12130 0.00104
R41142 DVSS.n12023 DVSS.n12022 0.00104
R41143 DVSS.n20634 DVSS.n20633 0.00104
R41144 DVSS.n11 DVSS.n10 0.00104
R41145 DVSS.n21347 DVSS.n21346 0.00104
R41146 DVSS.n21380 DVSS.n21376 0.00104
R41147 DVSS.n20874 DVSS.n20873 0.00104
R41148 DVSS.n21100 DVSS.n21099 0.00104
R41149 DVSS.n21349 DVSS.n21348 0.00104
R41150 DVSS.n21379 DVSS.n21378 0.00104
R41151 DVSS.n20328 DVSS.n20114 0.00104
R41152 DVSS.n20613 DVSS.n20600 0.00104
R41153 DVSS.n20635 DVSS.n20627 0.00104
R41154 DVSS.n12 DVSS.n5 0.00104
R41155 DVSS.n13483 DVSS.n13467 0.00104
R41156 DVSS.n7929 DVSS.n7915 0.00104
R41157 DVSS.n12121 DVSS.n12120 0.00104
R41158 DVSS.n12025 DVSS.n12024 0.00104
R41159 DVSS.n18919 DVSS.n18918 0.00103333
R41160 DVSS.n19594 DVSS.n19593 0.00103333
R41161 DVSS.n1302 DVSS.n1301 0.00103333
R41162 DVSS.n10058 DVSS.n10057 0.00103214
R41163 DVSS.n10122 DVSS.n10121 0.00103214
R41164 DVSS.n10170 DVSS.n10169 0.00103214
R41165 DVSS.n10171 DVSS.n10170 0.00103214
R41166 DVSS.n10057 DVSS.n10056 0.00103214
R41167 DVSS.n10123 DVSS.n10122 0.00103214
R41168 DVSS.n5560 DVSS.n5559 0.0010315
R41169 DVSS.n5776 DVSS.n5775 0.0010315
R41170 DVSS.n5750 DVSS.n5749 0.0010315
R41171 DVSS.n4050 DVSS.n4049 0.0010315
R41172 DVSS.n7107 DVSS.n7106 0.0010315
R41173 DVSS.n7149 DVSS.n7148 0.0010315
R41174 DVSS.n7176 DVSS.n7175 0.0010315
R41175 DVSS.n7199 DVSS.n7198 0.0010315
R41176 DVSS.n10201 DVSS.n10200 0.0010315
R41177 DVSS.n11281 DVSS.n11280 0.0010315
R41178 DVSS.n13133 DVSS.n13132 0.0010315
R41179 DVSS.n12925 DVSS.n12924 0.0010315
R41180 DVSS.n12697 DVSS.n12696 0.0010315
R41181 DVSS.n12478 DVSS.n12477 0.0010315
R41182 DVSS.n12211 DVSS.n12210 0.0010315
R41183 DVSS.n12197 DVSS.n12196 0.0010315
R41184 DVSS.n21277 DVSS.n21276 0.0010315
R41185 DVSS.n21283 DVSS.n21282 0.0010315
R41186 DVSS.n16946 DVSS.n16945 0.0010315
R41187 DVSS.n17584 DVSS.n17583 0.0010315
R41188 DVSS.n15028 DVSS.n15027 0.0010315
R41189 DVSS.n13574 DVSS.n13573 0.0010315
R41190 DVSS.n13544 DVSS.n13543 0.0010315
R41191 DVSS.n13531 DVSS.n13530 0.0010315
R41192 DVSS.n13521 DVSS.n13520 0.0010315
R41193 DVSS.n10605 DVSS.n10604 0.0010315
R41194 DVSS.n10781 DVSS.n10780 0.0010315
R41195 DVSS.n11381 DVSS.n11380 0.0010315
R41196 DVSS.n11408 DVSS.n11407 0.0010315
R41197 DVSS.n11444 DVSS.n11443 0.0010315
R41198 DVSS.n13068 DVSS.n13067 0.0010315
R41199 DVSS.n12047 DVSS.n12046 0.0010315
R41200 DVSS.n5213 DVSS.n5212 0.0010315
R41201 DVSS.n3985 DVSS.n3984 0.0010315
R41202 DVSS.n3749 DVSS.n3748 0.0010315
R41203 DVSS.n3320 DVSS.n3319 0.0010315
R41204 DVSS.n3104 DVSS.n3103 0.0010315
R41205 DVSS.n2841 DVSS.n2840 0.0010315
R41206 DVSS.n2826 DVSS.n2825 0.0010315
R41207 DVSS.n654 DVSS.n653 0.0010315
R41208 DVSS.n660 DVSS.n659 0.0010315
R41209 DVSS.n9902 DVSS.n9901 0.0010315
R41210 DVSS.n11107 DVSS.n11106 0.0010315
R41211 DVSS.n9057 DVSS.n9056 0.0010315
R41212 DVSS.n13258 DVSS.n13257 0.0010315
R41213 DVSS.n13370 DVSS.n13369 0.0010315
R41214 DVSS.n13386 DVSS.n13385 0.0010315
R41215 DVSS.n13403 DVSS.n13402 0.0010315
R41216 DVSS.n17255 DVSS.n17254 0.0010315
R41217 DVSS.n16397 DVSS.n16396 0.0010315
R41218 DVSS.n16371 DVSS.n16370 0.0010315
R41219 DVSS.n7515 DVSS.n7514 0.0010315
R41220 DVSS.n18786 DVSS.n18785 0.0010315
R41221 DVSS.n18831 DVSS.n18830 0.0010315
R41222 DVSS.n18844 DVSS.n18843 0.0010315
R41223 DVSS.n18859 DVSS.n18858 0.0010315
R41224 DVSS.n5318 DVSS.n5317 0.0010315
R41225 DVSS.n5483 DVSS.n5482 0.0010315
R41226 DVSS.n6066 DVSS.n6065 0.0010315
R41227 DVSS.n6331 DVSS.n6330 0.0010315
R41228 DVSS.n6455 DVSS.n6454 0.0010315
R41229 DVSS.n6833 DVSS.n6832 0.0010315
R41230 DVSS.n3642 DVSS.n3641 0.0010315
R41231 DVSS.n13471 DVSS.n13470 0.00103
R41232 DVSS.n7917 DVSS.n7916 0.00103
R41233 DVSS.n12136 DVSS.n12135 0.00103
R41234 DVSS.n12135 DVSS.n12134 0.00103
R41235 DVSS.n13470 DVSS.n13469 0.00103
R41236 DVSS.n2057 VSS 0.00101429
R41237 DVSS.n4989 DVSS.n4988 0.00101429
R41238 DVSS.n4754 DVSS.n4753 0.00101429
R41239 DVSS.n10084 DVSS.n10083 0.00101429
R41240 DVSS.n10151 DVSS.n10150 0.00101429
R41241 DVSS.n10702 DVSS.n10701 0.00101429
R41242 DVSS.n10721 DVSS.n10720 0.00101429
R41243 DVSS.n6039 DVSS.n6038 0.00101429
R41244 DVSS.n11302 DVSS.n11301 0.00101429
R41245 DVSS.n6287 DVSS.n6286 0.00101429
R41246 DVSS.n8656 DVSS.n8655 0.00101429
R41247 DVSS.n8720 DVSS.n8719 0.00101429
R41248 DVSS.n8781 DVSS.n8780 0.00101429
R41249 DVSS.n8876 DVSS.n8875 0.00101429
R41250 DVSS.n8894 DVSS.n8893 0.00101429
R41251 DVSS.n9275 DVSS.n9274 0.00101
R41252 DVSS.n9328 DVSS.n9327 0.00101
R41253 DVSS.n9457 DVSS.n9456 0.00101
R41254 DVSS.n9435 DVSS.n9434 0.00101
R41255 DVSS.n14125 DVSS.n14124 0.00101
R41256 DVSS.n12130 DVSS.n12129 0.00101
R41257 DVSS.n12022 DVSS.n12021 0.00101
R41258 DVSS.n19629 DVSS.n19628 0.00101
R41259 DVSS.n20325 DVSS.n20324 0.00101
R41260 DVSS.n20610 DVSS.n20609 0.00101
R41261 DVSS.n20633 DVSS.n20632 0.00101
R41262 DVSS.n10 DVSS.n9 0.00101
R41263 DVSS.n116 DVSS.n115 0.00101
R41264 DVSS.n20870 DVSS.n20869 0.00101
R41265 DVSS.n21096 DVSS.n21095 0.00101
R41266 DVSS.n21346 DVSS.n21345 0.00101
R41267 DVSS.n21376 DVSS.n21375 0.00101
R41268 DVSS.n10362 DVSS.n10361 0.000992958
R41269 DVSS.n10366 DVSS.n10365 0.000992958
R41270 DVSS.n9211 DVSS.n9210 0.00098
R41271 DVSS.n1382 DVSS.n1381 0.00098
R41272 DVSS.n4140 DVSS.n4139 0.00098
R41273 DVSS.n4221 DVSS.n4220 0.00098
R41274 DVSS.n4175 DVSS.n4174 0.00098
R41275 DVSS.n9213 DVSS.n9212 0.00098
R41276 DVSS.n9214 DVSS.n9213 0.00098
R41277 DVSS.n3523 DVSS.n3522 0.00098
R41278 DVSS.n3691 DVSS.n3690 0.00098
R41279 DVSS.n7244 DVSS.n7243 0.00098
R41280 DVSS.n18903 DVSS.n18902 0.00098
R41281 DVSS.n18925 DVSS.n18924 0.00098
R41282 DVSS.n19045 DVSS.n19044 0.00098
R41283 DVSS.n19096 DVSS.n19095 0.00098
R41284 DVSS.n19362 DVSS.n19361 0.00098
R41285 DVSS.n20322 DVSS.n20321 0.00098
R41286 DVSS.n20607 DVSS.n20606 0.00098
R41287 DVSS.n510 DVSS.n509 0.00098
R41288 DVSS.n680 DVSS.n679 0.00098
R41289 DVSS.n833 DVSS.n832 0.00098
R41290 DVSS.n1120 DVSS.n1119 0.00098
R41291 DVSS.n20867 DVSS.n20866 0.00098
R41292 DVSS.n21093 DVSS.n21092 0.00098
R41293 DVSS.n285 DVSS.n277 0.00098
R41294 DVSS.n19849 DVSS.n19848 0.00098
R41295 DVSS.n14591 DVSS.n14590 0.00098
R41296 DVSS DVSS.n11334 0.000957143
R41297 DVSS.n7722 DVSS.n7721 0.00095
R41298 DVSS.n16053 DVSS.n16052 0.00095
R41299 DVSS.n4751 DVSS.n4750 0.00095
R41300 DVSS.n4752 DVSS.n4748 0.00095
R41301 DVSS.n1385 DVSS.n1383 0.00095
R41302 DVSS.n4143 DVSS.n4141 0.00095
R41303 DVSS.n4218 DVSS.n4216 0.00095
R41304 DVSS.n4172 DVSS.n4170 0.00095
R41305 DVSS.n1386 DVSS.n1382 0.00095
R41306 DVSS.n4144 DVSS.n4140 0.00095
R41307 DVSS.n4220 DVSS.n4219 0.00095
R41308 DVSS.n4174 DVSS.n4173 0.00095
R41309 DVSS.n8114 DVSS.n8113 0.00095
R41310 DVSS.n8116 DVSS.n8115 0.00095
R41311 DVSS.n8117 DVSS.n8116 0.00095
R41312 DVSS.n11791 DVSS.n11790 0.00095
R41313 DVSS.n11795 DVSS.n11794 0.00095
R41314 DVSS.n8406 DVSS.n8405 0.00095
R41315 DVSS.n8408 DVSS.n8407 0.00095
R41316 DVSS.n8409 DVSS.n8408 0.00095
R41317 DVSS.n8661 DVSS.n8660 0.00095
R41318 DVSS.n8662 DVSS.n8661 0.00095
R41319 DVSS.n8659 DVSS.n8658 0.00095
R41320 DVSS.n3525 DVSS.n3523 0.00095
R41321 DVSS.n3693 DVSS.n3691 0.00095
R41322 DVSS.n3729 DVSS.n3728 0.00095
R41323 DVSS.n7242 DVSS.n7241 0.00095
R41324 DVSS.n18901 DVSS.n18900 0.00095
R41325 DVSS.n14569 DVSS.n14568 0.00095
R41326 DVSS.n7893 DVSS.n7892 0.00095
R41327 DVSS.n13502 DVSS.n13501 0.00095
R41328 DVSS.n7950 DVSS.n7949 0.00095
R41329 DVSS.n13422 DVSS.n13421 0.00095
R41330 DVSS.n12136 DVSS.n12127 0.00095
R41331 DVSS.n18927 DVSS.n18925 0.00095
R41332 DVSS.n19047 DVSS.n19045 0.00095
R41333 DVSS.n19054 DVSS.n19053 0.00095
R41334 DVSS.n19094 DVSS.n19093 0.00095
R41335 DVSS.n19360 DVSS.n19359 0.00095
R41336 DVSS.n20039 DVSS.n20038 0.00095
R41337 DVSS.n20644 DVSS.n20643 0.00095
R41338 DVSS.n512 DVSS.n510 0.00095
R41339 DVSS.n682 DVSS.n680 0.00095
R41340 DVSS.n719 DVSS.n718 0.00095
R41341 DVSS.n831 DVSS.n830 0.00095
R41342 DVSS.n1118 DVSS.n1117 0.00095
R41343 DVSS.n463 DVSS.n462 0.00095
R41344 DVSS.n21270 DVSS.n21269 0.00095
R41345 DVSS.n513 DVSS.n506 0.00095
R41346 DVSS.n683 DVSS.n649 0.00095
R41347 DVSS.n827 DVSS.n825 0.00095
R41348 DVSS.n1114 DVSS.n1112 0.00095
R41349 DVSS.n18928 DVSS.n18921 0.00095
R41350 DVSS.n19048 DVSS.n19040 0.00095
R41351 DVSS.n19090 DVSS.n19088 0.00095
R41352 DVSS.n19356 DVSS.n19354 0.00095
R41353 DVSS.n3527 DVSS.n3519 0.00095
R41354 DVSS.n3695 DVSS.n3687 0.00095
R41355 DVSS.n1305 DVSS.n1303 0.00095
R41356 DVSS.n7287 DVSS.n7285 0.00095
R41357 DVSS.n14540 DVSS.n81 0.000926667
R41358 DVSS.n20079 DVSS.n20078 0.000926667
R41359 DVSS.n504 DVSS.n503 0.000926667
R41360 DVSS.n10364 DVSS.n10363 0.000922535
R41361 DVSS.n16643 DVSS.n16642 0.000922535
R41362 DVSS.n16653 DVSS.n16652 0.000922535
R41363 DVSS.n16659 DVSS.n16658 0.000922535
R41364 DVSS.n16663 DVSS.n16662 0.000922535
R41365 DVSS.n17467 DVSS.n17466 0.000922535
R41366 DVSS.n16105 DVSS.n16104 0.000922535
R41367 DVSS.n16062 DVSS.n16061 0.000922535
R41368 DVSS.n17731 DVSS.n17730 0.000922535
R41369 DVSS.n17732 DVSS.n17731 0.000922535
R41370 DVSS.n17742 DVSS.n17741 0.000922535
R41371 DVSS.n17796 DVSS.n17795 0.000922535
R41372 DVSS.n18139 DVSS.n18138 0.000922535
R41373 DVSS.n18251 DVSS.n18250 0.000922535
R41374 DVSS.n18435 DVSS.n18434 0.000922535
R41375 DVSS.n18473 DVSS.n18472 0.000922535
R41376 DVSS.n18478 DVSS.n18477 0.000922535
R41377 DVSS.n14375 DVSS.n14374 0.000922535
R41378 DVSS.n14396 DVSS.n14395 0.000922535
R41379 DVSS.n19725 DVSS.n19724 0.000922535
R41380 DVSS.n179 DVSS.n178 0.000922535
R41381 DVSS.n17180 DVSS.n17179 0.000922535
R41382 DVSS.n17170 DVSS.n17169 0.000922535
R41383 DVSS.n17164 DVSS.n17163 0.000922535
R41384 DVSS.n17160 DVSS.n17159 0.000922535
R41385 DVSS.n16808 DVSS.n16807 0.000922535
R41386 DVSS.n15986 DVSS.n15985 0.000922535
R41387 DVSS.n15954 DVSS.n15953 0.000922535
R41388 DVSS.n15932 DVSS.n15931 0.000922535
R41389 DVSS.n15931 DVSS.n15930 0.000922535
R41390 DVSS.n15921 DVSS.n15920 0.000922535
R41391 DVSS.n17670 DVSS.n17669 0.000922535
R41392 DVSS.n15444 DVSS.n15443 0.000922535
R41393 DVSS.n15489 DVSS.n15488 0.000922535
R41394 DVSS.n15194 DVSS.n15193 0.000922535
R41395 DVSS.n15129 DVSS.n15128 0.000922535
R41396 DVSS.n15124 DVSS.n15123 0.000922535
R41397 DVSS.n14775 DVSS.n14774 0.000922535
R41398 DVSS.n14754 DVSS.n14753 0.000922535
R41399 DVSS.n19944 DVSS.n19943 0.000922535
R41400 DVSS.n387 DVSS.n386 0.000922535
R41401 DVSS.n9183 DVSS.n9181 0.00092
R41402 DVSS.n9183 DVSS.n9182 0.00092
R41403 DVSS.n9180 DVSS.n9179 0.00092
R41404 DVSS.n9184 DVSS.n9180 0.00092
R41405 DVSS.n9185 DVSS.n9184 0.00092
R41406 DVSS.n14129 DVSS.n14128 0.00092
R41407 DVSS.n14130 DVSS.n14129 0.00092
R41408 DVSS.n19812 DVSS.n19635 0.00092
R41409 DVSS.n19813 DVSS.n19812 0.00092
R41410 DVSS.n253 DVSS.n127 0.00092
R41411 DVSS.n254 DVSS.n253 0.00092
R41412 DVSS.n257 DVSS.n256 0.00092
R41413 DVSS.n121 DVSS.n119 0.00092
R41414 DVSS.n121 DVSS.n120 0.00092
R41415 DVSS.n19817 DVSS.n19632 0.00092
R41416 DVSS.n19817 DVSS.n19816 0.00092
R41417 DVSS.n14133 DVSS.n14116 0.00092
R41418 DVSS.n14133 DVSS.n14117 0.00092
R41419 DVSS.n1385 DVSS.n1384 0.00089
R41420 DVSS.n4143 DVSS.n4142 0.00089
R41421 DVSS.n4218 DVSS.n4217 0.00089
R41422 DVSS.n4172 DVSS.n4171 0.00089
R41423 DVSS.n1387 DVSS.n1386 0.00089
R41424 DVSS.n4145 DVSS.n4144 0.00089
R41425 DVSS.n4219 DVSS.n4215 0.00089
R41426 DVSS.n4173 DVSS.n4169 0.00089
R41427 DVSS.n3525 DVSS.n3524 0.00089
R41428 DVSS.n3693 DVSS.n3692 0.00089
R41429 DVSS.n7220 DVSS.n7219 0.00089
R41430 DVSS.n18880 DVSS.n18879 0.00089
R41431 DVSS.n14128 DVSS.n14127 0.00089
R41432 DVSS.n14131 DVSS.n14130 0.00089
R41433 DVSS.n14579 DVSS.n14571 0.00089
R41434 DVSS.n18927 DVSS.n18926 0.00089
R41435 DVSS.n19047 DVSS.n19046 0.00089
R41436 DVSS.n19099 DVSS.n19098 0.00089
R41437 DVSS.n19365 DVSS.n19364 0.00089
R41438 DVSS.n19635 DVSS.n19634 0.00089
R41439 DVSS.n19814 DVSS.n19813 0.00089
R41440 DVSS.n20047 DVSS.n20041 0.00089
R41441 DVSS.n512 DVSS.n511 0.00089
R41442 DVSS.n682 DVSS.n681 0.00089
R41443 DVSS.n836 DVSS.n835 0.00089
R41444 DVSS.n1123 DVSS.n1122 0.00089
R41445 DVSS.n127 DVSS.n126 0.00089
R41446 DVSS.n255 DVSS.n254 0.00089
R41447 DVSS.n471 DVSS.n465 0.00089
R41448 DVSS.n513 DVSS.n507 0.00089
R41449 DVSS.n683 DVSS.n650 0.00089
R41450 DVSS.n827 DVSS.n826 0.00089
R41451 DVSS.n1114 DVSS.n1113 0.00089
R41452 DVSS.n18928 DVSS.n18922 0.00089
R41453 DVSS.n19048 DVSS.n19041 0.00089
R41454 DVSS.n19090 DVSS.n19089 0.00089
R41455 DVSS.n19356 DVSS.n19355 0.00089
R41456 DVSS.n3527 DVSS.n3526 0.00089
R41457 DVSS.n3695 DVSS.n3694 0.00089
R41458 DVSS.n1305 DVSS.n1304 0.00089
R41459 DVSS.n7287 DVSS.n7286 0.00089
R41460 DVSS.n4803 DVSS.n4802 0.000885714
R41461 DVSS.n4745 DVSS.n4744 0.000885714
R41462 DVSS.n11793 DVSS.n11792 0.000885714
R41463 DVSS.n8609 DVSS.n8608 0.000885714
R41464 DVSS.n8664 DVSS.n8663 0.000885714
R41465 DVSS.n9211 DVSS.n9209 0.00086
R41466 DVSS.n1381 DVSS.n1380 0.00086
R41467 DVSS.n4139 DVSS.n4138 0.00086
R41468 DVSS.n4176 DVSS.n4175 0.00086
R41469 DVSS.n9212 DVSS.n9208 0.00086
R41470 DVSS.n7215 DVSS.n1310 0.00086
R41471 DVSS.n7216 DVSS.n7215 0.00086
R41472 DVSS.n7243 DVSS.n7242 0.00086
R41473 DVSS.n18875 DVSS.n7293 0.00086
R41474 DVSS.n18876 DVSS.n18875 0.00086
R41475 DVSS.n18902 DVSS.n18901 0.00086
R41476 DVSS.n14589 DVSS.n14586 0.00086
R41477 DVSS.n14568 DVSS.n14567 0.00086
R41478 DVSS.n13503 DVSS.n13502 0.00086
R41479 DVSS.n13479 DVSS.n13478 0.00086
R41480 DVSS.n13421 DVSS.n13420 0.00086
R41481 DVSS.n7925 DVSS.n7924 0.00086
R41482 DVSS.n18924 DVSS.n18923 0.00086
R41483 DVSS.n19095 DVSS.n19094 0.00086
R41484 DVSS.n19361 DVSS.n19360 0.00086
R41485 DVSS.n19847 DVSS.n19844 0.00086
R41486 DVSS.n20038 DVSS.n20037 0.00086
R41487 DVSS.n509 DVSS.n508 0.00086
R41488 DVSS.n832 DVSS.n831 0.00086
R41489 DVSS.n1119 DVSS.n1118 0.00086
R41490 DVSS.n284 DVSS.n281 0.00086
R41491 DVSS.n462 DVSS.n461 0.00086
R41492 DVSS.n285 DVSS.n276 0.00086
R41493 DVSS.n19849 DVSS.n19840 0.00086
R41494 DVSS.n14591 DVSS.n14582 0.00086
R41495 DVSS.n5634 DVSS.n5633 0.000854331
R41496 DVSS.n5711 DVSS.n5710 0.000854331
R41497 DVSS.n5765 DVSS.n5764 0.000854331
R41498 DVSS.n5714 DVSS.n5713 0.000854331
R41499 DVSS.n4076 DVSS.n4075 0.000854331
R41500 DVSS.n6976 DVSS.n6975 0.000854331
R41501 DVSS.n6996 DVSS.n6995 0.000854331
R41502 DVSS.n19210 DVSS.n19209 0.000854331
R41503 DVSS.n10925 DVSS.n10924 0.000854331
R41504 DVSS.n11001 DVSS.n11000 0.000854331
R41505 DVSS.n11268 DVSS.n11267 0.000854331
R41506 DVSS.n11218 DVSS.n11217 0.000854331
R41507 DVSS.n8995 DVSS.n8994 0.000854331
R41508 DVSS.n12956 DVSS.n12955 0.000854331
R41509 DVSS.n12485 DVSS.n12484 0.000854331
R41510 DVSS.n12410 DVSS.n12409 0.000854331
R41511 DVSS.n12406 DVSS.n12405 0.000854331
R41512 DVSS.n21282 DVSS.n21281 0.000854331
R41513 DVSS.n21251 DVSS.n21250 0.000854331
R41514 DVSS.n21343 DVSS.n21342 0.000854331
R41515 DVSS.n17058 DVSS.n17057 0.000854331
R41516 DVSS.n16906 DVSS.n16905 0.000854331
R41517 DVSS.n17597 DVSS.n17596 0.000854331
R41518 DVSS.n17651 DVSS.n17650 0.000854331
R41519 DVSS.n15000 DVSS.n14999 0.000854331
R41520 DVSS.n13662 DVSS.n13661 0.000854331
R41521 DVSS.n13642 DVSS.n13641 0.000854331
R41522 DVSS.n20220 DVSS.n20219 0.000854331
R41523 DVSS.n10837 DVSS.n10836 0.000854331
R41524 DVSS.n10813 DVSS.n10812 0.000854331
R41525 DVSS.n10761 DVSS.n10760 0.000854331
R41526 DVSS.n11394 DVSS.n11393 0.000854331
R41527 DVSS.n11697 DVSS.n11696 0.000854331
R41528 DVSS.n13036 DVSS.n13035 0.000854331
R41529 DVSS.n4704 DVSS.n4703 0.000854331
R41530 DVSS.n3797 DVSS.n3796 0.000854331
R41531 DVSS.n3775 DVSS.n3774 0.000854331
R41532 DVSS.n3110 DVSS.n3109 0.000854331
R41533 DVSS.n3037 DVSS.n3036 0.000854331
R41534 DVSS.n3032 DVSS.n3031 0.000854331
R41535 DVSS.n659 DVSS.n658 0.000854331
R41536 DVSS.n734 DVSS.n733 0.000854331
R41537 DVSS.n730 DVSS.n729 0.000854331
R41538 DVSS.n9947 DVSS.n9946 0.000854331
R41539 DVSS.n9862 DVSS.n9861 0.000854331
R41540 DVSS.n11120 DVSS.n11119 0.000854331
R41541 DVSS.n9835 DVSS.n9834 0.000854331
R41542 DVSS.n9085 DVSS.n9084 0.000854331
R41543 DVSS.n13213 DVSS.n13212 0.000854331
R41544 DVSS.n13233 DVSS.n13232 0.000854331
R41545 DVSS.n20491 DVSS.n20490 0.000854331
R41546 DVSS.n17353 DVSS.n17352 0.000854331
R41547 DVSS.n17430 DVSS.n17429 0.000854331
R41548 DVSS.n16386 DVSS.n16385 0.000854331
R41549 DVSS.n16326 DVSS.n16325 0.000854331
R41550 DVSS.n7541 DVSS.n7540 0.000854331
R41551 DVSS.n18743 DVSS.n18742 0.000854331
R41552 DVSS.n18763 DVSS.n18762 0.000854331
R41553 DVSS.n19481 DVSS.n19480 0.000854331
R41554 DVSS.n5429 DVSS.n5428 0.000854331
R41555 DVSS.n5450 DVSS.n5449 0.000854331
R41556 DVSS.n5487 DVSS.n5486 0.000854331
R41557 DVSS.n6077 DVSS.n6076 0.000854331
R41558 DVSS.n6778 DVSS.n6777 0.000854331
R41559 DVSS.n3586 DVSS.n3585 0.000854331
R41560 DVSS.n10313 DVSS.n10312 0.000852113
R41561 DVSS.n10310 DVSS.n10309 0.000852113
R41562 DVSS.n10328 DVSS.n10327 0.000852113
R41563 DVSS.n10332 DVSS.n10331 0.000852113
R41564 DVSS.n10336 DVSS.n10335 0.000852113
R41565 DVSS.n10344 DVSS.n10343 0.000852113
R41566 DVSS.n10348 DVSS.n10347 0.000852113
R41567 DVSS.n10423 DVSS.n10422 0.000852113
R41568 DVSS.n10426 DVSS.n10425 0.000852113
R41569 DVSS.n10482 DVSS.n10481 0.000852113
R41570 DVSS.n10485 DVSS.n10484 0.000852113
R41571 DVSS.n10578 DVSS.n10577 0.000852113
R41572 DVSS.n10581 DVSS.n10580 0.000852113
R41573 DVSS.n9329 DVSS.n9328 0.00083
R41574 DVSS.n1309 DVSS.n1308 0.00083
R41575 DVSS.n7218 DVSS.n7217 0.00083
R41576 DVSS.n7245 DVSS.n7244 0.00083
R41577 DVSS.n7292 DVSS.n7291 0.00083
R41578 DVSS.n18878 DVSS.n18877 0.00083
R41579 DVSS.n18904 DVSS.n18903 0.00083
R41580 DVSS.n14588 DVSS.n14587 0.00083
R41581 DVSS.n7892 DVSS.n7891 0.00083
R41582 DVSS.n13478 DVSS.n13477 0.00083
R41583 DVSS.n13476 DVSS.n13475 0.00083
R41584 DVSS.n7949 DVSS.n7948 0.00083
R41585 DVSS.n7924 DVSS.n7923 0.00083
R41586 DVSS.n7922 DVSS.n7921 0.00083
R41587 DVSS.n12127 DVSS.n12126 0.00083
R41588 DVSS.n12134 DVSS.n12133 0.00083
R41589 DVSS.n12129 DVSS.n12128 0.00083
R41590 DVSS.n12021 DVSS.n12020 0.00083
R41591 DVSS.n19097 DVSS.n19096 0.00083
R41592 DVSS.n19363 DVSS.n19362 0.00083
R41593 DVSS.n19846 DVSS.n19845 0.00083
R41594 DVSS.n20645 DVSS.n20644 0.00083
R41595 DVSS.n834 DVSS.n833 0.00083
R41596 DVSS.n1121 DVSS.n1120 0.00083
R41597 DVSS.n283 DVSS.n282 0.00083
R41598 DVSS.n21271 DVSS.n21270 0.00083
R41599 DVSS.n21265 DVSS.n21264 0.00083
R41600 DVSS.n4806 DVSS.n4804 0.000821429
R41601 DVSS.n4780 DVSS.n4779 0.000821429
R41602 DVSS.n4808 DVSS.n4807 0.000821429
R41603 DVSS.n4781 DVSS.n4775 0.000821429
R41604 DVSS.n4764 DVSS.n4760 0.000821429
R41605 DVSS.n8069 DVSS.n8068 0.000821429
R41606 DVSS.n8067 DVSS.n8066 0.000821429
R41607 DVSS.n8070 DVSS.n8067 0.000821429
R41608 DVSS.n8083 DVSS.n8082 0.000821429
R41609 DVSS.n8086 DVSS.n8085 0.000821429
R41610 DVSS.n8090 DVSS.n8089 0.000821429
R41611 DVSS.n11748 DVSS.n11747 0.000821429
R41612 DVSS.n11745 DVSS.n11744 0.000821429
R41613 DVSS.n11762 DVSS.n11761 0.000821429
R41614 DVSS.n11768 DVSS.n11767 0.000821429
R41615 DVSS.n11775 DVSS.n11774 0.000821429
R41616 DVSS.n11778 DVSS.n11777 0.000821429
R41617 DVSS.n11852 DVSS.n11851 0.000821429
R41618 DVSS.n11855 DVSS.n11854 0.000821429
R41619 DVSS.n11911 DVSS.n11910 0.000821429
R41620 DVSS.n11914 DVSS.n11913 0.000821429
R41621 DVSS.n8361 DVSS.n8360 0.000821429
R41622 DVSS.n8359 DVSS.n8358 0.000821429
R41623 DVSS.n8362 DVSS.n8359 0.000821429
R41624 DVSS.n8375 DVSS.n8374 0.000821429
R41625 DVSS.n8378 DVSS.n8377 0.000821429
R41626 DVSS.n8382 DVSS.n8381 0.000821429
R41627 DVSS.n8604 DVSS.n8603 0.000821429
R41628 DVSS.n8607 DVSS.n8604 0.000821429
R41629 DVSS.n8624 DVSS.n8623 0.000821429
R41630 DVSS.n8632 DVSS.n8631 0.000821429
R41631 DVSS.n8650 DVSS.n8649 0.000821429
R41632 DVSS.n8606 DVSS.n8605 0.000821429
R41633 DVSS.n7913 DVSS.n80 0.00082
R41634 DVSS.n20673 DVSS.n20619 0.00082
R41635 DVSS.n21107 DVSS.n21106 0.00082
R41636 DVSS.n9272 DVSS.n9270 0.0008
R41637 DVSS.n9325 DVSS.n9323 0.0008
R41638 DVSS.n9454 DVSS.n9452 0.0008
R41639 DVSS.n9439 DVSS.n9436 0.0008
R41640 DVSS.n9273 DVSS.n9269 0.0008
R41641 DVSS.n9326 DVSS.n9322 0.0008
R41642 DVSS.n9455 DVSS.n9451 0.0008
R41643 DVSS.n9441 DVSS.n9440 0.0008
R41644 DVSS.n3514 DVSS.n3513 0.0008
R41645 DVSS.n3728 DVSS.n3727 0.0008
R41646 DVSS.n13482 DVSS.n13474 0.0008
R41647 DVSS.n13481 DVSS.n13480 0.0008
R41648 DVSS.n7928 DVSS.n7920 0.0008
R41649 DVSS.n7927 DVSS.n7926 0.0008
R41650 DVSS.n12132 DVSS.n12131 0.0008
R41651 DVSS.n12023 DVSS.n12019 0.0008
R41652 DVSS.n19052 DVSS.n19051 0.0008
R41653 DVSS.n19055 DVSS.n19054 0.0008
R41654 DVSS.n20327 DVSS.n20320 0.0008
R41655 DVSS.n20326 DVSS.n20325 0.0008
R41656 DVSS.n20612 DVSS.n20605 0.0008
R41657 DVSS.n20611 DVSS.n20610 0.0008
R41658 DVSS.n20634 DVSS.n20629 0.0008
R41659 DVSS.n11 DVSS.n6 0.0008
R41660 DVSS.n687 DVSS.n686 0.0008
R41661 DVSS.n720 DVSS.n719 0.0008
R41662 DVSS.n20872 DVSS.n20865 0.0008
R41663 DVSS.n20871 DVSS.n20870 0.0008
R41664 DVSS.n21098 DVSS.n21091 0.0008
R41665 DVSS.n21097 DVSS.n21096 0.0008
R41666 DVSS.n21381 DVSS.n21380 0.0008
R41667 DVSS.n20874 DVSS.n20708 0.0008
R41668 DVSS.n21100 DVSS.n20937 0.0008
R41669 DVSS.n21349 DVSS.n21275 0.0008
R41670 DVSS.n21379 DVSS.n21377 0.0008
R41671 DVSS.n20328 DVSS.n20113 0.0008
R41672 DVSS.n20613 DVSS.n20599 0.0008
R41673 DVSS.n20635 DVSS.n20626 0.0008
R41674 DVSS.n12 DVSS.n4 0.0008
R41675 DVSS.n13483 DVSS.n13466 0.0008
R41676 DVSS.n7929 DVSS.n7914 0.0008
R41677 DVSS.n12121 DVSS.n12119 0.0008
R41678 DVSS.n12025 DVSS.n12018 0.0008
R41679 DVSS.n5307 DVSS.n5270 0.00078169
R41680 DVSS.n5187 DVSS.n5186 0.00078169
R41681 DVSS.n5149 DVSS.n5148 0.00078169
R41682 DVSS.n5095 DVSS.n5094 0.00078169
R41683 DVSS.n5308 DVSS.n5268 0.00078169
R41684 DVSS.n5248 DVSS.n5247 0.00078169
R41685 DVSS.n5245 DVSS.n5244 0.00078169
R41686 DVSS.n5236 DVSS.n5190 0.00078169
R41687 DVSS.n5188 DVSS.n5185 0.00078169
R41688 DVSS.n5184 DVSS.n5183 0.00078169
R41689 DVSS.n5165 DVSS.n5164 0.00078169
R41690 DVSS.n5162 DVSS.n5161 0.00078169
R41691 DVSS.n5153 DVSS.n5152 0.00078169
R41692 DVSS.n5150 DVSS.n5147 0.00078169
R41693 DVSS.n5146 DVSS.n5145 0.00078169
R41694 DVSS.n5111 DVSS.n5110 0.00078169
R41695 DVSS.n5108 DVSS.n5107 0.00078169
R41696 DVSS.n5099 DVSS.n5098 0.00078169
R41697 DVSS.n5096 DVSS.n5093 0.00078169
R41698 DVSS.n5092 DVSS.n5091 0.00078169
R41699 DVSS.n10407 DVSS.n10406 0.00078169
R41700 DVSS.n10414 DVSS.n10413 0.00078169
R41701 DVSS.n10466 DVSS.n10465 0.00078169
R41702 DVSS.n10473 DVSS.n10472 0.00078169
R41703 DVSS.n10900 DVSS.n10899 0.00078169
R41704 DVSS.n10569 DVSS.n10568 0.00078169
R41705 DVSS.n4643 DVSS.n4640 0.000757143
R41706 DVSS.n4957 DVSS.n4956 0.000757143
R41707 DVSS.n4913 DVSS.n4912 0.000757143
R41708 DVSS.n4853 DVSS.n4852 0.000757143
R41709 DVSS.n4645 DVSS.n4644 0.000757143
R41710 DVSS.n4971 DVSS.n4970 0.000757143
R41711 DVSS.n4958 DVSS.n4954 0.000757143
R41712 DVSS.n4927 DVSS.n4926 0.000757143
R41713 DVSS.n4914 DVSS.n4910 0.000757143
R41714 DVSS.n4867 DVSS.n4866 0.000757143
R41715 DVSS.n4854 DVSS.n4851 0.000757143
R41716 DVSS.n4812 DVSS.n4811 0.000757143
R41717 DVSS.n4784 DVSS.n4783 0.000757143
R41718 DVSS.n6813 DVSS.n6809 0.000757143
R41719 DVSS.n3965 DVSS.n3931 0.000757143
R41720 DVSS.n3901 DVSS.n3900 0.000757143
R41721 DVSS.n3855 DVSS.n3854 0.000757143
R41722 DVSS.n6814 DVSS.n6807 0.000757143
R41723 DVSS.n3966 DVSS.n3929 0.000757143
R41724 DVSS.n3902 DVSS.n3899 0.000757143
R41725 DVSS.n3856 DVSS.n3853 0.000757143
R41726 DVSS.n3612 DVSS.n3611 0.000757143
R41727 DVSS.n2604 DVSS.n2598 0.000757143
R41728 DVSS.n2693 DVSS.n2692 0.000757143
R41729 DVSS.n2639 DVSS.n2638 0.000757143
R41730 DVSS.n3614 DVSS.n3613 0.000757143
R41731 DVSS.n2606 DVSS.n2605 0.000757143
R41732 DVSS.n2710 DVSS.n2709 0.000757143
R41733 DVSS.n2707 DVSS.n2706 0.000757143
R41734 DVSS.n2697 DVSS.n2696 0.000757143
R41735 DVSS.n2694 DVSS.n2691 0.000757143
R41736 DVSS.n2690 DVSS.n2689 0.000757143
R41737 DVSS.n2656 DVSS.n2655 0.000757143
R41738 DVSS.n2653 DVSS.n2652 0.000757143
R41739 DVSS.n2643 DVSS.n2642 0.000757143
R41740 DVSS.n2640 DVSS.n2637 0.000757143
R41741 DVSS.n2636 DVSS.n2635 0.000757143
R41742 DVSS.n11836 DVSS.n11835 0.000757143
R41743 DVSS.n11843 DVSS.n11842 0.000757143
R41744 DVSS.n11895 DVSS.n11894 0.000757143
R41745 DVSS.n11902 DVSS.n11901 0.000757143
R41746 DVSS.n5910 DVSS.n5873 0.000757143
R41747 DVSS.n5979 DVSS.n5978 0.000757143
R41748 DVSS.n5933 DVSS.n5932 0.000757143
R41749 DVSS.n6046 DVSS.n6045 0.000757143
R41750 DVSS.n5980 DVSS.n5977 0.000757143
R41751 DVSS.n5934 DVSS.n5931 0.000757143
R41752 DVSS.n6107 DVSS.n6106 0.000757143
R41753 DVSS.n6243 DVSS.n6242 0.000757143
R41754 DVSS.n6231 DVSS.n6227 0.000757143
R41755 DVSS.n6185 DVSS.n6184 0.000757143
R41756 DVSS.n6173 DVSS.n6169 0.000757143
R41757 DVSS.n8602 DVSS.n8601 0.000757143
R41758 DVSS.n8627 DVSS.n8626 0.000757143
R41759 DVSS.n6105 DVSS.n6103 0.000757143
R41760 DVSS.n6230 DVSS.n6229 0.000757143
R41761 DVSS.n6172 DVSS.n6171 0.000757143
R41762 DVSS.n5403 DVSS.n5402 0.000751397
R41763 DVSS.n10624 DVSS.n10621 0.000751397
R41764 DVSS.n8029 DVSS.n8026 0.000751397
R41765 DVSS.n1374 DVSS.n1372 0.000751397
R41766 DVSS.n14571 DVSS.n14570 0.00074
R41767 DVSS.n13482 DVSS.n13481 0.00074
R41768 DVSS.n7928 DVSS.n7927 0.00074
R41769 DVSS.n20041 DVSS.n20040 0.00074
R41770 DVSS.n20327 DVSS.n20326 0.00074
R41771 DVSS.n20612 DVSS.n20611 0.00074
R41772 DVSS.n465 DVSS.n464 0.00074
R41773 DVSS.n20872 DVSS.n20871 0.00074
R41774 DVSS.n21098 DVSS.n21097 0.00074
R41775 DVSS.n16596 DVSS.n16595 0.000725
R41776 DVSS.n16607 DVSS.n16606 0.000725
R41777 DVSS DVSS.n15105 0.000725
R41778 DVSS.n18309 DVSS.n18308 0.000725
R41779 DVSS.n18320 DVSS.n18319 0.000725
R41780 DVSS.n10340 DVSS.n10339 0.000711268
R41781 DVSS.n5311 DVSS.n5070 0.000711268
R41782 DVSS.n5237 DVSS.n5236 0.000711268
R41783 DVSS.n5154 DVSS.n5153 0.000711268
R41784 DVSS.n5100 DVSS.n5099 0.000711268
R41785 DVSS.n10308 DVSS.n10307 0.000711268
R41786 DVSS.n10311 DVSS.n10310 0.000711268
R41787 DVSS.n10327 DVSS.n10326 0.000711268
R41788 DVSS.n10331 DVSS.n10330 0.000711268
R41789 DVSS.n10341 DVSS.n10337 0.000711268
R41790 DVSS.n10347 DVSS.n10346 0.000711268
R41791 DVSS.n16561 DVSS.n16560 0.000711268
R41792 DVSS.n16566 DVSS.n16565 0.000711268
R41793 DVSS.n16587 DVSS.n16586 0.000711268
R41794 DVSS.n16080 DVSS.n16079 0.000711268
R41795 DVSS.n16077 DVSS.n16076 0.000711268
R41796 DVSS.n17739 DVSS.n17738 0.000711268
R41797 DVSS.n18117 DVSS.n18116 0.000711268
R41798 DVSS.n18133 DVSS.n18132 0.000711268
R41799 DVSS.n18148 DVSS.n18147 0.000711268
R41800 DVSS.n18254 DVSS.n18253 0.000711268
R41801 DVSS.n18252 DVSS.n18251 0.000711268
R41802 DVSS.n18245 DVSS.n18244 0.000711268
R41803 DVSS.n18231 DVSS.n18230 0.000711268
R41804 DVSS.n18171 DVSS.n18170 0.000711268
R41805 DVSS.n18460 DVSS.n18459 0.000711268
R41806 DVSS.n14462 DVSS.n14461 0.000711268
R41807 DVSS.n14511 DVSS.n14510 0.000711268
R41808 DVSS.n19673 DVSS.n19672 0.000711268
R41809 DVSS.n19801 DVSS.n19800 0.000711268
R41810 DVSS.n153 DVSS.n152 0.000711268
R41811 DVSS.n242 DVSS.n241 0.000711268
R41812 DVSS.n16748 DVSS.n16747 0.000711268
R41813 DVSS.n16753 DVSS.n16752 0.000711268
R41814 DVSS.n16774 DVSS.n16773 0.000711268
R41815 DVSS.n15972 DVSS.n15971 0.000711268
R41816 DVSS.n15969 DVSS.n15968 0.000711268
R41817 DVSS.n15924 DVSS.n15923 0.000711268
R41818 DVSS.n15407 DVSS.n15406 0.000711268
R41819 DVSS.n15438 DVSS.n15422 0.000711268
R41820 DVSS.n15453 DVSS.n15452 0.000711268
R41821 DVSS.n15486 DVSS.n15485 0.000711268
R41822 DVSS.n15488 DVSS.n15487 0.000711268
R41823 DVSS.n15495 DVSS.n15494 0.000711268
R41824 DVSS.n15509 DVSS.n15508 0.000711268
R41825 DVSS.n15569 DVSS.n15568 0.000711268
R41826 DVSS.n15157 DVSS.n15141 0.000711268
R41827 DVSS.n14660 DVSS.n14659 0.000711268
R41828 DVSS.n14608 DVSS.n14607 0.000711268
R41829 DVSS.n19888 DVSS.n19887 0.000711268
R41830 DVSS.n20026 DVSS.n20025 0.000711268
R41831 DVSS.n313 DVSS.n312 0.000711268
R41832 DVSS.n450 DVSS.n449 0.000711268
R41833 DVSS.n9220 DVSS.n9219 0.00071
R41834 DVSS.n9222 DVSS.n9221 0.00071
R41835 DVSS.n9223 DVSS.n9222 0.00071
R41836 DVSS.n3720 DVSS.n3719 0.00071
R41837 DVSS.n12007 DVSS.n12006 0.00071
R41838 DVSS.n19063 DVSS.n19062 0.00071
R41839 DVSS.n20047 DVSS.n20046 0.00071
R41840 DVSS.n20046 DVSS.n20045 0.00071
R41841 DVSS.n20639 DVSS.n20638 0.00071
R41842 DVSS.n792 DVSS.n791 0.00071
R41843 DVSS.n471 DVSS.n470 0.00071
R41844 DVSS.n470 DVSS.n469 0.00071
R41845 DVSS.n21254 DVSS.n21253 0.00071
R41846 DVSS.n473 DVSS.n472 0.00071
R41847 DVSS.n20048 DVSS.n19852 0.00071
R41848 DVSS.n14580 DVSS.n14566 0.00071
R41849 DVSS.n4778 DVSS.n4777 0.000692857
R41850 DVSS.n4636 DVSS.n4635 0.000692857
R41851 DVSS.n4774 DVSS.n4773 0.000692857
R41852 DVSS.n8094 DVSS.n8093 0.000692857
R41853 DVSS.n6816 DVSS.n6798 0.000692857
R41854 DVSS.n3968 DVSS.n3826 0.000692857
R41855 DVSS.n3905 DVSS.n3904 0.000692857
R41856 DVSS.n3859 DVSS.n3858 0.000692857
R41857 DVSS.n8095 DVSS.n8091 0.000692857
R41858 DVSS.n8100 DVSS.n8099 0.000692857
R41859 DVSS.n11772 DVSS.n11771 0.000692857
R41860 DVSS.n3606 DVSS.n3605 0.000692857
R41861 DVSS.n2595 DVSS.n2594 0.000692857
R41862 DVSS.n2698 DVSS.n2697 0.000692857
R41863 DVSS.n2644 DVSS.n2643 0.000692857
R41864 DVSS.n11743 DVSS.n11742 0.000692857
R41865 DVSS.n11746 DVSS.n11745 0.000692857
R41866 DVSS.n11761 DVSS.n11760 0.000692857
R41867 DVSS.n11764 DVSS.n11763 0.000692857
R41868 DVSS.n11773 DVSS.n11769 0.000692857
R41869 DVSS.n11777 DVSS.n11776 0.000692857
R41870 DVSS.n8386 DVSS.n8385 0.000692857
R41871 DVSS.n6049 DVSS.n5871 0.000692857
R41872 DVSS.n5983 DVSS.n5982 0.000692857
R41873 DVSS.n5937 DVSS.n5936 0.000692857
R41874 DVSS.n8387 DVSS.n8383 0.000692857
R41875 DVSS.n8392 DVSS.n8391 0.000692857
R41876 DVSS.n6099 DVSS.n6098 0.000692857
R41877 DVSS.n6235 DVSS.n6234 0.000692857
R41878 DVSS.n6177 DVSS.n6176 0.000692857
R41879 DVSS.n8637 DVSS.n8633 0.000692857
R41880 DVSS.n8642 DVSS.n8641 0.000692857
R41881 DVSS.n8636 DVSS.n8635 0.000692857
R41882 DVSS.n12771 DVSS.n12766 0.000692308
R41883 DVSS.n12743 DVSS.n12742 0.000692308
R41884 DVSS.n12616 DVSS.n12611 0.000692308
R41885 DVSS.n12593 DVSS.n12592 0.000692308
R41886 DVSS.n12328 DVSS.n12323 0.000692308
R41887 DVSS.n12305 DVSS.n12304 0.000692308
R41888 DVSS.n12236 DVSS.n12231 0.000692308
R41889 DVSS.n21341 DVSS.n21340 0.000692308
R41890 DVSS.n3383 DVSS.n3378 0.000692308
R41891 DVSS.n2781 DVSS.n2780 0.000692308
R41892 DVSS.n3240 DVSS.n3235 0.000692308
R41893 DVSS.n3217 DVSS.n3216 0.000692308
R41894 DVSS.n2955 DVSS.n2950 0.000692308
R41895 DVSS.n2932 DVSS.n2931 0.000692308
R41896 DVSS.n2863 DVSS.n2858 0.000692308
R41897 DVSS.n890 DVSS.n885 0.000692308
R41898 DVSS.n3406 DVSS.n3405 0.000692308
R41899 DVSS.n12780 DVSS.n12779 0.000692308
R41900 DVSS.n14126 DVSS.n14125 0.00068
R41901 DVSS.n14579 DVSS.n14578 0.00068
R41902 DVSS.n14573 DVSS.n14572 0.00068
R41903 DVSS.n20043 DVSS.n20042 0.00068
R41904 DVSS.n467 DVSS.n466 0.00068
R41905 DVSS.n21363 DVSS 0.00068
R41906 DVSS DVSS.n21364 0.00068
R41907 DVSS.n4446 DVSS.n4445 0.000677165
R41908 DVSS.n4390 DVSS.n4389 0.000677165
R41909 DVSS.n7204 DVSS.n7203 0.000677165
R41910 DVSS.n19134 DVSS.n19133 0.000677165
R41911 DVSS.n19151 DVSS.n19150 0.000677165
R41912 DVSS.n19209 DVSS.n19208 0.000677165
R41913 DVSS.n19290 DVSS.n19289 0.000677165
R41914 DVSS.n862 DVSS.n861 0.000677165
R41915 DVSS.n1045 DVSS.n1044 0.000677165
R41916 DVSS.n986 DVSS.n985 0.000677165
R41917 DVSS.n9513 DVSS.n9512 0.000677165
R41918 DVSS.n9576 DVSS.n9575 0.000677165
R41919 DVSS.n12896 DVSS.n12895 0.000677165
R41920 DVSS.n12832 DVSS.n12831 0.000677165
R41921 DVSS.n12822 DVSS.n12821 0.000677165
R41922 DVSS.n12819 DVSS.n12818 0.000677165
R41923 DVSS.n12764 DVSS.n12763 0.000677165
R41924 DVSS.n12744 DVSS.n12734 0.000677165
R41925 DVSS.n12711 DVSS.n12710 0.000677165
R41926 DVSS.n12690 DVSS.n12689 0.000677165
R41927 DVSS.n12675 DVSS.n12674 0.000677165
R41928 DVSS.n12442 DVSS.n12441 0.000677165
R41929 DVSS.n12441 DVSS.n12440 0.000677165
R41930 DVSS.n12437 DVSS.n12436 0.000677165
R41931 DVSS.n12420 DVSS.n12419 0.000677165
R41932 DVSS.n12398 DVSS.n12397 0.000677165
R41933 DVSS.n12387 DVSS.n12386 0.000677165
R41934 DVSS.n12168 DVSS.n12167 0.000677165
R41935 DVSS.n12167 DVSS.n12166 0.000677165
R41936 DVSS.n12166 DVSS.n12165 0.000677165
R41937 DVSS.n12159 DVSS.n12158 0.000677165
R41938 DVSS.n21230 DVSS.n21229 0.000677165
R41939 DVSS.n21278 DVSS.n21277 0.000677165
R41940 DVSS.n21303 DVSS.n21302 0.000677165
R41941 DVSS.n21227 DVSS.n21226 0.000677165
R41942 DVSS.n21194 DVSS.n21193 0.000677165
R41943 DVSS.n21342 DVSS.n21330 0.000677165
R41944 DVSS.n21144 DVSS.n21143 0.000677165
R41945 DVSS.n15684 DVSS.n15683 0.000677165
R41946 DVSS.n15621 DVSS.n15620 0.000677165
R41947 DVSS.n13507 DVSS.n13506 0.000677165
R41948 DVSS.n20162 DVSS.n20161 0.000677165
R41949 DVSS.n20306 DVSS.n20305 0.000677165
R41950 DVSS.n20847 DVSS.n20846 0.000677165
R41951 DVSS.n20812 DVSS.n20811 0.000677165
R41952 DVSS.n10793 DVSS.n10792 0.000677165
R41953 DVSS.n10738 DVSS.n10737 0.000677165
R41954 DVSS.n11551 DVSS.n11550 0.000677165
R41955 DVSS.n11614 DVSS.n11613 0.000677165
R41956 DVSS.n12081 DVSS.n12080 0.000677165
R41957 DVSS.n63 DVSS.n62 0.000677165
R41958 DVSS.n21545 DVSS.n21544 0.000677165
R41959 DVSS.n21482 DVSS.n21481 0.000677165
R41960 DVSS.n21457 DVSS.n21456 0.000677165
R41961 DVSS.n21394 DVSS.n21393 0.000677165
R41962 DVSS.n4284 DVSS.n4283 0.000677165
R41963 DVSS.n4340 DVSS.n4339 0.000677165
R41964 DVSS.n3503 DVSS.n3502 0.000677165
R41965 DVSS.n3444 DVSS.n3443 0.000677165
R41966 DVSS.n3434 DVSS.n3433 0.000677165
R41967 DVSS.n3431 DVSS.n3430 0.000677165
R41968 DVSS.n3376 DVSS.n3375 0.000677165
R41969 DVSS.n3357 DVSS.n3356 0.000677165
R41970 DVSS.n3334 DVSS.n3333 0.000677165
R41971 DVSS.n3313 DVSS.n3312 0.000677165
R41972 DVSS.n3299 DVSS.n3298 0.000677165
R41973 DVSS.n3069 DVSS.n3068 0.000677165
R41974 DVSS.n3068 DVSS.n3067 0.000677165
R41975 DVSS.n3063 DVSS.n3062 0.000677165
R41976 DVSS.n3047 DVSS.n3046 0.000677165
R41977 DVSS.n3024 DVSS.n3023 0.000677165
R41978 DVSS.n3014 DVSS.n3013 0.000677165
R41979 DVSS.n2796 DVSS.n2795 0.000677165
R41980 DVSS.n2795 DVSS.n2794 0.000677165
R41981 DVSS.n2794 DVSS.n2793 0.000677165
R41982 DVSS.n2787 DVSS.n2786 0.000677165
R41983 DVSS.n760 DVSS.n759 0.000677165
R41984 DVSS.n655 DVSS.n654 0.000677165
R41985 DVSS.n666 DVSS.n665 0.000677165
R41986 DVSS.n757 DVSS.n756 0.000677165
R41987 DVSS.n801 DVSS.n800 0.000677165
R41988 DVSS.n729 DVSS.n728 0.000677165
R41989 DVSS.n697 DVSS.n696 0.000677165
R41990 DVSS.n9681 DVSS.n9680 0.000677165
R41991 DVSS.n9618 DVSS.n9617 0.000677165
R41992 DVSS.n13409 DVSS.n13408 0.000677165
R41993 DVSS.n20433 DVSS.n20432 0.000677165
R41994 DVSS.n20580 DVSS.n20579 0.000677165
R41995 DVSS.n21073 DVSS.n21072 0.000677165
R41996 DVSS.n21038 DVSS.n21037 0.000677165
R41997 DVSS.n16196 DVSS.n16195 0.000677165
R41998 DVSS.n16139 DVSS.n16138 0.000677165
R41999 DVSS.n18864 DVSS.n18863 0.000677165
R42000 DVSS.n19408 DVSS.n19407 0.000677165
R42001 DVSS.n19425 DVSS.n19424 0.000677165
R42002 DVSS.n19480 DVSS.n19479 0.000677165
R42003 DVSS.n19561 DVSS.n19560 0.000677165
R42004 DVSS.n1149 DVSS.n1148 0.000677165
R42005 DVSS.n1260 DVSS.n1259 0.000677165
R42006 DVSS.n1202 DVSS.n1201 0.000677165
R42007 DVSS.n5471 DVSS.n5470 0.000677165
R42008 DVSS.n5855 DVSS.n5854 0.000677165
R42009 DVSS.n6598 DVSS.n6597 0.000677165
R42010 DVSS.n6655 DVSS.n6654 0.000677165
R42011 DVSS.n3565 DVSS.n3564 0.000677165
R42012 DVSS.n18962 DVSS.n18961 0.000677165
R42013 DVSS.n19009 DVSS.n19008 0.000677165
R42014 DVSS.n540 DVSS.n539 0.000677165
R42015 DVSS.n611 DVSS.n610 0.000677165
R42016 DVSS.n555 DVSS.n554 0.000677165
R42017 DVSS.n9174 DVSS.n9172 0.00065
R42018 DVSS.n9171 DVSS.n9170 0.00065
R42019 DVSS.n9175 DVSS.n9171 0.00065
R42020 DVSS.n9188 DVSS.n9187 0.00065
R42021 DVSS.n9191 DVSS.n9190 0.00065
R42022 DVSS.n9195 DVSS.n9194 0.00065
R42023 DVSS.n14122 DVSS.n14121 0.00065
R42024 DVSS.n14532 DVSS.n14531 0.00065
R42025 DVSS.n14598 DVSS.n14597 0.00065
R42026 DVSS.n14584 DVSS.n14583 0.00065
R42027 DVSS.n14589 DVSS.n14588 0.00065
R42028 DVSS.n13480 DVSS.n13479 0.00065
R42029 DVSS.n13477 DVSS.n13476 0.00065
R42030 DVSS.n7926 DVSS.n7925 0.00065
R42031 DVSS.n7923 DVSS.n7922 0.00065
R42032 DVSS.n19627 DVSS.n19626 0.00065
R42033 DVSS.n19629 DVSS.n19627 0.00065
R42034 DVSS.n19829 DVSS.n19828 0.00065
R42035 DVSS.n19847 DVSS.n19846 0.00065
R42036 DVSS.n114 DVSS.n113 0.00065
R42037 DVSS.n116 DVSS.n114 0.00065
R42038 DVSS.n265 DVSS.n264 0.00065
R42039 DVSS.n284 DVSS.n283 0.00065
R42040 DVSS.n117 DVSS.n109 0.00065
R42041 DVSS.n266 DVSS.n124 0.00065
R42042 DVSS.n19630 DVSS.n19622 0.00065
R42043 DVSS.n19830 DVSS.n19820 0.00065
R42044 DVSS.n14114 DVSS.n14112 0.00065
R42045 DVSS.n14534 DVSS.n14533 0.00065
R42046 DVSS.n10402 DVSS.n10401 0.000640845
R42047 DVSS.n10461 DVSS.n10460 0.000640845
R42048 DVSS.n10559 DVSS.n10503 0.000640845
R42049 DVSS.n10887 DVSS.n10567 0.000640845
R42050 DVSS.n5266 DVSS.n5265 0.000640845
R42051 DVSS.n10314 DVSS.n10311 0.000640845
R42052 DVSS.n10343 DVSS.n10342 0.000640845
R42053 DVSS.n10404 DVSS.n10403 0.000640845
R42054 DVSS.n10415 DVSS.n10414 0.000640845
R42055 DVSS.n10463 DVSS.n10462 0.000640845
R42056 DVSS.n10474 DVSS.n10473 0.000640845
R42057 DVSS.n10561 DVSS.n10560 0.000640845
R42058 DVSS.n10570 DVSS.n10569 0.000640845
R42059 DVSS.n10886 DVSS.n10885 0.000640845
R42060 DVSS.n10884 DVSS.n10883 0.000640845
R42061 DVSS.n10872 DVSS.n10871 0.000640845
R42062 DVSS.n4577 DVSS.n4575 0.000638889
R42063 DVSS.n11015 DVSS.n11012 0.000638889
R42064 DVSS.n6762 DVSS.n6760 0.000638889
R42065 DVSS.n11675 DVSS.n11672 0.000638889
R42066 DVSS.n6707 DVSS.n6705 0.000638889
R42067 DVSS.n11638 DVSS.n11635 0.000638889
R42068 DVSS.n2539 DVSS.n2537 0.000638889
R42069 DVSS.n11513 DVSS.n11510 0.000638889
R42070 DVSS.n4523 DVSS.n4521 0.000638889
R42071 DVSS.n11185 DVSS.n11182 0.000638889
R42072 DVSS.n6400 DVSS.n6398 0.000638889
R42073 DVSS.n11476 DVSS.n11472 0.000638889
R42074 DVSS.n6889 DVSS.n6887 0.000638889
R42075 DVSS.n11724 DVSS.n11721 0.000638889
R42076 DVSS.n5507 DVSS.n5505 0.000638889
R42077 DVSS.n10025 DVSS.n10022 0.000638889
R42078 DVSS.n10725 DVSS.n10694 0.000628571
R42079 DVSS.n5058 DVSS.n5057 0.000628571
R42080 DVSS.n4960 DVSS.n4959 0.000628571
R42081 DVSS.n4916 DVSS.n4915 0.000628571
R42082 DVSS.n4856 DVSS.n4855 0.000628571
R42083 DVSS.n4772 DVSS.n4771 0.000628571
R42084 DVSS.n10065 DVSS.n10064 0.000628571
R42085 DVSS.n10129 DVSS.n10128 0.000628571
R42086 DVSS.n10141 DVSS.n10140 0.000628571
R42087 DVSS.n10177 DVSS.n10176 0.000628571
R42088 DVSS.n10695 DVSS.n10192 0.000628571
R42089 DVSS.n10724 DVSS.n10723 0.000628571
R42090 DVSS.n10733 DVSS.n10644 0.000628571
R42091 DVSS.n10656 DVSS.n10655 0.000628571
R42092 DVSS.n8286 DVSS.n8235 0.000628571
R42093 DVSS.n8320 DVSS.n8319 0.000628571
R42094 DVSS.n8097 DVSS.n8096 0.000628571
R42095 DVSS.n8151 DVSS.n8150 0.000628571
R42096 DVSS.n8160 DVSS.n8159 0.000628571
R42097 DVSS.n8202 DVSS.n8201 0.000628571
R42098 DVSS.n8211 DVSS.n8210 0.000628571
R42099 DVSS.n8288 DVSS.n8287 0.000628571
R42100 DVSS.n8296 DVSS.n8295 0.000628571
R42101 DVSS.n8322 DVSS.n8321 0.000628571
R42102 DVSS.n13098 DVSS.n13097 0.000628571
R42103 DVSS.n11831 DVSS.n11830 0.000628571
R42104 DVSS.n11890 DVSS.n11889 0.000628571
R42105 DVSS.n11981 DVSS.n11930 0.000628571
R42106 DVSS.n13002 DVSS.n11735 0.000628571
R42107 DVSS.n11749 DVSS.n11746 0.000628571
R42108 DVSS.n11833 DVSS.n11832 0.000628571
R42109 DVSS.n11844 DVSS.n11843 0.000628571
R42110 DVSS.n11892 DVSS.n11891 0.000628571
R42111 DVSS.n11903 DVSS.n11902 0.000628571
R42112 DVSS.n11983 DVSS.n11982 0.000628571
R42113 DVSS.n12990 DVSS.n12989 0.000628571
R42114 DVSS.n13004 DVSS.n13003 0.000628571
R42115 DVSS.n13015 DVSS.n13014 0.000628571
R42116 DVSS.n8583 DVSS.n8527 0.000628571
R42117 DVSS.n11336 DVSS.n8340 0.000628571
R42118 DVSS.n6043 DVSS.n6042 0.000628571
R42119 DVSS.n8389 DVSS.n8388 0.000628571
R42120 DVSS.n8443 DVSS.n8442 0.000628571
R42121 DVSS.n8452 DVSS.n8451 0.000628571
R42122 DVSS.n8494 DVSS.n8493 0.000628571
R42123 DVSS.n8503 DVSS.n8502 0.000628571
R42124 DVSS.n8585 DVSS.n8584 0.000628571
R42125 DVSS.n11324 DVSS.n11323 0.000628571
R42126 DVSS.n11338 DVSS.n11337 0.000628571
R42127 DVSS.n11362 DVSS.n11339 0.000628571
R42128 DVSS.n11351 DVSS.n11350 0.000628571
R42129 DVSS.n6326 DVSS.n6325 0.000628571
R42130 DVSS.n6233 DVSS.n6232 0.000628571
R42131 DVSS.n6175 DVSS.n6174 0.000628571
R42132 DVSS.n8639 DVSS.n8638 0.000628571
R42133 DVSS.n8697 DVSS.n8696 0.000628571
R42134 DVSS.n8713 DVSS.n8712 0.000628571
R42135 DVSS.n8760 DVSS.n8759 0.000628571
R42136 DVSS.n8774 DVSS.n8773 0.000628571
R42137 DVSS.n8861 DVSS.n8860 0.000628571
R42138 DVSS.n8869 DVSS.n8868 0.000628571
R42139 DVSS.n8900 DVSS.n8899 0.000628571
R42140 DVSS.n8902 DVSS.n8901 0.000628571
R42141 DVSS.n8336 DVSS.n8335 0.000628571
R42142 DVSS.n8706 DVSS.n8705 0.000628571
R42143 DVSS.n8859 DVSS.n8803 0.000628571
R42144 DVSS.n8898 DVSS.n8897 0.000628571
R42145 DVSS.n1398 DVSS.n1397 0.00062
R42146 DVSS.n4256 DVSS.n4240 0.00062
R42147 DVSS.n4210 DVSS.n4209 0.00062
R42148 DVSS.n4164 DVSS.n4163 0.00062
R42149 DVSS.n1399 DVSS.n1395 0.00062
R42150 DVSS.n4257 DVSS.n4238 0.00062
R42151 DVSS.n4211 DVSS.n4207 0.00062
R42152 DVSS.n4165 DVSS.n4160 0.00062
R42153 DVSS.n3664 DVSS.n3663 0.00062
R42154 DVSS.n3726 DVSS.n3515 0.00062
R42155 DVSS.n1310 DVSS.n1309 0.00062
R42156 DVSS.n7217 DVSS.n7216 0.00062
R42157 DVSS.n7219 DVSS.n7218 0.00062
R42158 DVSS.n7225 DVSS.n7224 0.00062
R42159 DVSS.n7229 DVSS.n7228 0.00062
R42160 DVSS.n7237 DVSS.n7236 0.00062
R42161 DVSS.n7293 DVSS.n7292 0.00062
R42162 DVSS.n18877 DVSS.n18876 0.00062
R42163 DVSS.n18879 DVSS.n18878 0.00062
R42164 DVSS.n18885 DVSS.n18884 0.00062
R42165 DVSS.n18889 DVSS.n18888 0.00062
R42166 DVSS.n18896 DVSS.n18895 0.00062
R42167 DVSS.n14119 DVSS.n14118 0.00062
R42168 DVSS.n14530 DVSS.n14529 0.00062
R42169 DVSS.n13489 DVSS.n13488 0.00062
R42170 DVSS.n13469 DVSS.n13468 0.00062
R42171 DVSS.n7935 DVSS.n7934 0.00062
R42172 DVSS.n7939 DVSS.n7938 0.00062
R42173 DVSS.n18935 DVSS.n18934 0.00062
R42174 DVSS.n19057 DVSS.n19056 0.00062
R42175 DVSS.n19098 DVSS.n19097 0.00062
R42176 DVSS.n19304 DVSS.n19303 0.00062
R42177 DVSS.n19364 DVSS.n19363 0.00062
R42178 DVSS.n19373 DVSS.n19372 0.00062
R42179 DVSS.n19625 DVSS.n19624 0.00062
R42180 DVSS.n19827 DVSS.n19826 0.00062
R42181 DVSS.n625 DVSS.n624 0.00062
R42182 DVSS.n722 DVSS.n721 0.00062
R42183 DVSS.n835 DVSS.n834 0.00062
R42184 DVSS.n1060 DVSS.n1059 0.00062
R42185 DVSS.n1122 DVSS.n1121 0.00062
R42186 DVSS.n1275 DVSS.n1274 0.00062
R42187 DVSS.n112 DVSS.n111 0.00062
R42188 DVSS.n263 DVSS.n262 0.00062
R42189 DVSS.n627 DVSS.n626 0.00062
R42190 DVSS.n724 DVSS.n723 0.00062
R42191 DVSS.n1062 DVSS.n1061 0.00062
R42192 DVSS.n1277 DVSS.n1276 0.00062
R42193 DVSS.n18937 DVSS.n18936 0.00062
R42194 DVSS.n19059 DVSS.n19058 0.00062
R42195 DVSS.n19306 DVSS.n19305 0.00062
R42196 DVSS.n19375 DVSS.n19374 0.00062
R42197 DVSS.n3665 DVSS.n3530 0.00062
R42198 DVSS.n3725 DVSS.n3517 0.00062
R42199 DVSS.n7231 DVSS.n7230 0.00062
R42200 DVSS.n18890 DVSS.n7290 0.00062
R42201 DVSS DVSS.n2 0.00062
R42202 DVSS.n9200 DVSS.n9198 0.00059
R42203 DVSS.n1401 DVSS.n1388 0.00059
R42204 DVSS.n4259 DVSS.n4146 0.00059
R42205 DVSS.n4214 DVSS.n4213 0.00059
R42206 DVSS.n4168 DVSS.n4167 0.00059
R42207 DVSS.n9201 DVSS.n9196 0.00059
R42208 DVSS.n9206 DVSS.n9205 0.00059
R42209 DVSS.n3661 DVSS.n3531 0.00059
R42210 DVSS.n3729 DVSS.n3514 0.00059
R42211 DVSS.n3713 DVSS.n3712 0.00059
R42212 DVSS.n7222 DVSS.n7221 0.00059
R42213 DVSS.n7224 DVSS.n7223 0.00059
R42214 DVSS.n7239 DVSS.n7238 0.00059
R42215 DVSS.n18882 DVSS.n18881 0.00059
R42216 DVSS.n18884 DVSS.n18883 0.00059
R42217 DVSS.n18898 DVSS.n18897 0.00059
R42218 DVSS.n14120 DVSS.n14119 0.00059
R42219 DVSS.n14123 DVSS.n14122 0.00059
R42220 DVSS.n14525 DVSS.n14524 0.00059
R42221 DVSS.n14529 DVSS.n14528 0.00059
R42222 DVSS.n14595 DVSS.n14082 0.00059
R42223 DVSS.n13487 DVSS.n13486 0.00059
R42224 DVSS.n13473 DVSS.n13472 0.00059
R42225 DVSS.n7933 DVSS.n7932 0.00059
R42226 DVSS.n7919 DVSS.n7918 0.00059
R42227 DVSS.n18932 DVSS.n18931 0.00059
R42228 DVSS.n19053 DVSS.n19052 0.00059
R42229 DVSS.n19068 DVSS.n19067 0.00059
R42230 DVSS.n19102 DVSS.n19101 0.00059
R42231 DVSS.n19368 DVSS.n19367 0.00059
R42232 DVSS.n19836 DVSS.n19833 0.00059
R42233 DVSS.n19842 DVSS.n19841 0.00059
R42234 DVSS.n20655 DVSS.n20654 0.00059
R42235 DVSS.n622 DVSS.n516 0.00059
R42236 DVSS.n718 DVSS.n687 0.00059
R42237 DVSS.n805 DVSS.n796 0.00059
R42238 DVSS.n1056 DVSS.n838 0.00059
R42239 DVSS.n1271 DVSS.n1125 0.00059
R42240 DVSS.n272 DVSS.n269 0.00059
R42241 DVSS.n279 DVSS.n278 0.00059
R42242 DVSS.n21191 DVSS.n21190 0.00059
R42243 DVSS.n274 DVSS.n268 0.00059
R42244 DVSS.n19838 DVSS.n19832 0.00059
R42245 DVSS.n14594 DVSS.n14083 0.00059
R42246 DVSS.n13103 DVSS 0.000585714
R42247 DVSS.n10410 DVSS.n10409 0.000570422
R42248 DVSS.n10469 DVSS.n10468 0.000570422
R42249 DVSS.n10896 DVSS.n10564 0.000570422
R42250 DVSS.n10879 DVSS.n10875 0.000570422
R42251 DVSS.n10329 DVSS.n10328 0.000570422
R42252 DVSS.n10346 DVSS.n10345 0.000570422
R42253 DVSS.n10365 DVSS.n10364 0.000570422
R42254 DVSS.n10368 DVSS.n10367 0.000570422
R42255 DVSS.n10397 DVSS.n10396 0.000570422
R42256 DVSS.n10411 DVSS.n10408 0.000570422
R42257 DVSS.n10456 DVSS.n10455 0.000570422
R42258 DVSS.n10470 DVSS.n10467 0.000570422
R42259 DVSS.n10499 DVSS.n10498 0.000570422
R42260 DVSS.n10898 DVSS.n10897 0.000570422
R42261 DVSS.n10594 DVSS.n10593 0.000570422
R42262 DVSS.n10881 DVSS.n10880 0.000570422
R42263 DVSS.n1997 DVSS.n1996 0.000564286
R42264 DVSS.n2065 DVSS.n2064 0.000564286
R42265 DVSS.n2067 DVSS.n2066 0.000564286
R42266 DVSS.n1998 DVSS.n1995 0.000564286
R42267 DVSS.n10074 DVSS.n10073 0.000564286
R42268 DVSS.n10146 DVSS.n10145 0.000564286
R42269 DVSS.n10187 DVSS.n10185 0.000564286
R42270 DVSS.n10729 DVSS.n10659 0.000564286
R42271 DVSS.n4797 DVSS.n4796 0.000564286
R42272 DVSS.n4790 DVSS.n4789 0.000564286
R42273 DVSS.n4786 DVSS.n4785 0.000564286
R42274 DVSS.n4783 DVSS.n4782 0.000564286
R42275 DVSS.n4770 DVSS.n4769 0.000564286
R42276 DVSS.n10075 DVSS.n10071 0.000564286
R42277 DVSS.n10077 DVSS.n10076 0.000564286
R42278 DVSS.n10136 DVSS.n10135 0.000564286
R42279 DVSS.n10138 DVSS.n10137 0.000564286
R42280 DVSS.n10188 DVSS.n10183 0.000564286
R42281 DVSS.n10190 DVSS.n10189 0.000564286
R42282 DVSS.n10720 DVSS.n10719 0.000564286
R42283 DVSS.n10731 DVSS.n10730 0.000564286
R42284 DVSS.n8156 DVSS.n8155 0.000564286
R42285 DVSS.n8207 DVSS.n8206 0.000564286
R42286 DVSS.n13111 DVSS.n8290 0.000564286
R42287 DVSS.n13101 DVSS.n8293 0.000564286
R42288 DVSS.n8084 DVSS.n8083 0.000564286
R42289 DVSS.n8099 DVSS.n8098 0.000564286
R42290 DVSS.n8146 DVSS.n8145 0.000564286
R42291 DVSS.n8157 DVSS.n8153 0.000564286
R42292 DVSS.n8197 DVSS.n8196 0.000564286
R42293 DVSS.n8208 DVSS.n8204 0.000564286
R42294 DVSS.n8232 DVSS.n8231 0.000564286
R42295 DVSS.n13113 DVSS.n13112 0.000564286
R42296 DVSS.n8316 DVSS.n8315 0.000564286
R42297 DVSS.n13100 DVSS.n13087 0.000564286
R42298 DVSS.n11839 DVSS.n11838 0.000564286
R42299 DVSS.n11898 DVSS.n11897 0.000564286
R42300 DVSS.n12993 DVSS.n11736 0.000564286
R42301 DVSS.n13021 DVSS.n13017 0.000564286
R42302 DVSS.n11794 DVSS.n11793 0.000564286
R42303 DVSS.n11797 DVSS.n11796 0.000564286
R42304 DVSS.n11826 DVSS.n11825 0.000564286
R42305 DVSS.n11840 DVSS.n11837 0.000564286
R42306 DVSS.n11885 DVSS.n11884 0.000564286
R42307 DVSS.n11899 DVSS.n11896 0.000564286
R42308 DVSS.n11927 DVSS.n11926 0.000564286
R42309 DVSS.n12992 DVSS.n12968 0.000564286
R42310 DVSS.n12970 DVSS.n12969 0.000564286
R42311 DVSS.n13023 DVSS.n13022 0.000564286
R42312 DVSS.n8448 DVSS.n8447 0.000564286
R42313 DVSS.n8499 DVSS.n8498 0.000564286
R42314 DVSS.n11327 DVSS.n8341 0.000564286
R42315 DVSS.n11358 DVSS.n11354 0.000564286
R42316 DVSS.n8376 DVSS.n8375 0.000564286
R42317 DVSS.n8391 DVSS.n8390 0.000564286
R42318 DVSS.n8438 DVSS.n8437 0.000564286
R42319 DVSS.n8449 DVSS.n8445 0.000564286
R42320 DVSS.n8489 DVSS.n8488 0.000564286
R42321 DVSS.n8500 DVSS.n8496 0.000564286
R42322 DVSS.n8524 DVSS.n8523 0.000564286
R42323 DVSS.n11326 DVSS.n11300 0.000564286
R42324 DVSS.n11303 DVSS.n11302 0.000564286
R42325 DVSS.n11360 DVSS.n11359 0.000564286
R42326 DVSS.n8619 DVSS.n8614 0.000564286
R42327 DVSS.n8622 DVSS.n8621 0.000564286
R42328 DVSS.n8625 DVSS.n8624 0.000564286
R42329 DVSS.n8628 DVSS.n8627 0.000564286
R42330 DVSS.n8641 DVSS.n8640 0.000564286
R42331 DVSS.n8693 DVSS.n8692 0.000564286
R42332 DVSS.n8709 DVSS.n8703 0.000564286
R42333 DVSS.n8711 DVSS.n8710 0.000564286
R42334 DVSS.n8754 DVSS.n8753 0.000564286
R42335 DVSS.n8770 DVSS.n8766 0.000564286
R42336 DVSS.n8772 DVSS.n8771 0.000564286
R42337 DVSS.n8799 DVSS.n8798 0.000564286
R42338 DVSS.n8922 DVSS.n8921 0.000564286
R42339 DVSS.n8867 DVSS.n8864 0.000564286
R42340 DVSS.n8893 DVSS.n8892 0.000564286
R42341 DVSS.n8907 DVSS.n8904 0.000564286
R42342 DVSS.n8708 DVSS.n8707 0.000564286
R42343 DVSS.n8769 DVSS.n8768 0.000564286
R42344 DVSS.n8920 DVSS.n8865 0.000564286
R42345 DVSS.n8909 DVSS.n8866 0.000564286
R42346 DVSS.n9422 DVSS.n9344 0.00056
R42347 DVSS.n9469 DVSS.n9468 0.00056
R42348 DVSS.n9203 DVSS.n9202 0.00056
R42349 DVSS.n9258 DVSS.n9257 0.00056
R42350 DVSS.n9268 DVSS.n9267 0.00056
R42351 DVSS.n9311 DVSS.n9310 0.00056
R42352 DVSS.n9321 DVSS.n9320 0.00056
R42353 DVSS.n9424 DVSS.n9423 0.00056
R42354 DVSS.n9450 DVSS.n9449 0.00056
R42355 DVSS.n9470 DVSS.n9466 0.00056
R42356 DVSS.n9443 DVSS.n9442 0.00056
R42357 DVSS.n7227 DVSS.n7226 0.00056
R42358 DVSS.n18887 DVSS.n18886 0.00056
R42359 DVSS.n14124 DVSS.n14123 0.00056
R42360 DVSS.n14597 DVSS.n14596 0.00056
R42361 DVSS.n13500 DVSS.n7894 0.00056
R42362 DVSS.n13424 DVSS.n13423 0.00056
R42363 DVSS.n12009 DVSS.n12008 0.00056
R42364 DVSS.n12104 DVSS.n12103 0.00056
R42365 DVSS.n12092 DVSS.n12030 0.00056
R42366 DVSS.n19104 DVSS.n19103 0.00056
R42367 DVSS.n19370 DVSS.n19369 0.00056
R42368 DVSS.n19835 DVSS.n19834 0.00056
R42369 DVSS.n20100 DVSS.n20099 0.00056
R42370 DVSS.n20318 DVSS.n20317 0.00056
R42371 DVSS.n20377 DVSS.n20376 0.00056
R42372 DVSS.n20603 DVSS.n20602 0.00056
R42373 DVSS.n20658 DVSS.n20657 0.00056
R42374 DVSS.n20643 DVSS.n20642 0.00056
R42375 DVSS.n21571 DVSS.n21570 0.00056
R42376 DVSS.n21557 DVSS.n21556 0.00056
R42377 DVSS.n1058 DVSS.n1057 0.00056
R42378 DVSS.n1273 DVSS.n1272 0.00056
R42379 DVSS.n271 DVSS.n270 0.00056
R42380 DVSS.n20693 DVSS.n20692 0.00056
R42381 DVSS.n20863 DVSS.n20862 0.00056
R42382 DVSS.n20922 DVSS.n20921 0.00056
R42383 DVSS.n21089 DVSS.n21088 0.00056
R42384 DVSS.n21256 DVSS.n21255 0.00056
R42385 DVSS.n21269 DVSS.n21265 0.00056
R42386 DVSS.n21371 DVSS.n21370 0.00056
R42387 DVSS.n21383 DVSS.n21382 0.00056
R42388 DVSS.n20695 DVSS.n20694 0.00056
R42389 DVSS.n20924 DVSS.n20923 0.00056
R42390 DVSS.n21258 DVSS.n21257 0.00056
R42391 DVSS.n21369 DVSS.n79 0.00056
R42392 DVSS.n20101 DVSS.n20093 0.00056
R42393 DVSS.n20378 DVSS.n20369 0.00056
R42394 DVSS.n20659 DVSS.n20651 0.00056
R42395 DVSS.n21572 DVSS.n21565 0.00056
R42396 DVSS.n13499 DVSS.n7896 0.00056
R42397 DVSS.n13425 DVSS.n7947 0.00056
R42398 DVSS.n12011 DVSS.n12010 0.00056
R42399 DVSS.n12106 DVSS.n12105 0.00056
R42400 VSS DVSS.n1718 0.000557143
R42401 DVSS.n9264 DVSS.n9262 0.00053
R42402 DVSS.n9317 DVSS.n9315 0.00053
R42403 DVSS.n9485 DVSS.n9426 0.00053
R42404 DVSS.n9446 DVSS.n9429 0.00053
R42405 DVSS.n9189 DVSS.n9188 0.00053
R42406 DVSS.n9205 DVSS.n9204 0.00053
R42407 DVSS.n9253 DVSS.n9252 0.00053
R42408 DVSS.n9265 DVSS.n9260 0.00053
R42409 DVSS.n9305 DVSS.n9304 0.00053
R42410 DVSS.n9318 DVSS.n9313 0.00053
R42411 DVSS.n9341 DVSS.n9340 0.00053
R42412 DVSS.n9487 DVSS.n9486 0.00053
R42413 DVSS.n9473 DVSS.n9472 0.00053
R42414 DVSS.n9445 DVSS.n9431 0.00053
R42415 DVSS.n14132 DVSS.n14131 0.00053
R42416 DVSS.n14578 DVSS.n14577 0.00053
R42417 DVSS.n14574 DVSS.n14573 0.00053
R42418 DVSS.n13503 DVSS.n7893 0.00053
R42419 DVSS.n13494 DVSS.n13491 0.00053
R42420 DVSS.n13493 DVSS.n13492 0.00053
R42421 DVSS.n13420 DVSS.n7950 0.00053
R42422 DVSS.n7942 DVSS.n7937 0.00053
R42423 DVSS.n7941 DVSS.n7940 0.00053
R42424 DVSS.n11997 DVSS.n11996 0.00053
R42425 DVSS.n12125 DVSS.n11984 0.00053
R42426 DVSS.n12100 DVSS.n12099 0.00053
R42427 DVSS.n12095 DVSS.n12029 0.00053
R42428 DVSS.n19815 DVSS.n19814 0.00053
R42429 DVSS.n20096 DVSS.n20095 0.00053
R42430 DVSS.n20109 DVSS.n20107 0.00053
R42431 DVSS.n20373 DVSS.n20372 0.00053
R42432 DVSS.n20595 DVSS.n20593 0.00053
R42433 DVSS.n20654 DVSS.n20653 0.00053
R42434 DVSS.n20646 DVSS.n20641 0.00053
R42435 DVSS.n21567 DVSS.n21566 0.00053
R42436 DVSS.n21559 DVSS.n15 0.00053
R42437 DVSS.n256 DVSS.n255 0.00053
R42438 DVSS.n20689 DVSS.n20688 0.00053
R42439 DVSS.n20705 DVSS.n20702 0.00053
R42440 DVSS.n20704 DVSS.n20703 0.00053
R42441 DVSS.n20918 DVSS.n20917 0.00053
R42442 DVSS.n20934 DVSS.n20931 0.00053
R42443 DVSS.n20933 DVSS.n20932 0.00053
R42444 DVSS.n21272 DVSS.n21262 0.00053
R42445 DVSS.n21362 DVSS.n21361 0.00053
R42446 DVSS.n21391 DVSS.n21390 0.00053
R42447 DVSS.n20706 DVSS.n20697 0.00053
R42448 DVSS.n20935 DVSS.n20926 0.00053
R42449 DVSS.n21273 DVSS.n21260 0.00053
R42450 DVSS.n21389 DVSS.n21385 0.00053
R42451 DVSS.n20111 DVSS.n20103 0.00053
R42452 DVSS.n20597 DVSS.n20380 0.00053
R42453 DVSS.n20648 DVSS.n20637 0.00053
R42454 DVSS.n21561 DVSS.n14 0.00053
R42455 DVSS.n13496 DVSS.n13485 0.00053
R42456 DVSS.n7944 DVSS.n7931 0.00053
R42457 DVSS.n12124 DVSS.n11985 0.00053
R42458 DVSS.n12096 DVSS.n12027 0.00053
R42459 DVSS.n9448 DVSS 0.000526667
R42460 ASIG5V.n9783 ASIG5V 7.62481
R42461 ASIG5V.n10340 ASIG5V 7.62056
R42462 ASIG5V.n12966 ASIG5V 7.61152
R42463 ASIG5V.n13052 ASIG5V 7.60922
R42464 ASIG5V.n12999 ASIG5V 7.60798
R42465 ASIG5V.n1975 ASIG5V 7.60674
R42466 ASIG5V.n1434 ASIG5V 7.60674
R42467 ASIG5V.n2264 ASIG5V 7.60674
R42468 ASIG5V.n11486 ASIG5V.n8859 2.2505
R42469 ASIG5V.n11486 ASIG5V.n11423 2.2505
R42470 ASIG5V.n11486 ASIG5V.n8858 2.2505
R42471 ASIG5V.n11486 ASIG5V.n11424 2.2505
R42472 ASIG5V.n11486 ASIG5V.n8857 2.2505
R42473 ASIG5V.n11324 ASIG5V.n11320 2.24164
R42474 ASIG5V.n11324 ASIG5V.n8864 2.24164
R42475 ASIG5V.n11324 ASIG5V.n11321 2.24164
R42476 ASIG5V.n11324 ASIG5V.n8863 2.24164
R42477 ASIG5V.n11324 ASIG5V.n11322 2.24164
R42478 ASIG5V.n11324 ASIG5V.n8862 2.24164
R42479 ASIG5V.n8975 ASIG5V.n8883 1.49791
R42480 ASIG5V.n12862 ASIG5V.n12861 1.49652
R42481 ASIG5V.n12891 ASIG5V.n12890 1.49652
R42482 ASIG5V.n10033 ASIG5V.n9973 1.49652
R42483 ASIG5V.n10005 ASIG5V.n9978 1.49652
R42484 ASIG5V.n10061 ASIG5V.n10060 1.49652
R42485 ASIG5V.n13123 ASIG5V.n13121 1.49652
R42486 ASIG5V.n13192 ASIG5V.n7173 1.49652
R42487 ASIG5V.n13161 ASIG5V.n7175 1.49652
R42488 ASIG5V.n13130 ASIG5V.n7181 1.49652
R42489 ASIG5V.n13220 ASIG5V.n13219 1.49652
R42490 ASIG5V.n13253 ASIG5V.n13252 1.49652
R42491 ASIG5V.n13262 ASIG5V.n398 1.49652
R42492 ASIG5V.n12808 ASIG5V.n12807 1.49652
R42493 ASIG5V.n13046 ASIG5V.n13045 1.49652
R42494 ASIG5V.n13093 ASIG5V.n13051 1.49652
R42495 ASIG5V.n1574 ASIG5V.n1403 1.49652
R42496 ASIG5V.n1544 ASIG5V.n1412 1.49652
R42497 ASIG5V.n1514 ASIG5V.n1421 1.49652
R42498 ASIG5V.n1484 ASIG5V.n1426 1.49652
R42499 ASIG5V.n1602 ASIG5V.n1601 1.49652
R42500 ASIG5V.n1634 ASIG5V.n1385 1.49652
R42501 ASIG5V.n12779 ASIG5V.n12778 1.49652
R42502 ASIG5V.n1664 ASIG5V.n1376 1.49652
R42503 ASIG5V.n2163 ASIG5V.n1974 1.49652
R42504 ASIG5V.n7145 ASIG5V.n7144 1.49652
R42505 ASIG5V.n10453 ASIG5V.n10304 1.49652
R42506 ASIG5V.n10428 ASIG5V.n10313 1.49652
R42507 ASIG5V.n10403 ASIG5V.n10326 1.49652
R42508 ASIG5V.n10378 ASIG5V.n10339 1.49652
R42509 ASIG5V.n10485 ASIG5V.n10484 1.49652
R42510 ASIG5V.n10487 ASIG5V.n10295 1.49652
R42511 ASIG5V.n10516 ASIG5V.n10515 1.49652
R42512 ASIG5V.n12982 ASIG5V.n12981 1.49652
R42513 ASIG5V.n13014 ASIG5V.n12998 1.49652
R42514 ASIG5V.n1452 ASIG5V.n1433 1.49652
R42515 ASIG5V.n10070 ASIG5V.n10069 1.49652
R42516 ASIG5V.n9925 ASIG5V.n9758 1.49652
R42517 ASIG5V.n9897 ASIG5V.n9766 1.49652
R42518 ASIG5V.n9869 ASIG5V.n9774 1.49652
R42519 ASIG5V.n9841 ASIG5V.n9782 1.49652
R42520 ASIG5V.n10100 ASIG5V.n10099 1.49652
R42521 ASIG5V.n2378 ASIG5V.n2224 1.49652
R42522 ASIG5V.n2353 ASIG5V.n2233 1.49652
R42523 ASIG5V.n2328 ASIG5V.n2242 1.49652
R42524 ASIG5V.n2303 ASIG5V.n2252 1.49652
R42525 ASIG5V.n2428 ASIG5V.n2205 1.49652
R42526 ASIG5V.n2277 ASIG5V.n2263 1.49652
R42527 ASIG5V.n2453 ASIG5V.n2195 1.49652
R42528 ASIG5V.n10031 ASIG5V.n10030 1.49641
R42529 ASIG5V.n10003 ASIG5V.n10002 1.49641
R42530 ASIG5V.n10066 ASIG5V.n10063 1.49641
R42531 ASIG5V.n13119 ASIG5V.n13118 1.49641
R42532 ASIG5V.n13159 ASIG5V.n13158 1.49641
R42533 ASIG5V.n13190 ASIG5V.n13189 1.49641
R42534 ASIG5V.n13128 ASIG5V.n13127 1.49641
R42535 ASIG5V.n13222 ASIG5V.n7171 1.49641
R42536 ASIG5V.n13250 ASIG5V.n13249 1.49641
R42537 ASIG5V.n13260 ASIG5V.n13259 1.49641
R42538 ASIG5V.n13043 ASIG5V.n13042 1.49641
R42539 ASIG5V.n13091 ASIG5V.n13090 1.49641
R42540 ASIG5V.n1512 ASIG5V.n1511 1.49641
R42541 ASIG5V.n1542 ASIG5V.n1541 1.49641
R42542 ASIG5V.n1572 ASIG5V.n1571 1.49641
R42543 ASIG5V.n1632 ASIG5V.n1631 1.49641
R42544 ASIG5V.n1482 ASIG5V.n1481 1.49641
R42545 ASIG5V.n1604 ASIG5V.n1394 1.49641
R42546 ASIG5V.n1662 ASIG5V.n1661 1.49641
R42547 ASIG5V.n7147 ASIG5V.n404 1.49641
R42548 ASIG5V.n13289 ASIG5V.n13288 1.49641
R42549 ASIG5V.n13291 ASIG5V.n396 1.49641
R42550 ASIG5V.n12781 ASIG5V.n7209 1.49641
R42551 ASIG5V.n10549 ASIG5V.n10548 1.49641
R42552 ASIG5V.n10561 ASIG5V.n10560 1.49641
R42553 ASIG5V.n1450 ASIG5V.n1449 1.49641
R42554 ASIG5V.n12979 ASIG5V.n12978 1.49641
R42555 ASIG5V.n13012 ASIG5V.n13011 1.49641
R42556 ASIG5V.n10072 ASIG5V.n9750 1.49641
R42557 ASIG5V.n9923 ASIG5V.n9922 1.49641
R42558 ASIG5V.n9895 ASIG5V.n9894 1.49641
R42559 ASIG5V.n9867 ASIG5V.n9866 1.49641
R42560 ASIG5V.n9839 ASIG5V.n9838 1.49641
R42561 ASIG5V.n9808 ASIG5V.n9807 1.49641
R42562 ASIG5V.n9813 ASIG5V.n9812 1.49641
R42563 ASIG5V.n10102 ASIG5V.n9742 1.49641
R42564 ASIG5V.n2301 ASIG5V.n2300 1.49641
R42565 ASIG5V.n2403 ASIG5V.n2215 1.49641
R42566 ASIG5V.n3512 ASIG5V.n3511 1.1255
R42567 ASIG5V.n3663 ASIG5V.n3662 1.1255
R42568 ASIG5V.n3516 ASIG5V.n3515 1.1255
R42569 ASIG5V.n3987 ASIG5V.n3986 1.1255
R42570 ASIG5V.n3776 ASIG5V.n3775 1.1255
R42571 ASIG5V.n3983 ASIG5V.n3982 1.1255
R42572 ASIG5V.n3780 ASIG5V.n3779 1.1255
R42573 ASIG5V.n3927 ASIG5V.n3926 1.1255
R42574 ASIG5V.n3784 ASIG5V.n3783 1.1255
R42575 ASIG5V.n4038 ASIG5V.n4037 1.1255
R42576 ASIG5V.n4203 ASIG5V.n4202 1.1255
R42577 ASIG5V.n4042 ASIG5V.n4041 1.1255
R42578 ASIG5V.n4258 ASIG5V.n4257 1.1255
R42579 ASIG5V.n4046 ASIG5V.n4045 1.1255
R42580 ASIG5V.n4254 ASIG5V.n4253 1.1255
R42581 ASIG5V.n4050 ASIG5V.n4049 1.1255
R42582 ASIG5V.n4199 ASIG5V.n4198 1.1255
R42583 ASIG5V.n4054 ASIG5V.n4053 1.1255
R42584 ASIG5V.n4250 ASIG5V.n4249 1.1255
R42585 ASIG5V.n4559 ASIG5V.n4558 1.1255
R42586 ASIG5V.n4309 ASIG5V.n4308 1.1255
R42587 ASIG5V.n4487 ASIG5V.n4486 1.1255
R42588 ASIG5V.n4313 ASIG5V.n4312 1.1255
R42589 ASIG5V.n4483 ASIG5V.n4482 1.1255
R42590 ASIG5V.n4317 ASIG5V.n4316 1.1255
R42591 ASIG5V.n4541 ASIG5V.n4540 1.1255
R42592 ASIG5V.n4321 ASIG5V.n4320 1.1255
R42593 ASIG5V.n4537 ASIG5V.n4536 1.1255
R42594 ASIG5V.n4325 ASIG5V.n4324 1.1255
R42595 ASIG5V.n4479 ASIG5V.n4478 1.1255
R42596 ASIG5V.n4329 ASIG5V.n4328 1.1255
R42597 ASIG5V.n4533 ASIG5V.n4532 1.1255
R42598 ASIG5V.n4529 ASIG5V.n4528 1.1255
R42599 ASIG5V.n4526 ASIG5V.n4525 1.1255
R42600 ASIG5V.n4573 ASIG5V.n4572 1.1255
R42601 ASIG5V.n4584 ASIG5V.n4583 1.1255
R42602 ASIG5V.n4828 ASIG5V.n4827 1.1255
R42603 ASIG5V.n4588 ASIG5V.n4587 1.1255
R42604 ASIG5V.n4750 ASIG5V.n4749 1.1255
R42605 ASIG5V.n4746 ASIG5V.n4745 1.1255
R42606 ASIG5V.n4743 ASIG5V.n4742 1.1255
R42607 ASIG5V.n4824 ASIG5V.n4823 1.1255
R42608 ASIG5V.n4821 ASIG5V.n4820 1.1255
R42609 ASIG5V.n4817 ASIG5V.n4816 1.1255
R42610 ASIG5V.n4814 ASIG5V.n4813 1.1255
R42611 ASIG5V.n4595 ASIG5V.n4594 1.1255
R42612 ASIG5V.n4602 ASIG5V.n4601 1.1255
R42613 ASIG5V.n4599 ASIG5V.n4598 1.1255
R42614 ASIG5V.n4810 ASIG5V.n4809 1.1255
R42615 ASIG5V.n4806 ASIG5V.n4805 1.1255
R42616 ASIG5V.n4803 ASIG5V.n4802 1.1255
R42617 ASIG5V.n4607 ASIG5V.n4606 1.1255
R42618 ASIG5V.n4859 ASIG5V.n4858 1.1255
R42619 ASIG5V.n5043 ASIG5V.n5042 1.1255
R42620 ASIG5V.n4871 ASIG5V.n4870 1.1255
R42621 ASIG5V.n5130 ASIG5V.n5129 1.1255
R42622 ASIG5V.n5126 ASIG5V.n5125 1.1255
R42623 ASIG5V.n5123 ASIG5V.n5122 1.1255
R42624 ASIG5V.n5039 ASIG5V.n5038 1.1255
R42625 ASIG5V.n5036 ASIG5V.n5035 1.1255
R42626 ASIG5V.n5032 ASIG5V.n5031 1.1255
R42627 ASIG5V.n5029 ASIG5V.n5028 1.1255
R42628 ASIG5V.n5119 ASIG5V.n5118 1.1255
R42629 ASIG5V.n5116 ASIG5V.n5115 1.1255
R42630 ASIG5V.n5112 ASIG5V.n5111 1.1255
R42631 ASIG5V.n5109 ASIG5V.n5108 1.1255
R42632 ASIG5V.n5025 ASIG5V.n5024 1.1255
R42633 ASIG5V.n5022 ASIG5V.n5021 1.1255
R42634 ASIG5V.n5105 ASIG5V.n5104 1.1255
R42635 ASIG5V.n5102 ASIG5V.n5101 1.1255
R42636 ASIG5V.n5098 ASIG5V.n5097 1.1255
R42637 ASIG5V.n5095 ASIG5V.n5094 1.1255
R42638 ASIG5V.n5018 ASIG5V.n5017 1.1255
R42639 ASIG5V.n5015 ASIG5V.n5014 1.1255
R42640 ASIG5V.n5011 ASIG5V.n5010 1.1255
R42641 ASIG5V.n5440 ASIG5V.n5439 1.1255
R42642 ASIG5V.n5180 ASIG5V.n5179 1.1255
R42643 ASIG5V.n5177 ASIG5V.n5176 1.1255
R42644 ASIG5V.n5187 ASIG5V.n5186 1.1255
R42645 ASIG5V.n5184 ASIG5V.n5183 1.1255
R42646 ASIG5V.n5194 ASIG5V.n5193 1.1255
R42647 ASIG5V.n5191 ASIG5V.n5190 1.1255
R42648 ASIG5V.n5201 ASIG5V.n5200 1.1255
R42649 ASIG5V.n5198 ASIG5V.n5197 1.1255
R42650 ASIG5V.n5208 ASIG5V.n5207 1.1255
R42651 ASIG5V.n5205 ASIG5V.n5204 1.1255
R42652 ASIG5V.n5215 ASIG5V.n5214 1.1255
R42653 ASIG5V.n5212 ASIG5V.n5211 1.1255
R42654 ASIG5V.n5222 ASIG5V.n5221 1.1255
R42655 ASIG5V.n5219 ASIG5V.n5218 1.1255
R42656 ASIG5V.n5229 ASIG5V.n5228 1.1255
R42657 ASIG5V.n5226 ASIG5V.n5225 1.1255
R42658 ASIG5V.n5236 ASIG5V.n5235 1.1255
R42659 ASIG5V.n5233 ASIG5V.n5232 1.1255
R42660 ASIG5V.n5243 ASIG5V.n5242 1.1255
R42661 ASIG5V.n5240 ASIG5V.n5239 1.1255
R42662 ASIG5V.n5250 ASIG5V.n5249 1.1255
R42663 ASIG5V.n5247 ASIG5V.n5246 1.1255
R42664 ASIG5V.n5257 ASIG5V.n5256 1.1255
R42665 ASIG5V.n5254 ASIG5V.n5253 1.1255
R42666 ASIG5V.n5263 ASIG5V.n5262 1.1255
R42667 ASIG5V.n5457 ASIG5V.n5456 1.1255
R42668 ASIG5V.n5468 ASIG5V.n5467 1.1255
R42669 ASIG5V.n5465 ASIG5V.n5464 1.1255
R42670 ASIG5V.n5786 ASIG5V.n5785 1.1255
R42671 ASIG5V.n5472 ASIG5V.n5471 1.1255
R42672 ASIG5V.n5723 ASIG5V.n5722 1.1255
R42673 ASIG5V.n5476 ASIG5V.n5475 1.1255
R42674 ASIG5V.n5782 ASIG5V.n5781 1.1255
R42675 ASIG5V.n5480 ASIG5V.n5479 1.1255
R42676 ASIG5V.n5487 ASIG5V.n5486 1.1255
R42677 ASIG5V.n5484 ASIG5V.n5483 1.1255
R42678 ASIG5V.n5719 ASIG5V.n5718 1.1255
R42679 ASIG5V.n5491 ASIG5V.n5490 1.1255
R42680 ASIG5V.n5715 ASIG5V.n5714 1.1255
R42681 ASIG5V.n5777 ASIG5V.n5776 1.1255
R42682 ASIG5V.n5774 ASIG5V.n5773 1.1255
R42683 ASIG5V.n5770 ASIG5V.n5769 1.1255
R42684 ASIG5V.n5767 ASIG5V.n5766 1.1255
R42685 ASIG5V.n5497 ASIG5V.n5496 1.1255
R42686 ASIG5V.n5711 ASIG5V.n5710 1.1255
R42687 ASIG5V.n5501 ASIG5V.n5500 1.1255
R42688 ASIG5V.n5763 ASIG5V.n5762 1.1255
R42689 ASIG5V.n5505 ASIG5V.n5504 1.1255
R42690 ASIG5V.n5759 ASIG5V.n5758 1.1255
R42691 ASIG5V.n5509 ASIG5V.n5508 1.1255
R42692 ASIG5V.n5707 ASIG5V.n5706 1.1255
R42693 ASIG5V.n5513 ASIG5V.n5512 1.1255
R42694 ASIG5V.n5703 ASIG5V.n5702 1.1255
R42695 ASIG5V.n5517 ASIG5V.n5516 1.1255
R42696 ASIG5V.n6147 ASIG5V.n6146 1.1255
R42697 ASIG5V.n6055 ASIG5V.n6054 1.1255
R42698 ASIG5V.n6052 ASIG5V.n6051 1.1255
R42699 ASIG5V.n5813 ASIG5V.n5812 1.1255
R42700 ASIG5V.n5817 ASIG5V.n5816 1.1255
R42701 ASIG5V.n6140 ASIG5V.n6139 1.1255
R42702 ASIG5V.n6137 ASIG5V.n6136 1.1255
R42703 ASIG5V.n6048 ASIG5V.n6047 1.1255
R42704 ASIG5V.n6045 ASIG5V.n6044 1.1255
R42705 ASIG5V.n5822 ASIG5V.n5821 1.1255
R42706 ASIG5V.n5826 ASIG5V.n5825 1.1255
R42707 ASIG5V.n6132 ASIG5V.n6131 1.1255
R42708 ASIG5V.n6129 ASIG5V.n6128 1.1255
R42709 ASIG5V.n6041 ASIG5V.n6040 1.1255
R42710 ASIG5V.n6038 ASIG5V.n6037 1.1255
R42711 ASIG5V.n6034 ASIG5V.n6033 1.1255
R42712 ASIG5V.n6031 ASIG5V.n6030 1.1255
R42713 ASIG5V.n6125 ASIG5V.n6124 1.1255
R42714 ASIG5V.n6122 ASIG5V.n6121 1.1255
R42715 ASIG5V.n6118 ASIG5V.n6117 1.1255
R42716 ASIG5V.n6115 ASIG5V.n6114 1.1255
R42717 ASIG5V.n6027 ASIG5V.n6026 1.1255
R42718 ASIG5V.n6024 ASIG5V.n6023 1.1255
R42719 ASIG5V.n6111 ASIG5V.n6110 1.1255
R42720 ASIG5V.n6108 ASIG5V.n6107 1.1255
R42721 ASIG5V.n6104 ASIG5V.n6103 1.1255
R42722 ASIG5V.n6101 ASIG5V.n6100 1.1255
R42723 ASIG5V.n6020 ASIG5V.n6019 1.1255
R42724 ASIG5V.n6017 ASIG5V.n6016 1.1255
R42725 ASIG5V.n6013 ASIG5V.n6012 1.1255
R42726 ASIG5V.n6010 ASIG5V.n6009 1.1255
R42727 ASIG5V.n6097 ASIG5V.n6096 1.1255
R42728 ASIG5V.n6165 ASIG5V.n6164 1.1255
R42729 ASIG5V.n6168 ASIG5V.n6167 1.1255
R42730 ASIG5V.n7094 ASIG5V.n7093 1.1255
R42731 ASIG5V.n6172 ASIG5V.n6171 1.1255
R42732 ASIG5V.n7090 ASIG5V.n7089 1.1255
R42733 ASIG5V.n6176 ASIG5V.n6175 1.1255
R42734 ASIG5V.n6183 ASIG5V.n6182 1.1255
R42735 ASIG5V.n6180 ASIG5V.n6179 1.1255
R42736 ASIG5V.n6187 ASIG5V.n6186 1.1255
R42737 ASIG5V.n7086 ASIG5V.n7085 1.1255
R42738 ASIG5V.n7083 ASIG5V.n7082 1.1255
R42739 ASIG5V.n6191 ASIG5V.n6190 1.1255
R42740 ASIG5V.n7115 ASIG5V.n7114 1.1255
R42741 ASIG5V.n6195 ASIG5V.n6194 1.1255
R42742 ASIG5V.n7111 ASIG5V.n7110 1.1255
R42743 ASIG5V.n7079 ASIG5V.n7078 1.1255
R42744 ASIG5V.n6203 ASIG5V.n6202 1.1255
R42745 ASIG5V.n6200 ASIG5V.n6199 1.1255
R42746 ASIG5V.n6210 ASIG5V.n6209 1.1255
R42747 ASIG5V.n6207 ASIG5V.n6206 1.1255
R42748 ASIG5V.n6217 ASIG5V.n6216 1.1255
R42749 ASIG5V.n6214 ASIG5V.n6213 1.1255
R42750 ASIG5V.n6224 ASIG5V.n6223 1.1255
R42751 ASIG5V.n6221 ASIG5V.n6220 1.1255
R42752 ASIG5V.n6231 ASIG5V.n6230 1.1255
R42753 ASIG5V.n6228 ASIG5V.n6227 1.1255
R42754 ASIG5V.n6238 ASIG5V.n6237 1.1255
R42755 ASIG5V.n6235 ASIG5V.n6234 1.1255
R42756 ASIG5V.n6245 ASIG5V.n6244 1.1255
R42757 ASIG5V.n6242 ASIG5V.n6241 1.1255
R42758 ASIG5V.n6252 ASIG5V.n6251 1.1255
R42759 ASIG5V.n6249 ASIG5V.n6248 1.1255
R42760 ASIG5V.n6259 ASIG5V.n6258 1.1255
R42761 ASIG5V.n6256 ASIG5V.n6255 1.1255
R42762 ASIG5V.n6420 ASIG5V.n6419 1.1255
R42763 ASIG5V.n6926 ASIG5V.n6925 1.1255
R42764 ASIG5V.n6925 ASIG5V.n6924 1.1255
R42765 ASIG5V.n6922 ASIG5V.n6921 1.1255
R42766 ASIG5V.n6340 ASIG5V.n6339 1.1255
R42767 ASIG5V.n6826 ASIG5V.n6825 1.1255
R42768 ASIG5V.n6344 ASIG5V.n6343 1.1255
R42769 ASIG5V.n6822 ASIG5V.n6821 1.1255
R42770 ASIG5V.n6918 ASIG5V.n6917 1.1255
R42771 ASIG5V.n6915 ASIG5V.n6914 1.1255
R42772 ASIG5V.n6911 ASIG5V.n6910 1.1255
R42773 ASIG5V.n6908 ASIG5V.n6907 1.1255
R42774 ASIG5V.n6350 ASIG5V.n6349 1.1255
R42775 ASIG5V.n6354 ASIG5V.n6353 1.1255
R42776 ASIG5V.n6904 ASIG5V.n6903 1.1255
R42777 ASIG5V.n6901 ASIG5V.n6900 1.1255
R42778 ASIG5V.n6897 ASIG5V.n6896 1.1255
R42779 ASIG5V.n6894 ASIG5V.n6893 1.1255
R42780 ASIG5V.n6359 ASIG5V.n6358 1.1255
R42781 ASIG5V.n6366 ASIG5V.n6365 1.1255
R42782 ASIG5V.n6363 ASIG5V.n6362 1.1255
R42783 ASIG5V.n6816 ASIG5V.n6815 1.1255
R42784 ASIG5V.n6890 ASIG5V.n6889 1.1255
R42785 ASIG5V.n6887 ASIG5V.n6886 1.1255
R42786 ASIG5V.n6883 ASIG5V.n6882 1.1255
R42787 ASIG5V.n6880 ASIG5V.n6879 1.1255
R42788 ASIG5V.n6372 ASIG5V.n6371 1.1255
R42789 ASIG5V.n6812 ASIG5V.n6811 1.1255
R42790 ASIG5V.n6876 ASIG5V.n6875 1.1255
R42791 ASIG5V.n6873 ASIG5V.n6872 1.1255
R42792 ASIG5V.n6869 ASIG5V.n6868 1.1255
R42793 ASIG5V.n6866 ASIG5V.n6865 1.1255
R42794 ASIG5V.n6378 ASIG5V.n6377 1.1255
R42795 ASIG5V.n6808 ASIG5V.n6807 1.1255
R42796 ASIG5V.n6382 ASIG5V.n6381 1.1255
R42797 ASIG5V.n6804 ASIG5V.n6803 1.1255
R42798 ASIG5V.n6427 ASIG5V.n6426 1.1255
R42799 ASIG5V.n6425 ASIG5V.n6424 1.1255
R42800 ASIG5V.n6424 ASIG5V.n6423 1.1255
R42801 ASIG5V.n6431 ASIG5V.n6430 1.1255
R42802 ASIG5V.n6613 ASIG5V.n6612 1.1255
R42803 ASIG5V.n6435 ASIG5V.n6434 1.1255
R42804 ASIG5V.n6609 ASIG5V.n6608 1.1255
R42805 ASIG5V.n6606 ASIG5V.n6605 1.1255
R42806 ASIG5V.n6439 ASIG5V.n6438 1.1255
R42807 ASIG5V.n6446 ASIG5V.n6445 1.1255
R42808 ASIG5V.n6443 ASIG5V.n6442 1.1255
R42809 ASIG5V.n6450 ASIG5V.n6449 1.1255
R42810 ASIG5V.n6602 ASIG5V.n6601 1.1255
R42811 ASIG5V.n6599 ASIG5V.n6598 1.1255
R42812 ASIG5V.n6454 ASIG5V.n6453 1.1255
R42813 ASIG5V.n6461 ASIG5V.n6460 1.1255
R42814 ASIG5V.n6458 ASIG5V.n6457 1.1255
R42815 ASIG5V.n6465 ASIG5V.n6464 1.1255
R42816 ASIG5V.n6595 ASIG5V.n6594 1.1255
R42817 ASIG5V.n6592 ASIG5V.n6591 1.1255
R42818 ASIG5V.n6588 ASIG5V.n6587 1.1255
R42819 ASIG5V.n6585 ASIG5V.n6584 1.1255
R42820 ASIG5V.n6470 ASIG5V.n6469 1.1255
R42821 ASIG5V.n6477 ASIG5V.n6476 1.1255
R42822 ASIG5V.n6474 ASIG5V.n6473 1.1255
R42823 ASIG5V.n6643 ASIG5V.n6642 1.1255
R42824 ASIG5V.n6581 ASIG5V.n6580 1.1255
R42825 ASIG5V.n6578 ASIG5V.n6577 1.1255
R42826 ASIG5V.n6482 ASIG5V.n6481 1.1255
R42827 ASIG5V.n6489 ASIG5V.n6488 1.1255
R42828 ASIG5V.n6486 ASIG5V.n6485 1.1255
R42829 ASIG5V.n6496 ASIG5V.n6495 1.1255
R42830 ASIG5V.n6493 ASIG5V.n6492 1.1255
R42831 ASIG5V.n6574 ASIG5V.n6573 1.1255
R42832 ASIG5V.n6500 ASIG5V.n6499 1.1255
R42833 ASIG5V.n6570 ASIG5V.n6569 1.1255
R42834 ASIG5V.n6504 ASIG5V.n6503 1.1255
R42835 ASIG5V.n6771 ASIG5V.n6770 1.1255
R42836 ASIG5V.n6774 ASIG5V.n6773 1.1255
R42837 ASIG5V.n5 ASIG5V.n4 1.1255
R42838 ASIG5V.n13493 ASIG5V.n13492 1.1255
R42839 ASIG5V.n13492 ASIG5V.n13491 1.1255
R42840 ASIG5V.n13489 ASIG5V.n13488 1.1255
R42841 ASIG5V.n9 ASIG5V.n8 1.1255
R42842 ASIG5V.n13406 ASIG5V.n13405 1.1255
R42843 ASIG5V.n13 ASIG5V.n12 1.1255
R42844 ASIG5V.n17 ASIG5V.n16 1.1255
R42845 ASIG5V.n13485 ASIG5V.n13484 1.1255
R42846 ASIG5V.n13482 ASIG5V.n13481 1.1255
R42847 ASIG5V.n13478 ASIG5V.n13477 1.1255
R42848 ASIG5V.n13475 ASIG5V.n13474 1.1255
R42849 ASIG5V.n22 ASIG5V.n21 1.1255
R42850 ASIG5V.n26 ASIG5V.n25 1.1255
R42851 ASIG5V.n13471 ASIG5V.n13470 1.1255
R42852 ASIG5V.n13468 ASIG5V.n13467 1.1255
R42853 ASIG5V.n13464 ASIG5V.n13463 1.1255
R42854 ASIG5V.n13461 ASIG5V.n13460 1.1255
R42855 ASIG5V.n31 ASIG5V.n30 1.1255
R42856 ASIG5V.n13400 ASIG5V.n13399 1.1255
R42857 ASIG5V.n13396 ASIG5V.n13395 1.1255
R42858 ASIG5V.n13393 ASIG5V.n13392 1.1255
R42859 ASIG5V.n13457 ASIG5V.n13456 1.1255
R42860 ASIG5V.n13454 ASIG5V.n13453 1.1255
R42861 ASIG5V.n13450 ASIG5V.n13449 1.1255
R42862 ASIG5V.n13447 ASIG5V.n13446 1.1255
R42863 ASIG5V.n38 ASIG5V.n37 1.1255
R42864 ASIG5V.n42 ASIG5V.n41 1.1255
R42865 ASIG5V.n13443 ASIG5V.n13442 1.1255
R42866 ASIG5V.n13440 ASIG5V.n13439 1.1255
R42867 ASIG5V.n13436 ASIG5V.n13435 1.1255
R42868 ASIG5V.n13433 ASIG5V.n13432 1.1255
R42869 ASIG5V.n47 ASIG5V.n46 1.1255
R42870 ASIG5V.n13388 ASIG5V.n13387 1.1255
R42871 ASIG5V.n51 ASIG5V.n50 1.1255
R42872 ASIG5V.n55 ASIG5V.n54 1.1255
R42873 ASIG5V.n13429 ASIG5V.n13428 1.1255
R42874 ASIG5V.n329 ASIG5V.n328 1.1255
R42875 ASIG5V.n326 ASIG5V.n325 1.1255
R42876 ASIG5V.n229 ASIG5V.n228 1.1255
R42877 ASIG5V.n226 ASIG5V.n225 1.1255
R42878 ASIG5V.n222 ASIG5V.n221 1.1255
R42879 ASIG5V.n219 ASIG5V.n218 1.1255
R42880 ASIG5V.n322 ASIG5V.n321 1.1255
R42881 ASIG5V.n319 ASIG5V.n318 1.1255
R42882 ASIG5V.n315 ASIG5V.n314 1.1255
R42883 ASIG5V.n312 ASIG5V.n311 1.1255
R42884 ASIG5V.n215 ASIG5V.n214 1.1255
R42885 ASIG5V.n212 ASIG5V.n211 1.1255
R42886 ASIG5V.n308 ASIG5V.n307 1.1255
R42887 ASIG5V.n305 ASIG5V.n304 1.1255
R42888 ASIG5V.n301 ASIG5V.n300 1.1255
R42889 ASIG5V.n298 ASIG5V.n297 1.1255
R42890 ASIG5V.n208 ASIG5V.n207 1.1255
R42891 ASIG5V.n205 ASIG5V.n204 1.1255
R42892 ASIG5V.n201 ASIG5V.n200 1.1255
R42893 ASIG5V.n198 ASIG5V.n197 1.1255
R42894 ASIG5V.n294 ASIG5V.n293 1.1255
R42895 ASIG5V.n291 ASIG5V.n290 1.1255
R42896 ASIG5V.n287 ASIG5V.n286 1.1255
R42897 ASIG5V.n284 ASIG5V.n283 1.1255
R42898 ASIG5V.n194 ASIG5V.n193 1.1255
R42899 ASIG5V.n191 ASIG5V.n190 1.1255
R42900 ASIG5V.n280 ASIG5V.n279 1.1255
R42901 ASIG5V.n277 ASIG5V.n276 1.1255
R42902 ASIG5V.n273 ASIG5V.n272 1.1255
R42903 ASIG5V.n270 ASIG5V.n269 1.1255
R42904 ASIG5V.n187 ASIG5V.n186 1.1255
R42905 ASIG5V.n184 ASIG5V.n183 1.1255
R42906 ASIG5V.n180 ASIG5V.n179 1.1255
R42907 ASIG5V.n177 ASIG5V.n176 1.1255
R42908 ASIG5V.n266 ASIG5V.n265 1.1255
R42909 ASIG5V.n7287 ASIG5V.n7286 1.1255
R42910 ASIG5V.n7293 ASIG5V.n7292 1.1255
R42911 ASIG5V.n7559 ASIG5V.n7558 1.1255
R42912 ASIG5V.n7297 ASIG5V.n7296 1.1255
R42913 ASIG5V.n7304 ASIG5V.n7303 1.1255
R42914 ASIG5V.n7301 ASIG5V.n7300 1.1255
R42915 ASIG5V.n7619 ASIG5V.n7618 1.1255
R42916 ASIG5V.n7308 ASIG5V.n7307 1.1255
R42917 ASIG5V.n7555 ASIG5V.n7554 1.1255
R42918 ASIG5V.n7312 ASIG5V.n7311 1.1255
R42919 ASIG5V.n7615 ASIG5V.n7614 1.1255
R42920 ASIG5V.n7316 ASIG5V.n7315 1.1255
R42921 ASIG5V.n7611 ASIG5V.n7610 1.1255
R42922 ASIG5V.n7320 ASIG5V.n7319 1.1255
R42923 ASIG5V.n7551 ASIG5V.n7550 1.1255
R42924 ASIG5V.n7324 ASIG5V.n7323 1.1255
R42925 ASIG5V.n7331 ASIG5V.n7330 1.1255
R42926 ASIG5V.n7328 ASIG5V.n7327 1.1255
R42927 ASIG5V.n7607 ASIG5V.n7606 1.1255
R42928 ASIG5V.n7335 ASIG5V.n7334 1.1255
R42929 ASIG5V.n7603 ASIG5V.n7602 1.1255
R42930 ASIG5V.n7339 ASIG5V.n7338 1.1255
R42931 ASIG5V.n7343 ASIG5V.n7342 1.1255
R42932 ASIG5V.n7599 ASIG5V.n7598 1.1255
R42933 ASIG5V.n7596 ASIG5V.n7595 1.1255
R42934 ASIG5V.n7347 ASIG5V.n7346 1.1255
R42935 ASIG5V.n7592 ASIG5V.n7591 1.1255
R42936 ASIG5V.n7351 ASIG5V.n7350 1.1255
R42937 ASIG5V.n7545 ASIG5V.n7544 1.1255
R42938 ASIG5V.n7355 ASIG5V.n7354 1.1255
R42939 ASIG5V.n7541 ASIG5V.n7540 1.1255
R42940 ASIG5V.n7642 ASIG5V.n7641 1.1255
R42941 ASIG5V.n7657 ASIG5V.n7656 1.1255
R42942 ASIG5V.n7666 ASIG5V.n7665 1.1255
R42943 ASIG5V.n7663 ASIG5V.n7662 1.1255
R42944 ASIG5V.n7673 ASIG5V.n7672 1.1255
R42945 ASIG5V.n7670 ASIG5V.n7669 1.1255
R42946 ASIG5V.n7680 ASIG5V.n7679 1.1255
R42947 ASIG5V.n7677 ASIG5V.n7676 1.1255
R42948 ASIG5V.n7687 ASIG5V.n7686 1.1255
R42949 ASIG5V.n7684 ASIG5V.n7683 1.1255
R42950 ASIG5V.n7694 ASIG5V.n7693 1.1255
R42951 ASIG5V.n7691 ASIG5V.n7690 1.1255
R42952 ASIG5V.n7701 ASIG5V.n7700 1.1255
R42953 ASIG5V.n7698 ASIG5V.n7697 1.1255
R42954 ASIG5V.n7708 ASIG5V.n7707 1.1255
R42955 ASIG5V.n7705 ASIG5V.n7704 1.1255
R42956 ASIG5V.n7715 ASIG5V.n7714 1.1255
R42957 ASIG5V.n7712 ASIG5V.n7711 1.1255
R42958 ASIG5V.n7722 ASIG5V.n7721 1.1255
R42959 ASIG5V.n7719 ASIG5V.n7718 1.1255
R42960 ASIG5V.n7729 ASIG5V.n7728 1.1255
R42961 ASIG5V.n7726 ASIG5V.n7725 1.1255
R42962 ASIG5V.n7736 ASIG5V.n7735 1.1255
R42963 ASIG5V.n7733 ASIG5V.n7732 1.1255
R42964 ASIG5V.n7743 ASIG5V.n7742 1.1255
R42965 ASIG5V.n7740 ASIG5V.n7739 1.1255
R42966 ASIG5V.n7750 ASIG5V.n7749 1.1255
R42967 ASIG5V.n7747 ASIG5V.n7746 1.1255
R42968 ASIG5V.n7756 ASIG5V.n7755 1.1255
R42969 ASIG5V.n7995 ASIG5V.n7994 1.1255
R42970 ASIG5V.n8011 ASIG5V.n8010 1.1255
R42971 ASIG5V.n12743 ASIG5V.n12742 1.1255
R42972 ASIG5V.n8015 ASIG5V.n8014 1.1255
R42973 ASIG5V.n8022 ASIG5V.n8021 1.1255
R42974 ASIG5V.n8019 ASIG5V.n8018 1.1255
R42975 ASIG5V.n12739 ASIG5V.n12738 1.1255
R42976 ASIG5V.n8026 ASIG5V.n8025 1.1255
R42977 ASIG5V.n12735 ASIG5V.n12734 1.1255
R42978 ASIG5V.n8030 ASIG5V.n8029 1.1255
R42979 ASIG5V.n8037 ASIG5V.n8036 1.1255
R42980 ASIG5V.n8034 ASIG5V.n8033 1.1255
R42981 ASIG5V.n8044 ASIG5V.n8043 1.1255
R42982 ASIG5V.n8041 ASIG5V.n8040 1.1255
R42983 ASIG5V.n12731 ASIG5V.n12730 1.1255
R42984 ASIG5V.n8048 ASIG5V.n8047 1.1255
R42985 ASIG5V.n12727 ASIG5V.n12726 1.1255
R42986 ASIG5V.n8052 ASIG5V.n8051 1.1255
R42987 ASIG5V.n12696 ASIG5V.n12695 1.1255
R42988 ASIG5V.n8056 ASIG5V.n8055 1.1255
R42989 ASIG5V.n8063 ASIG5V.n8062 1.1255
R42990 ASIG5V.n8060 ASIG5V.n8059 1.1255
R42991 ASIG5V.n8070 ASIG5V.n8069 1.1255
R42992 ASIG5V.n8067 ASIG5V.n8066 1.1255
R42993 ASIG5V.n12692 ASIG5V.n12691 1.1255
R42994 ASIG5V.n8074 ASIG5V.n8073 1.1255
R42995 ASIG5V.n12688 ASIG5V.n12687 1.1255
R42996 ASIG5V.n12579 ASIG5V.n12578 1.1255
R42997 ASIG5V.n12473 ASIG5V.n12472 1.1255
R42998 ASIG5V.n12563 ASIG5V.n12562 1.1255
R42999 ASIG5V.n12560 ASIG5V.n12559 1.1255
R43000 ASIG5V.n12556 ASIG5V.n12555 1.1255
R43001 ASIG5V.n12553 ASIG5V.n12552 1.1255
R43002 ASIG5V.n8138 ASIG5V.n8137 1.1255
R43003 ASIG5V.n12469 ASIG5V.n12468 1.1255
R43004 ASIG5V.n8142 ASIG5V.n8141 1.1255
R43005 ASIG5V.n8146 ASIG5V.n8145 1.1255
R43006 ASIG5V.n12549 ASIG5V.n12548 1.1255
R43007 ASIG5V.n12546 ASIG5V.n12545 1.1255
R43008 ASIG5V.n12542 ASIG5V.n12541 1.1255
R43009 ASIG5V.n12539 ASIG5V.n12538 1.1255
R43010 ASIG5V.n8151 ASIG5V.n8150 1.1255
R43011 ASIG5V.n12464 ASIG5V.n12463 1.1255
R43012 ASIG5V.n12535 ASIG5V.n12534 1.1255
R43013 ASIG5V.n12532 ASIG5V.n12531 1.1255
R43014 ASIG5V.n12528 ASIG5V.n12527 1.1255
R43015 ASIG5V.n12525 ASIG5V.n12524 1.1255
R43016 ASIG5V.n8157 ASIG5V.n8156 1.1255
R43017 ASIG5V.n12460 ASIG5V.n12459 1.1255
R43018 ASIG5V.n12456 ASIG5V.n12455 1.1255
R43019 ASIG5V.n8197 ASIG5V.n8196 1.1255
R43020 ASIG5V.n8235 ASIG5V.n8234 1.1255
R43021 ASIG5V.n8232 ASIG5V.n8231 1.1255
R43022 ASIG5V.n8242 ASIG5V.n8241 1.1255
R43023 ASIG5V.n8239 ASIG5V.n8238 1.1255
R43024 ASIG5V.n8249 ASIG5V.n8248 1.1255
R43025 ASIG5V.n8246 ASIG5V.n8245 1.1255
R43026 ASIG5V.n8256 ASIG5V.n8255 1.1255
R43027 ASIG5V.n8253 ASIG5V.n8252 1.1255
R43028 ASIG5V.n8263 ASIG5V.n8262 1.1255
R43029 ASIG5V.n8260 ASIG5V.n8259 1.1255
R43030 ASIG5V.n8270 ASIG5V.n8269 1.1255
R43031 ASIG5V.n8267 ASIG5V.n8266 1.1255
R43032 ASIG5V.n8277 ASIG5V.n8276 1.1255
R43033 ASIG5V.n8274 ASIG5V.n8273 1.1255
R43034 ASIG5V.n8284 ASIG5V.n8283 1.1255
R43035 ASIG5V.n8281 ASIG5V.n8280 1.1255
R43036 ASIG5V.n8291 ASIG5V.n8290 1.1255
R43037 ASIG5V.n8288 ASIG5V.n8287 1.1255
R43038 ASIG5V.n8297 ASIG5V.n8296 1.1255
R43039 ASIG5V.n8368 ASIG5V.n8367 1.1255
R43040 ASIG5V.n12225 ASIG5V.n12224 1.1255
R43041 ASIG5V.n8399 ASIG5V.n8398 1.1255
R43042 ASIG5V.n8406 ASIG5V.n8405 1.1255
R43043 ASIG5V.n8403 ASIG5V.n8402 1.1255
R43044 ASIG5V.n12185 ASIG5V.n12184 1.1255
R43045 ASIG5V.n8410 ASIG5V.n8409 1.1255
R43046 ASIG5V.n12221 ASIG5V.n12220 1.1255
R43047 ASIG5V.n8414 ASIG5V.n8413 1.1255
R43048 ASIG5V.n12217 ASIG5V.n12216 1.1255
R43049 ASIG5V.n8418 ASIG5V.n8417 1.1255
R43050 ASIG5V.n8425 ASIG5V.n8424 1.1255
R43051 ASIG5V.n8422 ASIG5V.n8421 1.1255
R43052 ASIG5V.n8432 ASIG5V.n8431 1.1255
R43053 ASIG5V.n8429 ASIG5V.n8428 1.1255
R43054 ASIG5V.n12212 ASIG5V.n12211 1.1255
R43055 ASIG5V.n8527 ASIG5V.n8526 1.1255
R43056 ASIG5V.n8534 ASIG5V.n8533 1.1255
R43057 ASIG5V.n8531 ASIG5V.n8530 1.1255
R43058 ASIG5V.n12070 ASIG5V.n12069 1.1255
R43059 ASIG5V.n8538 ASIG5V.n8537 1.1255
R43060 ASIG5V.n12066 ASIG5V.n12065 1.1255
R43061 ASIG5V.n8542 ASIG5V.n8541 1.1255
R43062 ASIG5V.n8549 ASIG5V.n8548 1.1255
R43063 ASIG5V.n8546 ASIG5V.n8545 1.1255
R43064 ASIG5V.n12062 ASIG5V.n12061 1.1255
R43065 ASIG5V.n8553 ASIG5V.n8552 1.1255
R43066 ASIG5V.n8642 ASIG5V.n8641 1.1255
R43067 ASIG5V.n11907 ASIG5V.n11906 1.1255
R43068 ASIG5V.n8646 ASIG5V.n8645 1.1255
R43069 ASIG5V.n11903 ASIG5V.n11902 1.1255
R43070 ASIG5V.n8650 ASIG5V.n8649 1.1255
R43071 ASIG5V.n11863 ASIG5V.n11862 1.1255
R43072 ASIG5V.n8654 ASIG5V.n8653 1.1255
R43073 ASIG5V.n11740 ASIG5V.n11739 1.1255
R43074 ASIG5V.n8754 ASIG5V.n8753 1.1255
R43075 ASIG5V.n11697 ASIG5V.n11696 1.1255
R43076 ASIG5V.n3088 ASIG5V.n3087 1.1255
R43077 ASIG5V.n3159 ASIG5V.n3158 1.1255
R43078 ASIG5V.n3161 ASIG5V.n3160 1.1255
R43079 ASIG5V.n3208 ASIG5V.n3207 1.1255
R43080 ASIG5V.n3084 ASIG5V.n3083 1.1255
R43081 ASIG5V.n3211 ASIG5V.n3210 1.1255
R43082 ASIG5V.n3213 ASIG5V.n3212 1.1255
R43083 ASIG5V.n3164 ASIG5V.n3163 1.1255
R43084 ASIG5V.n3166 ASIG5V.n3165 1.1255
R43085 ASIG5V.n3216 ASIG5V.n3215 1.1255
R43086 ASIG5V.n3218 ASIG5V.n3217 1.1255
R43087 ASIG5V.n3221 ASIG5V.n3220 1.1255
R43088 ASIG5V.n3078 ASIG5V.n3077 1.1255
R43089 ASIG5V.n3169 ASIG5V.n3168 1.1255
R43090 ASIG5V.n3075 ASIG5V.n3074 1.1255
R43091 ASIG5V.n3172 ASIG5V.n3171 1.1255
R43092 ASIG5V.n3174 ASIG5V.n3173 1.1255
R43093 ASIG5V.n3224 ASIG5V.n3223 1.1255
R43094 ASIG5V.n3071 ASIG5V.n3070 1.1255
R43095 ASIG5V.n3227 ASIG5V.n3226 1.1255
R43096 ASIG5V.n3068 ASIG5V.n3067 1.1255
R43097 ASIG5V.n3177 ASIG5V.n3176 1.1255
R43098 ASIG5V.n3065 ASIG5V.n3064 1.1255
R43099 ASIG5V.n3230 ASIG5V.n3229 1.1255
R43100 ASIG5V.n3062 ASIG5V.n3061 1.1255
R43101 ASIG5V.n3233 ASIG5V.n3232 1.1255
R43102 ASIG5V.n3235 ASIG5V.n3234 1.1255
R43103 ASIG5V.n3180 ASIG5V.n3179 1.1255
R43104 ASIG5V.n3058 ASIG5V.n3057 1.1255
R43105 ASIG5V.n3183 ASIG5V.n3182 1.1255
R43106 ASIG5V.n3185 ASIG5V.n3184 1.1255
R43107 ASIG5V.n3238 ASIG5V.n3237 1.1255
R43108 ASIG5V.n3054 ASIG5V.n3053 1.1255
R43109 ASIG5V.n3241 ASIG5V.n3240 1.1255
R43110 ASIG5V.n3243 ASIG5V.n3242 1.1255
R43111 ASIG5V.n3188 ASIG5V.n3187 1.1255
R43112 ASIG5V.n3350 ASIG5V.n3349 1.1255
R43113 ASIG5V.n3352 ASIG5V.n3351 1.1255
R43114 ASIG5V.n3355 ASIG5V.n3354 1.1255
R43115 ASIG5V.n3357 ASIG5V.n3356 1.1255
R43116 ASIG5V.n3416 ASIG5V.n3415 1.1255
R43117 ASIG5V.n3418 ASIG5V.n3417 1.1255
R43118 ASIG5V.n3421 ASIG5V.n3420 1.1255
R43119 ASIG5V.n3423 ASIG5V.n3422 1.1255
R43120 ASIG5V.n3360 ASIG5V.n3359 1.1255
R43121 ASIG5V.n3362 ASIG5V.n3361 1.1255
R43122 ASIG5V.n3426 ASIG5V.n3425 1.1255
R43123 ASIG5V.n3428 ASIG5V.n3427 1.1255
R43124 ASIG5V.n3431 ASIG5V.n3430 1.1255
R43125 ASIG5V.n3433 ASIG5V.n3432 1.1255
R43126 ASIG5V.n3365 ASIG5V.n3364 1.1255
R43127 ASIG5V.n3367 ASIG5V.n3366 1.1255
R43128 ASIG5V.n3370 ASIG5V.n3369 1.1255
R43129 ASIG5V.n3372 ASIG5V.n3371 1.1255
R43130 ASIG5V.n3436 ASIG5V.n3435 1.1255
R43131 ASIG5V.n3438 ASIG5V.n3437 1.1255
R43132 ASIG5V.n3441 ASIG5V.n3440 1.1255
R43133 ASIG5V.n3443 ASIG5V.n3442 1.1255
R43134 ASIG5V.n3375 ASIG5V.n3374 1.1255
R43135 ASIG5V.n3377 ASIG5V.n3376 1.1255
R43136 ASIG5V.n3446 ASIG5V.n3445 1.1255
R43137 ASIG5V.n3448 ASIG5V.n3447 1.1255
R43138 ASIG5V.n3451 ASIG5V.n3450 1.1255
R43139 ASIG5V.n3453 ASIG5V.n3452 1.1255
R43140 ASIG5V.n3380 ASIG5V.n3379 1.1255
R43141 ASIG5V.n3382 ASIG5V.n3381 1.1255
R43142 ASIG5V.n3385 ASIG5V.n3384 1.1255
R43143 ASIG5V.n3387 ASIG5V.n3386 1.1255
R43144 ASIG5V.n3456 ASIG5V.n3455 1.1255
R43145 ASIG5V.n3458 ASIG5V.n3457 1.1255
R43146 ASIG5V.n3461 ASIG5V.n3460 1.1255
R43147 ASIG5V.n3463 ASIG5V.n3462 1.1255
R43148 ASIG5V.n3390 ASIG5V.n3389 1.1255
R43149 ASIG5V.n3392 ASIG5V.n3391 1.1255
R43150 ASIG5V.n3466 ASIG5V.n3465 1.1255
R43151 ASIG5V.n3468 ASIG5V.n3467 1.1255
R43152 ASIG5V.n3689 ASIG5V.n3688 1.1255
R43153 ASIG5V.n3640 ASIG5V.n3639 1.1255
R43154 ASIG5V.n3642 ASIG5V.n3641 1.1255
R43155 ASIG5V.n3645 ASIG5V.n3644 1.1255
R43156 ASIG5V.n3647 ASIG5V.n3646 1.1255
R43157 ASIG5V.n3692 ASIG5V.n3691 1.1255
R43158 ASIG5V.n3533 ASIG5V.n3532 1.1255
R43159 ASIG5V.n3535 ASIG5V.n3534 1.1255
R43160 ASIG5V.n3695 ASIG5V.n3694 1.1255
R43161 ASIG5V.n3530 ASIG5V.n3529 1.1255
R43162 ASIG5V.n3650 ASIG5V.n3649 1.1255
R43163 ASIG5V.n3698 ASIG5V.n3697 1.1255
R43164 ASIG5V.n3700 ASIG5V.n3699 1.1255
R43165 ASIG5V.n3526 ASIG5V.n3525 1.1255
R43166 ASIG5V.n3703 ASIG5V.n3702 1.1255
R43167 ASIG5V.n3653 ASIG5V.n3652 1.1255
R43168 ASIG5V.n3655 ASIG5V.n3654 1.1255
R43169 ASIG5V.n3658 ASIG5V.n3657 1.1255
R43170 ASIG5V.n3660 ASIG5V.n3659 1.1255
R43171 ASIG5V.n3521 ASIG5V.n3520 1.1255
R43172 ASIG5V.n3706 ASIG5V.n3705 1.1255
R43173 ASIG5V.n3709 ASIG5V.n3708 1.1255
R43174 ASIG5V.n3711 ASIG5V.n3710 1.1255
R43175 ASIG5V.n3517 ASIG5V.n3516 1.1255
R43176 ASIG5V.n3664 ASIG5V.n3663 1.1255
R43177 ASIG5V.n3513 ASIG5V.n3512 1.1255
R43178 ASIG5V.n3714 ASIG5V.n3713 1.1255
R43179 ASIG5V.n3717 ASIG5V.n3716 1.1255
R43180 ASIG5V.n3719 ASIG5V.n3718 1.1255
R43181 ASIG5V.n3667 ASIG5V.n3666 1.1255
R43182 ASIG5V.n3669 ASIG5V.n3668 1.1255
R43183 ASIG5V.n3507 ASIG5V.n3506 1.1255
R43184 ASIG5V.n3504 ASIG5V.n3503 1.1255
R43185 ASIG5V.n3722 ASIG5V.n3721 1.1255
R43186 ASIG5V.n3724 ASIG5V.n3723 1.1255
R43187 ASIG5V.n3501 ASIG5V.n3500 1.1255
R43188 ASIG5V.n3727 ASIG5V.n3726 1.1255
R43189 ASIG5V.n3498 ASIG5V.n3497 1.1255
R43190 ASIG5V.n3673 ASIG5V.n3672 1.1255
R43191 ASIG5V.n3495 ASIG5V.n3494 1.1255
R43192 ASIG5V.n3730 ASIG5V.n3729 1.1255
R43193 ASIG5V.n3492 ASIG5V.n3491 1.1255
R43194 ASIG5V.n3733 ASIG5V.n3732 1.1255
R43195 ASIG5V.n3960 ASIG5V.n3959 1.1255
R43196 ASIG5V.n3912 ASIG5V.n3911 1.1255
R43197 ASIG5V.n3914 ASIG5V.n3913 1.1255
R43198 ASIG5V.n3917 ASIG5V.n3916 1.1255
R43199 ASIG5V.n3812 ASIG5V.n3811 1.1255
R43200 ASIG5V.n3963 ASIG5V.n3962 1.1255
R43201 ASIG5V.n3965 ASIG5V.n3964 1.1255
R43202 ASIG5V.n3968 ASIG5V.n3967 1.1255
R43203 ASIG5V.n3806 ASIG5V.n3805 1.1255
R43204 ASIG5V.n3808 ASIG5V.n3807 1.1255
R43205 ASIG5V.n3803 ASIG5V.n3802 1.1255
R43206 ASIG5V.n3971 ASIG5V.n3970 1.1255
R43207 ASIG5V.n3800 ASIG5V.n3799 1.1255
R43208 ASIG5V.n3974 ASIG5V.n3973 1.1255
R43209 ASIG5V.n3797 ASIG5V.n3796 1.1255
R43210 ASIG5V.n3921 ASIG5V.n3920 1.1255
R43211 ASIG5V.n3794 ASIG5V.n3793 1.1255
R43212 ASIG5V.n3924 ASIG5V.n3923 1.1255
R43213 ASIG5V.n3791 ASIG5V.n3790 1.1255
R43214 ASIG5V.n3977 ASIG5V.n3976 1.1255
R43215 ASIG5V.n3788 ASIG5V.n3787 1.1255
R43216 ASIG5V.n3980 ASIG5V.n3979 1.1255
R43217 ASIG5V.n3785 ASIG5V.n3784 1.1255
R43218 ASIG5V.n3928 ASIG5V.n3927 1.1255
R43219 ASIG5V.n3781 ASIG5V.n3780 1.1255
R43220 ASIG5V.n3984 ASIG5V.n3983 1.1255
R43221 ASIG5V.n3777 ASIG5V.n3776 1.1255
R43222 ASIG5V.n3988 ASIG5V.n3987 1.1255
R43223 ASIG5V.n3773 ASIG5V.n3772 1.1255
R43224 ASIG5V.n3931 ASIG5V.n3930 1.1255
R43225 ASIG5V.n3770 ASIG5V.n3769 1.1255
R43226 ASIG5V.n3934 ASIG5V.n3933 1.1255
R43227 ASIG5V.n3936 ASIG5V.n3935 1.1255
R43228 ASIG5V.n3767 ASIG5V.n3766 1.1255
R43229 ASIG5V.n3991 ASIG5V.n3990 1.1255
R43230 ASIG5V.n3994 ASIG5V.n3993 1.1255
R43231 ASIG5V.n3763 ASIG5V.n3762 1.1255
R43232 ASIG5V.n3939 ASIG5V.n3938 1.1255
R43233 ASIG5V.n3941 ASIG5V.n3940 1.1255
R43234 ASIG5V.n3760 ASIG5V.n3759 1.1255
R43235 ASIG5V.n3757 ASIG5V.n3756 1.1255
R43236 ASIG5V.n3998 ASIG5V.n3997 1.1255
R43237 ASIG5V.n4000 ASIG5V.n3999 1.1255
R43238 ASIG5V.n3944 ASIG5V.n3943 1.1255
R43239 ASIG5V.n3753 ASIG5V.n3752 1.1255
R43240 ASIG5V.n4084 ASIG5V.n4083 1.1255
R43241 ASIG5V.n4182 ASIG5V.n4181 1.1255
R43242 ASIG5V.n4081 ASIG5V.n4080 1.1255
R43243 ASIG5V.n4185 ASIG5V.n4184 1.1255
R43244 ASIG5V.n4187 ASIG5V.n4186 1.1255
R43245 ASIG5V.n4233 ASIG5V.n4232 1.1255
R43246 ASIG5V.n4077 ASIG5V.n4076 1.1255
R43247 ASIG5V.n4236 ASIG5V.n4235 1.1255
R43248 ASIG5V.n4238 ASIG5V.n4237 1.1255
R43249 ASIG5V.n4190 ASIG5V.n4189 1.1255
R43250 ASIG5V.n4073 ASIG5V.n4072 1.1255
R43251 ASIG5V.n4241 ASIG5V.n4240 1.1255
R43252 ASIG5V.n4070 ASIG5V.n4069 1.1255
R43253 ASIG5V.n4244 ASIG5V.n4243 1.1255
R43254 ASIG5V.n4067 ASIG5V.n4066 1.1255
R43255 ASIG5V.n4193 ASIG5V.n4192 1.1255
R43256 ASIG5V.n4064 ASIG5V.n4063 1.1255
R43257 ASIG5V.n4196 ASIG5V.n4195 1.1255
R43258 ASIG5V.n4061 ASIG5V.n4060 1.1255
R43259 ASIG5V.n4247 ASIG5V.n4246 1.1255
R43260 ASIG5V.n4058 ASIG5V.n4057 1.1255
R43261 ASIG5V.n4251 ASIG5V.n4250 1.1255
R43262 ASIG5V.n4055 ASIG5V.n4054 1.1255
R43263 ASIG5V.n4200 ASIG5V.n4199 1.1255
R43264 ASIG5V.n4051 ASIG5V.n4050 1.1255
R43265 ASIG5V.n4255 ASIG5V.n4254 1.1255
R43266 ASIG5V.n4047 ASIG5V.n4046 1.1255
R43267 ASIG5V.n4259 ASIG5V.n4258 1.1255
R43268 ASIG5V.n4043 ASIG5V.n4042 1.1255
R43269 ASIG5V.n4204 ASIG5V.n4203 1.1255
R43270 ASIG5V.n4039 ASIG5V.n4038 1.1255
R43271 ASIG5V.n4207 ASIG5V.n4206 1.1255
R43272 ASIG5V.n4035 ASIG5V.n4034 1.1255
R43273 ASIG5V.n4262 ASIG5V.n4261 1.1255
R43274 ASIG5V.n4032 ASIG5V.n4031 1.1255
R43275 ASIG5V.n4265 ASIG5V.n4264 1.1255
R43276 ASIG5V.n4029 ASIG5V.n4028 1.1255
R43277 ASIG5V.n4210 ASIG5V.n4209 1.1255
R43278 ASIG5V.n4026 ASIG5V.n4025 1.1255
R43279 ASIG5V.n4268 ASIG5V.n4267 1.1255
R43280 ASIG5V.n4270 ASIG5V.n4269 1.1255
R43281 ASIG5V.n4273 ASIG5V.n4272 1.1255
R43282 ASIG5V.n4022 ASIG5V.n4021 1.1255
R43283 ASIG5V.n4213 ASIG5V.n4212 1.1255
R43284 ASIG5V.n4019 ASIG5V.n4018 1.1255
R43285 ASIG5V.n4216 ASIG5V.n4215 1.1255
R43286 ASIG5V.n4016 ASIG5V.n4015 1.1255
R43287 ASIG5V.n4359 ASIG5V.n4358 1.1255
R43288 ASIG5V.n4462 ASIG5V.n4461 1.1255
R43289 ASIG5V.n4356 ASIG5V.n4355 1.1255
R43290 ASIG5V.n4465 ASIG5V.n4464 1.1255
R43291 ASIG5V.n4467 ASIG5V.n4466 1.1255
R43292 ASIG5V.n4514 ASIG5V.n4513 1.1255
R43293 ASIG5V.n4352 ASIG5V.n4351 1.1255
R43294 ASIG5V.n4517 ASIG5V.n4516 1.1255
R43295 ASIG5V.n4349 ASIG5V.n4348 1.1255
R43296 ASIG5V.n4470 ASIG5V.n4469 1.1255
R43297 ASIG5V.n4346 ASIG5V.n4345 1.1255
R43298 ASIG5V.n4520 ASIG5V.n4519 1.1255
R43299 ASIG5V.n4343 ASIG5V.n4342 1.1255
R43300 ASIG5V.n4523 ASIG5V.n4522 1.1255
R43301 ASIG5V.n4340 ASIG5V.n4339 1.1255
R43302 ASIG5V.n4473 ASIG5V.n4472 1.1255
R43303 ASIG5V.n4337 ASIG5V.n4336 1.1255
R43304 ASIG5V.n4476 ASIG5V.n4475 1.1255
R43305 ASIG5V.n4334 ASIG5V.n4333 1.1255
R43306 ASIG5V.n4527 ASIG5V.n4526 1.1255
R43307 ASIG5V.n4530 ASIG5V.n4529 1.1255
R43308 ASIG5V.n4534 ASIG5V.n4533 1.1255
R43309 ASIG5V.n4330 ASIG5V.n4329 1.1255
R43310 ASIG5V.n4480 ASIG5V.n4479 1.1255
R43311 ASIG5V.n4326 ASIG5V.n4325 1.1255
R43312 ASIG5V.n4538 ASIG5V.n4537 1.1255
R43313 ASIG5V.n4322 ASIG5V.n4321 1.1255
R43314 ASIG5V.n4542 ASIG5V.n4541 1.1255
R43315 ASIG5V.n4318 ASIG5V.n4317 1.1255
R43316 ASIG5V.n4484 ASIG5V.n4483 1.1255
R43317 ASIG5V.n4314 ASIG5V.n4313 1.1255
R43318 ASIG5V.n4488 ASIG5V.n4487 1.1255
R43319 ASIG5V.n4310 ASIG5V.n4309 1.1255
R43320 ASIG5V.n4545 ASIG5V.n4544 1.1255
R43321 ASIG5V.n4306 ASIG5V.n4305 1.1255
R43322 ASIG5V.n4548 ASIG5V.n4547 1.1255
R43323 ASIG5V.n4303 ASIG5V.n4302 1.1255
R43324 ASIG5V.n4491 ASIG5V.n4490 1.1255
R43325 ASIG5V.n4300 ASIG5V.n4299 1.1255
R43326 ASIG5V.n4551 ASIG5V.n4550 1.1255
R43327 ASIG5V.n4297 ASIG5V.n4296 1.1255
R43328 ASIG5V.n4554 ASIG5V.n4553 1.1255
R43329 ASIG5V.n4294 ASIG5V.n4293 1.1255
R43330 ASIG5V.n4494 ASIG5V.n4493 1.1255
R43331 ASIG5V.n4496 ASIG5V.n4495 1.1255
R43332 ASIG5V.n4499 ASIG5V.n4498 1.1255
R43333 ASIG5V.n4290 ASIG5V.n4289 1.1255
R43334 ASIG5V.n4557 ASIG5V.n4556 1.1255
R43335 ASIG5V.n4782 ASIG5V.n4781 1.1255
R43336 ASIG5V.n4719 ASIG5V.n4718 1.1255
R43337 ASIG5V.n4721 ASIG5V.n4720 1.1255
R43338 ASIG5V.n4724 ASIG5V.n4723 1.1255
R43339 ASIG5V.n4726 ASIG5V.n4725 1.1255
R43340 ASIG5V.n4785 ASIG5V.n4784 1.1255
R43341 ASIG5V.n4787 ASIG5V.n4786 1.1255
R43342 ASIG5V.n4790 ASIG5V.n4789 1.1255
R43343 ASIG5V.n4792 ASIG5V.n4791 1.1255
R43344 ASIG5V.n4729 ASIG5V.n4728 1.1255
R43345 ASIG5V.n4731 ASIG5V.n4730 1.1255
R43346 ASIG5V.n4795 ASIG5V.n4794 1.1255
R43347 ASIG5V.n4613 ASIG5V.n4612 1.1255
R43348 ASIG5V.n4798 ASIG5V.n4797 1.1255
R43349 ASIG5V.n4800 ASIG5V.n4799 1.1255
R43350 ASIG5V.n4734 ASIG5V.n4733 1.1255
R43351 ASIG5V.n4736 ASIG5V.n4735 1.1255
R43352 ASIG5V.n4739 ASIG5V.n4738 1.1255
R43353 ASIG5V.n4608 ASIG5V.n4607 1.1255
R43354 ASIG5V.n4804 ASIG5V.n4803 1.1255
R43355 ASIG5V.n4807 ASIG5V.n4806 1.1255
R43356 ASIG5V.n4811 ASIG5V.n4810 1.1255
R43357 ASIG5V.n4600 ASIG5V.n4599 1.1255
R43358 ASIG5V.n4603 ASIG5V.n4602 1.1255
R43359 ASIG5V.n4596 ASIG5V.n4595 1.1255
R43360 ASIG5V.n4815 ASIG5V.n4814 1.1255
R43361 ASIG5V.n4818 ASIG5V.n4817 1.1255
R43362 ASIG5V.n4822 ASIG5V.n4821 1.1255
R43363 ASIG5V.n4825 ASIG5V.n4824 1.1255
R43364 ASIG5V.n4744 ASIG5V.n4743 1.1255
R43365 ASIG5V.n4747 ASIG5V.n4746 1.1255
R43366 ASIG5V.n4751 ASIG5V.n4750 1.1255
R43367 ASIG5V.n4589 ASIG5V.n4588 1.1255
R43368 ASIG5V.n4829 ASIG5V.n4828 1.1255
R43369 ASIG5V.n4585 ASIG5V.n4584 1.1255
R43370 ASIG5V.n4832 ASIG5V.n4831 1.1255
R43371 ASIG5V.n4834 ASIG5V.n4833 1.1255
R43372 ASIG5V.n4754 ASIG5V.n4753 1.1255
R43373 ASIG5V.n4756 ASIG5V.n4755 1.1255
R43374 ASIG5V.n4837 ASIG5V.n4836 1.1255
R43375 ASIG5V.n4839 ASIG5V.n4838 1.1255
R43376 ASIG5V.n4842 ASIG5V.n4841 1.1255
R43377 ASIG5V.n4578 ASIG5V.n4577 1.1255
R43378 ASIG5V.n4759 ASIG5V.n4758 1.1255
R43379 ASIG5V.n4761 ASIG5V.n4760 1.1255
R43380 ASIG5V.n4764 ASIG5V.n4763 1.1255
R43381 ASIG5V.n4766 ASIG5V.n4765 1.1255
R43382 ASIG5V.n4845 ASIG5V.n4844 1.1255
R43383 ASIG5V.n4703 ASIG5V.n4702 1.1255
R43384 ASIG5V.n5072 ASIG5V.n5071 1.1255
R43385 ASIG5V.n4994 ASIG5V.n4993 1.1255
R43386 ASIG5V.n4996 ASIG5V.n4995 1.1255
R43387 ASIG5V.n4999 ASIG5V.n4998 1.1255
R43388 ASIG5V.n5001 ASIG5V.n5000 1.1255
R43389 ASIG5V.n5075 ASIG5V.n5074 1.1255
R43390 ASIG5V.n5077 ASIG5V.n5076 1.1255
R43391 ASIG5V.n5080 ASIG5V.n5079 1.1255
R43392 ASIG5V.n5082 ASIG5V.n5081 1.1255
R43393 ASIG5V.n5004 ASIG5V.n5003 1.1255
R43394 ASIG5V.n5006 ASIG5V.n5005 1.1255
R43395 ASIG5V.n5085 ASIG5V.n5084 1.1255
R43396 ASIG5V.n5087 ASIG5V.n5086 1.1255
R43397 ASIG5V.n5090 ASIG5V.n5089 1.1255
R43398 ASIG5V.n5092 ASIG5V.n5091 1.1255
R43399 ASIG5V.n5009 ASIG5V.n5008 1.1255
R43400 ASIG5V.n5012 ASIG5V.n5011 1.1255
R43401 ASIG5V.n5016 ASIG5V.n5015 1.1255
R43402 ASIG5V.n5019 ASIG5V.n5018 1.1255
R43403 ASIG5V.n5096 ASIG5V.n5095 1.1255
R43404 ASIG5V.n5099 ASIG5V.n5098 1.1255
R43405 ASIG5V.n5103 ASIG5V.n5102 1.1255
R43406 ASIG5V.n5106 ASIG5V.n5105 1.1255
R43407 ASIG5V.n5023 ASIG5V.n5022 1.1255
R43408 ASIG5V.n5026 ASIG5V.n5025 1.1255
R43409 ASIG5V.n5110 ASIG5V.n5109 1.1255
R43410 ASIG5V.n5113 ASIG5V.n5112 1.1255
R43411 ASIG5V.n5117 ASIG5V.n5116 1.1255
R43412 ASIG5V.n5120 ASIG5V.n5119 1.1255
R43413 ASIG5V.n5030 ASIG5V.n5029 1.1255
R43414 ASIG5V.n5033 ASIG5V.n5032 1.1255
R43415 ASIG5V.n5037 ASIG5V.n5036 1.1255
R43416 ASIG5V.n5040 ASIG5V.n5039 1.1255
R43417 ASIG5V.n5124 ASIG5V.n5123 1.1255
R43418 ASIG5V.n5127 ASIG5V.n5126 1.1255
R43419 ASIG5V.n5131 ASIG5V.n5130 1.1255
R43420 ASIG5V.n4872 ASIG5V.n4871 1.1255
R43421 ASIG5V.n5044 ASIG5V.n5043 1.1255
R43422 ASIG5V.n5046 ASIG5V.n5045 1.1255
R43423 ASIG5V.n5134 ASIG5V.n5133 1.1255
R43424 ASIG5V.n4867 ASIG5V.n4866 1.1255
R43425 ASIG5V.n5137 ASIG5V.n5136 1.1255
R43426 ASIG5V.n4864 ASIG5V.n4863 1.1255
R43427 ASIG5V.n5049 ASIG5V.n5048 1.1255
R43428 ASIG5V.n5051 ASIG5V.n5050 1.1255
R43429 ASIG5V.n5054 ASIG5V.n5053 1.1255
R43430 ASIG5V.n5056 ASIG5V.n5055 1.1255
R43431 ASIG5V.n5140 ASIG5V.n5139 1.1255
R43432 ASIG5V.n4978 ASIG5V.n4977 1.1255
R43433 ASIG5V.n5295 ASIG5V.n5294 1.1255
R43434 ASIG5V.n5297 ASIG5V.n5296 1.1255
R43435 ASIG5V.n5290 ASIG5V.n5289 1.1255
R43436 ASIG5V.n5292 ASIG5V.n5291 1.1255
R43437 ASIG5V.n5287 ASIG5V.n5286 1.1255
R43438 ASIG5V.n5426 ASIG5V.n5425 1.1255
R43439 ASIG5V.n5282 ASIG5V.n5281 1.1255
R43440 ASIG5V.n5284 ASIG5V.n5283 1.1255
R43441 ASIG5V.n5277 ASIG5V.n5276 1.1255
R43442 ASIG5V.n5279 ASIG5V.n5278 1.1255
R43443 ASIG5V.n5272 ASIG5V.n5271 1.1255
R43444 ASIG5V.n5274 ASIG5V.n5273 1.1255
R43445 ASIG5V.n5267 ASIG5V.n5266 1.1255
R43446 ASIG5V.n5269 ASIG5V.n5268 1.1255
R43447 ASIG5V.n5261 ASIG5V.n5260 1.1255
R43448 ASIG5V.n5264 ASIG5V.n5263 1.1255
R43449 ASIG5V.n5255 ASIG5V.n5254 1.1255
R43450 ASIG5V.n5258 ASIG5V.n5257 1.1255
R43451 ASIG5V.n5248 ASIG5V.n5247 1.1255
R43452 ASIG5V.n5251 ASIG5V.n5250 1.1255
R43453 ASIG5V.n5241 ASIG5V.n5240 1.1255
R43454 ASIG5V.n5244 ASIG5V.n5243 1.1255
R43455 ASIG5V.n5234 ASIG5V.n5233 1.1255
R43456 ASIG5V.n5237 ASIG5V.n5236 1.1255
R43457 ASIG5V.n5227 ASIG5V.n5226 1.1255
R43458 ASIG5V.n5230 ASIG5V.n5229 1.1255
R43459 ASIG5V.n5220 ASIG5V.n5219 1.1255
R43460 ASIG5V.n5223 ASIG5V.n5222 1.1255
R43461 ASIG5V.n5213 ASIG5V.n5212 1.1255
R43462 ASIG5V.n5216 ASIG5V.n5215 1.1255
R43463 ASIG5V.n5206 ASIG5V.n5205 1.1255
R43464 ASIG5V.n5209 ASIG5V.n5208 1.1255
R43465 ASIG5V.n5199 ASIG5V.n5198 1.1255
R43466 ASIG5V.n5202 ASIG5V.n5201 1.1255
R43467 ASIG5V.n5192 ASIG5V.n5191 1.1255
R43468 ASIG5V.n5195 ASIG5V.n5194 1.1255
R43469 ASIG5V.n5185 ASIG5V.n5184 1.1255
R43470 ASIG5V.n5188 ASIG5V.n5187 1.1255
R43471 ASIG5V.n5178 ASIG5V.n5177 1.1255
R43472 ASIG5V.n5181 ASIG5V.n5180 1.1255
R43473 ASIG5V.n5172 ASIG5V.n5171 1.1255
R43474 ASIG5V.n5174 ASIG5V.n5173 1.1255
R43475 ASIG5V.n5167 ASIG5V.n5166 1.1255
R43476 ASIG5V.n5169 ASIG5V.n5168 1.1255
R43477 ASIG5V.n5162 ASIG5V.n5161 1.1255
R43478 ASIG5V.n5164 ASIG5V.n5163 1.1255
R43479 ASIG5V.n5157 ASIG5V.n5156 1.1255
R43480 ASIG5V.n5159 ASIG5V.n5158 1.1255
R43481 ASIG5V.n5403 ASIG5V.n5402 1.1255
R43482 ASIG5V.n5539 ASIG5V.n5538 1.1255
R43483 ASIG5V.n5694 ASIG5V.n5693 1.1255
R43484 ASIG5V.n5536 ASIG5V.n5535 1.1255
R43485 ASIG5V.n5697 ASIG5V.n5696 1.1255
R43486 ASIG5V.n5533 ASIG5V.n5532 1.1255
R43487 ASIG5V.n5747 ASIG5V.n5746 1.1255
R43488 ASIG5V.n5530 ASIG5V.n5529 1.1255
R43489 ASIG5V.n5750 ASIG5V.n5749 1.1255
R43490 ASIG5V.n5527 ASIG5V.n5526 1.1255
R43491 ASIG5V.n5700 ASIG5V.n5699 1.1255
R43492 ASIG5V.n5524 ASIG5V.n5523 1.1255
R43493 ASIG5V.n5753 ASIG5V.n5752 1.1255
R43494 ASIG5V.n5521 ASIG5V.n5520 1.1255
R43495 ASIG5V.n5756 ASIG5V.n5755 1.1255
R43496 ASIG5V.n5518 ASIG5V.n5517 1.1255
R43497 ASIG5V.n5704 ASIG5V.n5703 1.1255
R43498 ASIG5V.n5514 ASIG5V.n5513 1.1255
R43499 ASIG5V.n5708 ASIG5V.n5707 1.1255
R43500 ASIG5V.n5510 ASIG5V.n5509 1.1255
R43501 ASIG5V.n5760 ASIG5V.n5759 1.1255
R43502 ASIG5V.n5506 ASIG5V.n5505 1.1255
R43503 ASIG5V.n5764 ASIG5V.n5763 1.1255
R43504 ASIG5V.n5502 ASIG5V.n5501 1.1255
R43505 ASIG5V.n5712 ASIG5V.n5711 1.1255
R43506 ASIG5V.n5498 ASIG5V.n5497 1.1255
R43507 ASIG5V.n5768 ASIG5V.n5767 1.1255
R43508 ASIG5V.n5771 ASIG5V.n5770 1.1255
R43509 ASIG5V.n5775 ASIG5V.n5774 1.1255
R43510 ASIG5V.n5778 ASIG5V.n5777 1.1255
R43511 ASIG5V.n5716 ASIG5V.n5715 1.1255
R43512 ASIG5V.n5492 ASIG5V.n5491 1.1255
R43513 ASIG5V.n5720 ASIG5V.n5719 1.1255
R43514 ASIG5V.n5485 ASIG5V.n5484 1.1255
R43515 ASIG5V.n5488 ASIG5V.n5487 1.1255
R43516 ASIG5V.n5481 ASIG5V.n5480 1.1255
R43517 ASIG5V.n5783 ASIG5V.n5782 1.1255
R43518 ASIG5V.n5477 ASIG5V.n5476 1.1255
R43519 ASIG5V.n5724 ASIG5V.n5723 1.1255
R43520 ASIG5V.n5473 ASIG5V.n5472 1.1255
R43521 ASIG5V.n5787 ASIG5V.n5786 1.1255
R43522 ASIG5V.n5466 ASIG5V.n5465 1.1255
R43523 ASIG5V.n5469 ASIG5V.n5468 1.1255
R43524 ASIG5V.n5462 ASIG5V.n5461 1.1255
R43525 ASIG5V.n5727 ASIG5V.n5726 1.1255
R43526 ASIG5V.n5729 ASIG5V.n5728 1.1255
R43527 ASIG5V.n5732 ASIG5V.n5731 1.1255
R43528 ASIG5V.n5734 ASIG5V.n5733 1.1255
R43529 ASIG5V.n5791 ASIG5V.n5790 1.1255
R43530 ASIG5V.n5683 ASIG5V.n5682 1.1255
R43531 ASIG5V.n6077 ASIG5V.n6076 1.1255
R43532 ASIG5V.n5995 ASIG5V.n5994 1.1255
R43533 ASIG5V.n5997 ASIG5V.n5996 1.1255
R43534 ASIG5V.n6000 ASIG5V.n5999 1.1255
R43535 ASIG5V.n6002 ASIG5V.n6001 1.1255
R43536 ASIG5V.n6080 ASIG5V.n6079 1.1255
R43537 ASIG5V.n6082 ASIG5V.n6081 1.1255
R43538 ASIG5V.n6085 ASIG5V.n6084 1.1255
R43539 ASIG5V.n6087 ASIG5V.n6086 1.1255
R43540 ASIG5V.n6005 ASIG5V.n6004 1.1255
R43541 ASIG5V.n6007 ASIG5V.n6006 1.1255
R43542 ASIG5V.n6090 ASIG5V.n6089 1.1255
R43543 ASIG5V.n6092 ASIG5V.n6091 1.1255
R43544 ASIG5V.n6095 ASIG5V.n6094 1.1255
R43545 ASIG5V.n6098 ASIG5V.n6097 1.1255
R43546 ASIG5V.n6011 ASIG5V.n6010 1.1255
R43547 ASIG5V.n6014 ASIG5V.n6013 1.1255
R43548 ASIG5V.n6018 ASIG5V.n6017 1.1255
R43549 ASIG5V.n6021 ASIG5V.n6020 1.1255
R43550 ASIG5V.n6102 ASIG5V.n6101 1.1255
R43551 ASIG5V.n6105 ASIG5V.n6104 1.1255
R43552 ASIG5V.n6109 ASIG5V.n6108 1.1255
R43553 ASIG5V.n6112 ASIG5V.n6111 1.1255
R43554 ASIG5V.n6025 ASIG5V.n6024 1.1255
R43555 ASIG5V.n6028 ASIG5V.n6027 1.1255
R43556 ASIG5V.n6116 ASIG5V.n6115 1.1255
R43557 ASIG5V.n6119 ASIG5V.n6118 1.1255
R43558 ASIG5V.n6123 ASIG5V.n6122 1.1255
R43559 ASIG5V.n6126 ASIG5V.n6125 1.1255
R43560 ASIG5V.n6032 ASIG5V.n6031 1.1255
R43561 ASIG5V.n6035 ASIG5V.n6034 1.1255
R43562 ASIG5V.n6039 ASIG5V.n6038 1.1255
R43563 ASIG5V.n6042 ASIG5V.n6041 1.1255
R43564 ASIG5V.n6130 ASIG5V.n6129 1.1255
R43565 ASIG5V.n6133 ASIG5V.n6132 1.1255
R43566 ASIG5V.n5827 ASIG5V.n5826 1.1255
R43567 ASIG5V.n5823 ASIG5V.n5822 1.1255
R43568 ASIG5V.n6046 ASIG5V.n6045 1.1255
R43569 ASIG5V.n6049 ASIG5V.n6048 1.1255
R43570 ASIG5V.n6138 ASIG5V.n6137 1.1255
R43571 ASIG5V.n6141 ASIG5V.n6140 1.1255
R43572 ASIG5V.n5818 ASIG5V.n5817 1.1255
R43573 ASIG5V.n5814 ASIG5V.n5813 1.1255
R43574 ASIG5V.n6053 ASIG5V.n6052 1.1255
R43575 ASIG5V.n6056 ASIG5V.n6055 1.1255
R43576 ASIG5V.n6059 ASIG5V.n6058 1.1255
R43577 ASIG5V.n6061 ASIG5V.n6060 1.1255
R43578 ASIG5V.n6145 ASIG5V.n6144 1.1255
R43579 ASIG5V.n5979 ASIG5V.n5978 1.1255
R43580 ASIG5V.n6293 ASIG5V.n6292 1.1255
R43581 ASIG5V.n6295 ASIG5V.n6294 1.1255
R43582 ASIG5V.n6288 ASIG5V.n6287 1.1255
R43583 ASIG5V.n6290 ASIG5V.n6289 1.1255
R43584 ASIG5V.n6283 ASIG5V.n6282 1.1255
R43585 ASIG5V.n6285 ASIG5V.n6284 1.1255
R43586 ASIG5V.n6278 ASIG5V.n6277 1.1255
R43587 ASIG5V.n6280 ASIG5V.n6279 1.1255
R43588 ASIG5V.n6273 ASIG5V.n6272 1.1255
R43589 ASIG5V.n6275 ASIG5V.n6274 1.1255
R43590 ASIG5V.n6268 ASIG5V.n6267 1.1255
R43591 ASIG5V.n6270 ASIG5V.n6269 1.1255
R43592 ASIG5V.n6263 ASIG5V.n6262 1.1255
R43593 ASIG5V.n6265 ASIG5V.n6264 1.1255
R43594 ASIG5V.n6257 ASIG5V.n6256 1.1255
R43595 ASIG5V.n6260 ASIG5V.n6259 1.1255
R43596 ASIG5V.n6250 ASIG5V.n6249 1.1255
R43597 ASIG5V.n6253 ASIG5V.n6252 1.1255
R43598 ASIG5V.n6243 ASIG5V.n6242 1.1255
R43599 ASIG5V.n6246 ASIG5V.n6245 1.1255
R43600 ASIG5V.n6236 ASIG5V.n6235 1.1255
R43601 ASIG5V.n6239 ASIG5V.n6238 1.1255
R43602 ASIG5V.n6229 ASIG5V.n6228 1.1255
R43603 ASIG5V.n6232 ASIG5V.n6231 1.1255
R43604 ASIG5V.n6222 ASIG5V.n6221 1.1255
R43605 ASIG5V.n6225 ASIG5V.n6224 1.1255
R43606 ASIG5V.n6215 ASIG5V.n6214 1.1255
R43607 ASIG5V.n6218 ASIG5V.n6217 1.1255
R43608 ASIG5V.n6208 ASIG5V.n6207 1.1255
R43609 ASIG5V.n6211 ASIG5V.n6210 1.1255
R43610 ASIG5V.n6201 ASIG5V.n6200 1.1255
R43611 ASIG5V.n6204 ASIG5V.n6203 1.1255
R43612 ASIG5V.n7080 ASIG5V.n7079 1.1255
R43613 ASIG5V.n7112 ASIG5V.n7111 1.1255
R43614 ASIG5V.n6196 ASIG5V.n6195 1.1255
R43615 ASIG5V.n7116 ASIG5V.n7115 1.1255
R43616 ASIG5V.n6192 ASIG5V.n6191 1.1255
R43617 ASIG5V.n7084 ASIG5V.n7083 1.1255
R43618 ASIG5V.n7087 ASIG5V.n7086 1.1255
R43619 ASIG5V.n6188 ASIG5V.n6187 1.1255
R43620 ASIG5V.n6181 ASIG5V.n6180 1.1255
R43621 ASIG5V.n6184 ASIG5V.n6183 1.1255
R43622 ASIG5V.n6177 ASIG5V.n6176 1.1255
R43623 ASIG5V.n7091 ASIG5V.n7090 1.1255
R43624 ASIG5V.n6173 ASIG5V.n6172 1.1255
R43625 ASIG5V.n7095 ASIG5V.n7094 1.1255
R43626 ASIG5V.n6169 ASIG5V.n6168 1.1255
R43627 ASIG5V.n7121 ASIG5V.n7120 1.1255
R43628 ASIG5V.n6336 ASIG5V.n6335 1.1255
R43629 ASIG5V.n6843 ASIG5V.n6842 1.1255
R43630 ASIG5V.n6401 ASIG5V.n6400 1.1255
R43631 ASIG5V.n6398 ASIG5V.n6397 1.1255
R43632 ASIG5V.n6800 ASIG5V.n6799 1.1255
R43633 ASIG5V.n6395 ASIG5V.n6394 1.1255
R43634 ASIG5V.n6846 ASIG5V.n6845 1.1255
R43635 ASIG5V.n6848 ASIG5V.n6847 1.1255
R43636 ASIG5V.n6851 ASIG5V.n6850 1.1255
R43637 ASIG5V.n6853 ASIG5V.n6852 1.1255
R43638 ASIG5V.n6391 ASIG5V.n6390 1.1255
R43639 ASIG5V.n6388 ASIG5V.n6387 1.1255
R43640 ASIG5V.n6856 ASIG5V.n6855 1.1255
R43641 ASIG5V.n6858 ASIG5V.n6857 1.1255
R43642 ASIG5V.n6861 ASIG5V.n6860 1.1255
R43643 ASIG5V.n6863 ASIG5V.n6862 1.1255
R43644 ASIG5V.n6805 ASIG5V.n6804 1.1255
R43645 ASIG5V.n6383 ASIG5V.n6382 1.1255
R43646 ASIG5V.n6809 ASIG5V.n6808 1.1255
R43647 ASIG5V.n6379 ASIG5V.n6378 1.1255
R43648 ASIG5V.n6867 ASIG5V.n6866 1.1255
R43649 ASIG5V.n6870 ASIG5V.n6869 1.1255
R43650 ASIG5V.n6874 ASIG5V.n6873 1.1255
R43651 ASIG5V.n6877 ASIG5V.n6876 1.1255
R43652 ASIG5V.n6813 ASIG5V.n6812 1.1255
R43653 ASIG5V.n6373 ASIG5V.n6372 1.1255
R43654 ASIG5V.n6881 ASIG5V.n6880 1.1255
R43655 ASIG5V.n6884 ASIG5V.n6883 1.1255
R43656 ASIG5V.n6888 ASIG5V.n6887 1.1255
R43657 ASIG5V.n6891 ASIG5V.n6890 1.1255
R43658 ASIG5V.n6817 ASIG5V.n6816 1.1255
R43659 ASIG5V.n6364 ASIG5V.n6363 1.1255
R43660 ASIG5V.n6367 ASIG5V.n6366 1.1255
R43661 ASIG5V.n6360 ASIG5V.n6359 1.1255
R43662 ASIG5V.n6895 ASIG5V.n6894 1.1255
R43663 ASIG5V.n6898 ASIG5V.n6897 1.1255
R43664 ASIG5V.n6902 ASIG5V.n6901 1.1255
R43665 ASIG5V.n6905 ASIG5V.n6904 1.1255
R43666 ASIG5V.n6355 ASIG5V.n6354 1.1255
R43667 ASIG5V.n6351 ASIG5V.n6350 1.1255
R43668 ASIG5V.n6909 ASIG5V.n6908 1.1255
R43669 ASIG5V.n6912 ASIG5V.n6911 1.1255
R43670 ASIG5V.n6916 ASIG5V.n6915 1.1255
R43671 ASIG5V.n6919 ASIG5V.n6918 1.1255
R43672 ASIG5V.n6823 ASIG5V.n6822 1.1255
R43673 ASIG5V.n6345 ASIG5V.n6344 1.1255
R43674 ASIG5V.n6827 ASIG5V.n6826 1.1255
R43675 ASIG5V.n6341 ASIG5V.n6340 1.1255
R43676 ASIG5V.n6923 ASIG5V.n6922 1.1255
R43677 ASIG5V.n6421 ASIG5V.n6420 1.1255
R43678 ASIG5V.n6530 ASIG5V.n6529 1.1255
R43679 ASIG5V.n6563 ASIG5V.n6562 1.1255
R43680 ASIG5V.n6525 ASIG5V.n6524 1.1255
R43681 ASIG5V.n6527 ASIG5V.n6526 1.1255
R43682 ASIG5V.n6522 ASIG5V.n6521 1.1255
R43683 ASIG5V.n6631 ASIG5V.n6630 1.1255
R43684 ASIG5V.n6519 ASIG5V.n6518 1.1255
R43685 ASIG5V.n6634 ASIG5V.n6633 1.1255
R43686 ASIG5V.n6516 ASIG5V.n6515 1.1255
R43687 ASIG5V.n6567 ASIG5V.n6566 1.1255
R43688 ASIG5V.n6513 ASIG5V.n6512 1.1255
R43689 ASIG5V.n6637 ASIG5V.n6636 1.1255
R43690 ASIG5V.n6508 ASIG5V.n6507 1.1255
R43691 ASIG5V.n6510 ASIG5V.n6509 1.1255
R43692 ASIG5V.n6505 ASIG5V.n6504 1.1255
R43693 ASIG5V.n6571 ASIG5V.n6570 1.1255
R43694 ASIG5V.n6501 ASIG5V.n6500 1.1255
R43695 ASIG5V.n6575 ASIG5V.n6574 1.1255
R43696 ASIG5V.n6494 ASIG5V.n6493 1.1255
R43697 ASIG5V.n6497 ASIG5V.n6496 1.1255
R43698 ASIG5V.n6487 ASIG5V.n6486 1.1255
R43699 ASIG5V.n6490 ASIG5V.n6489 1.1255
R43700 ASIG5V.n6483 ASIG5V.n6482 1.1255
R43701 ASIG5V.n6579 ASIG5V.n6578 1.1255
R43702 ASIG5V.n6582 ASIG5V.n6581 1.1255
R43703 ASIG5V.n6644 ASIG5V.n6643 1.1255
R43704 ASIG5V.n6475 ASIG5V.n6474 1.1255
R43705 ASIG5V.n6478 ASIG5V.n6477 1.1255
R43706 ASIG5V.n6471 ASIG5V.n6470 1.1255
R43707 ASIG5V.n6586 ASIG5V.n6585 1.1255
R43708 ASIG5V.n6589 ASIG5V.n6588 1.1255
R43709 ASIG5V.n6593 ASIG5V.n6592 1.1255
R43710 ASIG5V.n6596 ASIG5V.n6595 1.1255
R43711 ASIG5V.n6466 ASIG5V.n6465 1.1255
R43712 ASIG5V.n6459 ASIG5V.n6458 1.1255
R43713 ASIG5V.n6462 ASIG5V.n6461 1.1255
R43714 ASIG5V.n6455 ASIG5V.n6454 1.1255
R43715 ASIG5V.n6600 ASIG5V.n6599 1.1255
R43716 ASIG5V.n6603 ASIG5V.n6602 1.1255
R43717 ASIG5V.n6451 ASIG5V.n6450 1.1255
R43718 ASIG5V.n6444 ASIG5V.n6443 1.1255
R43719 ASIG5V.n6447 ASIG5V.n6446 1.1255
R43720 ASIG5V.n6440 ASIG5V.n6439 1.1255
R43721 ASIG5V.n6607 ASIG5V.n6606 1.1255
R43722 ASIG5V.n6610 ASIG5V.n6609 1.1255
R43723 ASIG5V.n6436 ASIG5V.n6435 1.1255
R43724 ASIG5V.n6614 ASIG5V.n6613 1.1255
R43725 ASIG5V.n6432 ASIG5V.n6431 1.1255
R43726 ASIG5V.n6428 ASIG5V.n6427 1.1255
R43727 ASIG5V.n13415 ASIG5V.n13414 1.1255
R43728 ASIG5V.n13378 ASIG5V.n13377 1.1255
R43729 ASIG5V.n74 ASIG5V.n73 1.1255
R43730 ASIG5V.n13381 ASIG5V.n13380 1.1255
R43731 ASIG5V.n71 ASIG5V.n70 1.1255
R43732 ASIG5V.n13418 ASIG5V.n13417 1.1255
R43733 ASIG5V.n68 ASIG5V.n67 1.1255
R43734 ASIG5V.n13421 ASIG5V.n13420 1.1255
R43735 ASIG5V.n65 ASIG5V.n64 1.1255
R43736 ASIG5V.n13384 ASIG5V.n13383 1.1255
R43737 ASIG5V.n62 ASIG5V.n61 1.1255
R43738 ASIG5V.n13424 ASIG5V.n13423 1.1255
R43739 ASIG5V.n59 ASIG5V.n58 1.1255
R43740 ASIG5V.n13427 ASIG5V.n13426 1.1255
R43741 ASIG5V.n13430 ASIG5V.n13429 1.1255
R43742 ASIG5V.n56 ASIG5V.n55 1.1255
R43743 ASIG5V.n52 ASIG5V.n51 1.1255
R43744 ASIG5V.n13389 ASIG5V.n13388 1.1255
R43745 ASIG5V.n48 ASIG5V.n47 1.1255
R43746 ASIG5V.n13434 ASIG5V.n13433 1.1255
R43747 ASIG5V.n13437 ASIG5V.n13436 1.1255
R43748 ASIG5V.n13441 ASIG5V.n13440 1.1255
R43749 ASIG5V.n13444 ASIG5V.n13443 1.1255
R43750 ASIG5V.n43 ASIG5V.n42 1.1255
R43751 ASIG5V.n39 ASIG5V.n38 1.1255
R43752 ASIG5V.n13448 ASIG5V.n13447 1.1255
R43753 ASIG5V.n13451 ASIG5V.n13450 1.1255
R43754 ASIG5V.n13455 ASIG5V.n13454 1.1255
R43755 ASIG5V.n13458 ASIG5V.n13457 1.1255
R43756 ASIG5V.n13394 ASIG5V.n13393 1.1255
R43757 ASIG5V.n13397 ASIG5V.n13396 1.1255
R43758 ASIG5V.n13401 ASIG5V.n13400 1.1255
R43759 ASIG5V.n32 ASIG5V.n31 1.1255
R43760 ASIG5V.n13462 ASIG5V.n13461 1.1255
R43761 ASIG5V.n13465 ASIG5V.n13464 1.1255
R43762 ASIG5V.n13469 ASIG5V.n13468 1.1255
R43763 ASIG5V.n13472 ASIG5V.n13471 1.1255
R43764 ASIG5V.n27 ASIG5V.n26 1.1255
R43765 ASIG5V.n23 ASIG5V.n22 1.1255
R43766 ASIG5V.n13476 ASIG5V.n13475 1.1255
R43767 ASIG5V.n13479 ASIG5V.n13478 1.1255
R43768 ASIG5V.n13483 ASIG5V.n13482 1.1255
R43769 ASIG5V.n13486 ASIG5V.n13485 1.1255
R43770 ASIG5V.n18 ASIG5V.n17 1.1255
R43771 ASIG5V.n14 ASIG5V.n13 1.1255
R43772 ASIG5V.n13407 ASIG5V.n13406 1.1255
R43773 ASIG5V.n10 ASIG5V.n9 1.1255
R43774 ASIG5V.n13490 ASIG5V.n13489 1.1255
R43775 ASIG5V.n6 ASIG5V.n5 1.1255
R43776 ASIG5V.n246 ASIG5V.n245 1.1255
R43777 ASIG5V.n162 ASIG5V.n161 1.1255
R43778 ASIG5V.n164 ASIG5V.n163 1.1255
R43779 ASIG5V.n167 ASIG5V.n166 1.1255
R43780 ASIG5V.n169 ASIG5V.n168 1.1255
R43781 ASIG5V.n249 ASIG5V.n248 1.1255
R43782 ASIG5V.n251 ASIG5V.n250 1.1255
R43783 ASIG5V.n254 ASIG5V.n253 1.1255
R43784 ASIG5V.n256 ASIG5V.n255 1.1255
R43785 ASIG5V.n172 ASIG5V.n171 1.1255
R43786 ASIG5V.n174 ASIG5V.n173 1.1255
R43787 ASIG5V.n259 ASIG5V.n258 1.1255
R43788 ASIG5V.n261 ASIG5V.n260 1.1255
R43789 ASIG5V.n264 ASIG5V.n263 1.1255
R43790 ASIG5V.n267 ASIG5V.n266 1.1255
R43791 ASIG5V.n178 ASIG5V.n177 1.1255
R43792 ASIG5V.n181 ASIG5V.n180 1.1255
R43793 ASIG5V.n185 ASIG5V.n184 1.1255
R43794 ASIG5V.n188 ASIG5V.n187 1.1255
R43795 ASIG5V.n271 ASIG5V.n270 1.1255
R43796 ASIG5V.n274 ASIG5V.n273 1.1255
R43797 ASIG5V.n278 ASIG5V.n277 1.1255
R43798 ASIG5V.n281 ASIG5V.n280 1.1255
R43799 ASIG5V.n192 ASIG5V.n191 1.1255
R43800 ASIG5V.n195 ASIG5V.n194 1.1255
R43801 ASIG5V.n285 ASIG5V.n284 1.1255
R43802 ASIG5V.n288 ASIG5V.n287 1.1255
R43803 ASIG5V.n292 ASIG5V.n291 1.1255
R43804 ASIG5V.n295 ASIG5V.n294 1.1255
R43805 ASIG5V.n199 ASIG5V.n198 1.1255
R43806 ASIG5V.n202 ASIG5V.n201 1.1255
R43807 ASIG5V.n206 ASIG5V.n205 1.1255
R43808 ASIG5V.n209 ASIG5V.n208 1.1255
R43809 ASIG5V.n299 ASIG5V.n298 1.1255
R43810 ASIG5V.n302 ASIG5V.n301 1.1255
R43811 ASIG5V.n306 ASIG5V.n305 1.1255
R43812 ASIG5V.n309 ASIG5V.n308 1.1255
R43813 ASIG5V.n213 ASIG5V.n212 1.1255
R43814 ASIG5V.n216 ASIG5V.n215 1.1255
R43815 ASIG5V.n313 ASIG5V.n312 1.1255
R43816 ASIG5V.n316 ASIG5V.n315 1.1255
R43817 ASIG5V.n320 ASIG5V.n319 1.1255
R43818 ASIG5V.n323 ASIG5V.n322 1.1255
R43819 ASIG5V.n220 ASIG5V.n219 1.1255
R43820 ASIG5V.n223 ASIG5V.n222 1.1255
R43821 ASIG5V.n227 ASIG5V.n226 1.1255
R43822 ASIG5V.n230 ASIG5V.n229 1.1255
R43823 ASIG5V.n327 ASIG5V.n326 1.1255
R43824 ASIG5V.n146 ASIG5V.n145 1.1255
R43825 ASIG5V.n7376 ASIG5V.n7375 1.1255
R43826 ASIG5V.n7532 ASIG5V.n7531 1.1255
R43827 ASIG5V.n7373 ASIG5V.n7372 1.1255
R43828 ASIG5V.n7535 ASIG5V.n7534 1.1255
R43829 ASIG5V.n7370 ASIG5V.n7369 1.1255
R43830 ASIG5V.n7576 ASIG5V.n7575 1.1255
R43831 ASIG5V.n7367 ASIG5V.n7366 1.1255
R43832 ASIG5V.n7579 ASIG5V.n7578 1.1255
R43833 ASIG5V.n7581 ASIG5V.n7580 1.1255
R43834 ASIG5V.n7538 ASIG5V.n7537 1.1255
R43835 ASIG5V.n7363 ASIG5V.n7362 1.1255
R43836 ASIG5V.n7584 ASIG5V.n7583 1.1255
R43837 ASIG5V.n7360 ASIG5V.n7359 1.1255
R43838 ASIG5V.n7587 ASIG5V.n7586 1.1255
R43839 ASIG5V.n7589 ASIG5V.n7588 1.1255
R43840 ASIG5V.n7542 ASIG5V.n7541 1.1255
R43841 ASIG5V.n7356 ASIG5V.n7355 1.1255
R43842 ASIG5V.n7546 ASIG5V.n7545 1.1255
R43843 ASIG5V.n7352 ASIG5V.n7351 1.1255
R43844 ASIG5V.n7593 ASIG5V.n7592 1.1255
R43845 ASIG5V.n7348 ASIG5V.n7347 1.1255
R43846 ASIG5V.n7597 ASIG5V.n7596 1.1255
R43847 ASIG5V.n7600 ASIG5V.n7599 1.1255
R43848 ASIG5V.n7344 ASIG5V.n7343 1.1255
R43849 ASIG5V.n7340 ASIG5V.n7339 1.1255
R43850 ASIG5V.n7604 ASIG5V.n7603 1.1255
R43851 ASIG5V.n7336 ASIG5V.n7335 1.1255
R43852 ASIG5V.n7608 ASIG5V.n7607 1.1255
R43853 ASIG5V.n7329 ASIG5V.n7328 1.1255
R43854 ASIG5V.n7332 ASIG5V.n7331 1.1255
R43855 ASIG5V.n7325 ASIG5V.n7324 1.1255
R43856 ASIG5V.n7552 ASIG5V.n7551 1.1255
R43857 ASIG5V.n7321 ASIG5V.n7320 1.1255
R43858 ASIG5V.n7612 ASIG5V.n7611 1.1255
R43859 ASIG5V.n7317 ASIG5V.n7316 1.1255
R43860 ASIG5V.n7616 ASIG5V.n7615 1.1255
R43861 ASIG5V.n7313 ASIG5V.n7312 1.1255
R43862 ASIG5V.n7556 ASIG5V.n7555 1.1255
R43863 ASIG5V.n7309 ASIG5V.n7308 1.1255
R43864 ASIG5V.n7620 ASIG5V.n7619 1.1255
R43865 ASIG5V.n7302 ASIG5V.n7301 1.1255
R43866 ASIG5V.n7305 ASIG5V.n7304 1.1255
R43867 ASIG5V.n7298 ASIG5V.n7297 1.1255
R43868 ASIG5V.n7560 ASIG5V.n7559 1.1255
R43869 ASIG5V.n7294 ASIG5V.n7293 1.1255
R43870 ASIG5V.n7563 ASIG5V.n7562 1.1255
R43871 ASIG5V.n7290 ASIG5V.n7289 1.1255
R43872 ASIG5V.n7624 ASIG5V.n7623 1.1255
R43873 ASIG5V.n7524 ASIG5V.n7523 1.1255
R43874 ASIG5V.n7790 ASIG5V.n7789 1.1255
R43875 ASIG5V.n7792 ASIG5V.n7791 1.1255
R43876 ASIG5V.n7785 ASIG5V.n7784 1.1255
R43877 ASIG5V.n7787 ASIG5V.n7786 1.1255
R43878 ASIG5V.n7780 ASIG5V.n7779 1.1255
R43879 ASIG5V.n7782 ASIG5V.n7781 1.1255
R43880 ASIG5V.n7775 ASIG5V.n7774 1.1255
R43881 ASIG5V.n7777 ASIG5V.n7776 1.1255
R43882 ASIG5V.n7770 ASIG5V.n7769 1.1255
R43883 ASIG5V.n7772 ASIG5V.n7771 1.1255
R43884 ASIG5V.n7765 ASIG5V.n7764 1.1255
R43885 ASIG5V.n7767 ASIG5V.n7766 1.1255
R43886 ASIG5V.n7760 ASIG5V.n7759 1.1255
R43887 ASIG5V.n7762 ASIG5V.n7761 1.1255
R43888 ASIG5V.n7754 ASIG5V.n7753 1.1255
R43889 ASIG5V.n7757 ASIG5V.n7756 1.1255
R43890 ASIG5V.n7748 ASIG5V.n7747 1.1255
R43891 ASIG5V.n7751 ASIG5V.n7750 1.1255
R43892 ASIG5V.n7741 ASIG5V.n7740 1.1255
R43893 ASIG5V.n7744 ASIG5V.n7743 1.1255
R43894 ASIG5V.n7734 ASIG5V.n7733 1.1255
R43895 ASIG5V.n7737 ASIG5V.n7736 1.1255
R43896 ASIG5V.n7727 ASIG5V.n7726 1.1255
R43897 ASIG5V.n7730 ASIG5V.n7729 1.1255
R43898 ASIG5V.n7720 ASIG5V.n7719 1.1255
R43899 ASIG5V.n7723 ASIG5V.n7722 1.1255
R43900 ASIG5V.n7713 ASIG5V.n7712 1.1255
R43901 ASIG5V.n7716 ASIG5V.n7715 1.1255
R43902 ASIG5V.n7706 ASIG5V.n7705 1.1255
R43903 ASIG5V.n7709 ASIG5V.n7708 1.1255
R43904 ASIG5V.n7699 ASIG5V.n7698 1.1255
R43905 ASIG5V.n7702 ASIG5V.n7701 1.1255
R43906 ASIG5V.n7692 ASIG5V.n7691 1.1255
R43907 ASIG5V.n7695 ASIG5V.n7694 1.1255
R43908 ASIG5V.n7685 ASIG5V.n7684 1.1255
R43909 ASIG5V.n7688 ASIG5V.n7687 1.1255
R43910 ASIG5V.n7678 ASIG5V.n7677 1.1255
R43911 ASIG5V.n7681 ASIG5V.n7680 1.1255
R43912 ASIG5V.n7671 ASIG5V.n7670 1.1255
R43913 ASIG5V.n7674 ASIG5V.n7673 1.1255
R43914 ASIG5V.n7664 ASIG5V.n7663 1.1255
R43915 ASIG5V.n7667 ASIG5V.n7666 1.1255
R43916 ASIG5V.n7658 ASIG5V.n7657 1.1255
R43917 ASIG5V.n7660 ASIG5V.n7659 1.1255
R43918 ASIG5V.n7652 ASIG5V.n7651 1.1255
R43919 ASIG5V.n7654 ASIG5V.n7653 1.1255
R43920 ASIG5V.n7647 ASIG5V.n7646 1.1255
R43921 ASIG5V.n7649 ASIG5V.n7648 1.1255
R43922 ASIG5V.n7644 ASIG5V.n7643 1.1255
R43923 ASIG5V.n8097 ASIG5V.n8096 1.1255
R43924 ASIG5V.n12677 ASIG5V.n12676 1.1255
R43925 ASIG5V.n8094 ASIG5V.n8093 1.1255
R43926 ASIG5V.n12680 ASIG5V.n12679 1.1255
R43927 ASIG5V.n12682 ASIG5V.n12681 1.1255
R43928 ASIG5V.n12713 ASIG5V.n12712 1.1255
R43929 ASIG5V.n8090 ASIG5V.n8089 1.1255
R43930 ASIG5V.n12716 ASIG5V.n12715 1.1255
R43931 ASIG5V.n8087 ASIG5V.n8086 1.1255
R43932 ASIG5V.n12685 ASIG5V.n12684 1.1255
R43933 ASIG5V.n8084 ASIG5V.n8083 1.1255
R43934 ASIG5V.n12719 ASIG5V.n12718 1.1255
R43935 ASIG5V.n8081 ASIG5V.n8080 1.1255
R43936 ASIG5V.n12722 ASIG5V.n12721 1.1255
R43937 ASIG5V.n8078 ASIG5V.n8077 1.1255
R43938 ASIG5V.n12689 ASIG5V.n12688 1.1255
R43939 ASIG5V.n8075 ASIG5V.n8074 1.1255
R43940 ASIG5V.n12693 ASIG5V.n12692 1.1255
R43941 ASIG5V.n8068 ASIG5V.n8067 1.1255
R43942 ASIG5V.n8071 ASIG5V.n8070 1.1255
R43943 ASIG5V.n8061 ASIG5V.n8060 1.1255
R43944 ASIG5V.n8064 ASIG5V.n8063 1.1255
R43945 ASIG5V.n8057 ASIG5V.n8056 1.1255
R43946 ASIG5V.n12697 ASIG5V.n12696 1.1255
R43947 ASIG5V.n8053 ASIG5V.n8052 1.1255
R43948 ASIG5V.n12728 ASIG5V.n12727 1.1255
R43949 ASIG5V.n8049 ASIG5V.n8048 1.1255
R43950 ASIG5V.n12732 ASIG5V.n12731 1.1255
R43951 ASIG5V.n8042 ASIG5V.n8041 1.1255
R43952 ASIG5V.n8045 ASIG5V.n8044 1.1255
R43953 ASIG5V.n8035 ASIG5V.n8034 1.1255
R43954 ASIG5V.n8038 ASIG5V.n8037 1.1255
R43955 ASIG5V.n8031 ASIG5V.n8030 1.1255
R43956 ASIG5V.n12736 ASIG5V.n12735 1.1255
R43957 ASIG5V.n8027 ASIG5V.n8026 1.1255
R43958 ASIG5V.n12740 ASIG5V.n12739 1.1255
R43959 ASIG5V.n8020 ASIG5V.n8019 1.1255
R43960 ASIG5V.n8023 ASIG5V.n8022 1.1255
R43961 ASIG5V.n8016 ASIG5V.n8015 1.1255
R43962 ASIG5V.n12744 ASIG5V.n12743 1.1255
R43963 ASIG5V.n8012 ASIG5V.n8011 1.1255
R43964 ASIG5V.n12747 ASIG5V.n12746 1.1255
R43965 ASIG5V.n8006 ASIG5V.n8005 1.1255
R43966 ASIG5V.n8008 ASIG5V.n8007 1.1255
R43967 ASIG5V.n8001 ASIG5V.n8000 1.1255
R43968 ASIG5V.n8003 ASIG5V.n8002 1.1255
R43969 ASIG5V.n7998 ASIG5V.n7997 1.1255
R43970 ASIG5V.n12750 ASIG5V.n12749 1.1255
R43971 ASIG5V.n8127 ASIG5V.n8126 1.1255
R43972 ASIG5V.n12502 ASIG5V.n12501 1.1255
R43973 ASIG5V.n12445 ASIG5V.n12444 1.1255
R43974 ASIG5V.n8172 ASIG5V.n8171 1.1255
R43975 ASIG5V.n12448 ASIG5V.n12447 1.1255
R43976 ASIG5V.n8169 ASIG5V.n8168 1.1255
R43977 ASIG5V.n12505 ASIG5V.n12504 1.1255
R43978 ASIG5V.n12507 ASIG5V.n12506 1.1255
R43979 ASIG5V.n12510 ASIG5V.n12509 1.1255
R43980 ASIG5V.n12512 ASIG5V.n12511 1.1255
R43981 ASIG5V.n12451 ASIG5V.n12450 1.1255
R43982 ASIG5V.n8164 ASIG5V.n8163 1.1255
R43983 ASIG5V.n12515 ASIG5V.n12514 1.1255
R43984 ASIG5V.n12517 ASIG5V.n12516 1.1255
R43985 ASIG5V.n12520 ASIG5V.n12519 1.1255
R43986 ASIG5V.n12522 ASIG5V.n12521 1.1255
R43987 ASIG5V.n12454 ASIG5V.n12453 1.1255
R43988 ASIG5V.n12457 ASIG5V.n12456 1.1255
R43989 ASIG5V.n12461 ASIG5V.n12460 1.1255
R43990 ASIG5V.n8158 ASIG5V.n8157 1.1255
R43991 ASIG5V.n12526 ASIG5V.n12525 1.1255
R43992 ASIG5V.n12529 ASIG5V.n12528 1.1255
R43993 ASIG5V.n12533 ASIG5V.n12532 1.1255
R43994 ASIG5V.n12536 ASIG5V.n12535 1.1255
R43995 ASIG5V.n12465 ASIG5V.n12464 1.1255
R43996 ASIG5V.n8152 ASIG5V.n8151 1.1255
R43997 ASIG5V.n12540 ASIG5V.n12539 1.1255
R43998 ASIG5V.n12543 ASIG5V.n12542 1.1255
R43999 ASIG5V.n12547 ASIG5V.n12546 1.1255
R44000 ASIG5V.n12550 ASIG5V.n12549 1.1255
R44001 ASIG5V.n8147 ASIG5V.n8146 1.1255
R44002 ASIG5V.n8143 ASIG5V.n8142 1.1255
R44003 ASIG5V.n12470 ASIG5V.n12469 1.1255
R44004 ASIG5V.n8139 ASIG5V.n8138 1.1255
R44005 ASIG5V.n12554 ASIG5V.n12553 1.1255
R44006 ASIG5V.n12557 ASIG5V.n12556 1.1255
R44007 ASIG5V.n12561 ASIG5V.n12560 1.1255
R44008 ASIG5V.n12564 ASIG5V.n12563 1.1255
R44009 ASIG5V.n12474 ASIG5V.n12473 1.1255
R44010 ASIG5V.n12476 ASIG5V.n12475 1.1255
R44011 ASIG5V.n12567 ASIG5V.n12566 1.1255
R44012 ASIG5V.n12569 ASIG5V.n12568 1.1255
R44013 ASIG5V.n12572 ASIG5V.n12571 1.1255
R44014 ASIG5V.n12574 ASIG5V.n12573 1.1255
R44015 ASIG5V.n12479 ASIG5V.n12478 1.1255
R44016 ASIG5V.n12481 ASIG5V.n12480 1.1255
R44017 ASIG5V.n12484 ASIG5V.n12483 1.1255
R44018 ASIG5V.n12486 ASIG5V.n12485 1.1255
R44019 ASIG5V.n12577 ASIG5V.n12576 1.1255
R44020 ASIG5V.n8192 ASIG5V.n8191 1.1255
R44021 ASIG5V.n8336 ASIG5V.n8335 1.1255
R44022 ASIG5V.n8338 ASIG5V.n8337 1.1255
R44023 ASIG5V.n8331 ASIG5V.n8330 1.1255
R44024 ASIG5V.n8333 ASIG5V.n8332 1.1255
R44025 ASIG5V.n8326 ASIG5V.n8325 1.1255
R44026 ASIG5V.n8328 ASIG5V.n8327 1.1255
R44027 ASIG5V.n8321 ASIG5V.n8320 1.1255
R44028 ASIG5V.n8323 ASIG5V.n8322 1.1255
R44029 ASIG5V.n8316 ASIG5V.n8315 1.1255
R44030 ASIG5V.n8318 ASIG5V.n8317 1.1255
R44031 ASIG5V.n8311 ASIG5V.n8310 1.1255
R44032 ASIG5V.n8313 ASIG5V.n8312 1.1255
R44033 ASIG5V.n8306 ASIG5V.n8305 1.1255
R44034 ASIG5V.n8308 ASIG5V.n8307 1.1255
R44035 ASIG5V.n8301 ASIG5V.n8300 1.1255
R44036 ASIG5V.n8303 ASIG5V.n8302 1.1255
R44037 ASIG5V.n8295 ASIG5V.n8294 1.1255
R44038 ASIG5V.n8298 ASIG5V.n8297 1.1255
R44039 ASIG5V.n8289 ASIG5V.n8288 1.1255
R44040 ASIG5V.n8292 ASIG5V.n8291 1.1255
R44041 ASIG5V.n8282 ASIG5V.n8281 1.1255
R44042 ASIG5V.n8285 ASIG5V.n8284 1.1255
R44043 ASIG5V.n8275 ASIG5V.n8274 1.1255
R44044 ASIG5V.n8278 ASIG5V.n8277 1.1255
R44045 ASIG5V.n8268 ASIG5V.n8267 1.1255
R44046 ASIG5V.n8271 ASIG5V.n8270 1.1255
R44047 ASIG5V.n8261 ASIG5V.n8260 1.1255
R44048 ASIG5V.n8264 ASIG5V.n8263 1.1255
R44049 ASIG5V.n8254 ASIG5V.n8253 1.1255
R44050 ASIG5V.n8257 ASIG5V.n8256 1.1255
R44051 ASIG5V.n8247 ASIG5V.n8246 1.1255
R44052 ASIG5V.n8250 ASIG5V.n8249 1.1255
R44053 ASIG5V.n8240 ASIG5V.n8239 1.1255
R44054 ASIG5V.n8243 ASIG5V.n8242 1.1255
R44055 ASIG5V.n8233 ASIG5V.n8232 1.1255
R44056 ASIG5V.n8236 ASIG5V.n8235 1.1255
R44057 ASIG5V.n8227 ASIG5V.n8226 1.1255
R44058 ASIG5V.n8229 ASIG5V.n8228 1.1255
R44059 ASIG5V.n8222 ASIG5V.n8221 1.1255
R44060 ASIG5V.n8224 ASIG5V.n8223 1.1255
R44061 ASIG5V.n8217 ASIG5V.n8216 1.1255
R44062 ASIG5V.n8219 ASIG5V.n8218 1.1255
R44063 ASIG5V.n8212 ASIG5V.n8211 1.1255
R44064 ASIG5V.n8214 ASIG5V.n8213 1.1255
R44065 ASIG5V.n8207 ASIG5V.n8206 1.1255
R44066 ASIG5V.n8209 ASIG5V.n8208 1.1255
R44067 ASIG5V.n8202 ASIG5V.n8201 1.1255
R44068 ASIG5V.n8204 ASIG5V.n8203 1.1255
R44069 ASIG5V.n8199 ASIG5V.n8198 1.1255
R44070 ASIG5V.n8467 ASIG5V.n8466 1.1255
R44071 ASIG5V.n8469 ASIG5V.n8468 1.1255
R44072 ASIG5V.n8464 ASIG5V.n8463 1.1255
R44073 ASIG5V.n12172 ASIG5V.n12171 1.1255
R44074 ASIG5V.n8461 ASIG5V.n8460 1.1255
R44075 ASIG5V.n12204 ASIG5V.n12203 1.1255
R44076 ASIG5V.n8456 ASIG5V.n8455 1.1255
R44077 ASIG5V.n8458 ASIG5V.n8457 1.1255
R44078 ASIG5V.n8453 ASIG5V.n8452 1.1255
R44079 ASIG5V.n12175 ASIG5V.n12174 1.1255
R44080 ASIG5V.n8448 ASIG5V.n8447 1.1255
R44081 ASIG5V.n8450 ASIG5V.n8449 1.1255
R44082 ASIG5V.n8445 ASIG5V.n8444 1.1255
R44083 ASIG5V.n12209 ASIG5V.n12208 1.1255
R44084 ASIG5V.n8442 ASIG5V.n8441 1.1255
R44085 ASIG5V.n12178 ASIG5V.n12177 1.1255
R44086 ASIG5V.n8439 ASIG5V.n8438 1.1255
R44087 ASIG5V.n12181 ASIG5V.n12180 1.1255
R44088 ASIG5V.n8436 ASIG5V.n8435 1.1255
R44089 ASIG5V.n12213 ASIG5V.n12212 1.1255
R44090 ASIG5V.n8430 ASIG5V.n8429 1.1255
R44091 ASIG5V.n8433 ASIG5V.n8432 1.1255
R44092 ASIG5V.n8423 ASIG5V.n8422 1.1255
R44093 ASIG5V.n8426 ASIG5V.n8425 1.1255
R44094 ASIG5V.n8419 ASIG5V.n8418 1.1255
R44095 ASIG5V.n12218 ASIG5V.n12217 1.1255
R44096 ASIG5V.n8415 ASIG5V.n8414 1.1255
R44097 ASIG5V.n12222 ASIG5V.n12221 1.1255
R44098 ASIG5V.n8411 ASIG5V.n8410 1.1255
R44099 ASIG5V.n12186 ASIG5V.n12185 1.1255
R44100 ASIG5V.n8404 ASIG5V.n8403 1.1255
R44101 ASIG5V.n8407 ASIG5V.n8406 1.1255
R44102 ASIG5V.n8400 ASIG5V.n8399 1.1255
R44103 ASIG5V.n12226 ASIG5V.n12225 1.1255
R44104 ASIG5V.n8396 ASIG5V.n8395 1.1255
R44105 ASIG5V.n12229 ASIG5V.n12228 1.1255
R44106 ASIG5V.n8393 ASIG5V.n8392 1.1255
R44107 ASIG5V.n12190 ASIG5V.n12189 1.1255
R44108 ASIG5V.n8388 ASIG5V.n8387 1.1255
R44109 ASIG5V.n8390 ASIG5V.n8389 1.1255
R44110 ASIG5V.n8385 ASIG5V.n8384 1.1255
R44111 ASIG5V.n12233 ASIG5V.n12232 1.1255
R44112 ASIG5V.n8380 ASIG5V.n8379 1.1255
R44113 ASIG5V.n8382 ASIG5V.n8381 1.1255
R44114 ASIG5V.n8375 ASIG5V.n8374 1.1255
R44115 ASIG5V.n8377 ASIG5V.n8376 1.1255
R44116 ASIG5V.n8372 ASIG5V.n8371 1.1255
R44117 ASIG5V.n12236 ASIG5V.n12235 1.1255
R44118 ASIG5V.n8590 ASIG5V.n8589 1.1255
R44119 ASIG5V.n12017 ASIG5V.n12016 1.1255
R44120 ASIG5V.n8587 ASIG5V.n8586 1.1255
R44121 ASIG5V.n12020 ASIG5V.n12019 1.1255
R44122 ASIG5V.n8584 ASIG5V.n8583 1.1255
R44123 ASIG5V.n12051 ASIG5V.n12050 1.1255
R44124 ASIG5V.n8579 ASIG5V.n8578 1.1255
R44125 ASIG5V.n8581 ASIG5V.n8580 1.1255
R44126 ASIG5V.n8574 ASIG5V.n8573 1.1255
R44127 ASIG5V.n8576 ASIG5V.n8575 1.1255
R44128 ASIG5V.n8571 ASIG5V.n8570 1.1255
R44129 ASIG5V.n12055 ASIG5V.n12054 1.1255
R44130 ASIG5V.n8566 ASIG5V.n8565 1.1255
R44131 ASIG5V.n8568 ASIG5V.n8567 1.1255
R44132 ASIG5V.n8563 ASIG5V.n8562 1.1255
R44133 ASIG5V.n12024 ASIG5V.n12023 1.1255
R44134 ASIG5V.n8560 ASIG5V.n8559 1.1255
R44135 ASIG5V.n12027 ASIG5V.n12026 1.1255
R44136 ASIG5V.n8557 ASIG5V.n8556 1.1255
R44137 ASIG5V.n12059 ASIG5V.n12058 1.1255
R44138 ASIG5V.n8554 ASIG5V.n8553 1.1255
R44139 ASIG5V.n12063 ASIG5V.n12062 1.1255
R44140 ASIG5V.n8547 ASIG5V.n8546 1.1255
R44141 ASIG5V.n8550 ASIG5V.n8549 1.1255
R44142 ASIG5V.n8543 ASIG5V.n8542 1.1255
R44143 ASIG5V.n12067 ASIG5V.n12066 1.1255
R44144 ASIG5V.n8539 ASIG5V.n8538 1.1255
R44145 ASIG5V.n12071 ASIG5V.n12070 1.1255
R44146 ASIG5V.n8532 ASIG5V.n8531 1.1255
R44147 ASIG5V.n8535 ASIG5V.n8534 1.1255
R44148 ASIG5V.n8528 ASIG5V.n8527 1.1255
R44149 ASIG5V.n12032 ASIG5V.n12031 1.1255
R44150 ASIG5V.n8524 ASIG5V.n8523 1.1255
R44151 ASIG5V.n12074 ASIG5V.n12073 1.1255
R44152 ASIG5V.n8519 ASIG5V.n8518 1.1255
R44153 ASIG5V.n8521 ASIG5V.n8520 1.1255
R44154 ASIG5V.n8516 ASIG5V.n8515 1.1255
R44155 ASIG5V.n12035 ASIG5V.n12034 1.1255
R44156 ASIG5V.n8513 ASIG5V.n8512 1.1255
R44157 ASIG5V.n12078 ASIG5V.n12077 1.1255
R44158 ASIG5V.n8508 ASIG5V.n8507 1.1255
R44159 ASIG5V.n8510 ASIG5V.n8509 1.1255
R44160 ASIG5V.n8505 ASIG5V.n8504 1.1255
R44161 ASIG5V.n12038 ASIG5V.n12037 1.1255
R44162 ASIG5V.n8500 ASIG5V.n8499 1.1255
R44163 ASIG5V.n8502 ASIG5V.n8501 1.1255
R44164 ASIG5V.n8496 ASIG5V.n8495 1.1255
R44165 ASIG5V.n8692 ASIG5V.n8691 1.1255
R44166 ASIG5V.n11850 ASIG5V.n11849 1.1255
R44167 ASIG5V.n8689 ASIG5V.n8688 1.1255
R44168 ASIG5V.n11853 ASIG5V.n11852 1.1255
R44169 ASIG5V.n8686 ASIG5V.n8685 1.1255
R44170 ASIG5V.n11887 ASIG5V.n11886 1.1255
R44171 ASIG5V.n8683 ASIG5V.n8682 1.1255
R44172 ASIG5V.n11890 ASIG5V.n11889 1.1255
R44173 ASIG5V.n8680 ASIG5V.n8679 1.1255
R44174 ASIG5V.n11856 ASIG5V.n11855 1.1255
R44175 ASIG5V.n8677 ASIG5V.n8676 1.1255
R44176 ASIG5V.n11893 ASIG5V.n11892 1.1255
R44177 ASIG5V.n8674 ASIG5V.n8673 1.1255
R44178 ASIG5V.n11896 ASIG5V.n11895 1.1255
R44179 ASIG5V.n8671 ASIG5V.n8670 1.1255
R44180 ASIG5V.n11859 ASIG5V.n11858 1.1255
R44181 ASIG5V.n8666 ASIG5V.n8665 1.1255
R44182 ASIG5V.n8668 ASIG5V.n8667 1.1255
R44183 ASIG5V.n8661 ASIG5V.n8660 1.1255
R44184 ASIG5V.n8663 ASIG5V.n8662 1.1255
R44185 ASIG5V.n8658 ASIG5V.n8657 1.1255
R44186 ASIG5V.n11900 ASIG5V.n11899 1.1255
R44187 ASIG5V.n8655 ASIG5V.n8654 1.1255
R44188 ASIG5V.n11864 ASIG5V.n11863 1.1255
R44189 ASIG5V.n8651 ASIG5V.n8650 1.1255
R44190 ASIG5V.n11904 ASIG5V.n11903 1.1255
R44191 ASIG5V.n8647 ASIG5V.n8646 1.1255
R44192 ASIG5V.n11908 ASIG5V.n11907 1.1255
R44193 ASIG5V.n8643 ASIG5V.n8642 1.1255
R44194 ASIG5V.n11867 ASIG5V.n11866 1.1255
R44195 ASIG5V.n8639 ASIG5V.n8638 1.1255
R44196 ASIG5V.n11870 ASIG5V.n11869 1.1255
R44197 ASIG5V.n8636 ASIG5V.n8635 1.1255
R44198 ASIG5V.n11911 ASIG5V.n11910 1.1255
R44199 ASIG5V.n8633 ASIG5V.n8632 1.1255
R44200 ASIG5V.n11914 ASIG5V.n11913 1.1255
R44201 ASIG5V.n11916 ASIG5V.n11915 1.1255
R44202 ASIG5V.n11873 ASIG5V.n11872 1.1255
R44203 ASIG5V.n8629 ASIG5V.n8628 1.1255
R44204 ASIG5V.n11919 ASIG5V.n11918 1.1255
R44205 ASIG5V.n8626 ASIG5V.n8625 1.1255
R44206 ASIG5V.n11922 ASIG5V.n11921 1.1255
R44207 ASIG5V.n8623 ASIG5V.n8622 1.1255
R44208 ASIG5V.n11876 ASIG5V.n11875 1.1255
R44209 ASIG5V.n8619 ASIG5V.n8618 1.1255
R44210 ASIG5V.n8795 ASIG5V.n8794 1.1255
R44211 ASIG5V.n11684 ASIG5V.n11683 1.1255
R44212 ASIG5V.n8790 ASIG5V.n8789 1.1255
R44213 ASIG5V.n8792 ASIG5V.n8791 1.1255
R44214 ASIG5V.n8787 ASIG5V.n8786 1.1255
R44215 ASIG5V.n11724 ASIG5V.n11723 1.1255
R44216 ASIG5V.n8784 ASIG5V.n8783 1.1255
R44217 ASIG5V.n11727 ASIG5V.n11726 1.1255
R44218 ASIG5V.n8781 ASIG5V.n8780 1.1255
R44219 ASIG5V.n11688 ASIG5V.n11687 1.1255
R44220 ASIG5V.n8778 ASIG5V.n8777 1.1255
R44221 ASIG5V.n11730 ASIG5V.n11729 1.1255
R44222 ASIG5V.n8775 ASIG5V.n8774 1.1255
R44223 ASIG5V.n11733 ASIG5V.n11732 1.1255
R44224 ASIG5V.n8772 ASIG5V.n8771 1.1255
R44225 ASIG5V.n11691 ASIG5V.n11690 1.1255
R44226 ASIG5V.n8769 ASIG5V.n8768 1.1255
R44227 ASIG5V.n11694 ASIG5V.n11693 1.1255
R44228 ASIG5V.n8766 ASIG5V.n8765 1.1255
R44229 ASIG5V.n11736 ASIG5V.n11735 1.1255
R44230 ASIG5V.n8761 ASIG5V.n8760 1.1255
R44231 ASIG5V.n8763 ASIG5V.n8762 1.1255
R44232 ASIG5V.n8758 ASIG5V.n8757 1.1255
R44233 ASIG5V.n11698 ASIG5V.n11697 1.1255
R44234 ASIG5V.n8755 ASIG5V.n8754 1.1255
R44235 ASIG5V.n11741 ASIG5V.n11740 1.1255
R44236 ASIG5V.n8751 ASIG5V.n8750 1.1255
R44237 ASIG5V.n11744 ASIG5V.n11743 1.1255
R44238 ASIG5V.n8748 ASIG5V.n8747 1.1255
R44239 ASIG5V.n11701 ASIG5V.n11700 1.1255
R44240 ASIG5V.n8745 ASIG5V.n8744 1.1255
R44241 ASIG5V.n11704 ASIG5V.n11703 1.1255
R44242 ASIG5V.n8742 ASIG5V.n8741 1.1255
R44243 ASIG5V.n11747 ASIG5V.n11746 1.1255
R44244 ASIG5V.n8739 ASIG5V.n8738 1.1255
R44245 ASIG5V.n11750 ASIG5V.n11749 1.1255
R44246 ASIG5V.n8736 ASIG5V.n8735 1.1255
R44247 ASIG5V.n11707 ASIG5V.n11706 1.1255
R44248 ASIG5V.n8733 ASIG5V.n8732 1.1255
R44249 ASIG5V.n11753 ASIG5V.n11752 1.1255
R44250 ASIG5V.n8730 ASIG5V.n8729 1.1255
R44251 ASIG5V.n11756 ASIG5V.n11755 1.1255
R44252 ASIG5V.n8727 ASIG5V.n8726 1.1255
R44253 ASIG5V.n11505 ASIG5V.n11504 1.1255
R44254 ASIG5V.n11507 ASIG5V.n11506 1.1255
R44255 ASIG5V.n11510 ASIG5V.n11509 1.1255
R44256 ASIG5V.n11512 ASIG5V.n11511 1.1255
R44257 ASIG5V.n11571 ASIG5V.n11570 1.1255
R44258 ASIG5V.n11573 ASIG5V.n11572 1.1255
R44259 ASIG5V.n11576 ASIG5V.n11575 1.1255
R44260 ASIG5V.n11578 ASIG5V.n11577 1.1255
R44261 ASIG5V.n11515 ASIG5V.n11514 1.1255
R44262 ASIG5V.n11517 ASIG5V.n11516 1.1255
R44263 ASIG5V.n11581 ASIG5V.n11580 1.1255
R44264 ASIG5V.n11583 ASIG5V.n11582 1.1255
R44265 ASIG5V.n11586 ASIG5V.n11585 1.1255
R44266 ASIG5V.n11588 ASIG5V.n11587 1.1255
R44267 ASIG5V.n11520 ASIG5V.n11519 1.1255
R44268 ASIG5V.n11522 ASIG5V.n11521 1.1255
R44269 ASIG5V.n11525 ASIG5V.n11524 1.1255
R44270 ASIG5V.n11527 ASIG5V.n11526 1.1255
R44271 ASIG5V.n11591 ASIG5V.n11590 1.1255
R44272 ASIG5V.n11593 ASIG5V.n11592 1.1255
R44273 ASIG5V.n11596 ASIG5V.n11595 1.1255
R44274 ASIG5V.n11598 ASIG5V.n11597 1.1255
R44275 ASIG5V.n11530 ASIG5V.n11529 1.1255
R44276 ASIG5V.n11532 ASIG5V.n11531 1.1255
R44277 ASIG5V.n11601 ASIG5V.n11600 1.1255
R44278 ASIG5V.n11603 ASIG5V.n11602 1.1255
R44279 ASIG5V.n11606 ASIG5V.n11605 1.1255
R44280 ASIG5V.n11608 ASIG5V.n11607 1.1255
R44281 ASIG5V.n11535 ASIG5V.n11534 1.1255
R44282 ASIG5V.n11537 ASIG5V.n11536 1.1255
R44283 ASIG5V.n11540 ASIG5V.n11539 1.1255
R44284 ASIG5V.n11542 ASIG5V.n11541 1.1255
R44285 ASIG5V.n11611 ASIG5V.n11610 1.1255
R44286 ASIG5V.n11613 ASIG5V.n11612 1.1255
R44287 ASIG5V.n11616 ASIG5V.n11615 1.1255
R44288 ASIG5V.n11618 ASIG5V.n11617 1.1255
R44289 ASIG5V.n11545 ASIG5V.n11544 1.1255
R44290 ASIG5V.n11547 ASIG5V.n11546 1.1255
R44291 ASIG5V.n11621 ASIG5V.n11620 1.1255
R44292 ASIG5V.n11623 ASIG5V.n11622 1.1255
R44293 ASIG5V.n12423 ASIG5V.n12422 1.1255
R44294 ASIG5V.n8187 ASIG5V.n8186 1.1255
R44295 ASIG5V.n8189 ASIG5V.n8188 1.1255
R44296 ASIG5V.n8194 ASIG5V.n8193 1.1255
R44297 ASIG5V.n8122 ASIG5V.n8121 1.1255
R44298 ASIG5V.n8124 ASIG5V.n8123 1.1255
R44299 ASIG5V.n8118 ASIG5V.n8117 1.1255
R44300 ASIG5V.n7819 ASIG5V.n7818 1.1255
R44301 ASIG5V.n7943 ASIG5V.n7942 1.1255
R44302 ASIG5V.n7821 ASIG5V.n7820 1.1255
R44303 ASIG5V.n7397 ASIG5V.n7396 1.1255
R44304 ASIG5V.n7521 ASIG5V.n7520 1.1255
R44305 ASIG5V.n7399 ASIG5V.n7398 1.1255
R44306 ASIG5V.n141 ASIG5V.n140 1.1255
R44307 ASIG5V.n143 ASIG5V.n142 1.1255
R44308 ASIG5V.n148 ASIG5V.n147 1.1255
R44309 ASIG5V.n100 ASIG5V.n99 1.1255
R44310 ASIG5V.n102 ASIG5V.n101 1.1255
R44311 ASIG5V.n105 ASIG5V.n104 1.1255
R44312 ASIG5V.n6772 ASIG5V.n6771 1.1255
R44313 ASIG5V.n6547 ASIG5V.n6546 1.1255
R44314 ASIG5V.n6775 ASIG5V.n6774 1.1255
R44315 ASIG5V.n6417 ASIG5V.n6416 1.1255
R44316 ASIG5V.n7050 ASIG5V.n7049 1.1255
R44317 ASIG5V.n6322 ASIG5V.n6321 1.1255
R44318 ASIG5V.n6333 ASIG5V.n6332 1.1255
R44319 ASIG5V.n6324 ASIG5V.n6323 1.1255
R44320 ASIG5V.n5974 ASIG5V.n5973 1.1255
R44321 ASIG5V.n5976 ASIG5V.n5975 1.1255
R44322 ASIG5V.n5981 ASIG5V.n5980 1.1255
R44323 ASIG5V.n5678 ASIG5V.n5677 1.1255
R44324 ASIG5V.n5680 ASIG5V.n5679 1.1255
R44325 ASIG5V.n5685 ASIG5V.n5684 1.1255
R44326 ASIG5V.n5324 ASIG5V.n5323 1.1255
R44327 ASIG5V.n5400 ASIG5V.n5399 1.1255
R44328 ASIG5V.n5326 ASIG5V.n5325 1.1255
R44329 ASIG5V.n4973 ASIG5V.n4972 1.1255
R44330 ASIG5V.n4975 ASIG5V.n4974 1.1255
R44331 ASIG5V.n4980 ASIG5V.n4979 1.1255
R44332 ASIG5V.n4705 ASIG5V.n4704 1.1255
R44333 ASIG5V.n1068 ASIG5V.n1067 1.1255
R44334 ASIG5V.n2823 ASIG5V.n2822 1.1255
R44335 ASIG5V.n2883 ASIG5V.n2882 1.1255
R44336 ASIG5V.n3034 ASIG5V.n3033 1.1255
R44337 ASIG5V.n3038 ASIG5V.n3037 1.1255
R44338 ASIG5V.n3139 ASIG5V.n3138 1.1255
R44339 ASIG5V.n3255 ASIG5V.n3254 1.1255
R44340 ASIG5V.n3259 ASIG5V.n3258 1.1255
R44341 ASIG5V.n3299 ASIG5V.n3298 1.1255
R44342 ASIG5V.n3477 ASIG5V.n3476 1.1255
R44343 ASIG5V.n3481 ASIG5V.n3480 1.1255
R44344 ASIG5V.n3626 ASIG5V.n3625 1.1255
R44345 ASIG5V.n3742 ASIG5V.n3741 1.1255
R44346 ASIG5V.n3747 ASIG5V.n3746 1.1255
R44347 ASIG5V.n3899 ASIG5V.n3898 1.1255
R44348 ASIG5V.n4009 ASIG5V.n4008 1.1255
R44349 ASIG5V.n4099 ASIG5V.n4098 1.1255
R44350 ASIG5V.n4279 ASIG5V.n4278 1.1255
R44351 ASIG5V.n4287 ASIG5V.n4286 1.1255
R44352 ASIG5V.n4443 ASIG5V.n4442 1.1255
R44353 ASIG5V.n4563 ASIG5V.n4562 1.1255
R44354 ASIG5V.n4568 ASIG5V.n4567 1.1255
R44355 ASIG5V.n4633 ASIG5V.n4632 1.1255
R44356 ASIG5V.n4849 ASIG5V.n4848 1.1255
R44357 ASIG5V.n4854 ASIG5V.n4853 1.1255
R44358 ASIG5V.n4971 ASIG5V.n4970 1.1255
R44359 ASIG5V.n5148 ASIG5V.n5147 1.1255
R44360 ASIG5V.n5154 ASIG5V.n5153 1.1255
R44361 ASIG5V.n5398 ASIG5V.n5397 1.1255
R44362 ASIG5V.n5448 ASIG5V.n5447 1.1255
R44363 ASIG5V.n5455 ASIG5V.n5454 1.1255
R44364 ASIG5V.n5676 ASIG5V.n5675 1.1255
R44365 ASIG5V.n5804 ASIG5V.n5803 1.1255
R44366 ASIG5V.n5860 ASIG5V.n5859 1.1255
R44367 ASIG5V.n6152 ASIG5V.n6151 1.1255
R44368 ASIG5V.n6159 ASIG5V.n6158 1.1255
R44369 ASIG5V.n6331 ASIG5V.n6330 1.1255
R44370 ASIG5V.n7066 ASIG5V.n7065 1.1255
R44371 ASIG5V.n7059 ASIG5V.n7058 1.1255
R44372 ASIG5V.n6935 ASIG5V.n6934 1.1255
R44373 ASIG5V.n6787 ASIG5V.n6786 1.1255
R44374 ASIG5V.n6780 ASIG5V.n6779 1.1255
R44375 ASIG5V.n6657 ASIG5V.n6656 1.1255
R44376 ASIG5V.n6552 ASIG5V.n6551 1.1255
R44377 ASIG5V.n13621 ASIG5V.n13620 1.1255
R44378 ASIG5V.n13612 ASIG5V.n13611 1.1255
R44379 ASIG5V.n13367 ASIG5V.n13366 1.1255
R44380 ASIG5V.n13358 ASIG5V.n13357 1.1255
R44381 ASIG5V.n7274 ASIG5V.n7273 1.1255
R44382 ASIG5V.n7281 ASIG5V.n7280 1.1255
R44383 ASIG5V.n7406 ASIG5V.n7405 1.1255
R44384 ASIG5V.n7629 ASIG5V.n7628 1.1255
R44385 ASIG5V.n7636 ASIG5V.n7635 1.1255
R44386 ASIG5V.n7941 ASIG5V.n7940 1.1255
R44387 ASIG5V.n7986 ASIG5V.n7985 1.1255
R44388 ASIG5V.n7993 ASIG5V.n7992 1.1255
R44389 ASIG5V.n12757 ASIG5V.n12756 1.1255
R44390 ASIG5V.n12665 ASIG5V.n12664 1.1255
R44391 ASIG5V.n12659 ASIG5V.n12658 1.1255
R44392 ASIG5V.n12651 ASIG5V.n12650 1.1255
R44393 ASIG5V.n12432 ASIG5V.n12431 1.1255
R44394 ASIG5V.n12427 ASIG5V.n12426 1.1255
R44395 ASIG5V.n12355 ASIG5V.n12354 1.1255
R44396 ASIG5V.n12315 ASIG5V.n12314 1.1255
R44397 ASIG5V.n12306 ASIG5V.n12305 1.1255
R44398 ASIG5V.n12164 ASIG5V.n12163 1.1255
R44399 ASIG5V.n12159 ASIG5V.n12158 1.1255
R44400 ASIG5V.n12085 ASIG5V.n12084 1.1255
R44401 ASIG5V.n12006 ASIG5V.n12005 1.1255
R44402 ASIG5V.n12001 ASIG5V.n12000 1.1255
R44403 ASIG5V.n11962 ASIG5V.n11961 1.1255
R44404 ASIG5V.n11841 ASIG5V.n11840 1.1255
R44405 ASIG5V.n11836 ASIG5V.n11835 1.1255
R44406 ASIG5V.n11763 ASIG5V.n11762 1.1255
R44407 ASIG5V.n11674 ASIG5V.n11673 1.1255
R44408 ASIG5V.n11670 ASIG5V.n11669 1.1255
R44409 ASIG5V.n11634 ASIG5V.n11633 1.1255
R44410 ASIG5V.n11490 ASIG5V.n11489 1.1255
R44411 ASIG5V.n11419 ASIG5V.n11418 1.1255
R44412 ASIG5V.n11319 ASIG5V.n11318 1.1255
R44413 ASIG5V.n11313 ASIG5V.n11312 1.1255
R44414 ASIG5V.n11157 ASIG5V.n11156 1.1255
R44415 ASIG5V.n11104 ASIG5V.n11103 1.1255
R44416 ASIG5V.n11100 ASIG5V.n11099 1.1255
R44417 ASIG5V.n9433 ASIG5V.n9432 1.1255
R44418 ASIG5V.n11292 ASIG5V.n11291 1.1255
R44419 ASIG5V.n11289 ASIG5V.n11288 1.1255
R44420 ASIG5V.n11287 ASIG5V.n11286 1.1255
R44421 ASIG5V.n11284 ASIG5V.n11283 1.1255
R44422 ASIG5V.n11282 ASIG5V.n11281 1.1255
R44423 ASIG5V.n11279 ASIG5V.n11278 1.1255
R44424 ASIG5V.n11277 ASIG5V.n11276 1.1255
R44425 ASIG5V.n11274 ASIG5V.n11273 1.1255
R44426 ASIG5V.n11272 ASIG5V.n11271 1.1255
R44427 ASIG5V.n11269 ASIG5V.n11268 1.1255
R44428 ASIG5V.n11267 ASIG5V.n11266 1.1255
R44429 ASIG5V.n11264 ASIG5V.n11263 1.1255
R44430 ASIG5V.n11136 ASIG5V.n11135 1.1255
R44431 ASIG5V.n11261 ASIG5V.n11260 1.1255
R44432 ASIG5V.n11259 ASIG5V.n11258 1.1255
R44433 ASIG5V.n11256 ASIG5V.n11255 1.1255
R44434 ASIG5V.n11254 ASIG5V.n11253 1.1255
R44435 ASIG5V.n11251 ASIG5V.n11250 1.1255
R44436 ASIG5V.n11249 ASIG5V.n11248 1.1255
R44437 ASIG5V.n11131 ASIG5V.n11130 1.1255
R44438 ASIG5V.n11128 ASIG5V.n11127 1.1255
R44439 ASIG5V.n11245 ASIG5V.n11244 1.1255
R44440 ASIG5V.n11243 ASIG5V.n11242 1.1255
R44441 ASIG5V.n11240 ASIG5V.n11239 1.1255
R44442 ASIG5V.n11238 ASIG5V.n11237 1.1255
R44443 ASIG5V.n11235 ASIG5V.n11234 1.1255
R44444 ASIG5V.n11233 ASIG5V.n11232 1.1255
R44445 ASIG5V.n11230 ASIG5V.n11229 1.1255
R44446 ASIG5V.n11228 ASIG5V.n11227 1.1255
R44447 ASIG5V.n11225 ASIG5V.n11224 1.1255
R44448 ASIG5V.n11223 ASIG5V.n11222 1.1255
R44449 ASIG5V.n11220 ASIG5V.n11219 1.1255
R44450 ASIG5V.n11218 ASIG5V.n11217 1.1255
R44451 ASIG5V.n11215 ASIG5V.n11214 1.1255
R44452 ASIG5V.n4970 ASIG5V.n4969 1.1255
R44453 ASIG5V.n5147 ASIG5V.n5146 1.1255
R44454 ASIG5V.n5153 ASIG5V.n5152 1.1255
R44455 ASIG5V.n5397 ASIG5V.n5396 1.1255
R44456 ASIG5V.n5447 ASIG5V.n5446 1.1255
R44457 ASIG5V.n5454 ASIG5V.n5453 1.1255
R44458 ASIG5V.n5675 ASIG5V.n5674 1.1255
R44459 ASIG5V.n5803 ASIG5V.n5802 1.1255
R44460 ASIG5V.n5859 ASIG5V.n5858 1.1255
R44461 ASIG5V.n6151 ASIG5V.n6150 1.1255
R44462 ASIG5V.n6158 ASIG5V.n6157 1.1255
R44463 ASIG5V.n6330 ASIG5V.n6329 1.1255
R44464 ASIG5V.n7065 ASIG5V.n7064 1.1255
R44465 ASIG5V.n7058 ASIG5V.n7057 1.1255
R44466 ASIG5V.n6934 ASIG5V.n6933 1.1255
R44467 ASIG5V.n6786 ASIG5V.n6785 1.1255
R44468 ASIG5V.n6779 ASIG5V.n6778 1.1255
R44469 ASIG5V.n6656 ASIG5V.n6655 1.1255
R44470 ASIG5V.n6551 ASIG5V.n6550 1.1255
R44471 ASIG5V.n13620 ASIG5V.n13619 1.1255
R44472 ASIG5V.n13611 ASIG5V.n13610 1.1255
R44473 ASIG5V.n13366 ASIG5V.n13365 1.1255
R44474 ASIG5V.n13357 ASIG5V.n13356 1.1255
R44475 ASIG5V.n7273 ASIG5V.n7272 1.1255
R44476 ASIG5V.n7280 ASIG5V.n7279 1.1255
R44477 ASIG5V.n7405 ASIG5V.n7404 1.1255
R44478 ASIG5V.n7628 ASIG5V.n7627 1.1255
R44479 ASIG5V.n7635 ASIG5V.n7634 1.1255
R44480 ASIG5V.n7940 ASIG5V.n7939 1.1255
R44481 ASIG5V.n7985 ASIG5V.n7984 1.1255
R44482 ASIG5V.n7992 ASIG5V.n7991 1.1255
R44483 ASIG5V.n12756 ASIG5V.n12755 1.1255
R44484 ASIG5V.n12664 ASIG5V.n12663 1.1255
R44485 ASIG5V.n12658 ASIG5V.n12657 1.1255
R44486 ASIG5V.n12650 ASIG5V.n12649 1.1255
R44487 ASIG5V.n2937 ASIG5V.n2936 1.1255
R44488 ASIG5V.n2940 ASIG5V.n2939 1.1255
R44489 ASIG5V.n2867 ASIG5V.n2866 1.1255
R44490 ASIG5V.n2943 ASIG5V.n2942 1.1255
R44491 ASIG5V.n2945 ASIG5V.n2944 1.1255
R44492 ASIG5V.n2948 ASIG5V.n2947 1.1255
R44493 ASIG5V.n2863 ASIG5V.n2862 1.1255
R44494 ASIG5V.n2951 ASIG5V.n2950 1.1255
R44495 ASIG5V.n2860 ASIG5V.n2859 1.1255
R44496 ASIG5V.n2954 ASIG5V.n2953 1.1255
R44497 ASIG5V.n2956 ASIG5V.n2955 1.1255
R44498 ASIG5V.n2959 ASIG5V.n2958 1.1255
R44499 ASIG5V.n2961 ASIG5V.n2960 1.1255
R44500 ASIG5V.n2964 ASIG5V.n2963 1.1255
R44501 ASIG5V.n2966 ASIG5V.n2965 1.1255
R44502 ASIG5V.n2969 ASIG5V.n2968 1.1255
R44503 ASIG5V.n2971 ASIG5V.n2970 1.1255
R44504 ASIG5V.n2854 ASIG5V.n2853 1.1255
R44505 ASIG5V.n2974 ASIG5V.n2973 1.1255
R44506 ASIG5V.n2977 ASIG5V.n2976 1.1255
R44507 ASIG5V.n2850 ASIG5V.n2849 1.1255
R44508 ASIG5V.n2980 ASIG5V.n2979 1.1255
R44509 ASIG5V.n2982 ASIG5V.n2981 1.1255
R44510 ASIG5V.n2985 ASIG5V.n2984 1.1255
R44511 ASIG5V.n2987 ASIG5V.n2986 1.1255
R44512 ASIG5V.n2990 ASIG5V.n2989 1.1255
R44513 ASIG5V.n2845 ASIG5V.n2844 1.1255
R44514 ASIG5V.n2993 ASIG5V.n2992 1.1255
R44515 ASIG5V.n2995 ASIG5V.n2994 1.1255
R44516 ASIG5V.n2998 ASIG5V.n2997 1.1255
R44517 ASIG5V.n3000 ASIG5V.n2999 1.1255
R44518 ASIG5V.n3003 ASIG5V.n3002 1.1255
R44519 ASIG5V.n2840 ASIG5V.n2839 1.1255
R44520 ASIG5V.n8975 ASIG5V.n8878 1.12271
R44521 ASIG5V.n621 ASIG5V.n521 1.12271
R44522 ASIG5V.n744 ASIG5V.n743 1.12271
R44523 ASIG5V.n9116 ASIG5V.n8986 1.12271
R44524 ASIG5V.n8981 ASIG5V.n8980 1.12271
R44525 ASIG5V.n8975 ASIG5V.n8974 1.12271
R44526 ASIG5V.n9116 ASIG5V.n8874 1.12271
R44527 ASIG5V.n621 ASIG5V.n620 1.12271
R44528 ASIG5V.n627 ASIG5V.n626 1.12271
R44529 ASIG5V.n741 ASIG5V.n740 1.12271
R44530 ASIG5V.n9116 ASIG5V.n9115 1.12271
R44531 ASIG5V.n3104 ASIG5V.n3103 1.11687
R44532 ASIG5V.n3558 ASIG5V.n3557 1.11687
R44533 ASIG5V.n3833 ASIG5V.n3832 1.11687
R44534 ASIG5V.n4096 ASIG5V.n4095 1.11687
R44535 ASIG5V.n4375 ASIG5V.n4374 1.11687
R44536 ASIG5V.n4630 ASIG5V.n4629 1.11687
R44537 ASIG5V.n4901 ASIG5V.n4900 1.11687
R44538 ASIG5V.n5328 ASIG5V.n5327 1.11687
R44539 ASIG5V.n5559 ASIG5V.n5558 1.11687
R44540 ASIG5V.n5855 ASIG5V.n5854 1.11687
R44541 ASIG5V.n6326 ASIG5V.n6325 1.11687
R44542 ASIG5V.n7052 ASIG5V.n7051 1.11687
R44543 ASIG5V.n6777 ASIG5V.n6776 1.11687
R44544 ASIG5V.n13618 ASIG5V.n13617 1.11687
R44545 ASIG5V.n13360 ASIG5V.n13359 1.11687
R44546 ASIG5V.n7401 ASIG5V.n7400 1.11687
R44547 ASIG5V.n7823 ASIG5V.n7822 1.11687
R44548 ASIG5V.n8120 ASIG5V.n8119 1.11687
R44549 ASIG5V.n12653 ASIG5V.n12652 1.11687
R44550 ASIG5V.n12425 ASIG5V.n12424 1.11687
R44551 ASIG5V.n12310 ASIG5V.n12309 1.11687
R44552 ASIG5V.n12154 ASIG5V.n12153 1.11687
R44553 ASIG5V.n11999 ASIG5V.n11998 1.11687
R44554 ASIG5V.n11831 ASIG5V.n11830 1.11687
R44555 ASIG5V.n11668 ASIG5V.n11667 1.11687
R44556 ASIG5V.n11486 ASIG5V.n11422 1.11687
R44557 ASIG5V.n11631 ASIG5V.n11494 1.11687
R44558 ASIG5V.n11760 ASIG5V.n11677 1.11687
R44559 ASIG5V.n11926 ASIG5V.n11842 1.11687
R44560 ASIG5V.n12082 ASIG5V.n12010 1.11687
R44561 ASIG5V.n12238 ASIG5V.n12165 1.11687
R44562 ASIG5V.n12352 ASIG5V.n12319 1.11687
R44563 ASIG5V.n12581 ASIG5V.n12436 1.11687
R44564 ASIG5V.n12752 ASIG5V.n12669 1.11687
R44565 ASIG5V.n7979 ASIG5V.n7946 1.11687
R44566 ASIG5V.n7626 ASIG5V.n7526 1.11687
R44567 ASIG5V.n331 ASIG5V.n151 1.11687
R44568 ASIG5V.n13495 ASIG5V.n13372 1.11687
R44569 ASIG5V.n6652 ASIG5V.n6557 1.11687
R44570 ASIG5V.n6928 ASIG5V.n6792 1.11687
R44571 ASIG5V.n7123 ASIG5V.n7067 1.11687
R44572 ASIG5V.n6149 ASIG5V.n5984 1.11687
R44573 ASIG5V.n5793 ASIG5V.n5687 1.11687
R44574 ASIG5V.n5442 ASIG5V.n5405 1.11687
R44575 ASIG5V.n5142 ASIG5V.n4983 1.11687
R44576 ASIG5V.n4847 ASIG5V.n4708 1.11687
R44577 ASIG5V.n4561 ASIG5V.n4454 1.11687
R44578 ASIG5V.n4277 ASIG5V.n4171 1.11687
R44579 ASIG5V.n4004 ASIG5V.n3904 1.11687
R44580 ASIG5V.n3737 ASIG5V.n3631 1.11687
R44581 ASIG5V.n3475 ASIG5V.n3339 1.11687
R44582 ASIG5V.n3251 ASIG5V.n3147 1.11687
R44583 ASIG5V.n3251 ASIG5V.n3150 1.11687
R44584 ASIG5V.n3475 ASIG5V.n3342 1.11687
R44585 ASIG5V.n3737 ASIG5V.n3632 1.11687
R44586 ASIG5V.n4004 ASIG5V.n3906 1.11687
R44587 ASIG5V.n4277 ASIG5V.n4174 1.11687
R44588 ASIG5V.n4561 ASIG5V.n4456 1.11687
R44589 ASIG5V.n4847 ASIG5V.n4711 1.11687
R44590 ASIG5V.n5142 ASIG5V.n4986 1.11687
R44591 ASIG5V.n5442 ASIG5V.n5406 1.11687
R44592 ASIG5V.n5793 ASIG5V.n5690 1.11687
R44593 ASIG5V.n6149 ASIG5V.n5987 1.11687
R44594 ASIG5V.n7123 ASIG5V.n7068 1.11687
R44595 ASIG5V.n6928 ASIG5V.n6793 1.11687
R44596 ASIG5V.n6652 ASIG5V.n6558 1.11687
R44597 ASIG5V.n13495 ASIG5V.n13373 1.11687
R44598 ASIG5V.n331 ASIG5V.n154 1.11687
R44599 ASIG5V.n7626 ASIG5V.n7528 1.11687
R44600 ASIG5V.n7979 ASIG5V.n7947 1.11687
R44601 ASIG5V.n12752 ASIG5V.n12671 1.11687
R44602 ASIG5V.n12581 ASIG5V.n12438 1.11687
R44603 ASIG5V.n12352 ASIG5V.n12320 1.11687
R44604 ASIG5V.n12238 ASIG5V.n12166 1.11687
R44605 ASIG5V.n12082 ASIG5V.n12012 1.11687
R44606 ASIG5V.n11926 ASIG5V.n11844 1.11687
R44607 ASIG5V.n11760 ASIG5V.n11679 1.11687
R44608 ASIG5V.n11631 ASIG5V.n11497 1.11687
R44609 ASIG5V.n3251 ASIG5V.n3153 1.11687
R44610 ASIG5V.n3475 ASIG5V.n3345 1.11687
R44611 ASIG5V.n3737 ASIG5V.n3635 1.11687
R44612 ASIG5V.n4004 ASIG5V.n3908 1.11687
R44613 ASIG5V.n4277 ASIG5V.n4177 1.11687
R44614 ASIG5V.n4561 ASIG5V.n4458 1.11687
R44615 ASIG5V.n4847 ASIG5V.n4714 1.11687
R44616 ASIG5V.n5142 ASIG5V.n4989 1.11687
R44617 ASIG5V.n5442 ASIG5V.n5407 1.11687
R44618 ASIG5V.n5793 ASIG5V.n5691 1.11687
R44619 ASIG5V.n6149 ASIG5V.n5990 1.11687
R44620 ASIG5V.n7123 ASIG5V.n7069 1.11687
R44621 ASIG5V.n6928 ASIG5V.n6795 1.11687
R44622 ASIG5V.n6652 ASIG5V.n6560 1.11687
R44623 ASIG5V.n13495 ASIG5V.n13374 1.11687
R44624 ASIG5V.n331 ASIG5V.n157 1.11687
R44625 ASIG5V.n7626 ASIG5V.n7529 1.11687
R44626 ASIG5V.n7979 ASIG5V.n7948 1.11687
R44627 ASIG5V.n12752 ASIG5V.n12673 1.11687
R44628 ASIG5V.n12581 ASIG5V.n12440 1.11687
R44629 ASIG5V.n12352 ASIG5V.n12321 1.11687
R44630 ASIG5V.n12238 ASIG5V.n12167 1.11687
R44631 ASIG5V.n12082 ASIG5V.n12013 1.11687
R44632 ASIG5V.n11926 ASIG5V.n11846 1.11687
R44633 ASIG5V.n11760 ASIG5V.n11681 1.11687
R44634 ASIG5V.n11631 ASIG5V.n11500 1.11687
R44635 ASIG5V.n11631 ASIG5V.n11503 1.11687
R44636 ASIG5V.n11760 ASIG5V.n11682 1.11687
R44637 ASIG5V.n11926 ASIG5V.n11848 1.11687
R44638 ASIG5V.n12082 ASIG5V.n12015 1.11687
R44639 ASIG5V.n12238 ASIG5V.n12169 1.11687
R44640 ASIG5V.n12352 ASIG5V.n12322 1.11687
R44641 ASIG5V.n12581 ASIG5V.n12443 1.11687
R44642 ASIG5V.n12752 ASIG5V.n12675 1.11687
R44643 ASIG5V.n7979 ASIG5V.n7949 1.11687
R44644 ASIG5V.n7626 ASIG5V.n7530 1.11687
R44645 ASIG5V.n331 ASIG5V.n160 1.11687
R44646 ASIG5V.n13495 ASIG5V.n13376 1.11687
R44647 ASIG5V.n6652 ASIG5V.n6561 1.11687
R44648 ASIG5V.n6928 ASIG5V.n6797 1.11687
R44649 ASIG5V.n7123 ASIG5V.n7070 1.11687
R44650 ASIG5V.n6149 ASIG5V.n5993 1.11687
R44651 ASIG5V.n5793 ASIG5V.n5692 1.11687
R44652 ASIG5V.n5442 ASIG5V.n5408 1.11687
R44653 ASIG5V.n5142 ASIG5V.n4992 1.11687
R44654 ASIG5V.n4847 ASIG5V.n4717 1.11687
R44655 ASIG5V.n4561 ASIG5V.n4460 1.11687
R44656 ASIG5V.n4277 ASIG5V.n4180 1.11687
R44657 ASIG5V.n4004 ASIG5V.n3910 1.11687
R44658 ASIG5V.n3737 ASIG5V.n3638 1.11687
R44659 ASIG5V.n3475 ASIG5V.n3348 1.11687
R44660 ASIG5V.n3251 ASIG5V.n3155 1.11687
R44661 ASIG5V.n3251 ASIG5V.n3157 1.11687
R44662 ASIG5V.n3475 ASIG5V.n3353 1.11687
R44663 ASIG5V.n3737 ASIG5V.n3643 1.11687
R44664 ASIG5V.n4004 ASIG5V.n3915 1.11687
R44665 ASIG5V.n4277 ASIG5V.n4183 1.11687
R44666 ASIG5V.n4561 ASIG5V.n4463 1.11687
R44667 ASIG5V.n4847 ASIG5V.n4722 1.11687
R44668 ASIG5V.n5142 ASIG5V.n4997 1.11687
R44669 ASIG5V.n5442 ASIG5V.n5409 1.11687
R44670 ASIG5V.n5793 ASIG5V.n5695 1.11687
R44671 ASIG5V.n6149 ASIG5V.n5998 1.11687
R44672 ASIG5V.n7123 ASIG5V.n7071 1.11687
R44673 ASIG5V.n6928 ASIG5V.n6798 1.11687
R44674 ASIG5V.n6652 ASIG5V.n6564 1.11687
R44675 ASIG5V.n13495 ASIG5V.n13379 1.11687
R44676 ASIG5V.n331 ASIG5V.n165 1.11687
R44677 ASIG5V.n7626 ASIG5V.n7533 1.11687
R44678 ASIG5V.n7979 ASIG5V.n7950 1.11687
R44679 ASIG5V.n12752 ASIG5V.n12678 1.11687
R44680 ASIG5V.n12581 ASIG5V.n12446 1.11687
R44681 ASIG5V.n12352 ASIG5V.n12323 1.11687
R44682 ASIG5V.n12238 ASIG5V.n12170 1.11687
R44683 ASIG5V.n12082 ASIG5V.n12018 1.11687
R44684 ASIG5V.n11926 ASIG5V.n11851 1.11687
R44685 ASIG5V.n11760 ASIG5V.n11685 1.11687
R44686 ASIG5V.n11631 ASIG5V.n11508 1.11687
R44687 ASIG5V.n11631 ASIG5V.n11513 1.11687
R44688 ASIG5V.n11760 ASIG5V.n11686 1.11687
R44689 ASIG5V.n11926 ASIG5V.n11854 1.11687
R44690 ASIG5V.n12082 ASIG5V.n12021 1.11687
R44691 ASIG5V.n12238 ASIG5V.n12173 1.11687
R44692 ASIG5V.n12352 ASIG5V.n12324 1.11687
R44693 ASIG5V.n12581 ASIG5V.n12449 1.11687
R44694 ASIG5V.n12752 ASIG5V.n12683 1.11687
R44695 ASIG5V.n7979 ASIG5V.n7951 1.11687
R44696 ASIG5V.n7626 ASIG5V.n7536 1.11687
R44697 ASIG5V.n331 ASIG5V.n170 1.11687
R44698 ASIG5V.n13495 ASIG5V.n13382 1.11687
R44699 ASIG5V.n6652 ASIG5V.n6565 1.11687
R44700 ASIG5V.n6928 ASIG5V.n6801 1.11687
R44701 ASIG5V.n7123 ASIG5V.n7072 1.11687
R44702 ASIG5V.n6149 ASIG5V.n6003 1.11687
R44703 ASIG5V.n5793 ASIG5V.n5698 1.11687
R44704 ASIG5V.n5442 ASIG5V.n5410 1.11687
R44705 ASIG5V.n5142 ASIG5V.n5002 1.11687
R44706 ASIG5V.n4847 ASIG5V.n4727 1.11687
R44707 ASIG5V.n4561 ASIG5V.n4468 1.11687
R44708 ASIG5V.n4277 ASIG5V.n4188 1.11687
R44709 ASIG5V.n4004 ASIG5V.n3918 1.11687
R44710 ASIG5V.n3737 ASIG5V.n3648 1.11687
R44711 ASIG5V.n3475 ASIG5V.n3358 1.11687
R44712 ASIG5V.n3251 ASIG5V.n3162 1.11687
R44713 ASIG5V.n3251 ASIG5V.n3167 1.11687
R44714 ASIG5V.n3475 ASIG5V.n3363 1.11687
R44715 ASIG5V.n3737 ASIG5V.n3651 1.11687
R44716 ASIG5V.n4004 ASIG5V.n3919 1.11687
R44717 ASIG5V.n4277 ASIG5V.n4191 1.11687
R44718 ASIG5V.n4561 ASIG5V.n4471 1.11687
R44719 ASIG5V.n4847 ASIG5V.n4732 1.11687
R44720 ASIG5V.n5142 ASIG5V.n5007 1.11687
R44721 ASIG5V.n5442 ASIG5V.n5411 1.11687
R44722 ASIG5V.n5793 ASIG5V.n5701 1.11687
R44723 ASIG5V.n6149 ASIG5V.n6008 1.11687
R44724 ASIG5V.n7123 ASIG5V.n7073 1.11687
R44725 ASIG5V.n6928 ASIG5V.n6802 1.11687
R44726 ASIG5V.n6652 ASIG5V.n6568 1.11687
R44727 ASIG5V.n13495 ASIG5V.n13385 1.11687
R44728 ASIG5V.n331 ASIG5V.n175 1.11687
R44729 ASIG5V.n7626 ASIG5V.n7539 1.11687
R44730 ASIG5V.n7979 ASIG5V.n7952 1.11687
R44731 ASIG5V.n12752 ASIG5V.n12686 1.11687
R44732 ASIG5V.n12581 ASIG5V.n12452 1.11687
R44733 ASIG5V.n12352 ASIG5V.n12325 1.11687
R44734 ASIG5V.n12238 ASIG5V.n12176 1.11687
R44735 ASIG5V.n12082 ASIG5V.n12022 1.11687
R44736 ASIG5V.n11926 ASIG5V.n11857 1.11687
R44737 ASIG5V.n11760 ASIG5V.n11689 1.11687
R44738 ASIG5V.n11631 ASIG5V.n11518 1.11687
R44739 ASIG5V.n3251 ASIG5V.n3170 1.11687
R44740 ASIG5V.n3475 ASIG5V.n3368 1.11687
R44741 ASIG5V.n3737 ASIG5V.n3656 1.11687
R44742 ASIG5V.n4004 ASIG5V.n3922 1.11687
R44743 ASIG5V.n4277 ASIG5V.n4194 1.11687
R44744 ASIG5V.n4561 ASIG5V.n4474 1.11687
R44745 ASIG5V.n4847 ASIG5V.n4737 1.11687
R44746 ASIG5V.n5142 ASIG5V.n5013 1.11687
R44747 ASIG5V.n5442 ASIG5V.n5412 1.11687
R44748 ASIG5V.n5793 ASIG5V.n5705 1.11687
R44749 ASIG5V.n6149 ASIG5V.n6015 1.11687
R44750 ASIG5V.n7123 ASIG5V.n7074 1.11687
R44751 ASIG5V.n6928 ASIG5V.n6806 1.11687
R44752 ASIG5V.n6652 ASIG5V.n6572 1.11687
R44753 ASIG5V.n13495 ASIG5V.n13386 1.11687
R44754 ASIG5V.n331 ASIG5V.n182 1.11687
R44755 ASIG5V.n7626 ASIG5V.n7543 1.11687
R44756 ASIG5V.n7979 ASIG5V.n7953 1.11687
R44757 ASIG5V.n12752 ASIG5V.n12690 1.11687
R44758 ASIG5V.n12581 ASIG5V.n12458 1.11687
R44759 ASIG5V.n12352 ASIG5V.n12326 1.11687
R44760 ASIG5V.n12238 ASIG5V.n12179 1.11687
R44761 ASIG5V.n12082 ASIG5V.n12025 1.11687
R44762 ASIG5V.n11926 ASIG5V.n11860 1.11687
R44763 ASIG5V.n11760 ASIG5V.n11692 1.11687
R44764 ASIG5V.n11631 ASIG5V.n11523 1.11687
R44765 ASIG5V.n11631 ASIG5V.n11528 1.11687
R44766 ASIG5V.n11760 ASIG5V.n11695 1.11687
R44767 ASIG5V.n11926 ASIG5V.n11861 1.11687
R44768 ASIG5V.n12082 ASIG5V.n12028 1.11687
R44769 ASIG5V.n12238 ASIG5V.n12182 1.11687
R44770 ASIG5V.n12352 ASIG5V.n12327 1.11687
R44771 ASIG5V.n12581 ASIG5V.n12462 1.11687
R44772 ASIG5V.n12752 ASIG5V.n12694 1.11687
R44773 ASIG5V.n7979 ASIG5V.n7954 1.11687
R44774 ASIG5V.n7626 ASIG5V.n7547 1.11687
R44775 ASIG5V.n331 ASIG5V.n189 1.11687
R44776 ASIG5V.n13495 ASIG5V.n13390 1.11687
R44777 ASIG5V.n6652 ASIG5V.n6576 1.11687
R44778 ASIG5V.n6928 ASIG5V.n6810 1.11687
R44779 ASIG5V.n7123 ASIG5V.n7075 1.11687
R44780 ASIG5V.n6149 ASIG5V.n6022 1.11687
R44781 ASIG5V.n5793 ASIG5V.n5709 1.11687
R44782 ASIG5V.n5442 ASIG5V.n5413 1.11687
R44783 ASIG5V.n5142 ASIG5V.n5020 1.11687
R44784 ASIG5V.n4847 ASIG5V.n4740 1.11687
R44785 ASIG5V.n4561 ASIG5V.n4477 1.11687
R44786 ASIG5V.n4277 ASIG5V.n4197 1.11687
R44787 ASIG5V.n4004 ASIG5V.n3925 1.11687
R44788 ASIG5V.n3737 ASIG5V.n3661 1.11687
R44789 ASIG5V.n3475 ASIG5V.n3373 1.11687
R44790 ASIG5V.n3251 ASIG5V.n3175 1.11687
R44791 ASIG5V.n3251 ASIG5V.n3178 1.11687
R44792 ASIG5V.n3475 ASIG5V.n3378 1.11687
R44793 ASIG5V.n3737 ASIG5V.n3665 1.11687
R44794 ASIG5V.n4004 ASIG5V.n3929 1.11687
R44795 ASIG5V.n4277 ASIG5V.n4201 1.11687
R44796 ASIG5V.n4561 ASIG5V.n4481 1.11687
R44797 ASIG5V.n4847 ASIG5V.n4741 1.11687
R44798 ASIG5V.n5142 ASIG5V.n5027 1.11687
R44799 ASIG5V.n5442 ASIG5V.n5414 1.11687
R44800 ASIG5V.n5793 ASIG5V.n5713 1.11687
R44801 ASIG5V.n6149 ASIG5V.n6029 1.11687
R44802 ASIG5V.n7123 ASIG5V.n7076 1.11687
R44803 ASIG5V.n6928 ASIG5V.n6814 1.11687
R44804 ASIG5V.n6652 ASIG5V.n6583 1.11687
R44805 ASIG5V.n13495 ASIG5V.n13391 1.11687
R44806 ASIG5V.n331 ASIG5V.n196 1.11687
R44807 ASIG5V.n7626 ASIG5V.n7548 1.11687
R44808 ASIG5V.n7979 ASIG5V.n7955 1.11687
R44809 ASIG5V.n12752 ASIG5V.n12698 1.11687
R44810 ASIG5V.n12581 ASIG5V.n12466 1.11687
R44811 ASIG5V.n12352 ASIG5V.n12328 1.11687
R44812 ASIG5V.n12238 ASIG5V.n12183 1.11687
R44813 ASIG5V.n12082 ASIG5V.n12029 1.11687
R44814 ASIG5V.n11926 ASIG5V.n11865 1.11687
R44815 ASIG5V.n11760 ASIG5V.n11699 1.11687
R44816 ASIG5V.n11631 ASIG5V.n11533 1.11687
R44817 ASIG5V.n3251 ASIG5V.n3181 1.11687
R44818 ASIG5V.n3475 ASIG5V.n3383 1.11687
R44819 ASIG5V.n3737 ASIG5V.n3670 1.11687
R44820 ASIG5V.n4004 ASIG5V.n3932 1.11687
R44821 ASIG5V.n4277 ASIG5V.n4205 1.11687
R44822 ASIG5V.n4561 ASIG5V.n4485 1.11687
R44823 ASIG5V.n4847 ASIG5V.n4748 1.11687
R44824 ASIG5V.n5142 ASIG5V.n5034 1.11687
R44825 ASIG5V.n5442 ASIG5V.n5415 1.11687
R44826 ASIG5V.n5793 ASIG5V.n5717 1.11687
R44827 ASIG5V.n6149 ASIG5V.n6036 1.11687
R44828 ASIG5V.n7123 ASIG5V.n7077 1.11687
R44829 ASIG5V.n6928 ASIG5V.n6818 1.11687
R44830 ASIG5V.n6652 ASIG5V.n6590 1.11687
R44831 ASIG5V.n13495 ASIG5V.n13398 1.11687
R44832 ASIG5V.n331 ASIG5V.n203 1.11687
R44833 ASIG5V.n7626 ASIG5V.n7549 1.11687
R44834 ASIG5V.n7979 ASIG5V.n7956 1.11687
R44835 ASIG5V.n12752 ASIG5V.n12699 1.11687
R44836 ASIG5V.n12581 ASIG5V.n12467 1.11687
R44837 ASIG5V.n12352 ASIG5V.n12329 1.11687
R44838 ASIG5V.n12238 ASIG5V.n12187 1.11687
R44839 ASIG5V.n12082 ASIG5V.n12030 1.11687
R44840 ASIG5V.n11926 ASIG5V.n11868 1.11687
R44841 ASIG5V.n11760 ASIG5V.n11702 1.11687
R44842 ASIG5V.n11631 ASIG5V.n11538 1.11687
R44843 ASIG5V.n11631 ASIG5V.n11543 1.11687
R44844 ASIG5V.n11760 ASIG5V.n11705 1.11687
R44845 ASIG5V.n11926 ASIG5V.n11871 1.11687
R44846 ASIG5V.n12082 ASIG5V.n12033 1.11687
R44847 ASIG5V.n12238 ASIG5V.n12188 1.11687
R44848 ASIG5V.n12352 ASIG5V.n12330 1.11687
R44849 ASIG5V.n12581 ASIG5V.n12471 1.11687
R44850 ASIG5V.n12752 ASIG5V.n12700 1.11687
R44851 ASIG5V.n7979 ASIG5V.n7957 1.11687
R44852 ASIG5V.n7626 ASIG5V.n7553 1.11687
R44853 ASIG5V.n331 ASIG5V.n210 1.11687
R44854 ASIG5V.n13495 ASIG5V.n13402 1.11687
R44855 ASIG5V.n6652 ASIG5V.n6597 1.11687
R44856 ASIG5V.n6928 ASIG5V.n6819 1.11687
R44857 ASIG5V.n7123 ASIG5V.n7081 1.11687
R44858 ASIG5V.n6149 ASIG5V.n6043 1.11687
R44859 ASIG5V.n5793 ASIG5V.n5721 1.11687
R44860 ASIG5V.n5442 ASIG5V.n5416 1.11687
R44861 ASIG5V.n5142 ASIG5V.n5041 1.11687
R44862 ASIG5V.n4847 ASIG5V.n4752 1.11687
R44863 ASIG5V.n4561 ASIG5V.n4489 1.11687
R44864 ASIG5V.n4277 ASIG5V.n4208 1.11687
R44865 ASIG5V.n4004 ASIG5V.n3937 1.11687
R44866 ASIG5V.n3737 ASIG5V.n3671 1.11687
R44867 ASIG5V.n3475 ASIG5V.n3388 1.11687
R44868 ASIG5V.n3251 ASIG5V.n3186 1.11687
R44869 ASIG5V.n3251 ASIG5V.n3189 1.11687
R44870 ASIG5V.n3475 ASIG5V.n3393 1.11687
R44871 ASIG5V.n3737 ASIG5V.n3674 1.11687
R44872 ASIG5V.n4004 ASIG5V.n3942 1.11687
R44873 ASIG5V.n4277 ASIG5V.n4211 1.11687
R44874 ASIG5V.n4561 ASIG5V.n4492 1.11687
R44875 ASIG5V.n4847 ASIG5V.n4757 1.11687
R44876 ASIG5V.n5142 ASIG5V.n5047 1.11687
R44877 ASIG5V.n5442 ASIG5V.n5417 1.11687
R44878 ASIG5V.n5793 ASIG5V.n5725 1.11687
R44879 ASIG5V.n6149 ASIG5V.n6050 1.11687
R44880 ASIG5V.n7123 ASIG5V.n7088 1.11687
R44881 ASIG5V.n6928 ASIG5V.n6820 1.11687
R44882 ASIG5V.n6652 ASIG5V.n6604 1.11687
R44883 ASIG5V.n13495 ASIG5V.n13403 1.11687
R44884 ASIG5V.n331 ASIG5V.n217 1.11687
R44885 ASIG5V.n7626 ASIG5V.n7557 1.11687
R44886 ASIG5V.n7979 ASIG5V.n7958 1.11687
R44887 ASIG5V.n12752 ASIG5V.n12701 1.11687
R44888 ASIG5V.n12581 ASIG5V.n12477 1.11687
R44889 ASIG5V.n12352 ASIG5V.n12331 1.11687
R44890 ASIG5V.n12238 ASIG5V.n12191 1.11687
R44891 ASIG5V.n12082 ASIG5V.n12036 1.11687
R44892 ASIG5V.n11926 ASIG5V.n11874 1.11687
R44893 ASIG5V.n11760 ASIG5V.n11708 1.11687
R44894 ASIG5V.n11631 ASIG5V.n11548 1.11687
R44895 ASIG5V.n3251 ASIG5V.n3192 1.11687
R44896 ASIG5V.n3475 ASIG5V.n3396 1.11687
R44897 ASIG5V.n3737 ASIG5V.n3677 1.11687
R44898 ASIG5V.n4004 ASIG5V.n3945 1.11687
R44899 ASIG5V.n4277 ASIG5V.n4214 1.11687
R44900 ASIG5V.n4561 ASIG5V.n4497 1.11687
R44901 ASIG5V.n4847 ASIG5V.n4762 1.11687
R44902 ASIG5V.n5142 ASIG5V.n5052 1.11687
R44903 ASIG5V.n5442 ASIG5V.n5418 1.11687
R44904 ASIG5V.n5793 ASIG5V.n5730 1.11687
R44905 ASIG5V.n6149 ASIG5V.n6057 1.11687
R44906 ASIG5V.n7123 ASIG5V.n7092 1.11687
R44907 ASIG5V.n6928 ASIG5V.n6824 1.11687
R44908 ASIG5V.n6652 ASIG5V.n6611 1.11687
R44909 ASIG5V.n13495 ASIG5V.n13404 1.11687
R44910 ASIG5V.n331 ASIG5V.n224 1.11687
R44911 ASIG5V.n7626 ASIG5V.n7561 1.11687
R44912 ASIG5V.n7979 ASIG5V.n7959 1.11687
R44913 ASIG5V.n12752 ASIG5V.n12702 1.11687
R44914 ASIG5V.n12581 ASIG5V.n12482 1.11687
R44915 ASIG5V.n12352 ASIG5V.n12332 1.11687
R44916 ASIG5V.n12238 ASIG5V.n12192 1.11687
R44917 ASIG5V.n12082 ASIG5V.n12039 1.11687
R44918 ASIG5V.n11926 ASIG5V.n11877 1.11687
R44919 ASIG5V.n11760 ASIG5V.n11710 1.11687
R44920 ASIG5V.n11631 ASIG5V.n11551 1.11687
R44921 ASIG5V.n11631 ASIG5V.n11554 1.11687
R44922 ASIG5V.n11760 ASIG5V.n11712 1.11687
R44923 ASIG5V.n11926 ASIG5V.n11878 1.11687
R44924 ASIG5V.n12082 ASIG5V.n12040 1.11687
R44925 ASIG5V.n12238 ASIG5V.n12193 1.11687
R44926 ASIG5V.n12352 ASIG5V.n12333 1.11687
R44927 ASIG5V.n12581 ASIG5V.n12487 1.11687
R44928 ASIG5V.n12752 ASIG5V.n12703 1.11687
R44929 ASIG5V.n7979 ASIG5V.n7960 1.11687
R44930 ASIG5V.n7626 ASIG5V.n7564 1.11687
R44931 ASIG5V.n331 ASIG5V.n231 1.11687
R44932 ASIG5V.n13495 ASIG5V.n13408 1.11687
R44933 ASIG5V.n6652 ASIG5V.n6615 1.11687
R44934 ASIG5V.n6928 ASIG5V.n6828 1.11687
R44935 ASIG5V.n7123 ASIG5V.n7096 1.11687
R44936 ASIG5V.n6149 ASIG5V.n6062 1.11687
R44937 ASIG5V.n5793 ASIG5V.n5735 1.11687
R44938 ASIG5V.n5442 ASIG5V.n5419 1.11687
R44939 ASIG5V.n5142 ASIG5V.n5057 1.11687
R44940 ASIG5V.n4847 ASIG5V.n4767 1.11687
R44941 ASIG5V.n4561 ASIG5V.n4500 1.11687
R44942 ASIG5V.n4277 ASIG5V.n4217 1.11687
R44943 ASIG5V.n4004 ASIG5V.n3948 1.11687
R44944 ASIG5V.n3737 ASIG5V.n3679 1.11687
R44945 ASIG5V.n3475 ASIG5V.n3399 1.11687
R44946 ASIG5V.n3251 ASIG5V.n3194 1.11687
R44947 ASIG5V.n3104 ASIG5V.n3102 1.11687
R44948 ASIG5V.n3251 ASIG5V.n3197 1.11687
R44949 ASIG5V.n3104 ASIG5V.n3101 1.11687
R44950 ASIG5V.n3251 ASIG5V.n3200 1.11687
R44951 ASIG5V.n3104 ASIG5V.n3100 1.11687
R44952 ASIG5V.n3104 ASIG5V.n3099 1.11687
R44953 ASIG5V.n3251 ASIG5V.n3202 1.11687
R44954 ASIG5V.n3104 ASIG5V.n3098 1.11687
R44955 ASIG5V.n3251 ASIG5V.n3204 1.11687
R44956 ASIG5V.n3104 ASIG5V.n3096 1.11687
R44957 ASIG5V.n3104 ASIG5V.n3094 1.11687
R44958 ASIG5V.n3104 ASIG5V.n3093 1.11687
R44959 ASIG5V.n3251 ASIG5V.n3206 1.11687
R44960 ASIG5V.n3104 ASIG5V.n3091 1.11687
R44961 ASIG5V.n3104 ASIG5V.n3089 1.11687
R44962 ASIG5V.n3104 ASIG5V.n3086 1.11687
R44963 ASIG5V.n3251 ASIG5V.n3209 1.11687
R44964 ASIG5V.n3104 ASIG5V.n3085 1.11687
R44965 ASIG5V.n3251 ASIG5V.n3214 1.11687
R44966 ASIG5V.n3104 ASIG5V.n3082 1.11687
R44967 ASIG5V.n3104 ASIG5V.n3081 1.11687
R44968 ASIG5V.n3251 ASIG5V.n3219 1.11687
R44969 ASIG5V.n3104 ASIG5V.n3080 1.11687
R44970 ASIG5V.n3251 ASIG5V.n3222 1.11687
R44971 ASIG5V.n3104 ASIG5V.n3079 1.11687
R44972 ASIG5V.n3104 ASIG5V.n3076 1.11687
R44973 ASIG5V.n3104 ASIG5V.n3073 1.11687
R44974 ASIG5V.n3251 ASIG5V.n3225 1.11687
R44975 ASIG5V.n3104 ASIG5V.n3072 1.11687
R44976 ASIG5V.n3251 ASIG5V.n3228 1.11687
R44977 ASIG5V.n3104 ASIG5V.n3069 1.11687
R44978 ASIG5V.n3104 ASIG5V.n3066 1.11687
R44979 ASIG5V.n3251 ASIG5V.n3231 1.11687
R44980 ASIG5V.n3104 ASIG5V.n3063 1.11687
R44981 ASIG5V.n3251 ASIG5V.n3236 1.11687
R44982 ASIG5V.n3104 ASIG5V.n3060 1.11687
R44983 ASIG5V.n3104 ASIG5V.n3059 1.11687
R44984 ASIG5V.n3104 ASIG5V.n3056 1.11687
R44985 ASIG5V.n3251 ASIG5V.n3239 1.11687
R44986 ASIG5V.n3104 ASIG5V.n3055 1.11687
R44987 ASIG5V.n3251 ASIG5V.n3244 1.11687
R44988 ASIG5V.n3104 ASIG5V.n3052 1.11687
R44989 ASIG5V.n3104 ASIG5V.n3051 1.11687
R44990 ASIG5V.n3251 ASIG5V.n3246 1.11687
R44991 ASIG5V.n3104 ASIG5V.n3049 1.11687
R44992 ASIG5V.n3251 ASIG5V.n3248 1.11687
R44993 ASIG5V.n3104 ASIG5V.n3047 1.11687
R44994 ASIG5V.n3104 ASIG5V.n3045 1.11687
R44995 ASIG5V.n3104 ASIG5V.n3044 1.11687
R44996 ASIG5V.n3251 ASIG5V.n3250 1.11687
R44997 ASIG5V.n3104 ASIG5V.n3042 1.11687
R44998 ASIG5V.n3296 ASIG5V.n3293 1.11687
R44999 ASIG5V.n3475 ASIG5V.n3402 1.11687
R45000 ASIG5V.n3296 ASIG5V.n3292 1.11687
R45001 ASIG5V.n3475 ASIG5V.n3405 1.11687
R45002 ASIG5V.n3296 ASIG5V.n3291 1.11687
R45003 ASIG5V.n3296 ASIG5V.n3290 1.11687
R45004 ASIG5V.n3475 ASIG5V.n3408 1.11687
R45005 ASIG5V.n3296 ASIG5V.n3289 1.11687
R45006 ASIG5V.n3475 ASIG5V.n3411 1.11687
R45007 ASIG5V.n3296 ASIG5V.n3288 1.11687
R45008 ASIG5V.n3296 ASIG5V.n3287 1.11687
R45009 ASIG5V.n3296 ASIG5V.n3286 1.11687
R45010 ASIG5V.n3475 ASIG5V.n3414 1.11687
R45011 ASIG5V.n3296 ASIG5V.n3285 1.11687
R45012 ASIG5V.n3296 ASIG5V.n3284 1.11687
R45013 ASIG5V.n3296 ASIG5V.n3283 1.11687
R45014 ASIG5V.n3475 ASIG5V.n3419 1.11687
R45015 ASIG5V.n3296 ASIG5V.n3282 1.11687
R45016 ASIG5V.n3475 ASIG5V.n3424 1.11687
R45017 ASIG5V.n3296 ASIG5V.n3281 1.11687
R45018 ASIG5V.n3296 ASIG5V.n3280 1.11687
R45019 ASIG5V.n3475 ASIG5V.n3429 1.11687
R45020 ASIG5V.n3296 ASIG5V.n3279 1.11687
R45021 ASIG5V.n3475 ASIG5V.n3434 1.11687
R45022 ASIG5V.n3296 ASIG5V.n3278 1.11687
R45023 ASIG5V.n3296 ASIG5V.n3277 1.11687
R45024 ASIG5V.n3296 ASIG5V.n3276 1.11687
R45025 ASIG5V.n3475 ASIG5V.n3439 1.11687
R45026 ASIG5V.n3296 ASIG5V.n3275 1.11687
R45027 ASIG5V.n3475 ASIG5V.n3444 1.11687
R45028 ASIG5V.n3296 ASIG5V.n3274 1.11687
R45029 ASIG5V.n3296 ASIG5V.n3273 1.11687
R45030 ASIG5V.n3475 ASIG5V.n3449 1.11687
R45031 ASIG5V.n3296 ASIG5V.n3272 1.11687
R45032 ASIG5V.n3475 ASIG5V.n3454 1.11687
R45033 ASIG5V.n3296 ASIG5V.n3271 1.11687
R45034 ASIG5V.n3296 ASIG5V.n3270 1.11687
R45035 ASIG5V.n3296 ASIG5V.n3269 1.11687
R45036 ASIG5V.n3475 ASIG5V.n3459 1.11687
R45037 ASIG5V.n3296 ASIG5V.n3268 1.11687
R45038 ASIG5V.n3475 ASIG5V.n3464 1.11687
R45039 ASIG5V.n3296 ASIG5V.n3267 1.11687
R45040 ASIG5V.n3296 ASIG5V.n3266 1.11687
R45041 ASIG5V.n3475 ASIG5V.n3469 1.11687
R45042 ASIG5V.n3296 ASIG5V.n3265 1.11687
R45043 ASIG5V.n3475 ASIG5V.n3472 1.11687
R45044 ASIG5V.n3296 ASIG5V.n3264 1.11687
R45045 ASIG5V.n3296 ASIG5V.n3263 1.11687
R45046 ASIG5V.n3296 ASIG5V.n3262 1.11687
R45047 ASIG5V.n3475 ASIG5V.n3474 1.11687
R45048 ASIG5V.n3296 ASIG5V.n3261 1.11687
R45049 ASIG5V.n3558 ASIG5V.n3554 1.11687
R45050 ASIG5V.n3737 ASIG5V.n3682 1.11687
R45051 ASIG5V.n3558 ASIG5V.n3553 1.11687
R45052 ASIG5V.n3737 ASIG5V.n3684 1.11687
R45053 ASIG5V.n3558 ASIG5V.n3552 1.11687
R45054 ASIG5V.n3558 ASIG5V.n3549 1.11687
R45055 ASIG5V.n3737 ASIG5V.n3685 1.11687
R45056 ASIG5V.n3558 ASIG5V.n3546 1.11687
R45057 ASIG5V.n3737 ASIG5V.n3687 1.11687
R45058 ASIG5V.n3558 ASIG5V.n3543 1.11687
R45059 ASIG5V.n3558 ASIG5V.n3542 1.11687
R45060 ASIG5V.n3558 ASIG5V.n3541 1.11687
R45061 ASIG5V.n3737 ASIG5V.n3690 1.11687
R45062 ASIG5V.n3558 ASIG5V.n3539 1.11687
R45063 ASIG5V.n3558 ASIG5V.n3538 1.11687
R45064 ASIG5V.n3558 ASIG5V.n3537 1.11687
R45065 ASIG5V.n3737 ASIG5V.n3693 1.11687
R45066 ASIG5V.n3558 ASIG5V.n3536 1.11687
R45067 ASIG5V.n3737 ASIG5V.n3696 1.11687
R45068 ASIG5V.n3558 ASIG5V.n3531 1.11687
R45069 ASIG5V.n3558 ASIG5V.n3528 1.11687
R45070 ASIG5V.n3737 ASIG5V.n3701 1.11687
R45071 ASIG5V.n3558 ASIG5V.n3527 1.11687
R45072 ASIG5V.n3737 ASIG5V.n3704 1.11687
R45073 ASIG5V.n3558 ASIG5V.n3524 1.11687
R45074 ASIG5V.n3558 ASIG5V.n3523 1.11687
R45075 ASIG5V.n3558 ASIG5V.n3522 1.11687
R45076 ASIG5V.n3737 ASIG5V.n3707 1.11687
R45077 ASIG5V.n3558 ASIG5V.n3519 1.11687
R45078 ASIG5V.n3737 ASIG5V.n3712 1.11687
R45079 ASIG5V.n3558 ASIG5V.n3518 1.11687
R45080 ASIG5V.n3558 ASIG5V.n3514 1.11687
R45081 ASIG5V.n3737 ASIG5V.n3715 1.11687
R45082 ASIG5V.n3558 ASIG5V.n3510 1.11687
R45083 ASIG5V.n3737 ASIG5V.n3720 1.11687
R45084 ASIG5V.n3558 ASIG5V.n3509 1.11687
R45085 ASIG5V.n3558 ASIG5V.n3508 1.11687
R45086 ASIG5V.n3558 ASIG5V.n3505 1.11687
R45087 ASIG5V.n3737 ASIG5V.n3725 1.11687
R45088 ASIG5V.n3558 ASIG5V.n3502 1.11687
R45089 ASIG5V.n3737 ASIG5V.n3728 1.11687
R45090 ASIG5V.n3558 ASIG5V.n3499 1.11687
R45091 ASIG5V.n3558 ASIG5V.n3496 1.11687
R45092 ASIG5V.n3737 ASIG5V.n3731 1.11687
R45093 ASIG5V.n3558 ASIG5V.n3493 1.11687
R45094 ASIG5V.n3737 ASIG5V.n3734 1.11687
R45095 ASIG5V.n3558 ASIG5V.n3490 1.11687
R45096 ASIG5V.n3558 ASIG5V.n3489 1.11687
R45097 ASIG5V.n3558 ASIG5V.n3487 1.11687
R45098 ASIG5V.n3737 ASIG5V.n3736 1.11687
R45099 ASIG5V.n3558 ASIG5V.n3485 1.11687
R45100 ASIG5V.n3833 ASIG5V.n3830 1.11687
R45101 ASIG5V.n4004 ASIG5V.n3950 1.11687
R45102 ASIG5V.n3833 ASIG5V.n3828 1.11687
R45103 ASIG5V.n4004 ASIG5V.n3953 1.11687
R45104 ASIG5V.n3833 ASIG5V.n3826 1.11687
R45105 ASIG5V.n3833 ASIG5V.n3825 1.11687
R45106 ASIG5V.n4004 ASIG5V.n3955 1.11687
R45107 ASIG5V.n3833 ASIG5V.n3823 1.11687
R45108 ASIG5V.n4004 ASIG5V.n3957 1.11687
R45109 ASIG5V.n3833 ASIG5V.n3821 1.11687
R45110 ASIG5V.n3833 ASIG5V.n3819 1.11687
R45111 ASIG5V.n3833 ASIG5V.n3817 1.11687
R45112 ASIG5V.n4004 ASIG5V.n3961 1.11687
R45113 ASIG5V.n3833 ASIG5V.n3815 1.11687
R45114 ASIG5V.n3833 ASIG5V.n3814 1.11687
R45115 ASIG5V.n3833 ASIG5V.n3813 1.11687
R45116 ASIG5V.n4004 ASIG5V.n3966 1.11687
R45117 ASIG5V.n3833 ASIG5V.n3810 1.11687
R45118 ASIG5V.n4004 ASIG5V.n3969 1.11687
R45119 ASIG5V.n3833 ASIG5V.n3809 1.11687
R45120 ASIG5V.n3833 ASIG5V.n3804 1.11687
R45121 ASIG5V.n4004 ASIG5V.n3972 1.11687
R45122 ASIG5V.n3833 ASIG5V.n3801 1.11687
R45123 ASIG5V.n4004 ASIG5V.n3975 1.11687
R45124 ASIG5V.n3833 ASIG5V.n3798 1.11687
R45125 ASIG5V.n3833 ASIG5V.n3795 1.11687
R45126 ASIG5V.n3833 ASIG5V.n3792 1.11687
R45127 ASIG5V.n4004 ASIG5V.n3978 1.11687
R45128 ASIG5V.n3833 ASIG5V.n3789 1.11687
R45129 ASIG5V.n4004 ASIG5V.n3981 1.11687
R45130 ASIG5V.n3833 ASIG5V.n3786 1.11687
R45131 ASIG5V.n3833 ASIG5V.n3782 1.11687
R45132 ASIG5V.n4004 ASIG5V.n3985 1.11687
R45133 ASIG5V.n3833 ASIG5V.n3778 1.11687
R45134 ASIG5V.n4004 ASIG5V.n3989 1.11687
R45135 ASIG5V.n3833 ASIG5V.n3774 1.11687
R45136 ASIG5V.n3833 ASIG5V.n3771 1.11687
R45137 ASIG5V.n3833 ASIG5V.n3768 1.11687
R45138 ASIG5V.n4004 ASIG5V.n3992 1.11687
R45139 ASIG5V.n3833 ASIG5V.n3765 1.11687
R45140 ASIG5V.n4004 ASIG5V.n3995 1.11687
R45141 ASIG5V.n3833 ASIG5V.n3764 1.11687
R45142 ASIG5V.n3833 ASIG5V.n3761 1.11687
R45143 ASIG5V.n4004 ASIG5V.n3996 1.11687
R45144 ASIG5V.n3833 ASIG5V.n3758 1.11687
R45145 ASIG5V.n4004 ASIG5V.n4001 1.11687
R45146 ASIG5V.n3833 ASIG5V.n3755 1.11687
R45147 ASIG5V.n3833 ASIG5V.n3754 1.11687
R45148 ASIG5V.n3833 ASIG5V.n3751 1.11687
R45149 ASIG5V.n4004 ASIG5V.n4003 1.11687
R45150 ASIG5V.n3833 ASIG5V.n3750 1.11687
R45151 ASIG5V.n4096 ASIG5V.n4093 1.11687
R45152 ASIG5V.n4277 ASIG5V.n4220 1.11687
R45153 ASIG5V.n4096 ASIG5V.n4092 1.11687
R45154 ASIG5V.n4277 ASIG5V.n4223 1.11687
R45155 ASIG5V.n4096 ASIG5V.n4091 1.11687
R45156 ASIG5V.n4096 ASIG5V.n4090 1.11687
R45157 ASIG5V.n4277 ASIG5V.n4226 1.11687
R45158 ASIG5V.n4096 ASIG5V.n4089 1.11687
R45159 ASIG5V.n4277 ASIG5V.n4229 1.11687
R45160 ASIG5V.n4096 ASIG5V.n4088 1.11687
R45161 ASIG5V.n4096 ASIG5V.n4087 1.11687
R45162 ASIG5V.n4096 ASIG5V.n4086 1.11687
R45163 ASIG5V.n4277 ASIG5V.n4231 1.11687
R45164 ASIG5V.n4096 ASIG5V.n4085 1.11687
R45165 ASIG5V.n4096 ASIG5V.n4082 1.11687
R45166 ASIG5V.n4096 ASIG5V.n4079 1.11687
R45167 ASIG5V.n4277 ASIG5V.n4234 1.11687
R45168 ASIG5V.n4096 ASIG5V.n4078 1.11687
R45169 ASIG5V.n4277 ASIG5V.n4239 1.11687
R45170 ASIG5V.n4096 ASIG5V.n4075 1.11687
R45171 ASIG5V.n4096 ASIG5V.n4074 1.11687
R45172 ASIG5V.n4277 ASIG5V.n4242 1.11687
R45173 ASIG5V.n4096 ASIG5V.n4071 1.11687
R45174 ASIG5V.n4277 ASIG5V.n4245 1.11687
R45175 ASIG5V.n4096 ASIG5V.n4068 1.11687
R45176 ASIG5V.n4096 ASIG5V.n4065 1.11687
R45177 ASIG5V.n4096 ASIG5V.n4062 1.11687
R45178 ASIG5V.n4277 ASIG5V.n4248 1.11687
R45179 ASIG5V.n4096 ASIG5V.n4059 1.11687
R45180 ASIG5V.n4277 ASIG5V.n4252 1.11687
R45181 ASIG5V.n4096 ASIG5V.n4056 1.11687
R45182 ASIG5V.n4096 ASIG5V.n4052 1.11687
R45183 ASIG5V.n4277 ASIG5V.n4256 1.11687
R45184 ASIG5V.n4096 ASIG5V.n4048 1.11687
R45185 ASIG5V.n4277 ASIG5V.n4260 1.11687
R45186 ASIG5V.n4096 ASIG5V.n4044 1.11687
R45187 ASIG5V.n4096 ASIG5V.n4040 1.11687
R45188 ASIG5V.n4096 ASIG5V.n4036 1.11687
R45189 ASIG5V.n4277 ASIG5V.n4263 1.11687
R45190 ASIG5V.n4096 ASIG5V.n4033 1.11687
R45191 ASIG5V.n4277 ASIG5V.n4266 1.11687
R45192 ASIG5V.n4096 ASIG5V.n4030 1.11687
R45193 ASIG5V.n4096 ASIG5V.n4027 1.11687
R45194 ASIG5V.n4277 ASIG5V.n4271 1.11687
R45195 ASIG5V.n4096 ASIG5V.n4024 1.11687
R45196 ASIG5V.n4277 ASIG5V.n4274 1.11687
R45197 ASIG5V.n4096 ASIG5V.n4023 1.11687
R45198 ASIG5V.n4096 ASIG5V.n4020 1.11687
R45199 ASIG5V.n4096 ASIG5V.n4017 1.11687
R45200 ASIG5V.n4277 ASIG5V.n4276 1.11687
R45201 ASIG5V.n4096 ASIG5V.n4014 1.11687
R45202 ASIG5V.n4375 ASIG5V.n4373 1.11687
R45203 ASIG5V.n4561 ASIG5V.n4503 1.11687
R45204 ASIG5V.n4375 ASIG5V.n4372 1.11687
R45205 ASIG5V.n4561 ASIG5V.n4506 1.11687
R45206 ASIG5V.n4375 ASIG5V.n4371 1.11687
R45207 ASIG5V.n4375 ASIG5V.n4370 1.11687
R45208 ASIG5V.n4561 ASIG5V.n4508 1.11687
R45209 ASIG5V.n4375 ASIG5V.n4368 1.11687
R45210 ASIG5V.n4561 ASIG5V.n4510 1.11687
R45211 ASIG5V.n4375 ASIG5V.n4366 1.11687
R45212 ASIG5V.n4375 ASIG5V.n4364 1.11687
R45213 ASIG5V.n4375 ASIG5V.n4362 1.11687
R45214 ASIG5V.n4561 ASIG5V.n4512 1.11687
R45215 ASIG5V.n4375 ASIG5V.n4360 1.11687
R45216 ASIG5V.n4375 ASIG5V.n4357 1.11687
R45217 ASIG5V.n4375 ASIG5V.n4354 1.11687
R45218 ASIG5V.n4561 ASIG5V.n4515 1.11687
R45219 ASIG5V.n4375 ASIG5V.n4353 1.11687
R45220 ASIG5V.n4561 ASIG5V.n4518 1.11687
R45221 ASIG5V.n4375 ASIG5V.n4350 1.11687
R45222 ASIG5V.n4375 ASIG5V.n4347 1.11687
R45223 ASIG5V.n4561 ASIG5V.n4521 1.11687
R45224 ASIG5V.n4375 ASIG5V.n4344 1.11687
R45225 ASIG5V.n4561 ASIG5V.n4524 1.11687
R45226 ASIG5V.n4375 ASIG5V.n4341 1.11687
R45227 ASIG5V.n4375 ASIG5V.n4338 1.11687
R45228 ASIG5V.n4375 ASIG5V.n4335 1.11687
R45229 ASIG5V.n4561 ASIG5V.n4531 1.11687
R45230 ASIG5V.n4375 ASIG5V.n4332 1.11687
R45231 ASIG5V.n4561 ASIG5V.n4535 1.11687
R45232 ASIG5V.n4375 ASIG5V.n4331 1.11687
R45233 ASIG5V.n4375 ASIG5V.n4327 1.11687
R45234 ASIG5V.n4561 ASIG5V.n4539 1.11687
R45235 ASIG5V.n4375 ASIG5V.n4323 1.11687
R45236 ASIG5V.n4561 ASIG5V.n4543 1.11687
R45237 ASIG5V.n4375 ASIG5V.n4319 1.11687
R45238 ASIG5V.n4375 ASIG5V.n4315 1.11687
R45239 ASIG5V.n4375 ASIG5V.n4311 1.11687
R45240 ASIG5V.n4561 ASIG5V.n4546 1.11687
R45241 ASIG5V.n4375 ASIG5V.n4307 1.11687
R45242 ASIG5V.n4561 ASIG5V.n4549 1.11687
R45243 ASIG5V.n4375 ASIG5V.n4304 1.11687
R45244 ASIG5V.n4375 ASIG5V.n4301 1.11687
R45245 ASIG5V.n4561 ASIG5V.n4552 1.11687
R45246 ASIG5V.n4375 ASIG5V.n4298 1.11687
R45247 ASIG5V.n4561 ASIG5V.n4555 1.11687
R45248 ASIG5V.n4375 ASIG5V.n4295 1.11687
R45249 ASIG5V.n4375 ASIG5V.n4292 1.11687
R45250 ASIG5V.n4375 ASIG5V.n4291 1.11687
R45251 ASIG5V.n4561 ASIG5V.n4560 1.11687
R45252 ASIG5V.n4375 ASIG5V.n4288 1.11687
R45253 ASIG5V.n4630 ASIG5V.n4628 1.11687
R45254 ASIG5V.n4847 ASIG5V.n4770 1.11687
R45255 ASIG5V.n4630 ASIG5V.n4627 1.11687
R45256 ASIG5V.n4847 ASIG5V.n4773 1.11687
R45257 ASIG5V.n4630 ASIG5V.n4626 1.11687
R45258 ASIG5V.n4630 ASIG5V.n4625 1.11687
R45259 ASIG5V.n4847 ASIG5V.n4776 1.11687
R45260 ASIG5V.n4630 ASIG5V.n4624 1.11687
R45261 ASIG5V.n4847 ASIG5V.n4779 1.11687
R45262 ASIG5V.n4630 ASIG5V.n4623 1.11687
R45263 ASIG5V.n4630 ASIG5V.n4622 1.11687
R45264 ASIG5V.n4630 ASIG5V.n4621 1.11687
R45265 ASIG5V.n4847 ASIG5V.n4783 1.11687
R45266 ASIG5V.n4630 ASIG5V.n4620 1.11687
R45267 ASIG5V.n4630 ASIG5V.n4619 1.11687
R45268 ASIG5V.n4630 ASIG5V.n4618 1.11687
R45269 ASIG5V.n4847 ASIG5V.n4788 1.11687
R45270 ASIG5V.n4630 ASIG5V.n4617 1.11687
R45271 ASIG5V.n4847 ASIG5V.n4793 1.11687
R45272 ASIG5V.n4630 ASIG5V.n4616 1.11687
R45273 ASIG5V.n4630 ASIG5V.n4615 1.11687
R45274 ASIG5V.n4847 ASIG5V.n4796 1.11687
R45275 ASIG5V.n4630 ASIG5V.n4614 1.11687
R45276 ASIG5V.n4847 ASIG5V.n4801 1.11687
R45277 ASIG5V.n4630 ASIG5V.n4611 1.11687
R45278 ASIG5V.n4630 ASIG5V.n4610 1.11687
R45279 ASIG5V.n4630 ASIG5V.n4609 1.11687
R45280 ASIG5V.n4847 ASIG5V.n4808 1.11687
R45281 ASIG5V.n4630 ASIG5V.n4605 1.11687
R45282 ASIG5V.n4847 ASIG5V.n4812 1.11687
R45283 ASIG5V.n4630 ASIG5V.n4604 1.11687
R45284 ASIG5V.n4630 ASIG5V.n4597 1.11687
R45285 ASIG5V.n4847 ASIG5V.n4819 1.11687
R45286 ASIG5V.n4630 ASIG5V.n4593 1.11687
R45287 ASIG5V.n4847 ASIG5V.n4826 1.11687
R45288 ASIG5V.n4630 ASIG5V.n4592 1.11687
R45289 ASIG5V.n4630 ASIG5V.n4591 1.11687
R45290 ASIG5V.n4630 ASIG5V.n4590 1.11687
R45291 ASIG5V.n4847 ASIG5V.n4830 1.11687
R45292 ASIG5V.n4630 ASIG5V.n4586 1.11687
R45293 ASIG5V.n4847 ASIG5V.n4835 1.11687
R45294 ASIG5V.n4630 ASIG5V.n4582 1.11687
R45295 ASIG5V.n4630 ASIG5V.n4581 1.11687
R45296 ASIG5V.n4847 ASIG5V.n4840 1.11687
R45297 ASIG5V.n4630 ASIG5V.n4580 1.11687
R45298 ASIG5V.n4847 ASIG5V.n4843 1.11687
R45299 ASIG5V.n4630 ASIG5V.n4579 1.11687
R45300 ASIG5V.n4630 ASIG5V.n4576 1.11687
R45301 ASIG5V.n4630 ASIG5V.n4575 1.11687
R45302 ASIG5V.n4847 ASIG5V.n4846 1.11687
R45303 ASIG5V.n4630 ASIG5V.n4574 1.11687
R45304 ASIG5V.n4901 ASIG5V.n4899 1.11687
R45305 ASIG5V.n5142 ASIG5V.n5060 1.11687
R45306 ASIG5V.n4901 ASIG5V.n4898 1.11687
R45307 ASIG5V.n5142 ASIG5V.n5063 1.11687
R45308 ASIG5V.n4901 ASIG5V.n4897 1.11687
R45309 ASIG5V.n4901 ASIG5V.n4896 1.11687
R45310 ASIG5V.n5142 ASIG5V.n5066 1.11687
R45311 ASIG5V.n4901 ASIG5V.n4895 1.11687
R45312 ASIG5V.n5142 ASIG5V.n5069 1.11687
R45313 ASIG5V.n4901 ASIG5V.n4894 1.11687
R45314 ASIG5V.n4901 ASIG5V.n4893 1.11687
R45315 ASIG5V.n4901 ASIG5V.n4892 1.11687
R45316 ASIG5V.n5142 ASIG5V.n5073 1.11687
R45317 ASIG5V.n4901 ASIG5V.n4891 1.11687
R45318 ASIG5V.n4901 ASIG5V.n4890 1.11687
R45319 ASIG5V.n4901 ASIG5V.n4889 1.11687
R45320 ASIG5V.n5142 ASIG5V.n5078 1.11687
R45321 ASIG5V.n4901 ASIG5V.n4888 1.11687
R45322 ASIG5V.n5142 ASIG5V.n5083 1.11687
R45323 ASIG5V.n4901 ASIG5V.n4887 1.11687
R45324 ASIG5V.n4901 ASIG5V.n4886 1.11687
R45325 ASIG5V.n5142 ASIG5V.n5088 1.11687
R45326 ASIG5V.n4901 ASIG5V.n4885 1.11687
R45327 ASIG5V.n5142 ASIG5V.n5093 1.11687
R45328 ASIG5V.n4901 ASIG5V.n4884 1.11687
R45329 ASIG5V.n4901 ASIG5V.n4883 1.11687
R45330 ASIG5V.n4901 ASIG5V.n4882 1.11687
R45331 ASIG5V.n5142 ASIG5V.n5100 1.11687
R45332 ASIG5V.n4901 ASIG5V.n4881 1.11687
R45333 ASIG5V.n5142 ASIG5V.n5107 1.11687
R45334 ASIG5V.n4901 ASIG5V.n4880 1.11687
R45335 ASIG5V.n4901 ASIG5V.n4879 1.11687
R45336 ASIG5V.n5142 ASIG5V.n5114 1.11687
R45337 ASIG5V.n4901 ASIG5V.n4878 1.11687
R45338 ASIG5V.n5142 ASIG5V.n5121 1.11687
R45339 ASIG5V.n4901 ASIG5V.n4877 1.11687
R45340 ASIG5V.n4901 ASIG5V.n4876 1.11687
R45341 ASIG5V.n4901 ASIG5V.n4875 1.11687
R45342 ASIG5V.n5142 ASIG5V.n5128 1.11687
R45343 ASIG5V.n4901 ASIG5V.n4874 1.11687
R45344 ASIG5V.n5142 ASIG5V.n5132 1.11687
R45345 ASIG5V.n4901 ASIG5V.n4873 1.11687
R45346 ASIG5V.n4901 ASIG5V.n4869 1.11687
R45347 ASIG5V.n5142 ASIG5V.n5135 1.11687
R45348 ASIG5V.n4901 ASIG5V.n4868 1.11687
R45349 ASIG5V.n5142 ASIG5V.n5138 1.11687
R45350 ASIG5V.n4901 ASIG5V.n4865 1.11687
R45351 ASIG5V.n4901 ASIG5V.n4862 1.11687
R45352 ASIG5V.n4901 ASIG5V.n4861 1.11687
R45353 ASIG5V.n5142 ASIG5V.n5141 1.11687
R45354 ASIG5V.n4901 ASIG5V.n4860 1.11687
R45355 ASIG5V.n5328 ASIG5V.n5322 1.11687
R45356 ASIG5V.n5442 ASIG5V.n5420 1.11687
R45357 ASIG5V.n5328 ASIG5V.n5319 1.11687
R45358 ASIG5V.n5442 ASIG5V.n5421 1.11687
R45359 ASIG5V.n5328 ASIG5V.n5316 1.11687
R45360 ASIG5V.n5328 ASIG5V.n5313 1.11687
R45361 ASIG5V.n5442 ASIG5V.n5422 1.11687
R45362 ASIG5V.n5328 ASIG5V.n5310 1.11687
R45363 ASIG5V.n5442 ASIG5V.n5423 1.11687
R45364 ASIG5V.n5328 ASIG5V.n5307 1.11687
R45365 ASIG5V.n5328 ASIG5V.n5304 1.11687
R45366 ASIG5V.n5328 ASIG5V.n5301 1.11687
R45367 ASIG5V.n5442 ASIG5V.n5424 1.11687
R45368 ASIG5V.n5328 ASIG5V.n5298 1.11687
R45369 ASIG5V.n5328 ASIG5V.n5293 1.11687
R45370 ASIG5V.n5328 ASIG5V.n5288 1.11687
R45371 ASIG5V.n5442 ASIG5V.n5427 1.11687
R45372 ASIG5V.n5328 ASIG5V.n5285 1.11687
R45373 ASIG5V.n5442 ASIG5V.n5428 1.11687
R45374 ASIG5V.n5328 ASIG5V.n5280 1.11687
R45375 ASIG5V.n5328 ASIG5V.n5275 1.11687
R45376 ASIG5V.n5442 ASIG5V.n5429 1.11687
R45377 ASIG5V.n5328 ASIG5V.n5270 1.11687
R45378 ASIG5V.n5442 ASIG5V.n5430 1.11687
R45379 ASIG5V.n5328 ASIG5V.n5265 1.11687
R45380 ASIG5V.n5328 ASIG5V.n5259 1.11687
R45381 ASIG5V.n5328 ASIG5V.n5252 1.11687
R45382 ASIG5V.n5442 ASIG5V.n5431 1.11687
R45383 ASIG5V.n5328 ASIG5V.n5245 1.11687
R45384 ASIG5V.n5442 ASIG5V.n5432 1.11687
R45385 ASIG5V.n5328 ASIG5V.n5238 1.11687
R45386 ASIG5V.n5328 ASIG5V.n5231 1.11687
R45387 ASIG5V.n5442 ASIG5V.n5433 1.11687
R45388 ASIG5V.n5328 ASIG5V.n5224 1.11687
R45389 ASIG5V.n5442 ASIG5V.n5434 1.11687
R45390 ASIG5V.n5328 ASIG5V.n5217 1.11687
R45391 ASIG5V.n5328 ASIG5V.n5210 1.11687
R45392 ASIG5V.n5328 ASIG5V.n5203 1.11687
R45393 ASIG5V.n5442 ASIG5V.n5435 1.11687
R45394 ASIG5V.n5328 ASIG5V.n5196 1.11687
R45395 ASIG5V.n5442 ASIG5V.n5436 1.11687
R45396 ASIG5V.n5328 ASIG5V.n5189 1.11687
R45397 ASIG5V.n5328 ASIG5V.n5182 1.11687
R45398 ASIG5V.n5442 ASIG5V.n5437 1.11687
R45399 ASIG5V.n5328 ASIG5V.n5175 1.11687
R45400 ASIG5V.n5442 ASIG5V.n5438 1.11687
R45401 ASIG5V.n5328 ASIG5V.n5170 1.11687
R45402 ASIG5V.n5328 ASIG5V.n5165 1.11687
R45403 ASIG5V.n5328 ASIG5V.n5160 1.11687
R45404 ASIG5V.n5442 ASIG5V.n5441 1.11687
R45405 ASIG5V.n5328 ASIG5V.n5155 1.11687
R45406 ASIG5V.n5559 ASIG5V.n5557 1.11687
R45407 ASIG5V.n5793 ASIG5V.n5737 1.11687
R45408 ASIG5V.n5559 ASIG5V.n5555 1.11687
R45409 ASIG5V.n5793 ASIG5V.n5739 1.11687
R45410 ASIG5V.n5559 ASIG5V.n5553 1.11687
R45411 ASIG5V.n5559 ASIG5V.n5551 1.11687
R45412 ASIG5V.n5793 ASIG5V.n5741 1.11687
R45413 ASIG5V.n5559 ASIG5V.n5550 1.11687
R45414 ASIG5V.n5793 ASIG5V.n5743 1.11687
R45415 ASIG5V.n5559 ASIG5V.n5548 1.11687
R45416 ASIG5V.n5559 ASIG5V.n5545 1.11687
R45417 ASIG5V.n5559 ASIG5V.n5542 1.11687
R45418 ASIG5V.n5793 ASIG5V.n5745 1.11687
R45419 ASIG5V.n5559 ASIG5V.n5540 1.11687
R45420 ASIG5V.n5559 ASIG5V.n5537 1.11687
R45421 ASIG5V.n5559 ASIG5V.n5534 1.11687
R45422 ASIG5V.n5793 ASIG5V.n5748 1.11687
R45423 ASIG5V.n5559 ASIG5V.n5531 1.11687
R45424 ASIG5V.n5793 ASIG5V.n5751 1.11687
R45425 ASIG5V.n5559 ASIG5V.n5528 1.11687
R45426 ASIG5V.n5559 ASIG5V.n5525 1.11687
R45427 ASIG5V.n5793 ASIG5V.n5754 1.11687
R45428 ASIG5V.n5559 ASIG5V.n5522 1.11687
R45429 ASIG5V.n5793 ASIG5V.n5757 1.11687
R45430 ASIG5V.n5559 ASIG5V.n5519 1.11687
R45431 ASIG5V.n5559 ASIG5V.n5515 1.11687
R45432 ASIG5V.n5559 ASIG5V.n5511 1.11687
R45433 ASIG5V.n5793 ASIG5V.n5761 1.11687
R45434 ASIG5V.n5559 ASIG5V.n5507 1.11687
R45435 ASIG5V.n5793 ASIG5V.n5765 1.11687
R45436 ASIG5V.n5559 ASIG5V.n5503 1.11687
R45437 ASIG5V.n5559 ASIG5V.n5499 1.11687
R45438 ASIG5V.n5793 ASIG5V.n5772 1.11687
R45439 ASIG5V.n5559 ASIG5V.n5495 1.11687
R45440 ASIG5V.n5793 ASIG5V.n5779 1.11687
R45441 ASIG5V.n5559 ASIG5V.n5494 1.11687
R45442 ASIG5V.n5559 ASIG5V.n5493 1.11687
R45443 ASIG5V.n5559 ASIG5V.n5489 1.11687
R45444 ASIG5V.n5793 ASIG5V.n5780 1.11687
R45445 ASIG5V.n5559 ASIG5V.n5482 1.11687
R45446 ASIG5V.n5793 ASIG5V.n5784 1.11687
R45447 ASIG5V.n5559 ASIG5V.n5478 1.11687
R45448 ASIG5V.n5559 ASIG5V.n5474 1.11687
R45449 ASIG5V.n5793 ASIG5V.n5788 1.11687
R45450 ASIG5V.n5559 ASIG5V.n5470 1.11687
R45451 ASIG5V.n5793 ASIG5V.n5789 1.11687
R45452 ASIG5V.n5559 ASIG5V.n5463 1.11687
R45453 ASIG5V.n5559 ASIG5V.n5460 1.11687
R45454 ASIG5V.n5559 ASIG5V.n5459 1.11687
R45455 ASIG5V.n5793 ASIG5V.n5792 1.11687
R45456 ASIG5V.n5559 ASIG5V.n5458 1.11687
R45457 ASIG5V.n5855 ASIG5V.n5853 1.11687
R45458 ASIG5V.n6149 ASIG5V.n6065 1.11687
R45459 ASIG5V.n5855 ASIG5V.n5852 1.11687
R45460 ASIG5V.n6149 ASIG5V.n6068 1.11687
R45461 ASIG5V.n5855 ASIG5V.n5851 1.11687
R45462 ASIG5V.n5855 ASIG5V.n5850 1.11687
R45463 ASIG5V.n6149 ASIG5V.n6071 1.11687
R45464 ASIG5V.n5855 ASIG5V.n5849 1.11687
R45465 ASIG5V.n6149 ASIG5V.n6074 1.11687
R45466 ASIG5V.n5855 ASIG5V.n5848 1.11687
R45467 ASIG5V.n5855 ASIG5V.n5847 1.11687
R45468 ASIG5V.n5855 ASIG5V.n5846 1.11687
R45469 ASIG5V.n6149 ASIG5V.n6078 1.11687
R45470 ASIG5V.n5855 ASIG5V.n5845 1.11687
R45471 ASIG5V.n5855 ASIG5V.n5844 1.11687
R45472 ASIG5V.n5855 ASIG5V.n5843 1.11687
R45473 ASIG5V.n6149 ASIG5V.n6083 1.11687
R45474 ASIG5V.n5855 ASIG5V.n5842 1.11687
R45475 ASIG5V.n6149 ASIG5V.n6088 1.11687
R45476 ASIG5V.n5855 ASIG5V.n5841 1.11687
R45477 ASIG5V.n5855 ASIG5V.n5840 1.11687
R45478 ASIG5V.n6149 ASIG5V.n6093 1.11687
R45479 ASIG5V.n5855 ASIG5V.n5839 1.11687
R45480 ASIG5V.n6149 ASIG5V.n6099 1.11687
R45481 ASIG5V.n5855 ASIG5V.n5838 1.11687
R45482 ASIG5V.n5855 ASIG5V.n5837 1.11687
R45483 ASIG5V.n5855 ASIG5V.n5836 1.11687
R45484 ASIG5V.n6149 ASIG5V.n6106 1.11687
R45485 ASIG5V.n5855 ASIG5V.n5835 1.11687
R45486 ASIG5V.n6149 ASIG5V.n6113 1.11687
R45487 ASIG5V.n5855 ASIG5V.n5834 1.11687
R45488 ASIG5V.n5855 ASIG5V.n5833 1.11687
R45489 ASIG5V.n6149 ASIG5V.n6120 1.11687
R45490 ASIG5V.n5855 ASIG5V.n5832 1.11687
R45491 ASIG5V.n6149 ASIG5V.n6127 1.11687
R45492 ASIG5V.n5855 ASIG5V.n5831 1.11687
R45493 ASIG5V.n5855 ASIG5V.n5830 1.11687
R45494 ASIG5V.n5855 ASIG5V.n5829 1.11687
R45495 ASIG5V.n6149 ASIG5V.n6134 1.11687
R45496 ASIG5V.n5855 ASIG5V.n5828 1.11687
R45497 ASIG5V.n6149 ASIG5V.n6135 1.11687
R45498 ASIG5V.n5855 ASIG5V.n5824 1.11687
R45499 ASIG5V.n5855 ASIG5V.n5820 1.11687
R45500 ASIG5V.n6149 ASIG5V.n6142 1.11687
R45501 ASIG5V.n5855 ASIG5V.n5819 1.11687
R45502 ASIG5V.n6149 ASIG5V.n6143 1.11687
R45503 ASIG5V.n5855 ASIG5V.n5815 1.11687
R45504 ASIG5V.n5855 ASIG5V.n5811 1.11687
R45505 ASIG5V.n5855 ASIG5V.n5810 1.11687
R45506 ASIG5V.n6149 ASIG5V.n6148 1.11687
R45507 ASIG5V.n5855 ASIG5V.n5809 1.11687
R45508 ASIG5V.n6326 ASIG5V.n6320 1.11687
R45509 ASIG5V.n7123 ASIG5V.n7097 1.11687
R45510 ASIG5V.n6326 ASIG5V.n6317 1.11687
R45511 ASIG5V.n7123 ASIG5V.n7098 1.11687
R45512 ASIG5V.n6326 ASIG5V.n6314 1.11687
R45513 ASIG5V.n6326 ASIG5V.n6311 1.11687
R45514 ASIG5V.n7123 ASIG5V.n7099 1.11687
R45515 ASIG5V.n6326 ASIG5V.n6308 1.11687
R45516 ASIG5V.n7123 ASIG5V.n7100 1.11687
R45517 ASIG5V.n6326 ASIG5V.n6305 1.11687
R45518 ASIG5V.n6326 ASIG5V.n6302 1.11687
R45519 ASIG5V.n6326 ASIG5V.n6299 1.11687
R45520 ASIG5V.n7123 ASIG5V.n7101 1.11687
R45521 ASIG5V.n6326 ASIG5V.n6296 1.11687
R45522 ASIG5V.n6326 ASIG5V.n6291 1.11687
R45523 ASIG5V.n6326 ASIG5V.n6286 1.11687
R45524 ASIG5V.n7123 ASIG5V.n7102 1.11687
R45525 ASIG5V.n6326 ASIG5V.n6281 1.11687
R45526 ASIG5V.n7123 ASIG5V.n7103 1.11687
R45527 ASIG5V.n6326 ASIG5V.n6276 1.11687
R45528 ASIG5V.n6326 ASIG5V.n6271 1.11687
R45529 ASIG5V.n7123 ASIG5V.n7104 1.11687
R45530 ASIG5V.n6326 ASIG5V.n6266 1.11687
R45531 ASIG5V.n7123 ASIG5V.n7105 1.11687
R45532 ASIG5V.n6326 ASIG5V.n6261 1.11687
R45533 ASIG5V.n6326 ASIG5V.n6254 1.11687
R45534 ASIG5V.n6326 ASIG5V.n6247 1.11687
R45535 ASIG5V.n7123 ASIG5V.n7106 1.11687
R45536 ASIG5V.n6326 ASIG5V.n6240 1.11687
R45537 ASIG5V.n7123 ASIG5V.n7107 1.11687
R45538 ASIG5V.n6326 ASIG5V.n6233 1.11687
R45539 ASIG5V.n6326 ASIG5V.n6226 1.11687
R45540 ASIG5V.n7123 ASIG5V.n7108 1.11687
R45541 ASIG5V.n6326 ASIG5V.n6219 1.11687
R45542 ASIG5V.n7123 ASIG5V.n7109 1.11687
R45543 ASIG5V.n6326 ASIG5V.n6212 1.11687
R45544 ASIG5V.n6326 ASIG5V.n6205 1.11687
R45545 ASIG5V.n6326 ASIG5V.n6198 1.11687
R45546 ASIG5V.n7123 ASIG5V.n7113 1.11687
R45547 ASIG5V.n6326 ASIG5V.n6197 1.11687
R45548 ASIG5V.n7123 ASIG5V.n7117 1.11687
R45549 ASIG5V.n6326 ASIG5V.n6193 1.11687
R45550 ASIG5V.n6326 ASIG5V.n6189 1.11687
R45551 ASIG5V.n7123 ASIG5V.n7118 1.11687
R45552 ASIG5V.n6326 ASIG5V.n6185 1.11687
R45553 ASIG5V.n7123 ASIG5V.n7119 1.11687
R45554 ASIG5V.n6326 ASIG5V.n6178 1.11687
R45555 ASIG5V.n6326 ASIG5V.n6174 1.11687
R45556 ASIG5V.n6326 ASIG5V.n6170 1.11687
R45557 ASIG5V.n7123 ASIG5V.n7122 1.11687
R45558 ASIG5V.n6326 ASIG5V.n6166 1.11687
R45559 ASIG5V.n7052 ASIG5V.n6415 1.11687
R45560 ASIG5V.n6928 ASIG5V.n6831 1.11687
R45561 ASIG5V.n7052 ASIG5V.n6413 1.11687
R45562 ASIG5V.n6928 ASIG5V.n6834 1.11687
R45563 ASIG5V.n7052 ASIG5V.n6412 1.11687
R45564 ASIG5V.n7052 ASIG5V.n6410 1.11687
R45565 ASIG5V.n6928 ASIG5V.n6837 1.11687
R45566 ASIG5V.n7052 ASIG5V.n6408 1.11687
R45567 ASIG5V.n6928 ASIG5V.n6840 1.11687
R45568 ASIG5V.n7052 ASIG5V.n6407 1.11687
R45569 ASIG5V.n7052 ASIG5V.n6406 1.11687
R45570 ASIG5V.n7052 ASIG5V.n6404 1.11687
R45571 ASIG5V.n6928 ASIG5V.n6844 1.11687
R45572 ASIG5V.n7052 ASIG5V.n6402 1.11687
R45573 ASIG5V.n7052 ASIG5V.n6399 1.11687
R45574 ASIG5V.n7052 ASIG5V.n6396 1.11687
R45575 ASIG5V.n6928 ASIG5V.n6849 1.11687
R45576 ASIG5V.n7052 ASIG5V.n6393 1.11687
R45577 ASIG5V.n6928 ASIG5V.n6854 1.11687
R45578 ASIG5V.n7052 ASIG5V.n6392 1.11687
R45579 ASIG5V.n7052 ASIG5V.n6389 1.11687
R45580 ASIG5V.n6928 ASIG5V.n6859 1.11687
R45581 ASIG5V.n7052 ASIG5V.n6386 1.11687
R45582 ASIG5V.n6928 ASIG5V.n6864 1.11687
R45583 ASIG5V.n7052 ASIG5V.n6385 1.11687
R45584 ASIG5V.n7052 ASIG5V.n6384 1.11687
R45585 ASIG5V.n7052 ASIG5V.n6380 1.11687
R45586 ASIG5V.n6928 ASIG5V.n6871 1.11687
R45587 ASIG5V.n7052 ASIG5V.n6376 1.11687
R45588 ASIG5V.n6928 ASIG5V.n6878 1.11687
R45589 ASIG5V.n7052 ASIG5V.n6375 1.11687
R45590 ASIG5V.n7052 ASIG5V.n6374 1.11687
R45591 ASIG5V.n6928 ASIG5V.n6885 1.11687
R45592 ASIG5V.n7052 ASIG5V.n6370 1.11687
R45593 ASIG5V.n6928 ASIG5V.n6892 1.11687
R45594 ASIG5V.n7052 ASIG5V.n6369 1.11687
R45595 ASIG5V.n7052 ASIG5V.n6368 1.11687
R45596 ASIG5V.n7052 ASIG5V.n6361 1.11687
R45597 ASIG5V.n6928 ASIG5V.n6899 1.11687
R45598 ASIG5V.n7052 ASIG5V.n6357 1.11687
R45599 ASIG5V.n6928 ASIG5V.n6906 1.11687
R45600 ASIG5V.n7052 ASIG5V.n6356 1.11687
R45601 ASIG5V.n7052 ASIG5V.n6352 1.11687
R45602 ASIG5V.n6928 ASIG5V.n6913 1.11687
R45603 ASIG5V.n7052 ASIG5V.n6348 1.11687
R45604 ASIG5V.n6928 ASIG5V.n6920 1.11687
R45605 ASIG5V.n7052 ASIG5V.n6347 1.11687
R45606 ASIG5V.n7052 ASIG5V.n6346 1.11687
R45607 ASIG5V.n7052 ASIG5V.n6342 1.11687
R45608 ASIG5V.n6928 ASIG5V.n6927 1.11687
R45609 ASIG5V.n7052 ASIG5V.n6338 1.11687
R45610 ASIG5V.n6777 ASIG5V.n6545 1.11687
R45611 ASIG5V.n6652 ASIG5V.n6618 1.11687
R45612 ASIG5V.n6777 ASIG5V.n6543 1.11687
R45613 ASIG5V.n6652 ASIG5V.n6621 1.11687
R45614 ASIG5V.n6777 ASIG5V.n6542 1.11687
R45615 ASIG5V.n6777 ASIG5V.n6540 1.11687
R45616 ASIG5V.n6652 ASIG5V.n6624 1.11687
R45617 ASIG5V.n6777 ASIG5V.n6538 1.11687
R45618 ASIG5V.n6652 ASIG5V.n6627 1.11687
R45619 ASIG5V.n6777 ASIG5V.n6537 1.11687
R45620 ASIG5V.n6777 ASIG5V.n6536 1.11687
R45621 ASIG5V.n6777 ASIG5V.n6533 1.11687
R45622 ASIG5V.n6652 ASIG5V.n6629 1.11687
R45623 ASIG5V.n6777 ASIG5V.n6531 1.11687
R45624 ASIG5V.n6777 ASIG5V.n6528 1.11687
R45625 ASIG5V.n6777 ASIG5V.n6523 1.11687
R45626 ASIG5V.n6652 ASIG5V.n6632 1.11687
R45627 ASIG5V.n6777 ASIG5V.n6520 1.11687
R45628 ASIG5V.n6652 ASIG5V.n6635 1.11687
R45629 ASIG5V.n6777 ASIG5V.n6517 1.11687
R45630 ASIG5V.n6777 ASIG5V.n6514 1.11687
R45631 ASIG5V.n6652 ASIG5V.n6638 1.11687
R45632 ASIG5V.n6777 ASIG5V.n6511 1.11687
R45633 ASIG5V.n6652 ASIG5V.n6639 1.11687
R45634 ASIG5V.n6777 ASIG5V.n6506 1.11687
R45635 ASIG5V.n6777 ASIG5V.n6502 1.11687
R45636 ASIG5V.n6777 ASIG5V.n6498 1.11687
R45637 ASIG5V.n6652 ASIG5V.n6640 1.11687
R45638 ASIG5V.n6777 ASIG5V.n6491 1.11687
R45639 ASIG5V.n6652 ASIG5V.n6641 1.11687
R45640 ASIG5V.n6777 ASIG5V.n6484 1.11687
R45641 ASIG5V.n6777 ASIG5V.n6480 1.11687
R45642 ASIG5V.n6652 ASIG5V.n6645 1.11687
R45643 ASIG5V.n6777 ASIG5V.n6479 1.11687
R45644 ASIG5V.n6652 ASIG5V.n6646 1.11687
R45645 ASIG5V.n6777 ASIG5V.n6472 1.11687
R45646 ASIG5V.n6777 ASIG5V.n6468 1.11687
R45647 ASIG5V.n6777 ASIG5V.n6467 1.11687
R45648 ASIG5V.n6652 ASIG5V.n6647 1.11687
R45649 ASIG5V.n6777 ASIG5V.n6463 1.11687
R45650 ASIG5V.n6652 ASIG5V.n6648 1.11687
R45651 ASIG5V.n6777 ASIG5V.n6456 1.11687
R45652 ASIG5V.n6777 ASIG5V.n6452 1.11687
R45653 ASIG5V.n6652 ASIG5V.n6649 1.11687
R45654 ASIG5V.n6777 ASIG5V.n6448 1.11687
R45655 ASIG5V.n6652 ASIG5V.n6650 1.11687
R45656 ASIG5V.n6777 ASIG5V.n6441 1.11687
R45657 ASIG5V.n6777 ASIG5V.n6437 1.11687
R45658 ASIG5V.n6777 ASIG5V.n6433 1.11687
R45659 ASIG5V.n6652 ASIG5V.n6651 1.11687
R45660 ASIG5V.n6777 ASIG5V.n6429 1.11687
R45661 ASIG5V.n13618 ASIG5V.n98 1.11687
R45662 ASIG5V.n13495 ASIG5V.n13409 1.11687
R45663 ASIG5V.n13618 ASIG5V.n95 1.11687
R45664 ASIG5V.n13495 ASIG5V.n13410 1.11687
R45665 ASIG5V.n13618 ASIG5V.n92 1.11687
R45666 ASIG5V.n13618 ASIG5V.n89 1.11687
R45667 ASIG5V.n13495 ASIG5V.n13411 1.11687
R45668 ASIG5V.n13618 ASIG5V.n86 1.11687
R45669 ASIG5V.n13495 ASIG5V.n13412 1.11687
R45670 ASIG5V.n13618 ASIG5V.n83 1.11687
R45671 ASIG5V.n13618 ASIG5V.n80 1.11687
R45672 ASIG5V.n13618 ASIG5V.n78 1.11687
R45673 ASIG5V.n13495 ASIG5V.n13416 1.11687
R45674 ASIG5V.n13618 ASIG5V.n76 1.11687
R45675 ASIG5V.n13618 ASIG5V.n75 1.11687
R45676 ASIG5V.n13618 ASIG5V.n72 1.11687
R45677 ASIG5V.n13495 ASIG5V.n13419 1.11687
R45678 ASIG5V.n13618 ASIG5V.n69 1.11687
R45679 ASIG5V.n13495 ASIG5V.n13422 1.11687
R45680 ASIG5V.n13618 ASIG5V.n66 1.11687
R45681 ASIG5V.n13618 ASIG5V.n63 1.11687
R45682 ASIG5V.n13495 ASIG5V.n13425 1.11687
R45683 ASIG5V.n13618 ASIG5V.n60 1.11687
R45684 ASIG5V.n13495 ASIG5V.n13431 1.11687
R45685 ASIG5V.n13618 ASIG5V.n57 1.11687
R45686 ASIG5V.n13618 ASIG5V.n53 1.11687
R45687 ASIG5V.n13618 ASIG5V.n49 1.11687
R45688 ASIG5V.n13495 ASIG5V.n13438 1.11687
R45689 ASIG5V.n13618 ASIG5V.n45 1.11687
R45690 ASIG5V.n13495 ASIG5V.n13445 1.11687
R45691 ASIG5V.n13618 ASIG5V.n44 1.11687
R45692 ASIG5V.n13618 ASIG5V.n40 1.11687
R45693 ASIG5V.n13495 ASIG5V.n13452 1.11687
R45694 ASIG5V.n13618 ASIG5V.n36 1.11687
R45695 ASIG5V.n13495 ASIG5V.n13459 1.11687
R45696 ASIG5V.n13618 ASIG5V.n35 1.11687
R45697 ASIG5V.n13618 ASIG5V.n34 1.11687
R45698 ASIG5V.n13618 ASIG5V.n33 1.11687
R45699 ASIG5V.n13495 ASIG5V.n13466 1.11687
R45700 ASIG5V.n13618 ASIG5V.n29 1.11687
R45701 ASIG5V.n13495 ASIG5V.n13473 1.11687
R45702 ASIG5V.n13618 ASIG5V.n28 1.11687
R45703 ASIG5V.n13618 ASIG5V.n24 1.11687
R45704 ASIG5V.n13495 ASIG5V.n13480 1.11687
R45705 ASIG5V.n13618 ASIG5V.n20 1.11687
R45706 ASIG5V.n13495 ASIG5V.n13487 1.11687
R45707 ASIG5V.n13618 ASIG5V.n19 1.11687
R45708 ASIG5V.n13618 ASIG5V.n15 1.11687
R45709 ASIG5V.n13618 ASIG5V.n11 1.11687
R45710 ASIG5V.n13495 ASIG5V.n13494 1.11687
R45711 ASIG5V.n13618 ASIG5V.n7 1.11687
R45712 ASIG5V.n13360 ASIG5V.n139 1.11687
R45713 ASIG5V.n331 ASIG5V.n234 1.11687
R45714 ASIG5V.n13360 ASIG5V.n138 1.11687
R45715 ASIG5V.n331 ASIG5V.n237 1.11687
R45716 ASIG5V.n13360 ASIG5V.n137 1.11687
R45717 ASIG5V.n13360 ASIG5V.n136 1.11687
R45718 ASIG5V.n331 ASIG5V.n240 1.11687
R45719 ASIG5V.n13360 ASIG5V.n135 1.11687
R45720 ASIG5V.n331 ASIG5V.n243 1.11687
R45721 ASIG5V.n13360 ASIG5V.n134 1.11687
R45722 ASIG5V.n13360 ASIG5V.n133 1.11687
R45723 ASIG5V.n13360 ASIG5V.n132 1.11687
R45724 ASIG5V.n331 ASIG5V.n247 1.11687
R45725 ASIG5V.n13360 ASIG5V.n131 1.11687
R45726 ASIG5V.n13360 ASIG5V.n130 1.11687
R45727 ASIG5V.n13360 ASIG5V.n129 1.11687
R45728 ASIG5V.n331 ASIG5V.n252 1.11687
R45729 ASIG5V.n13360 ASIG5V.n128 1.11687
R45730 ASIG5V.n331 ASIG5V.n257 1.11687
R45731 ASIG5V.n13360 ASIG5V.n127 1.11687
R45732 ASIG5V.n13360 ASIG5V.n126 1.11687
R45733 ASIG5V.n331 ASIG5V.n262 1.11687
R45734 ASIG5V.n13360 ASIG5V.n125 1.11687
R45735 ASIG5V.n331 ASIG5V.n268 1.11687
R45736 ASIG5V.n13360 ASIG5V.n124 1.11687
R45737 ASIG5V.n13360 ASIG5V.n123 1.11687
R45738 ASIG5V.n13360 ASIG5V.n122 1.11687
R45739 ASIG5V.n331 ASIG5V.n275 1.11687
R45740 ASIG5V.n13360 ASIG5V.n121 1.11687
R45741 ASIG5V.n331 ASIG5V.n282 1.11687
R45742 ASIG5V.n13360 ASIG5V.n120 1.11687
R45743 ASIG5V.n13360 ASIG5V.n119 1.11687
R45744 ASIG5V.n331 ASIG5V.n289 1.11687
R45745 ASIG5V.n13360 ASIG5V.n118 1.11687
R45746 ASIG5V.n331 ASIG5V.n296 1.11687
R45747 ASIG5V.n13360 ASIG5V.n117 1.11687
R45748 ASIG5V.n13360 ASIG5V.n116 1.11687
R45749 ASIG5V.n13360 ASIG5V.n115 1.11687
R45750 ASIG5V.n331 ASIG5V.n303 1.11687
R45751 ASIG5V.n13360 ASIG5V.n114 1.11687
R45752 ASIG5V.n331 ASIG5V.n310 1.11687
R45753 ASIG5V.n13360 ASIG5V.n113 1.11687
R45754 ASIG5V.n13360 ASIG5V.n112 1.11687
R45755 ASIG5V.n331 ASIG5V.n317 1.11687
R45756 ASIG5V.n13360 ASIG5V.n111 1.11687
R45757 ASIG5V.n331 ASIG5V.n324 1.11687
R45758 ASIG5V.n13360 ASIG5V.n110 1.11687
R45759 ASIG5V.n13360 ASIG5V.n109 1.11687
R45760 ASIG5V.n13360 ASIG5V.n108 1.11687
R45761 ASIG5V.n331 ASIG5V.n330 1.11687
R45762 ASIG5V.n13360 ASIG5V.n107 1.11687
R45763 ASIG5V.n7401 ASIG5V.n7395 1.11687
R45764 ASIG5V.n7626 ASIG5V.n7567 1.11687
R45765 ASIG5V.n7401 ASIG5V.n7393 1.11687
R45766 ASIG5V.n7626 ASIG5V.n7569 1.11687
R45767 ASIG5V.n7401 ASIG5V.n7392 1.11687
R45768 ASIG5V.n7401 ASIG5V.n7389 1.11687
R45769 ASIG5V.n7626 ASIG5V.n7570 1.11687
R45770 ASIG5V.n7401 ASIG5V.n7387 1.11687
R45771 ASIG5V.n7626 ASIG5V.n7572 1.11687
R45772 ASIG5V.n7401 ASIG5V.n7385 1.11687
R45773 ASIG5V.n7401 ASIG5V.n7382 1.11687
R45774 ASIG5V.n7401 ASIG5V.n7379 1.11687
R45775 ASIG5V.n7626 ASIG5V.n7574 1.11687
R45776 ASIG5V.n7401 ASIG5V.n7377 1.11687
R45777 ASIG5V.n7401 ASIG5V.n7374 1.11687
R45778 ASIG5V.n7401 ASIG5V.n7371 1.11687
R45779 ASIG5V.n7626 ASIG5V.n7577 1.11687
R45780 ASIG5V.n7401 ASIG5V.n7368 1.11687
R45781 ASIG5V.n7626 ASIG5V.n7582 1.11687
R45782 ASIG5V.n7401 ASIG5V.n7365 1.11687
R45783 ASIG5V.n7401 ASIG5V.n7364 1.11687
R45784 ASIG5V.n7626 ASIG5V.n7585 1.11687
R45785 ASIG5V.n7401 ASIG5V.n7361 1.11687
R45786 ASIG5V.n7626 ASIG5V.n7590 1.11687
R45787 ASIG5V.n7401 ASIG5V.n7358 1.11687
R45788 ASIG5V.n7401 ASIG5V.n7357 1.11687
R45789 ASIG5V.n7401 ASIG5V.n7353 1.11687
R45790 ASIG5V.n7626 ASIG5V.n7594 1.11687
R45791 ASIG5V.n7401 ASIG5V.n7349 1.11687
R45792 ASIG5V.n7626 ASIG5V.n7601 1.11687
R45793 ASIG5V.n7401 ASIG5V.n7345 1.11687
R45794 ASIG5V.n7401 ASIG5V.n7341 1.11687
R45795 ASIG5V.n7626 ASIG5V.n7605 1.11687
R45796 ASIG5V.n7401 ASIG5V.n7337 1.11687
R45797 ASIG5V.n7626 ASIG5V.n7609 1.11687
R45798 ASIG5V.n7401 ASIG5V.n7333 1.11687
R45799 ASIG5V.n7401 ASIG5V.n7326 1.11687
R45800 ASIG5V.n7401 ASIG5V.n7322 1.11687
R45801 ASIG5V.n7626 ASIG5V.n7613 1.11687
R45802 ASIG5V.n7401 ASIG5V.n7318 1.11687
R45803 ASIG5V.n7626 ASIG5V.n7617 1.11687
R45804 ASIG5V.n7401 ASIG5V.n7314 1.11687
R45805 ASIG5V.n7401 ASIG5V.n7310 1.11687
R45806 ASIG5V.n7626 ASIG5V.n7621 1.11687
R45807 ASIG5V.n7401 ASIG5V.n7306 1.11687
R45808 ASIG5V.n7626 ASIG5V.n7622 1.11687
R45809 ASIG5V.n7401 ASIG5V.n7299 1.11687
R45810 ASIG5V.n7401 ASIG5V.n7295 1.11687
R45811 ASIG5V.n7401 ASIG5V.n7291 1.11687
R45812 ASIG5V.n7626 ASIG5V.n7625 1.11687
R45813 ASIG5V.n7401 ASIG5V.n7288 1.11687
R45814 ASIG5V.n7823 ASIG5V.n7817 1.11687
R45815 ASIG5V.n7979 ASIG5V.n7961 1.11687
R45816 ASIG5V.n7823 ASIG5V.n7814 1.11687
R45817 ASIG5V.n7979 ASIG5V.n7962 1.11687
R45818 ASIG5V.n7823 ASIG5V.n7811 1.11687
R45819 ASIG5V.n7823 ASIG5V.n7808 1.11687
R45820 ASIG5V.n7979 ASIG5V.n7963 1.11687
R45821 ASIG5V.n7823 ASIG5V.n7805 1.11687
R45822 ASIG5V.n7979 ASIG5V.n7964 1.11687
R45823 ASIG5V.n7823 ASIG5V.n7802 1.11687
R45824 ASIG5V.n7823 ASIG5V.n7799 1.11687
R45825 ASIG5V.n7823 ASIG5V.n7796 1.11687
R45826 ASIG5V.n7979 ASIG5V.n7965 1.11687
R45827 ASIG5V.n7823 ASIG5V.n7793 1.11687
R45828 ASIG5V.n7823 ASIG5V.n7788 1.11687
R45829 ASIG5V.n7823 ASIG5V.n7783 1.11687
R45830 ASIG5V.n7979 ASIG5V.n7966 1.11687
R45831 ASIG5V.n7823 ASIG5V.n7778 1.11687
R45832 ASIG5V.n7979 ASIG5V.n7967 1.11687
R45833 ASIG5V.n7823 ASIG5V.n7773 1.11687
R45834 ASIG5V.n7823 ASIG5V.n7768 1.11687
R45835 ASIG5V.n7979 ASIG5V.n7968 1.11687
R45836 ASIG5V.n7823 ASIG5V.n7763 1.11687
R45837 ASIG5V.n7979 ASIG5V.n7969 1.11687
R45838 ASIG5V.n7823 ASIG5V.n7758 1.11687
R45839 ASIG5V.n7823 ASIG5V.n7752 1.11687
R45840 ASIG5V.n7823 ASIG5V.n7745 1.11687
R45841 ASIG5V.n7979 ASIG5V.n7970 1.11687
R45842 ASIG5V.n7823 ASIG5V.n7738 1.11687
R45843 ASIG5V.n7979 ASIG5V.n7971 1.11687
R45844 ASIG5V.n7823 ASIG5V.n7731 1.11687
R45845 ASIG5V.n7823 ASIG5V.n7724 1.11687
R45846 ASIG5V.n7979 ASIG5V.n7972 1.11687
R45847 ASIG5V.n7823 ASIG5V.n7717 1.11687
R45848 ASIG5V.n7979 ASIG5V.n7973 1.11687
R45849 ASIG5V.n7823 ASIG5V.n7710 1.11687
R45850 ASIG5V.n7823 ASIG5V.n7703 1.11687
R45851 ASIG5V.n7823 ASIG5V.n7696 1.11687
R45852 ASIG5V.n7979 ASIG5V.n7974 1.11687
R45853 ASIG5V.n7823 ASIG5V.n7689 1.11687
R45854 ASIG5V.n7979 ASIG5V.n7975 1.11687
R45855 ASIG5V.n7823 ASIG5V.n7682 1.11687
R45856 ASIG5V.n7823 ASIG5V.n7675 1.11687
R45857 ASIG5V.n7979 ASIG5V.n7976 1.11687
R45858 ASIG5V.n7823 ASIG5V.n7668 1.11687
R45859 ASIG5V.n7979 ASIG5V.n7977 1.11687
R45860 ASIG5V.n7823 ASIG5V.n7661 1.11687
R45861 ASIG5V.n7823 ASIG5V.n7655 1.11687
R45862 ASIG5V.n7823 ASIG5V.n7650 1.11687
R45863 ASIG5V.n7979 ASIG5V.n7978 1.11687
R45864 ASIG5V.n7823 ASIG5V.n7645 1.11687
R45865 ASIG5V.n8120 ASIG5V.n8116 1.11687
R45866 ASIG5V.n12752 ASIG5V.n12704 1.11687
R45867 ASIG5V.n8120 ASIG5V.n8113 1.11687
R45868 ASIG5V.n12752 ASIG5V.n12705 1.11687
R45869 ASIG5V.n8120 ASIG5V.n8110 1.11687
R45870 ASIG5V.n8120 ASIG5V.n8108 1.11687
R45871 ASIG5V.n12752 ASIG5V.n12707 1.11687
R45872 ASIG5V.n8120 ASIG5V.n8106 1.11687
R45873 ASIG5V.n12752 ASIG5V.n12709 1.11687
R45874 ASIG5V.n8120 ASIG5V.n8104 1.11687
R45875 ASIG5V.n8120 ASIG5V.n8102 1.11687
R45876 ASIG5V.n8120 ASIG5V.n8100 1.11687
R45877 ASIG5V.n12752 ASIG5V.n12711 1.11687
R45878 ASIG5V.n8120 ASIG5V.n8098 1.11687
R45879 ASIG5V.n8120 ASIG5V.n8095 1.11687
R45880 ASIG5V.n8120 ASIG5V.n8092 1.11687
R45881 ASIG5V.n12752 ASIG5V.n12714 1.11687
R45882 ASIG5V.n8120 ASIG5V.n8091 1.11687
R45883 ASIG5V.n12752 ASIG5V.n12717 1.11687
R45884 ASIG5V.n8120 ASIG5V.n8088 1.11687
R45885 ASIG5V.n8120 ASIG5V.n8085 1.11687
R45886 ASIG5V.n12752 ASIG5V.n12720 1.11687
R45887 ASIG5V.n8120 ASIG5V.n8082 1.11687
R45888 ASIG5V.n12752 ASIG5V.n12723 1.11687
R45889 ASIG5V.n8120 ASIG5V.n8079 1.11687
R45890 ASIG5V.n8120 ASIG5V.n8076 1.11687
R45891 ASIG5V.n8120 ASIG5V.n8072 1.11687
R45892 ASIG5V.n12752 ASIG5V.n12724 1.11687
R45893 ASIG5V.n8120 ASIG5V.n8065 1.11687
R45894 ASIG5V.n12752 ASIG5V.n12725 1.11687
R45895 ASIG5V.n8120 ASIG5V.n8058 1.11687
R45896 ASIG5V.n8120 ASIG5V.n8054 1.11687
R45897 ASIG5V.n12752 ASIG5V.n12729 1.11687
R45898 ASIG5V.n8120 ASIG5V.n8050 1.11687
R45899 ASIG5V.n12752 ASIG5V.n12733 1.11687
R45900 ASIG5V.n8120 ASIG5V.n8046 1.11687
R45901 ASIG5V.n8120 ASIG5V.n8039 1.11687
R45902 ASIG5V.n8120 ASIG5V.n8032 1.11687
R45903 ASIG5V.n12752 ASIG5V.n12737 1.11687
R45904 ASIG5V.n8120 ASIG5V.n8028 1.11687
R45905 ASIG5V.n12752 ASIG5V.n12741 1.11687
R45906 ASIG5V.n8120 ASIG5V.n8024 1.11687
R45907 ASIG5V.n8120 ASIG5V.n8017 1.11687
R45908 ASIG5V.n12752 ASIG5V.n12745 1.11687
R45909 ASIG5V.n8120 ASIG5V.n8013 1.11687
R45910 ASIG5V.n12752 ASIG5V.n12748 1.11687
R45911 ASIG5V.n8120 ASIG5V.n8009 1.11687
R45912 ASIG5V.n8120 ASIG5V.n8004 1.11687
R45913 ASIG5V.n8120 ASIG5V.n7999 1.11687
R45914 ASIG5V.n12752 ASIG5V.n12751 1.11687
R45915 ASIG5V.n8120 ASIG5V.n7996 1.11687
R45916 ASIG5V.n12653 ASIG5V.n8185 1.11687
R45917 ASIG5V.n12581 ASIG5V.n12490 1.11687
R45918 ASIG5V.n12653 ASIG5V.n8183 1.11687
R45919 ASIG5V.n12581 ASIG5V.n12493 1.11687
R45920 ASIG5V.n12653 ASIG5V.n8182 1.11687
R45921 ASIG5V.n12653 ASIG5V.n8181 1.11687
R45922 ASIG5V.n12581 ASIG5V.n12496 1.11687
R45923 ASIG5V.n12653 ASIG5V.n8179 1.11687
R45924 ASIG5V.n12581 ASIG5V.n12499 1.11687
R45925 ASIG5V.n12653 ASIG5V.n8178 1.11687
R45926 ASIG5V.n12653 ASIG5V.n8177 1.11687
R45927 ASIG5V.n12653 ASIG5V.n8175 1.11687
R45928 ASIG5V.n12581 ASIG5V.n12503 1.11687
R45929 ASIG5V.n12653 ASIG5V.n8174 1.11687
R45930 ASIG5V.n12653 ASIG5V.n8173 1.11687
R45931 ASIG5V.n12653 ASIG5V.n8170 1.11687
R45932 ASIG5V.n12581 ASIG5V.n12508 1.11687
R45933 ASIG5V.n12653 ASIG5V.n8167 1.11687
R45934 ASIG5V.n12581 ASIG5V.n12513 1.11687
R45935 ASIG5V.n12653 ASIG5V.n8166 1.11687
R45936 ASIG5V.n12653 ASIG5V.n8165 1.11687
R45937 ASIG5V.n12581 ASIG5V.n12518 1.11687
R45938 ASIG5V.n12653 ASIG5V.n8162 1.11687
R45939 ASIG5V.n12581 ASIG5V.n12523 1.11687
R45940 ASIG5V.n12653 ASIG5V.n8161 1.11687
R45941 ASIG5V.n12653 ASIG5V.n8160 1.11687
R45942 ASIG5V.n12653 ASIG5V.n8159 1.11687
R45943 ASIG5V.n12581 ASIG5V.n12530 1.11687
R45944 ASIG5V.n12653 ASIG5V.n8155 1.11687
R45945 ASIG5V.n12581 ASIG5V.n12537 1.11687
R45946 ASIG5V.n12653 ASIG5V.n8154 1.11687
R45947 ASIG5V.n12653 ASIG5V.n8153 1.11687
R45948 ASIG5V.n12581 ASIG5V.n12544 1.11687
R45949 ASIG5V.n12653 ASIG5V.n8149 1.11687
R45950 ASIG5V.n12581 ASIG5V.n12551 1.11687
R45951 ASIG5V.n12653 ASIG5V.n8148 1.11687
R45952 ASIG5V.n12653 ASIG5V.n8144 1.11687
R45953 ASIG5V.n12653 ASIG5V.n8140 1.11687
R45954 ASIG5V.n12581 ASIG5V.n12558 1.11687
R45955 ASIG5V.n12653 ASIG5V.n8136 1.11687
R45956 ASIG5V.n12581 ASIG5V.n12565 1.11687
R45957 ASIG5V.n12653 ASIG5V.n8135 1.11687
R45958 ASIG5V.n12653 ASIG5V.n8134 1.11687
R45959 ASIG5V.n12581 ASIG5V.n12570 1.11687
R45960 ASIG5V.n12653 ASIG5V.n8133 1.11687
R45961 ASIG5V.n12581 ASIG5V.n12575 1.11687
R45962 ASIG5V.n12653 ASIG5V.n8132 1.11687
R45963 ASIG5V.n12653 ASIG5V.n8131 1.11687
R45964 ASIG5V.n12653 ASIG5V.n8130 1.11687
R45965 ASIG5V.n12581 ASIG5V.n12580 1.11687
R45966 ASIG5V.n12653 ASIG5V.n8129 1.11687
R45967 ASIG5V.n12425 ASIG5V.n8363 1.11687
R45968 ASIG5V.n12352 ASIG5V.n12334 1.11687
R45969 ASIG5V.n12425 ASIG5V.n8360 1.11687
R45970 ASIG5V.n12352 ASIG5V.n12335 1.11687
R45971 ASIG5V.n12425 ASIG5V.n8357 1.11687
R45972 ASIG5V.n12425 ASIG5V.n8354 1.11687
R45973 ASIG5V.n12352 ASIG5V.n12336 1.11687
R45974 ASIG5V.n12425 ASIG5V.n8351 1.11687
R45975 ASIG5V.n12352 ASIG5V.n12337 1.11687
R45976 ASIG5V.n12425 ASIG5V.n8348 1.11687
R45977 ASIG5V.n12425 ASIG5V.n8345 1.11687
R45978 ASIG5V.n12425 ASIG5V.n8342 1.11687
R45979 ASIG5V.n12352 ASIG5V.n12338 1.11687
R45980 ASIG5V.n12425 ASIG5V.n8339 1.11687
R45981 ASIG5V.n12425 ASIG5V.n8334 1.11687
R45982 ASIG5V.n12425 ASIG5V.n8329 1.11687
R45983 ASIG5V.n12352 ASIG5V.n12339 1.11687
R45984 ASIG5V.n12425 ASIG5V.n8324 1.11687
R45985 ASIG5V.n12352 ASIG5V.n12340 1.11687
R45986 ASIG5V.n12425 ASIG5V.n8319 1.11687
R45987 ASIG5V.n12425 ASIG5V.n8314 1.11687
R45988 ASIG5V.n12352 ASIG5V.n12341 1.11687
R45989 ASIG5V.n12425 ASIG5V.n8309 1.11687
R45990 ASIG5V.n12352 ASIG5V.n12342 1.11687
R45991 ASIG5V.n12425 ASIG5V.n8304 1.11687
R45992 ASIG5V.n12425 ASIG5V.n8299 1.11687
R45993 ASIG5V.n12425 ASIG5V.n8293 1.11687
R45994 ASIG5V.n12352 ASIG5V.n12343 1.11687
R45995 ASIG5V.n12425 ASIG5V.n8286 1.11687
R45996 ASIG5V.n12352 ASIG5V.n12344 1.11687
R45997 ASIG5V.n12425 ASIG5V.n8279 1.11687
R45998 ASIG5V.n12425 ASIG5V.n8272 1.11687
R45999 ASIG5V.n12352 ASIG5V.n12345 1.11687
R46000 ASIG5V.n12425 ASIG5V.n8265 1.11687
R46001 ASIG5V.n12352 ASIG5V.n12346 1.11687
R46002 ASIG5V.n12425 ASIG5V.n8258 1.11687
R46003 ASIG5V.n12425 ASIG5V.n8251 1.11687
R46004 ASIG5V.n12425 ASIG5V.n8244 1.11687
R46005 ASIG5V.n12352 ASIG5V.n12347 1.11687
R46006 ASIG5V.n12425 ASIG5V.n8237 1.11687
R46007 ASIG5V.n12352 ASIG5V.n12348 1.11687
R46008 ASIG5V.n12425 ASIG5V.n8230 1.11687
R46009 ASIG5V.n12425 ASIG5V.n8225 1.11687
R46010 ASIG5V.n12352 ASIG5V.n12349 1.11687
R46011 ASIG5V.n12425 ASIG5V.n8220 1.11687
R46012 ASIG5V.n12352 ASIG5V.n12350 1.11687
R46013 ASIG5V.n12425 ASIG5V.n8215 1.11687
R46014 ASIG5V.n12425 ASIG5V.n8210 1.11687
R46015 ASIG5V.n12425 ASIG5V.n8205 1.11687
R46016 ASIG5V.n12352 ASIG5V.n12351 1.11687
R46017 ASIG5V.n12425 ASIG5V.n8200 1.11687
R46018 ASIG5V.n12310 ASIG5V.n8489 1.11687
R46019 ASIG5V.n12238 ASIG5V.n12195 1.11687
R46020 ASIG5V.n12310 ASIG5V.n8487 1.11687
R46021 ASIG5V.n12238 ASIG5V.n12197 1.11687
R46022 ASIG5V.n12310 ASIG5V.n8485 1.11687
R46023 ASIG5V.n12310 ASIG5V.n8482 1.11687
R46024 ASIG5V.n12238 ASIG5V.n12199 1.11687
R46025 ASIG5V.n12310 ASIG5V.n8480 1.11687
R46026 ASIG5V.n12238 ASIG5V.n12200 1.11687
R46027 ASIG5V.n12310 ASIG5V.n8477 1.11687
R46028 ASIG5V.n12310 ASIG5V.n8474 1.11687
R46029 ASIG5V.n12310 ASIG5V.n8472 1.11687
R46030 ASIG5V.n12238 ASIG5V.n12202 1.11687
R46031 ASIG5V.n12310 ASIG5V.n8470 1.11687
R46032 ASIG5V.n12310 ASIG5V.n8465 1.11687
R46033 ASIG5V.n12310 ASIG5V.n8462 1.11687
R46034 ASIG5V.n12238 ASIG5V.n12205 1.11687
R46035 ASIG5V.n12310 ASIG5V.n8459 1.11687
R46036 ASIG5V.n12238 ASIG5V.n12206 1.11687
R46037 ASIG5V.n12310 ASIG5V.n8454 1.11687
R46038 ASIG5V.n12310 ASIG5V.n8451 1.11687
R46039 ASIG5V.n12238 ASIG5V.n12207 1.11687
R46040 ASIG5V.n12310 ASIG5V.n8446 1.11687
R46041 ASIG5V.n12238 ASIG5V.n12210 1.11687
R46042 ASIG5V.n12310 ASIG5V.n8443 1.11687
R46043 ASIG5V.n12310 ASIG5V.n8440 1.11687
R46044 ASIG5V.n12310 ASIG5V.n8437 1.11687
R46045 ASIG5V.n12238 ASIG5V.n12214 1.11687
R46046 ASIG5V.n12310 ASIG5V.n8434 1.11687
R46047 ASIG5V.n12238 ASIG5V.n12215 1.11687
R46048 ASIG5V.n12310 ASIG5V.n8427 1.11687
R46049 ASIG5V.n12310 ASIG5V.n8420 1.11687
R46050 ASIG5V.n12238 ASIG5V.n12219 1.11687
R46051 ASIG5V.n12310 ASIG5V.n8416 1.11687
R46052 ASIG5V.n12238 ASIG5V.n12223 1.11687
R46053 ASIG5V.n12310 ASIG5V.n8412 1.11687
R46054 ASIG5V.n12310 ASIG5V.n8408 1.11687
R46055 ASIG5V.n12310 ASIG5V.n8401 1.11687
R46056 ASIG5V.n12238 ASIG5V.n12227 1.11687
R46057 ASIG5V.n12310 ASIG5V.n8397 1.11687
R46058 ASIG5V.n12238 ASIG5V.n12230 1.11687
R46059 ASIG5V.n12310 ASIG5V.n8394 1.11687
R46060 ASIG5V.n12310 ASIG5V.n8391 1.11687
R46061 ASIG5V.n12238 ASIG5V.n12231 1.11687
R46062 ASIG5V.n12310 ASIG5V.n8386 1.11687
R46063 ASIG5V.n12238 ASIG5V.n12234 1.11687
R46064 ASIG5V.n12310 ASIG5V.n8383 1.11687
R46065 ASIG5V.n12310 ASIG5V.n8378 1.11687
R46066 ASIG5V.n12310 ASIG5V.n8373 1.11687
R46067 ASIG5V.n12238 ASIG5V.n12237 1.11687
R46068 ASIG5V.n12310 ASIG5V.n8370 1.11687
R46069 ASIG5V.n12154 ASIG5V.n8609 1.11687
R46070 ASIG5V.n12082 ASIG5V.n12041 1.11687
R46071 ASIG5V.n12154 ASIG5V.n8606 1.11687
R46072 ASIG5V.n12082 ASIG5V.n12043 1.11687
R46073 ASIG5V.n12154 ASIG5V.n8604 1.11687
R46074 ASIG5V.n12154 ASIG5V.n8602 1.11687
R46075 ASIG5V.n12082 ASIG5V.n12045 1.11687
R46076 ASIG5V.n12154 ASIG5V.n8600 1.11687
R46077 ASIG5V.n12082 ASIG5V.n12047 1.11687
R46078 ASIG5V.n12154 ASIG5V.n8598 1.11687
R46079 ASIG5V.n12154 ASIG5V.n8595 1.11687
R46080 ASIG5V.n12154 ASIG5V.n8593 1.11687
R46081 ASIG5V.n12082 ASIG5V.n12049 1.11687
R46082 ASIG5V.n12154 ASIG5V.n8591 1.11687
R46083 ASIG5V.n12154 ASIG5V.n8588 1.11687
R46084 ASIG5V.n12154 ASIG5V.n8585 1.11687
R46085 ASIG5V.n12082 ASIG5V.n12052 1.11687
R46086 ASIG5V.n12154 ASIG5V.n8582 1.11687
R46087 ASIG5V.n12082 ASIG5V.n12053 1.11687
R46088 ASIG5V.n12154 ASIG5V.n8577 1.11687
R46089 ASIG5V.n12154 ASIG5V.n8572 1.11687
R46090 ASIG5V.n12082 ASIG5V.n12056 1.11687
R46091 ASIG5V.n12154 ASIG5V.n8569 1.11687
R46092 ASIG5V.n12082 ASIG5V.n12057 1.11687
R46093 ASIG5V.n12154 ASIG5V.n8564 1.11687
R46094 ASIG5V.n12154 ASIG5V.n8561 1.11687
R46095 ASIG5V.n12154 ASIG5V.n8558 1.11687
R46096 ASIG5V.n12082 ASIG5V.n12060 1.11687
R46097 ASIG5V.n12154 ASIG5V.n8555 1.11687
R46098 ASIG5V.n12082 ASIG5V.n12064 1.11687
R46099 ASIG5V.n12154 ASIG5V.n8551 1.11687
R46100 ASIG5V.n12154 ASIG5V.n8544 1.11687
R46101 ASIG5V.n12082 ASIG5V.n12068 1.11687
R46102 ASIG5V.n12154 ASIG5V.n8540 1.11687
R46103 ASIG5V.n12082 ASIG5V.n12072 1.11687
R46104 ASIG5V.n12154 ASIG5V.n8536 1.11687
R46105 ASIG5V.n12154 ASIG5V.n8529 1.11687
R46106 ASIG5V.n12154 ASIG5V.n8525 1.11687
R46107 ASIG5V.n12082 ASIG5V.n12075 1.11687
R46108 ASIG5V.n12154 ASIG5V.n8522 1.11687
R46109 ASIG5V.n12082 ASIG5V.n12076 1.11687
R46110 ASIG5V.n12154 ASIG5V.n8517 1.11687
R46111 ASIG5V.n12154 ASIG5V.n8514 1.11687
R46112 ASIG5V.n12082 ASIG5V.n12079 1.11687
R46113 ASIG5V.n12154 ASIG5V.n8511 1.11687
R46114 ASIG5V.n12082 ASIG5V.n12080 1.11687
R46115 ASIG5V.n12154 ASIG5V.n8506 1.11687
R46116 ASIG5V.n12154 ASIG5V.n8503 1.11687
R46117 ASIG5V.n12154 ASIG5V.n8498 1.11687
R46118 ASIG5V.n12082 ASIG5V.n12081 1.11687
R46119 ASIG5V.n12154 ASIG5V.n8494 1.11687
R46120 ASIG5V.n11999 ASIG5V.n8712 1.11687
R46121 ASIG5V.n11926 ASIG5V.n11879 1.11687
R46122 ASIG5V.n11999 ASIG5V.n8709 1.11687
R46123 ASIG5V.n11926 ASIG5V.n11880 1.11687
R46124 ASIG5V.n11999 ASIG5V.n8706 1.11687
R46125 ASIG5V.n11999 ASIG5V.n8704 1.11687
R46126 ASIG5V.n11926 ASIG5V.n11882 1.11687
R46127 ASIG5V.n11999 ASIG5V.n8702 1.11687
R46128 ASIG5V.n11926 ASIG5V.n11884 1.11687
R46129 ASIG5V.n11999 ASIG5V.n8700 1.11687
R46130 ASIG5V.n11999 ASIG5V.n8698 1.11687
R46131 ASIG5V.n11999 ASIG5V.n8696 1.11687
R46132 ASIG5V.n11926 ASIG5V.n11885 1.11687
R46133 ASIG5V.n11999 ASIG5V.n8693 1.11687
R46134 ASIG5V.n11999 ASIG5V.n8690 1.11687
R46135 ASIG5V.n11999 ASIG5V.n8687 1.11687
R46136 ASIG5V.n11926 ASIG5V.n11888 1.11687
R46137 ASIG5V.n11999 ASIG5V.n8684 1.11687
R46138 ASIG5V.n11926 ASIG5V.n11891 1.11687
R46139 ASIG5V.n11999 ASIG5V.n8681 1.11687
R46140 ASIG5V.n11999 ASIG5V.n8678 1.11687
R46141 ASIG5V.n11926 ASIG5V.n11894 1.11687
R46142 ASIG5V.n11999 ASIG5V.n8675 1.11687
R46143 ASIG5V.n11926 ASIG5V.n11897 1.11687
R46144 ASIG5V.n11999 ASIG5V.n8672 1.11687
R46145 ASIG5V.n11999 ASIG5V.n8669 1.11687
R46146 ASIG5V.n11999 ASIG5V.n8664 1.11687
R46147 ASIG5V.n11926 ASIG5V.n11898 1.11687
R46148 ASIG5V.n11999 ASIG5V.n8659 1.11687
R46149 ASIG5V.n11926 ASIG5V.n11901 1.11687
R46150 ASIG5V.n11999 ASIG5V.n8656 1.11687
R46151 ASIG5V.n11999 ASIG5V.n8652 1.11687
R46152 ASIG5V.n11926 ASIG5V.n11905 1.11687
R46153 ASIG5V.n11999 ASIG5V.n8648 1.11687
R46154 ASIG5V.n11926 ASIG5V.n11909 1.11687
R46155 ASIG5V.n11999 ASIG5V.n8644 1.11687
R46156 ASIG5V.n11999 ASIG5V.n8640 1.11687
R46157 ASIG5V.n11999 ASIG5V.n8637 1.11687
R46158 ASIG5V.n11926 ASIG5V.n11912 1.11687
R46159 ASIG5V.n11999 ASIG5V.n8634 1.11687
R46160 ASIG5V.n11926 ASIG5V.n11917 1.11687
R46161 ASIG5V.n11999 ASIG5V.n8631 1.11687
R46162 ASIG5V.n11999 ASIG5V.n8630 1.11687
R46163 ASIG5V.n11926 ASIG5V.n11920 1.11687
R46164 ASIG5V.n11999 ASIG5V.n8627 1.11687
R46165 ASIG5V.n11926 ASIG5V.n11923 1.11687
R46166 ASIG5V.n11999 ASIG5V.n8624 1.11687
R46167 ASIG5V.n11999 ASIG5V.n8621 1.11687
R46168 ASIG5V.n11999 ASIG5V.n8617 1.11687
R46169 ASIG5V.n11926 ASIG5V.n11925 1.11687
R46170 ASIG5V.n11999 ASIG5V.n8615 1.11687
R46171 ASIG5V.n11831 ASIG5V.n8813 1.11687
R46172 ASIG5V.n11760 ASIG5V.n11714 1.11687
R46173 ASIG5V.n11831 ASIG5V.n8811 1.11687
R46174 ASIG5V.n11760 ASIG5V.n11716 1.11687
R46175 ASIG5V.n11831 ASIG5V.n8809 1.11687
R46176 ASIG5V.n11831 ASIG5V.n8807 1.11687
R46177 ASIG5V.n11760 ASIG5V.n11718 1.11687
R46178 ASIG5V.n11831 ASIG5V.n8805 1.11687
R46179 ASIG5V.n11760 ASIG5V.n11720 1.11687
R46180 ASIG5V.n11831 ASIG5V.n8803 1.11687
R46181 ASIG5V.n11831 ASIG5V.n8801 1.11687
R46182 ASIG5V.n11831 ASIG5V.n8798 1.11687
R46183 ASIG5V.n11760 ASIG5V.n11722 1.11687
R46184 ASIG5V.n11831 ASIG5V.n8796 1.11687
R46185 ASIG5V.n11831 ASIG5V.n8793 1.11687
R46186 ASIG5V.n11831 ASIG5V.n8788 1.11687
R46187 ASIG5V.n11760 ASIG5V.n11725 1.11687
R46188 ASIG5V.n11831 ASIG5V.n8785 1.11687
R46189 ASIG5V.n11760 ASIG5V.n11728 1.11687
R46190 ASIG5V.n11831 ASIG5V.n8782 1.11687
R46191 ASIG5V.n11831 ASIG5V.n8779 1.11687
R46192 ASIG5V.n11760 ASIG5V.n11731 1.11687
R46193 ASIG5V.n11831 ASIG5V.n8776 1.11687
R46194 ASIG5V.n11760 ASIG5V.n11734 1.11687
R46195 ASIG5V.n11831 ASIG5V.n8773 1.11687
R46196 ASIG5V.n11831 ASIG5V.n8770 1.11687
R46197 ASIG5V.n11831 ASIG5V.n8767 1.11687
R46198 ASIG5V.n11760 ASIG5V.n11737 1.11687
R46199 ASIG5V.n11831 ASIG5V.n8764 1.11687
R46200 ASIG5V.n11760 ASIG5V.n11738 1.11687
R46201 ASIG5V.n11831 ASIG5V.n8759 1.11687
R46202 ASIG5V.n11831 ASIG5V.n8756 1.11687
R46203 ASIG5V.n11760 ASIG5V.n11742 1.11687
R46204 ASIG5V.n11831 ASIG5V.n8752 1.11687
R46205 ASIG5V.n11760 ASIG5V.n11745 1.11687
R46206 ASIG5V.n11831 ASIG5V.n8749 1.11687
R46207 ASIG5V.n11831 ASIG5V.n8746 1.11687
R46208 ASIG5V.n11831 ASIG5V.n8743 1.11687
R46209 ASIG5V.n11760 ASIG5V.n11748 1.11687
R46210 ASIG5V.n11831 ASIG5V.n8740 1.11687
R46211 ASIG5V.n11760 ASIG5V.n11751 1.11687
R46212 ASIG5V.n11831 ASIG5V.n8737 1.11687
R46213 ASIG5V.n11831 ASIG5V.n8734 1.11687
R46214 ASIG5V.n11760 ASIG5V.n11754 1.11687
R46215 ASIG5V.n11831 ASIG5V.n8731 1.11687
R46216 ASIG5V.n11760 ASIG5V.n11757 1.11687
R46217 ASIG5V.n11831 ASIG5V.n8728 1.11687
R46218 ASIG5V.n11831 ASIG5V.n8725 1.11687
R46219 ASIG5V.n11831 ASIG5V.n8723 1.11687
R46220 ASIG5V.n11760 ASIG5V.n11759 1.11687
R46221 ASIG5V.n11831 ASIG5V.n8720 1.11687
R46222 ASIG5V.n11668 ASIG5V.n8850 1.11687
R46223 ASIG5V.n11631 ASIG5V.n11557 1.11687
R46224 ASIG5V.n11668 ASIG5V.n8849 1.11687
R46225 ASIG5V.n11631 ASIG5V.n11560 1.11687
R46226 ASIG5V.n11668 ASIG5V.n8848 1.11687
R46227 ASIG5V.n11668 ASIG5V.n8847 1.11687
R46228 ASIG5V.n11631 ASIG5V.n11563 1.11687
R46229 ASIG5V.n11668 ASIG5V.n8846 1.11687
R46230 ASIG5V.n11631 ASIG5V.n11566 1.11687
R46231 ASIG5V.n11668 ASIG5V.n8845 1.11687
R46232 ASIG5V.n11668 ASIG5V.n8844 1.11687
R46233 ASIG5V.n11668 ASIG5V.n8843 1.11687
R46234 ASIG5V.n11631 ASIG5V.n11569 1.11687
R46235 ASIG5V.n11668 ASIG5V.n8842 1.11687
R46236 ASIG5V.n11668 ASIG5V.n8841 1.11687
R46237 ASIG5V.n11668 ASIG5V.n8840 1.11687
R46238 ASIG5V.n11631 ASIG5V.n11574 1.11687
R46239 ASIG5V.n11668 ASIG5V.n8839 1.11687
R46240 ASIG5V.n11631 ASIG5V.n11579 1.11687
R46241 ASIG5V.n11668 ASIG5V.n8838 1.11687
R46242 ASIG5V.n11668 ASIG5V.n8837 1.11687
R46243 ASIG5V.n11631 ASIG5V.n11584 1.11687
R46244 ASIG5V.n11668 ASIG5V.n8836 1.11687
R46245 ASIG5V.n11631 ASIG5V.n11589 1.11687
R46246 ASIG5V.n11668 ASIG5V.n8835 1.11687
R46247 ASIG5V.n11668 ASIG5V.n8834 1.11687
R46248 ASIG5V.n11668 ASIG5V.n8833 1.11687
R46249 ASIG5V.n11631 ASIG5V.n11594 1.11687
R46250 ASIG5V.n11668 ASIG5V.n8832 1.11687
R46251 ASIG5V.n11631 ASIG5V.n11599 1.11687
R46252 ASIG5V.n11668 ASIG5V.n8831 1.11687
R46253 ASIG5V.n11668 ASIG5V.n8830 1.11687
R46254 ASIG5V.n11631 ASIG5V.n11604 1.11687
R46255 ASIG5V.n11668 ASIG5V.n8829 1.11687
R46256 ASIG5V.n11631 ASIG5V.n11609 1.11687
R46257 ASIG5V.n11668 ASIG5V.n8828 1.11687
R46258 ASIG5V.n11668 ASIG5V.n8827 1.11687
R46259 ASIG5V.n11668 ASIG5V.n8826 1.11687
R46260 ASIG5V.n11631 ASIG5V.n11614 1.11687
R46261 ASIG5V.n11668 ASIG5V.n8825 1.11687
R46262 ASIG5V.n11631 ASIG5V.n11619 1.11687
R46263 ASIG5V.n11668 ASIG5V.n8824 1.11687
R46264 ASIG5V.n11668 ASIG5V.n8823 1.11687
R46265 ASIG5V.n11631 ASIG5V.n11624 1.11687
R46266 ASIG5V.n11668 ASIG5V.n8822 1.11687
R46267 ASIG5V.n11631 ASIG5V.n11627 1.11687
R46268 ASIG5V.n11668 ASIG5V.n8821 1.11687
R46269 ASIG5V.n11668 ASIG5V.n8820 1.11687
R46270 ASIG5V.n11668 ASIG5V.n8819 1.11687
R46271 ASIG5V.n11631 ASIG5V.n11630 1.11687
R46272 ASIG5V.n11668 ASIG5V.n8818 1.11687
R46273 ASIG5V.n11324 ASIG5V.n11323 1.11687
R46274 ASIG5V.n11631 ASIG5V.n8856 1.11687
R46275 ASIG5V.n11631 ASIG5V.n8853 1.11687
R46276 ASIG5V.n11760 ASIG5V.n8817 1.11687
R46277 ASIG5V.n11760 ASIG5V.n8816 1.11687
R46278 ASIG5V.n11926 ASIG5V.n8718 1.11687
R46279 ASIG5V.n11926 ASIG5V.n8715 1.11687
R46280 ASIG5V.n12082 ASIG5V.n8613 1.11687
R46281 ASIG5V.n12082 ASIG5V.n8611 1.11687
R46282 ASIG5V.n12238 ASIG5V.n8492 1.11687
R46283 ASIG5V.n12238 ASIG5V.n8491 1.11687
R46284 ASIG5V.n12352 ASIG5V.n8366 1.11687
R46285 ASIG5V.n12352 ASIG5V.n8365 1.11687
R46286 ASIG5V.n12581 ASIG5V.n8195 1.11687
R46287 ASIG5V.n12581 ASIG5V.n8190 1.11687
R46288 ASIG5V.n12752 ASIG5V.n8128 1.11687
R46289 ASIG5V.n12752 ASIG5V.n8125 1.11687
R46290 ASIG5V.n7979 ASIG5V.n7945 1.11687
R46291 ASIG5V.n7979 ASIG5V.n7944 1.11687
R46292 ASIG5V.n7626 ASIG5V.n7525 1.11687
R46293 ASIG5V.n7626 ASIG5V.n7522 1.11687
R46294 ASIG5V.n331 ASIG5V.n149 1.11687
R46295 ASIG5V.n331 ASIG5V.n144 1.11687
R46296 ASIG5V.n13495 ASIG5V.n106 1.11687
R46297 ASIG5V.n13495 ASIG5V.n103 1.11687
R46298 ASIG5V.n6652 ASIG5V.n6549 1.11687
R46299 ASIG5V.n6652 ASIG5V.n6548 1.11687
R46300 ASIG5V.n6928 ASIG5V.n6422 1.11687
R46301 ASIG5V.n6928 ASIG5V.n6418 1.11687
R46302 ASIG5V.n7123 ASIG5V.n6337 1.11687
R46303 ASIG5V.n7123 ASIG5V.n6334 1.11687
R46304 ASIG5V.n6149 ASIG5V.n5982 1.11687
R46305 ASIG5V.n6149 ASIG5V.n5977 1.11687
R46306 ASIG5V.n5793 ASIG5V.n5686 1.11687
R46307 ASIG5V.n5793 ASIG5V.n5681 1.11687
R46308 ASIG5V.n5442 ASIG5V.n5404 1.11687
R46309 ASIG5V.n5442 ASIG5V.n5401 1.11687
R46310 ASIG5V.n5142 ASIG5V.n4981 1.11687
R46311 ASIG5V.n5142 ASIG5V.n4976 1.11687
R46312 ASIG5V.n4847 ASIG5V.n4706 1.11687
R46313 ASIG5V.n4847 ASIG5V.n4701 1.11687
R46314 ASIG5V.n4561 ASIG5V.n4452 1.11687
R46315 ASIG5V.n4561 ASIG5V.n4449 1.11687
R46316 ASIG5V.n4277 ASIG5V.n4169 1.11687
R46317 ASIG5V.n4277 ASIG5V.n4166 1.11687
R46318 ASIG5V.n4004 ASIG5V.n3903 1.11687
R46319 ASIG5V.n4004 ASIG5V.n3901 1.11687
R46320 ASIG5V.n3737 ASIG5V.n3629 1.11687
R46321 ASIG5V.n3737 ASIG5V.n3628 1.11687
R46322 ASIG5V.n3475 ASIG5V.n3337 1.11687
R46323 ASIG5V.n3475 ASIG5V.n3334 1.11687
R46324 ASIG5V.n3296 ASIG5V.n3294 1.11687
R46325 ASIG5V.n3251 ASIG5V.n3145 1.11687
R46326 ASIG5V.n3251 ASIG5V.n3142 1.11687
R46327 ASIG5V.n11486 ASIG5V.n11485 1.11687
R46328 ASIG5V.n11324 ASIG5V.n8861 1.11687
R46329 ASIG5V.n2880 ASIG5V.n2827 1.11668
R46330 ASIG5V.n11311 ASIG5V.n8867 1.11668
R46331 ASIG5V.n11154 ASIG5V.n11107 1.11668
R46332 ASIG5V.n11311 ASIG5V.n11192 1.11668
R46333 ASIG5V.n3032 ASIG5V.n3031 1.11668
R46334 ASIG5V.n2880 ASIG5V.n2829 1.11668
R46335 ASIG5V.n11154 ASIG5V.n11108 1.11668
R46336 ASIG5V.n11311 ASIG5V.n11195 1.11668
R46337 ASIG5V.n3032 ASIG5V.n3030 1.11668
R46338 ASIG5V.n2880 ASIG5V.n2830 1.11668
R46339 ASIG5V.n2880 ASIG5V.n2831 1.11668
R46340 ASIG5V.n3032 ASIG5V.n3027 1.11668
R46341 ASIG5V.n11311 ASIG5V.n11198 1.11668
R46342 ASIG5V.n11154 ASIG5V.n11109 1.11668
R46343 ASIG5V.n2880 ASIG5V.n2832 1.11668
R46344 ASIG5V.n3032 ASIG5V.n3024 1.11668
R46345 ASIG5V.n11311 ASIG5V.n11201 1.11668
R46346 ASIG5V.n11154 ASIG5V.n11110 1.11668
R46347 ASIG5V.n11154 ASIG5V.n11111 1.11668
R46348 ASIG5V.n11311 ASIG5V.n11204 1.11668
R46349 ASIG5V.n3032 ASIG5V.n3021 1.11668
R46350 ASIG5V.n2880 ASIG5V.n2833 1.11668
R46351 ASIG5V.n2880 ASIG5V.n2834 1.11668
R46352 ASIG5V.n3032 ASIG5V.n3018 1.11668
R46353 ASIG5V.n11311 ASIG5V.n11206 1.11668
R46354 ASIG5V.n11154 ASIG5V.n11112 1.11668
R46355 ASIG5V.n2880 ASIG5V.n2836 1.11668
R46356 ASIG5V.n3032 ASIG5V.n3015 1.11668
R46357 ASIG5V.n11311 ASIG5V.n11208 1.11668
R46358 ASIG5V.n11154 ASIG5V.n11114 1.11668
R46359 ASIG5V.n11154 ASIG5V.n11116 1.11668
R46360 ASIG5V.n11311 ASIG5V.n11210 1.11668
R46361 ASIG5V.n3032 ASIG5V.n3012 1.11668
R46362 ASIG5V.n2880 ASIG5V.n2837 1.11668
R46363 ASIG5V.n11154 ASIG5V.n11119 1.11668
R46364 ASIG5V.n11311 ASIG5V.n11212 1.11668
R46365 ASIG5V.n3032 ASIG5V.n3010 1.11668
R46366 ASIG5V.n2880 ASIG5V.n2838 1.11668
R46367 ASIG5V.n2880 ASIG5V.n2841 1.11668
R46368 ASIG5V.n3032 ASIG5V.n3007 1.11668
R46369 ASIG5V.n11311 ASIG5V.n11216 1.11668
R46370 ASIG5V.n11154 ASIG5V.n11120 1.11668
R46371 ASIG5V.n11154 ASIG5V.n11121 1.11668
R46372 ASIG5V.n11311 ASIG5V.n11221 1.11668
R46373 ASIG5V.n3032 ASIG5V.n3004 1.11668
R46374 ASIG5V.n2880 ASIG5V.n2842 1.11668
R46375 ASIG5V.n11154 ASIG5V.n11122 1.11668
R46376 ASIG5V.n11311 ASIG5V.n11226 1.11668
R46377 ASIG5V.n3032 ASIG5V.n3001 1.11668
R46378 ASIG5V.n2880 ASIG5V.n2843 1.11668
R46379 ASIG5V.n2880 ASIG5V.n2846 1.11668
R46380 ASIG5V.n3032 ASIG5V.n2996 1.11668
R46381 ASIG5V.n11311 ASIG5V.n11231 1.11668
R46382 ASIG5V.n11154 ASIG5V.n11123 1.11668
R46383 ASIG5V.n2880 ASIG5V.n2847 1.11668
R46384 ASIG5V.n3032 ASIG5V.n2991 1.11668
R46385 ASIG5V.n11311 ASIG5V.n11236 1.11668
R46386 ASIG5V.n11154 ASIG5V.n11124 1.11668
R46387 ASIG5V.n11154 ASIG5V.n11125 1.11668
R46388 ASIG5V.n11311 ASIG5V.n11241 1.11668
R46389 ASIG5V.n3032 ASIG5V.n2988 1.11668
R46390 ASIG5V.n2880 ASIG5V.n2848 1.11668
R46391 ASIG5V.n11154 ASIG5V.n11126 1.11668
R46392 ASIG5V.n11311 ASIG5V.n11246 1.11668
R46393 ASIG5V.n3032 ASIG5V.n2983 1.11668
R46394 ASIG5V.n2880 ASIG5V.n2851 1.11668
R46395 ASIG5V.n2880 ASIG5V.n2852 1.11668
R46396 ASIG5V.n3032 ASIG5V.n2978 1.11668
R46397 ASIG5V.n11311 ASIG5V.n11247 1.11668
R46398 ASIG5V.n11154 ASIG5V.n11129 1.11668
R46399 ASIG5V.n11154 ASIG5V.n11132 1.11668
R46400 ASIG5V.n11311 ASIG5V.n11252 1.11668
R46401 ASIG5V.n3032 ASIG5V.n2975 1.11668
R46402 ASIG5V.n2880 ASIG5V.n2855 1.11668
R46403 ASIG5V.n11154 ASIG5V.n11133 1.11668
R46404 ASIG5V.n11311 ASIG5V.n11257 1.11668
R46405 ASIG5V.n3032 ASIG5V.n2972 1.11668
R46406 ASIG5V.n2880 ASIG5V.n2856 1.11668
R46407 ASIG5V.n2880 ASIG5V.n2857 1.11668
R46408 ASIG5V.n3032 ASIG5V.n2967 1.11668
R46409 ASIG5V.n11311 ASIG5V.n11262 1.11668
R46410 ASIG5V.n11154 ASIG5V.n11134 1.11668
R46411 ASIG5V.n2880 ASIG5V.n2858 1.11668
R46412 ASIG5V.n3032 ASIG5V.n2962 1.11668
R46413 ASIG5V.n11311 ASIG5V.n11265 1.11668
R46414 ASIG5V.n11154 ASIG5V.n11137 1.11668
R46415 ASIG5V.n11154 ASIG5V.n11138 1.11668
R46416 ASIG5V.n11311 ASIG5V.n11270 1.11668
R46417 ASIG5V.n3032 ASIG5V.n2957 1.11668
R46418 ASIG5V.n2880 ASIG5V.n2861 1.11668
R46419 ASIG5V.n11154 ASIG5V.n11139 1.11668
R46420 ASIG5V.n11311 ASIG5V.n11275 1.11668
R46421 ASIG5V.n3032 ASIG5V.n2952 1.11668
R46422 ASIG5V.n2880 ASIG5V.n2864 1.11668
R46423 ASIG5V.n2880 ASIG5V.n2865 1.11668
R46424 ASIG5V.n3032 ASIG5V.n2949 1.11668
R46425 ASIG5V.n11311 ASIG5V.n11280 1.11668
R46426 ASIG5V.n11154 ASIG5V.n11140 1.11668
R46427 ASIG5V.n11154 ASIG5V.n11141 1.11668
R46428 ASIG5V.n11311 ASIG5V.n11285 1.11668
R46429 ASIG5V.n3032 ASIG5V.n2946 1.11668
R46430 ASIG5V.n2880 ASIG5V.n2868 1.11668
R46431 ASIG5V.n11154 ASIG5V.n11142 1.11668
R46432 ASIG5V.n11311 ASIG5V.n11290 1.11668
R46433 ASIG5V.n3032 ASIG5V.n2941 1.11668
R46434 ASIG5V.n2880 ASIG5V.n2869 1.11668
R46435 ASIG5V.n2880 ASIG5V.n2871 1.11668
R46436 ASIG5V.n3032 ASIG5V.n2938 1.11668
R46437 ASIG5V.n11311 ASIG5V.n11293 1.11668
R46438 ASIG5V.n11154 ASIG5V.n11143 1.11668
R46439 ASIG5V.n2880 ASIG5V.n2872 1.11668
R46440 ASIG5V.n3032 ASIG5V.n2934 1.11668
R46441 ASIG5V.n11311 ASIG5V.n11296 1.11668
R46442 ASIG5V.n11154 ASIG5V.n11145 1.11668
R46443 ASIG5V.n11154 ASIG5V.n11146 1.11668
R46444 ASIG5V.n11311 ASIG5V.n11299 1.11668
R46445 ASIG5V.n3032 ASIG5V.n2932 1.11668
R46446 ASIG5V.n2880 ASIG5V.n2873 1.11668
R46447 ASIG5V.n11154 ASIG5V.n11147 1.11668
R46448 ASIG5V.n11311 ASIG5V.n11302 1.11668
R46449 ASIG5V.n3032 ASIG5V.n2929 1.11668
R46450 ASIG5V.n2880 ASIG5V.n2874 1.11668
R46451 ASIG5V.n2880 ASIG5V.n2875 1.11668
R46452 ASIG5V.n3032 ASIG5V.n2926 1.11668
R46453 ASIG5V.n11311 ASIG5V.n11305 1.11668
R46454 ASIG5V.n11154 ASIG5V.n11148 1.11668
R46455 ASIG5V.n11154 ASIG5V.n11149 1.11668
R46456 ASIG5V.n11311 ASIG5V.n11307 1.11668
R46457 ASIG5V.n3032 ASIG5V.n2923 1.11668
R46458 ASIG5V.n2880 ASIG5V.n2877 1.11668
R46459 ASIG5V.n11154 ASIG5V.n11151 1.11668
R46460 ASIG5V.n11311 ASIG5V.n11310 1.11668
R46461 ASIG5V.n3032 ASIG5V.n2921 1.11668
R46462 ASIG5V.n2880 ASIG5V.n2879 1.11668
R46463 ASIG5V.n11154 ASIG5V.n11153 1.11668
R46464 ASIG5V.n3032 ASIG5V.n2918 1.11668
R46465 ASIG5V.n2821 ASIG5V.n2820 0.563
R46466 ASIG5V.n2825 ASIG5V.n2824 0.563
R46467 ASIG5V.n2915 ASIG5V.n2914 0.563
R46468 ASIG5V.n3036 ASIG5V.n3035 0.563
R46469 ASIG5V.n3040 ASIG5V.n3039 0.563
R46470 ASIG5V.n3136 ASIG5V.n3135 0.563
R46471 ASIG5V.n3253 ASIG5V.n3252 0.563
R46472 ASIG5V.n3257 ASIG5V.n3256 0.563
R46473 ASIG5V.n3296 ASIG5V.n3295 0.563
R46474 ASIG5V.n3331 ASIG5V.n3330 0.563
R46475 ASIG5V.n3479 ASIG5V.n3478 0.563
R46476 ASIG5V.n3483 ASIG5V.n3482 0.563
R46477 ASIG5V.n3623 ASIG5V.n3622 0.563
R46478 ASIG5V.n3740 ASIG5V.n3739 0.563
R46479 ASIG5V.n3745 ASIG5V.n3744 0.563
R46480 ASIG5V.n3896 ASIG5V.n3895 0.563
R46481 ASIG5V.n4007 ASIG5V.n4006 0.563
R46482 ASIG5V.n4012 ASIG5V.n4011 0.563
R46483 ASIG5V.n4164 ASIG5V.n4163 0.563
R46484 ASIG5V.n4282 ASIG5V.n4281 0.563
R46485 ASIG5V.n4285 ASIG5V.n4284 0.563
R46486 ASIG5V.n4440 ASIG5V.n4439 0.563
R46487 ASIG5V.n4446 ASIG5V.n4445 0.563
R46488 ASIG5V.n4566 ASIG5V.n4565 0.563
R46489 ASIG5V.n4571 ASIG5V.n4570 0.563
R46490 ASIG5V.n4698 ASIG5V.n4697 0.563
R46491 ASIG5V.n4852 ASIG5V.n4851 0.563
R46492 ASIG5V.n4857 ASIG5V.n4856 0.563
R46493 ASIG5V.n4966 ASIG5V.n4965 0.563
R46494 ASIG5V.n5145 ASIG5V.n5144 0.563
R46495 ASIG5V.n5151 ASIG5V.n5150 0.563
R46496 ASIG5V.n5393 ASIG5V.n5392 0.563
R46497 ASIG5V.n5445 ASIG5V.n5444 0.563
R46498 ASIG5V.n5452 ASIG5V.n5451 0.563
R46499 ASIG5V.n5671 ASIG5V.n5670 0.563
R46500 ASIG5V.n5797 ASIG5V.n5796 0.563
R46501 ASIG5V.n5801 ASIG5V.n5800 0.563
R46502 ASIG5V.n5808 ASIG5V.n5807 0.563
R46503 ASIG5V.n5972 ASIG5V.n5971 0.563
R46504 ASIG5V.n6156 ASIG5V.n6155 0.563
R46505 ASIG5V.n6163 ASIG5V.n6162 0.563
R46506 ASIG5V.n7125 ASIG5V.n7124 0.563
R46507 ASIG5V.n7063 ASIG5V.n7062 0.563
R46508 ASIG5V.n7056 ASIG5V.n7055 0.563
R46509 ASIG5V.n7048 ASIG5V.n7047 0.563
R46510 ASIG5V.n6791 ASIG5V.n6790 0.563
R46511 ASIG5V.n6784 ASIG5V.n6783 0.563
R46512 ASIG5V.n6769 ASIG5V.n6768 0.563
R46513 ASIG5V.n6556 ASIG5V.n6555 0.563
R46514 ASIG5V.n3 ASIG5V.n2 0.563
R46515 ASIG5V.n13616 ASIG5V.n13615 0.563
R46516 ASIG5V.n13607 ASIG5V.n13606 0.563
R46517 ASIG5V.n13371 ASIG5V.n13370 0.563
R46518 ASIG5V.n13364 ASIG5V.n13363 0.563
R46519 ASIG5V.n13353 ASIG5V.n13352 0.563
R46520 ASIG5V.n7278 ASIG5V.n7277 0.563
R46521 ASIG5V.n7285 ASIG5V.n7284 0.563
R46522 ASIG5V.n7519 ASIG5V.n7518 0.563
R46523 ASIG5V.n7633 ASIG5V.n7632 0.563
R46524 ASIG5V.n7640 ASIG5V.n7639 0.563
R46525 ASIG5V.n7936 ASIG5V.n7935 0.563
R46526 ASIG5V.n7983 ASIG5V.n7982 0.563
R46527 ASIG5V.n7990 ASIG5V.n7989 0.563
R46528 ASIG5V.n12759 ASIG5V.n12758 0.563
R46529 ASIG5V.n12668 ASIG5V.n12667 0.563
R46530 ASIG5V.n12662 ASIG5V.n12661 0.563
R46531 ASIG5V.n12656 ASIG5V.n12655 0.563
R46532 ASIG5V.n12646 ASIG5V.n12645 0.563
R46533 ASIG5V.n12435 ASIG5V.n12434 0.563
R46534 ASIG5V.n12430 ASIG5V.n12429 0.563
R46535 ASIG5V.n12420 ASIG5V.n12419 0.563
R46536 ASIG5V.n12318 ASIG5V.n12317 0.563
R46537 ASIG5V.n12313 ASIG5V.n12312 0.563
R46538 ASIG5V.n12303 ASIG5V.n12302 0.563
R46539 ASIG5V.n12162 ASIG5V.n12161 0.563
R46540 ASIG5V.n12157 ASIG5V.n12156 0.563
R46541 ASIG5V.n12150 ASIG5V.n12149 0.563
R46542 ASIG5V.n12009 ASIG5V.n12008 0.563
R46543 ASIG5V.n12004 ASIG5V.n12003 0.563
R46544 ASIG5V.n11997 ASIG5V.n11996 0.563
R46545 ASIG5V.n11959 ASIG5V.n11958 0.563
R46546 ASIG5V.n11839 ASIG5V.n11838 0.563
R46547 ASIG5V.n11834 ASIG5V.n11833 0.563
R46548 ASIG5V.n11828 ASIG5V.n11827 0.563
R46549 ASIG5V.n11676 ASIG5V.n11675 0.563
R46550 ASIG5V.n11672 ASIG5V.n11671 0.563
R46551 ASIG5V.n11666 ASIG5V.n11665 0.563
R46552 ASIG5V.n11492 ASIG5V.n11491 0.563
R46553 ASIG5V.n11488 ASIG5V.n11487 0.563
R46554 ASIG5V.n11416 ASIG5V.n11415 0.563
R46555 ASIG5V.n11317 ASIG5V.n11316 0.563
R46556 ASIG5V.n11315 ASIG5V.n11314 0.563
R46557 ASIG5V.n11189 ASIG5V.n11188 0.563
R46558 ASIG5V.n11106 ASIG5V.n11105 0.563
R46559 ASIG5V.n11102 ASIG5V.n11101 0.563
R46560 ASIG5V.n11098 ASIG5V.n11097 0.563
R46561 ASIG5V.n3622 ASIG5V.n3621 0.563
R46562 ASIG5V.n3739 ASIG5V.n3738 0.563
R46563 ASIG5V.n3744 ASIG5V.n3743 0.563
R46564 ASIG5V.n3895 ASIG5V.n3894 0.563
R46565 ASIG5V.n4006 ASIG5V.n4005 0.563
R46566 ASIG5V.n4011 ASIG5V.n4010 0.563
R46567 ASIG5V.n4163 ASIG5V.n4162 0.563
R46568 ASIG5V.n4281 ASIG5V.n4280 0.563
R46569 ASIG5V.n4284 ASIG5V.n4283 0.563
R46570 ASIG5V.n4439 ASIG5V.n4438 0.563
R46571 ASIG5V.n4445 ASIG5V.n4444 0.563
R46572 ASIG5V.n4565 ASIG5V.n4564 0.563
R46573 ASIG5V.n4570 ASIG5V.n4569 0.563
R46574 ASIG5V.n4697 ASIG5V.n4696 0.563
R46575 ASIG5V.n4851 ASIG5V.n4850 0.563
R46576 ASIG5V.n4856 ASIG5V.n4855 0.563
R46577 ASIG5V.n4965 ASIG5V.n4964 0.563
R46578 ASIG5V.n5144 ASIG5V.n5143 0.563
R46579 ASIG5V.n5150 ASIG5V.n5149 0.563
R46580 ASIG5V.n5392 ASIG5V.n5391 0.563
R46581 ASIG5V.n5444 ASIG5V.n5443 0.563
R46582 ASIG5V.n5451 ASIG5V.n5450 0.563
R46583 ASIG5V.n5450 ASIG5V.n5449 0.563
R46584 ASIG5V.n5670 ASIG5V.n5669 0.563
R46585 ASIG5V.n5669 ASIG5V.n5668 0.563
R46586 ASIG5V.n5796 ASIG5V.n5795 0.563
R46587 ASIG5V.n5795 ASIG5V.n5794 0.563
R46588 ASIG5V.n5800 ASIG5V.n5799 0.563
R46589 ASIG5V.n5799 ASIG5V.n5798 0.563
R46590 ASIG5V.n5807 ASIG5V.n5806 0.563
R46591 ASIG5V.n5806 ASIG5V.n5805 0.563
R46592 ASIG5V.n5971 ASIG5V.n5970 0.563
R46593 ASIG5V.n5970 ASIG5V.n5969 0.563
R46594 ASIG5V.n6155 ASIG5V.n6154 0.563
R46595 ASIG5V.n6154 ASIG5V.n6153 0.563
R46596 ASIG5V.n6162 ASIG5V.n6161 0.563
R46597 ASIG5V.n6161 ASIG5V.n6160 0.563
R46598 ASIG5V.n7126 ASIG5V.n7125 0.563
R46599 ASIG5V.n7127 ASIG5V.n7126 0.563
R46600 ASIG5V.n7062 ASIG5V.n7061 0.563
R46601 ASIG5V.n7061 ASIG5V.n7060 0.563
R46602 ASIG5V.n7055 ASIG5V.n7054 0.563
R46603 ASIG5V.n7054 ASIG5V.n7053 0.563
R46604 ASIG5V.n7047 ASIG5V.n7046 0.563
R46605 ASIG5V.n7046 ASIG5V.n7045 0.563
R46606 ASIG5V.n6790 ASIG5V.n6789 0.563
R46607 ASIG5V.n6789 ASIG5V.n6788 0.563
R46608 ASIG5V.n6783 ASIG5V.n6782 0.563
R46609 ASIG5V.n6782 ASIG5V.n6781 0.563
R46610 ASIG5V.n6768 ASIG5V.n6767 0.563
R46611 ASIG5V.n6767 ASIG5V.n6766 0.563
R46612 ASIG5V.n6555 ASIG5V.n6554 0.563
R46613 ASIG5V.n6554 ASIG5V.n6553 0.563
R46614 ASIG5V.n2 ASIG5V.n1 0.563
R46615 ASIG5V.n1 ASIG5V.n0 0.563
R46616 ASIG5V.n13615 ASIG5V.n13614 0.563
R46617 ASIG5V.n13614 ASIG5V.n13613 0.563
R46618 ASIG5V.n13606 ASIG5V.n13605 0.563
R46619 ASIG5V.n13605 ASIG5V.n13604 0.563
R46620 ASIG5V.n13370 ASIG5V.n13369 0.563
R46621 ASIG5V.n13369 ASIG5V.n13368 0.563
R46622 ASIG5V.n13363 ASIG5V.n13362 0.563
R46623 ASIG5V.n13362 ASIG5V.n13361 0.563
R46624 ASIG5V.n13352 ASIG5V.n13351 0.563
R46625 ASIG5V.n13351 ASIG5V.n13350 0.563
R46626 ASIG5V.n7277 ASIG5V.n7276 0.563
R46627 ASIG5V.n7276 ASIG5V.n7275 0.563
R46628 ASIG5V.n7284 ASIG5V.n7283 0.563
R46629 ASIG5V.n7283 ASIG5V.n7282 0.563
R46630 ASIG5V.n7518 ASIG5V.n7517 0.563
R46631 ASIG5V.n7517 ASIG5V.n7516 0.563
R46632 ASIG5V.n7632 ASIG5V.n7631 0.563
R46633 ASIG5V.n7631 ASIG5V.n7630 0.563
R46634 ASIG5V.n7639 ASIG5V.n7638 0.563
R46635 ASIG5V.n7638 ASIG5V.n7637 0.563
R46636 ASIG5V.n7935 ASIG5V.n7934 0.563
R46637 ASIG5V.n7934 ASIG5V.n7933 0.563
R46638 ASIG5V.n7982 ASIG5V.n7981 0.563
R46639 ASIG5V.n7981 ASIG5V.n7980 0.563
R46640 ASIG5V.n7989 ASIG5V.n7988 0.563
R46641 ASIG5V.n7988 ASIG5V.n7987 0.563
R46642 ASIG5V.n12760 ASIG5V.n12759 0.563
R46643 ASIG5V.n12761 ASIG5V.n12760 0.563
R46644 ASIG5V.n12667 ASIG5V.n12666 0.563
R46645 ASIG5V.n12661 ASIG5V.n12660 0.563
R46646 ASIG5V.n12655 ASIG5V.n12654 0.563
R46647 ASIG5V.n12645 ASIG5V.n12644 0.563
R46648 ASIG5V.n12434 ASIG5V.n12433 0.563
R46649 ASIG5V.n12429 ASIG5V.n12428 0.563
R46650 ASIG5V.n12419 ASIG5V.n12418 0.563
R46651 ASIG5V.n12317 ASIG5V.n12316 0.563
R46652 ASIG5V.n12312 ASIG5V.n12311 0.563
R46653 ASIG5V.n12302 ASIG5V.n12301 0.563
R46654 ASIG5V.n12161 ASIG5V.n12160 0.563
R46655 ASIG5V.n12156 ASIG5V.n12155 0.563
R46656 ASIG5V.n12149 ASIG5V.n12148 0.563
R46657 ASIG5V.n12008 ASIG5V.n12007 0.563
R46658 ASIG5V.n12003 ASIG5V.n12002 0.563
R46659 ASIG5V.n11996 ASIG5V.n11995 0.563
R46660 ASIG5V.n11958 ASIG5V.n11957 0.563
R46661 ASIG5V.n11838 ASIG5V.n11837 0.563
R46662 ASIG5V.n11833 ASIG5V.n11832 0.563
R46663 ASIG5V.n11827 ASIG5V.n11826 0.563
R46664 ASIG5V.n12876 ASIG5V.n12875 0.475303
R46665 ASIG5V.n10017 ASIG5V.n10016 0.475303
R46666 ASIG5V.n13173 ASIG5V.n13172 0.475303
R46667 ASIG5V.n2075 ASIG5V.n2074 0.475303
R46668 ASIG5V.n1556 ASIG5V.n1555 0.475303
R46669 ASIG5V.n10440 ASIG5V.n10439 0.475303
R46670 ASIG5V.n9909 ASIG5V.n9908 0.475303
R46671 ASIG5V.n2365 ASIG5V.n2364 0.475303
R46672 ASIG5V.n1064 ASIG5V.n1063 0.452975
R46673 ASIG5V.n9429 ASIG5V.n9428 0.452975
R46674 ASIG5V.n9114 ASIG5V.n9113 0.4505
R46675 ASIG5V.n9113 ASIG5V.n9112 0.4505
R46676 ASIG5V.n8876 ASIG5V.n8875 0.4505
R46677 ASIG5V.n8984 ASIG5V.n8983 0.4505
R46678 ASIG5V.n8978 ASIG5V.n8977 0.4505
R46679 ASIG5V.n8872 ASIG5V.n8871 0.4505
R46680 ASIG5V.n8869 ASIG5V.n8868 0.4505
R46681 ASIG5V.n8972 ASIG5V.n8971 0.4505
R46682 ASIG5V.n8970 ASIG5V.n8969 0.4505
R46683 ASIG5V.n8962 ASIG5V.n8961 0.4505
R46684 ASIG5V.n8960 ASIG5V.n8959 0.4505
R46685 ASIG5V.n8958 ASIG5V.n8957 0.4505
R46686 ASIG5V.n8956 ASIG5V.n8955 0.4505
R46687 ASIG5V.n8952 ASIG5V.n8951 0.4505
R46688 ASIG5V.n8946 ASIG5V.n8945 0.4505
R46689 ASIG5V.n517 ASIG5V.n516 0.4505
R46690 ASIG5V.n516 ASIG5V.n515 0.4505
R46691 ASIG5V.n587 ASIG5V.n586 0.4505
R46692 ASIG5V.n589 ASIG5V.n588 0.4505
R46693 ASIG5V.n593 ASIG5V.n592 0.4505
R46694 ASIG5V.n599 ASIG5V.n598 0.4505
R46695 ASIG5V.n601 ASIG5V.n600 0.4505
R46696 ASIG5V.n611 ASIG5V.n610 0.4505
R46697 ASIG5V.n615 ASIG5V.n614 0.4505
R46698 ASIG5V.n618 ASIG5V.n617 0.4505
R46699 ASIG5V.n624 ASIG5V.n623 0.4505
R46700 ASIG5V.n519 ASIG5V.n518 0.4505
R46701 ASIG5V.n738 ASIG5V.n629 0.4505
R46702 ASIG5V.n1065 ASIG5V.n1064 0.4505
R46703 ASIG5V.n8985 ASIG5V.n8984 0.4505
R46704 ASIG5V.n8870 ASIG5V.n8869 0.4505
R46705 ASIG5V.n8973 ASIG5V.n8972 0.4505
R46706 ASIG5V.n8873 ASIG5V.n8872 0.4505
R46707 ASIG5V.n616 ASIG5V.n615 0.4505
R46708 ASIG5V.n619 ASIG5V.n618 0.4505
R46709 ASIG5V.n8877 ASIG5V.n8876 0.4505
R46710 ASIG5V.n8979 ASIG5V.n8978 0.4505
R46711 ASIG5V.n625 ASIG5V.n624 0.4505
R46712 ASIG5V.n520 ASIG5V.n519 0.4505
R46713 ASIG5V.n739 ASIG5V.n738 0.4505
R46714 ASIG5V.n9430 ASIG5V.n9429 0.4505
R46715 ASIG5V.n2500 ASIG5V.n2499 0.3755
R46716 ASIG5V.n10761 ASIG5V.n10760 0.3755
R46717 ASIG5V.n11095 ASIG5V.n11094 0.3755
R46718 ASIG5V.n2818 ASIG5V.n2817 0.3755
R46719 ASIG5V.n1508 ASIG5V.t0 0.327124
R46720 ASIG5V.n1423 ASIG5V.t1 0.327124
R46721 ASIG5V.n1446 ASIG5V.t4 0.32703
R46722 ASIG5V.n9893 ASIG5V.t6 0.326988
R46723 ASIG5V.t5 ASIG5V 0.3255
R46724 ASIG5V.n1628 ASIG5V.t3 0.301145
R46725 ASIG5V.n1658 ASIG5V.t2 0.301145
R46726 ASIG5V.n9921 ASIG5V.t7 0.30099
R46727 ASIG5V.n10068 ASIG5V.t5 0.30099
R46728 ASIG5V.n12763 ASIG5V.n12762 0.29424
R46729 ASIG5V.n13349 ASIG5V.n13302 0.29424
R46730 ASIG5V.n7129 ASIG5V.n7128 0.29424
R46731 ASIG5V.n2175 ASIG5V.n2174 0.29424
R46732 ASIG5V.n2478 ASIG5V.n1675 0.29424
R46733 ASIG5V.n10726 ASIG5V.n10572 0.29424
R46734 ASIG5V.n10739 ASIG5V.n10138 0.29424
R46735 ASIG5V.n2465 ASIG5V.n2464 0.29424
R46736 ASIG5V.n2498 ASIG5V.n2497 0.195812
R46737 ASIG5V.n10759 ASIG5V.n10758 0.195812
R46738 ASIG5V.n12955 ASIG5V.n12954 0.158
R46739 ASIG5V.n12930 ASIG5V.n12929 0.158
R46740 ASIG5V.n12905 ASIG5V.n12904 0.158
R46741 ASIG5V.n12847 ASIG5V.n12846 0.158
R46742 ASIG5V.n12822 ASIG5V.n12821 0.158
R46743 ASIG5V.n12793 ASIG5V.n12792 0.158
R46744 ASIG5V.n13077 ASIG5V.n13076 0.158
R46745 ASIG5V.n13105 ASIG5V.n13104 0.158
R46746 ASIG5V.n9989 ASIG5V.n9988 0.158
R46747 ASIG5V.n10045 ASIG5V.n10044 0.158
R46748 ASIG5V.n9958 ASIG5V.n9957 0.158
R46749 ASIG5V.n13274 ASIG5V.n13273 0.158
R46750 ASIG5V.n13026 ASIG5V.n13025 0.158
R46751 ASIG5V.n7196 ASIG5V.n7195 0.158
R46752 ASIG5V.n13142 ASIG5V.n13141 0.158
R46753 ASIG5V.n13204 ASIG5V.n13203 0.158
R46754 ASIG5V.n13234 ASIG5V.n13233 0.158
R46755 ASIG5V.n7159 ASIG5V.n7158 0.158
R46756 ASIG5V.n2000 ASIG5V.n1999 0.158
R46757 ASIG5V.n2025 ASIG5V.n2024 0.158
R46758 ASIG5V.n2050 ASIG5V.n2049 0.158
R46759 ASIG5V.n2100 ASIG5V.n2099 0.158
R46760 ASIG5V.n2125 ASIG5V.n2124 0.158
R46761 ASIG5V.n2150 ASIG5V.n2149 0.158
R46762 ASIG5V.n1464 ASIG5V.n1463 0.158
R46763 ASIG5V.n1496 ASIG5V.n1495 0.158
R46764 ASIG5V.n1526 ASIG5V.n1525 0.158
R46765 ASIG5V.n1586 ASIG5V.n1585 0.158
R46766 ASIG5V.n1616 ASIG5V.n1615 0.158
R46767 ASIG5V.n1646 ASIG5V.n1645 0.158
R46768 ASIG5V.n10365 ASIG5V.n10364 0.158
R46769 ASIG5V.n10390 ASIG5V.n10389 0.158
R46770 ASIG5V.n10415 ASIG5V.n10414 0.158
R46771 ASIG5V.n10465 ASIG5V.n10464 0.158
R46772 ASIG5V.n10499 ASIG5V.n10498 0.158
R46773 ASIG5V.n10530 ASIG5V.n10529 0.158
R46774 ASIG5V.n9825 ASIG5V.n9824 0.158
R46775 ASIG5V.n9853 ASIG5V.n9852 0.158
R46776 ASIG5V.n9881 ASIG5V.n9880 0.158
R46777 ASIG5V.n9937 ASIG5V.n9936 0.158
R46778 ASIG5V.n10084 ASIG5V.n10083 0.158
R46779 ASIG5V.n10114 ASIG5V.n10113 0.158
R46780 ASIG5V.n2289 ASIG5V.n2288 0.158
R46781 ASIG5V.n2315 ASIG5V.n2314 0.158
R46782 ASIG5V.n2340 ASIG5V.n2339 0.158
R46783 ASIG5V.n2390 ASIG5V.n2389 0.158
R46784 ASIG5V.n2415 ASIG5V.n2414 0.158
R46785 ASIG5V.n2440 ASIG5V.n2439 0.158
R46786 ASIG5V.n10322 ASIG5V.n10321 0.0910304
R46787 ASIG5V.n1480 ASIG5V.n1479 0.0910304
R46788 ASIG5V.n10335 ASIG5V.n10334 0.0910304
R46789 ASIG5V.n1433 ASIG5V.n1432 0.0910304
R46790 ASIG5V.n2260 ASIG5V.n2259 0.0910304
R46791 ASIG5V.n12986 ASIG5V.n12985 0.0910304
R46792 ASIG5V.n9795 ASIG5V.n9794 0.0910304
R46793 ASIG5V.n9803 ASIG5V.n9802 0.0910304
R46794 ASIG5V.n2195 ASIG5V.n2194 0.0890067
R46795 ASIG5V.n1394 ASIG5V.n1393 0.0883085
R46796 ASIG5V.n2214 ASIG5V.n2213 0.0883085
R46797 ASIG5V.n1385 ASIG5V.n1384 0.0883085
R46798 ASIG5V.n2204 ASIG5V.n2203 0.0883085
R46799 ASIG5V.n10483 ASIG5V.n10482 0.0883085
R46800 ASIG5V.n10514 ASIG5V.n10513 0.0883085
R46801 ASIG5V.n10543 ASIG5V.n10542 0.0883085
R46802 ASIG5V.n10559 ASIG5V.n10558 0.0883085
R46803 ASIG5V ASIG5V.n7173 0.0881
R46804 ASIG5V ASIG5V.n7175 0.0881
R46805 ASIG5V ASIG5V.n7171 0.0881
R46806 ASIG5V ASIG5V.n10066 0.0881
R46807 ASIG5V.n13127 ASIG5V 0.0881
R46808 ASIG5V ASIG5V.n13253 0.0881
R46809 ASIG5V ASIG5V.n13046 0.0881
R46810 ASIG5V.n402 ASIG5V 0.0881
R46811 ASIG5V.n12994 ASIG5V 0.0881
R46812 ASIG5V.n9970 ASIG5V.n9969 0.0659264
R46813 ASIG5V.n13255 ASIG5V.n13254 0.0659264
R46814 ASIG5V.n401 ASIG5V.n396 0.0659264
R46815 ASIG5V.n9975 ASIG5V.n9974 0.0631705
R46816 ASIG5V.n13126 ASIG5V.n13125 0.0631705
R46817 ASIG5V.n13048 ASIG5V.n13047 0.0631705
R46818 ASIG5V.n12993 ASIG5V.n12992 0.0631705
R46819 ASIG5V.n1403 ASIG5V.n1402 0.0578
R46820 ASIG5V.n1402 ASIG5V.n1401 0.0578
R46821 ASIG5V.n9754 ASIG5V.n9753 0.0578
R46822 ASIG5V.n9755 ASIG5V.n9754 0.0578
R46823 ASIG5V.n1412 ASIG5V.n1411 0.0578
R46824 ASIG5V.n1411 ASIG5V.n1410 0.0578
R46825 ASIG5V.n9762 ASIG5V.n9761 0.0578
R46826 ASIG5V.n9763 ASIG5V.n9762 0.0578
R46827 ASIG5V.n2207 ASIG5V.n2206 0.0578
R46828 ASIG5V.n10058 ASIG5V.n10057 0.0578
R46829 ASIG5V.n9746 ASIG5V.n9745 0.0578
R46830 ASIG5V.n9747 ASIG5V.n9746 0.0578
R46831 ASIG5V.n1421 ASIG5V.n1420 0.0578
R46832 ASIG5V.n1420 ASIG5V.n1419 0.0578
R46833 ASIG5V.n2197 ASIG5V.n2196 0.0578
R46834 ASIG5V.n1376 ASIG5V.n1375 0.0578
R46835 ASIG5V.n1375 ASIG5V.n1374 0.0578
R46836 ASIG5V.n2232 ASIG5V.n2231 0.0562034
R46837 ASIG5V.n2241 ASIG5V.n2240 0.0562034
R46838 ASIG5V.n2251 ASIG5V.n2250 0.0562034
R46839 ASIG5V.n10309 ASIG5V.n10308 0.0562034
R46840 ASIG5V.n9770 ASIG5V.n9769 0.0562034
R46841 ASIG5V.n9778 ASIG5V.n9777 0.0562034
R46842 ASIG5V.n2223 ASIG5V.n2222 0.0561949
R46843 ASIG5V.n10300 ASIG5V.n10299 0.0561949
R46844 ASIG5V.n9740 ASIG5V.n9739 0.0561949
R46845 ASIG5V.n10301 ASIG5V.n10300 0.0558048
R46846 ASIG5V.n9742 ASIG5V.n9740 0.0558048
R46847 ASIG5V.n2224 ASIG5V.n2223 0.0558048
R46848 ASIG5V.n2233 ASIG5V.n2232 0.0557963
R46849 ASIG5V.n2242 ASIG5V.n2241 0.0557963
R46850 ASIG5V.n2252 ASIG5V.n2251 0.0557963
R46851 ASIG5V.n10310 ASIG5V.n10309 0.0557963
R46852 ASIG5V.n9771 ASIG5V.n9770 0.0557963
R46853 ASIG5V.n9779 ASIG5V.n9778 0.0557963
R46854 ASIG5V.n9624 ASIG5V.n9623 0.0380882
R46855 ASIG5V.n9623 ASIG5V.n9622 0.0380882
R46856 ASIG5V.n9622 ASIG5V.n9621 0.0380882
R46857 ASIG5V.n9621 ASIG5V.n9620 0.0380882
R46858 ASIG5V.n9620 ASIG5V.n9619 0.0380882
R46859 ASIG5V.n9619 ASIG5V.n9618 0.0380882
R46860 ASIG5V.n9618 ASIG5V.n9617 0.0380882
R46861 ASIG5V.n9617 ASIG5V.n9616 0.0380882
R46862 ASIG5V.n9616 ASIG5V.n9615 0.0380882
R46863 ASIG5V.n9615 ASIG5V.n9614 0.0380882
R46864 ASIG5V.n9614 ASIG5V.n9613 0.0380882
R46865 ASIG5V.n9613 ASIG5V.n9612 0.0380882
R46866 ASIG5V.n9612 ASIG5V.n9611 0.0380882
R46867 ASIG5V.n9611 ASIG5V.n9610 0.0380882
R46868 ASIG5V.n9610 ASIG5V.n9609 0.0380882
R46869 ASIG5V.n9609 ASIG5V.n9608 0.0380882
R46870 ASIG5V.n9608 ASIG5V.n9607 0.0380882
R46871 ASIG5V.n9607 ASIG5V.n9606 0.0380882
R46872 ASIG5V.n9606 ASIG5V.n9605 0.0380882
R46873 ASIG5V.n9605 ASIG5V.n9604 0.0380882
R46874 ASIG5V.n9604 ASIG5V.n9603 0.0380882
R46875 ASIG5V.n9603 ASIG5V.n9602 0.0380882
R46876 ASIG5V.n9602 ASIG5V.n9601 0.0380882
R46877 ASIG5V.n9601 ASIG5V.n9600 0.0380882
R46878 ASIG5V.n9600 ASIG5V.n9599 0.0380882
R46879 ASIG5V.n9599 ASIG5V.n9598 0.0380882
R46880 ASIG5V.n9598 ASIG5V.n9597 0.0380882
R46881 ASIG5V.n9597 ASIG5V.n9596 0.0380882
R46882 ASIG5V.n9596 ASIG5V.n9595 0.0380882
R46883 ASIG5V.n9595 ASIG5V.n9594 0.0380882
R46884 ASIG5V.n9594 ASIG5V.n9593 0.0380882
R46885 ASIG5V.n9593 ASIG5V.n9592 0.0380882
R46886 ASIG5V.n9592 ASIG5V.n9591 0.0380882
R46887 ASIG5V.n9591 ASIG5V.n9590 0.0380882
R46888 ASIG5V.n9590 ASIG5V.n9589 0.0380882
R46889 ASIG5V.n9589 ASIG5V.n9588 0.0380882
R46890 ASIG5V.n9588 ASIG5V.n9587 0.0380882
R46891 ASIG5V.n9587 ASIG5V.n9586 0.0380882
R46892 ASIG5V.n9586 ASIG5V.n9585 0.0380882
R46893 ASIG5V.n9585 ASIG5V.n9584 0.0380882
R46894 ASIG5V.n9584 ASIG5V.n9583 0.0380882
R46895 ASIG5V.n9583 ASIG5V.n9582 0.0380882
R46896 ASIG5V.n9582 ASIG5V.n9581 0.0380882
R46897 ASIG5V.n9581 ASIG5V.n9580 0.0380882
R46898 ASIG5V.n9580 ASIG5V.n9579 0.0380882
R46899 ASIG5V.n9579 ASIG5V.n9578 0.0380882
R46900 ASIG5V.n9578 ASIG5V.n9577 0.0380882
R46901 ASIG5V.n9577 ASIG5V.n9576 0.0380882
R46902 ASIG5V.n9576 ASIG5V.n9575 0.0380882
R46903 ASIG5V.n9575 ASIG5V.n9574 0.0380882
R46904 ASIG5V.n9574 ASIG5V.n9573 0.0380882
R46905 ASIG5V.n9573 ASIG5V.n9572 0.0380882
R46906 ASIG5V.n9572 ASIG5V.n9571 0.0380882
R46907 ASIG5V.n9571 ASIG5V.n9570 0.0380882
R46908 ASIG5V.n9153 ASIG5V.n9152 0.0380882
R46909 ASIG5V.n9154 ASIG5V.n9153 0.0380882
R46910 ASIG5V.n9155 ASIG5V.n9154 0.0380882
R46911 ASIG5V.n9156 ASIG5V.n9155 0.0380882
R46912 ASIG5V.n9157 ASIG5V.n9156 0.0380882
R46913 ASIG5V.n9158 ASIG5V.n9157 0.0380882
R46914 ASIG5V.n9159 ASIG5V.n9158 0.0380882
R46915 ASIG5V.n9160 ASIG5V.n9159 0.0380882
R46916 ASIG5V.n9161 ASIG5V.n9160 0.0380882
R46917 ASIG5V.n9162 ASIG5V.n9161 0.0380882
R46918 ASIG5V.n9163 ASIG5V.n9162 0.0380882
R46919 ASIG5V.n9164 ASIG5V.n9163 0.0380882
R46920 ASIG5V.n9165 ASIG5V.n9164 0.0380882
R46921 ASIG5V.n9166 ASIG5V.n9165 0.0380882
R46922 ASIG5V.n9167 ASIG5V.n9166 0.0380882
R46923 ASIG5V.n9168 ASIG5V.n9167 0.0380882
R46924 ASIG5V.n9169 ASIG5V.n9168 0.0380882
R46925 ASIG5V.n9170 ASIG5V.n9169 0.0380882
R46926 ASIG5V.n9171 ASIG5V.n9170 0.0380882
R46927 ASIG5V.n9172 ASIG5V.n9171 0.0380882
R46928 ASIG5V.n9173 ASIG5V.n9172 0.0380882
R46929 ASIG5V.n9174 ASIG5V.n9173 0.0380882
R46930 ASIG5V.n9175 ASIG5V.n9174 0.0380882
R46931 ASIG5V.n9176 ASIG5V.n9175 0.0380882
R46932 ASIG5V.n9177 ASIG5V.n9176 0.0380882
R46933 ASIG5V.n9178 ASIG5V.n9177 0.0380882
R46934 ASIG5V.n9179 ASIG5V.n9178 0.0380882
R46935 ASIG5V.n9180 ASIG5V.n9179 0.0380882
R46936 ASIG5V.n1259 ASIG5V.n1258 0.0380882
R46937 ASIG5V.n1258 ASIG5V.n1257 0.0380882
R46938 ASIG5V.n1257 ASIG5V.n1256 0.0380882
R46939 ASIG5V.n1256 ASIG5V.n1255 0.0380882
R46940 ASIG5V.n1255 ASIG5V.n1254 0.0380882
R46941 ASIG5V.n1254 ASIG5V.n1253 0.0380882
R46942 ASIG5V.n1253 ASIG5V.n1252 0.0380882
R46943 ASIG5V.n1252 ASIG5V.n1251 0.0380882
R46944 ASIG5V.n1251 ASIG5V.n1250 0.0380882
R46945 ASIG5V.n1250 ASIG5V.n1249 0.0380882
R46946 ASIG5V.n1249 ASIG5V.n1248 0.0380882
R46947 ASIG5V.n1248 ASIG5V.n1247 0.0380882
R46948 ASIG5V.n1247 ASIG5V.n1246 0.0380882
R46949 ASIG5V.n1246 ASIG5V.n1245 0.0380882
R46950 ASIG5V.n1245 ASIG5V.n1244 0.0380882
R46951 ASIG5V.n1244 ASIG5V.n1243 0.0380882
R46952 ASIG5V.n1243 ASIG5V.n1242 0.0380882
R46953 ASIG5V.n1242 ASIG5V.n1241 0.0380882
R46954 ASIG5V.n1241 ASIG5V.n1240 0.0380882
R46955 ASIG5V.n1240 ASIG5V.n1239 0.0380882
R46956 ASIG5V.n1239 ASIG5V.n1238 0.0380882
R46957 ASIG5V.n1238 ASIG5V.n1237 0.0380882
R46958 ASIG5V.n1237 ASIG5V.n1236 0.0380882
R46959 ASIG5V.n1236 ASIG5V.n1235 0.0380882
R46960 ASIG5V.n1235 ASIG5V.n1234 0.0380882
R46961 ASIG5V.n1234 ASIG5V.n1233 0.0380882
R46962 ASIG5V.n1233 ASIG5V.n1232 0.0380882
R46963 ASIG5V.n1232 ASIG5V.n1231 0.0380882
R46964 ASIG5V.n1231 ASIG5V.n1230 0.0380882
R46965 ASIG5V.n1230 ASIG5V.n1229 0.0380882
R46966 ASIG5V.n1229 ASIG5V.n1228 0.0380882
R46967 ASIG5V.n1228 ASIG5V.n1227 0.0380882
R46968 ASIG5V.n1227 ASIG5V.n1226 0.0380882
R46969 ASIG5V.n1226 ASIG5V.n1225 0.0380882
R46970 ASIG5V.n1225 ASIG5V.n1224 0.0380882
R46971 ASIG5V.n1224 ASIG5V.n1223 0.0380882
R46972 ASIG5V.n1223 ASIG5V.n1222 0.0380882
R46973 ASIG5V.n1222 ASIG5V.n1221 0.0380882
R46974 ASIG5V.n1221 ASIG5V.n1220 0.0380882
R46975 ASIG5V.n1220 ASIG5V.n1219 0.0380882
R46976 ASIG5V.n1219 ASIG5V.n1218 0.0380882
R46977 ASIG5V.n1218 ASIG5V.n1217 0.0380882
R46978 ASIG5V.n1217 ASIG5V.n1216 0.0380882
R46979 ASIG5V.n1216 ASIG5V.n1215 0.0380882
R46980 ASIG5V.n1215 ASIG5V.n1214 0.0380882
R46981 ASIG5V.n1214 ASIG5V.n1213 0.0380882
R46982 ASIG5V.n1213 ASIG5V.n1212 0.0380882
R46983 ASIG5V.n1212 ASIG5V.n1211 0.0380882
R46984 ASIG5V.n1211 ASIG5V.n1210 0.0380882
R46985 ASIG5V.n1210 ASIG5V.n1209 0.0380882
R46986 ASIG5V.n1209 ASIG5V.n1208 0.0380882
R46987 ASIG5V.n1208 ASIG5V.n1207 0.0380882
R46988 ASIG5V.n1207 ASIG5V.n1206 0.0380882
R46989 ASIG5V.n1206 ASIG5V.n1205 0.0380882
R46990 ASIG5V.n749 ASIG5V.n748 0.0380882
R46991 ASIG5V.n750 ASIG5V.n749 0.0380882
R46992 ASIG5V.n751 ASIG5V.n750 0.0380882
R46993 ASIG5V.n752 ASIG5V.n751 0.0380882
R46994 ASIG5V.n753 ASIG5V.n752 0.0380882
R46995 ASIG5V.n754 ASIG5V.n753 0.0380882
R46996 ASIG5V.n755 ASIG5V.n754 0.0380882
R46997 ASIG5V.n756 ASIG5V.n755 0.0380882
R46998 ASIG5V.n757 ASIG5V.n756 0.0380882
R46999 ASIG5V.n758 ASIG5V.n757 0.0380882
R47000 ASIG5V.n759 ASIG5V.n758 0.0380882
R47001 ASIG5V.n760 ASIG5V.n759 0.0380882
R47002 ASIG5V.n761 ASIG5V.n760 0.0380882
R47003 ASIG5V.n762 ASIG5V.n761 0.0380882
R47004 ASIG5V.n763 ASIG5V.n762 0.0380882
R47005 ASIG5V.n764 ASIG5V.n763 0.0380882
R47006 ASIG5V.n765 ASIG5V.n764 0.0380882
R47007 ASIG5V.n766 ASIG5V.n765 0.0380882
R47008 ASIG5V.n767 ASIG5V.n766 0.0380882
R47009 ASIG5V.n768 ASIG5V.n767 0.0380882
R47010 ASIG5V.n769 ASIG5V.n768 0.0380882
R47011 ASIG5V.n770 ASIG5V.n769 0.0380882
R47012 ASIG5V.n771 ASIG5V.n770 0.0380882
R47013 ASIG5V.n772 ASIG5V.n771 0.0380882
R47014 ASIG5V.n773 ASIG5V.n772 0.0380882
R47015 ASIG5V.n774 ASIG5V.n773 0.0380882
R47016 ASIG5V.n775 ASIG5V.n774 0.0380882
R47017 ASIG5V.n776 ASIG5V.n775 0.0380882
R47018 ASIG5V.n2698 ASIG5V.n2697 0.0380882
R47019 ASIG5V.n2697 ASIG5V.n2696 0.0380882
R47020 ASIG5V.n2696 ASIG5V.n2695 0.0380882
R47021 ASIG5V.n2695 ASIG5V.n2694 0.0380882
R47022 ASIG5V.n2694 ASIG5V.n2693 0.0380882
R47023 ASIG5V.n2693 ASIG5V.n2692 0.0380882
R47024 ASIG5V.n2692 ASIG5V.n2691 0.0380882
R47025 ASIG5V.n2691 ASIG5V.n2690 0.0380882
R47026 ASIG5V.n2690 ASIG5V.n2689 0.0380882
R47027 ASIG5V.n2689 ASIG5V.n2688 0.0380882
R47028 ASIG5V.n2688 ASIG5V.n2687 0.0380882
R47029 ASIG5V.n2687 ASIG5V.n2686 0.0380882
R47030 ASIG5V.n2686 ASIG5V.n2685 0.0380882
R47031 ASIG5V.n2685 ASIG5V.n2684 0.0380882
R47032 ASIG5V.n2684 ASIG5V.n2683 0.0380882
R47033 ASIG5V.n2683 ASIG5V.n2682 0.0380882
R47034 ASIG5V.n2682 ASIG5V.n2681 0.0380882
R47035 ASIG5V.n2681 ASIG5V.n2680 0.0380882
R47036 ASIG5V.n2680 ASIG5V.n2679 0.0380882
R47037 ASIG5V.n2679 ASIG5V.n2678 0.0380882
R47038 ASIG5V.n2678 ASIG5V.n2677 0.0380882
R47039 ASIG5V.n2677 ASIG5V.n2676 0.0380882
R47040 ASIG5V.n2676 ASIG5V.n2675 0.0380882
R47041 ASIG5V.n2675 ASIG5V.n2674 0.0380882
R47042 ASIG5V.n2674 ASIG5V.n2673 0.0380882
R47043 ASIG5V.n2673 ASIG5V.n2672 0.0380882
R47044 ASIG5V.n2672 ASIG5V.n2671 0.0380882
R47045 ASIG5V.n2671 ASIG5V.n2670 0.0380882
R47046 ASIG5V.n2670 ASIG5V.n2669 0.0380882
R47047 ASIG5V.n2669 ASIG5V.n2668 0.0380882
R47048 ASIG5V.n2668 ASIG5V.n2667 0.0380882
R47049 ASIG5V.n2667 ASIG5V.n2666 0.0380882
R47050 ASIG5V.n648 ASIG5V.n647 0.0380882
R47051 ASIG5V.n649 ASIG5V.n648 0.0380882
R47052 ASIG5V.n650 ASIG5V.n649 0.0380882
R47053 ASIG5V.n651 ASIG5V.n650 0.0380882
R47054 ASIG5V.n652 ASIG5V.n651 0.0380882
R47055 ASIG5V.n653 ASIG5V.n652 0.0380882
R47056 ASIG5V.n654 ASIG5V.n653 0.0380882
R47057 ASIG5V.n655 ASIG5V.n654 0.0380882
R47058 ASIG5V.n656 ASIG5V.n655 0.0380882
R47059 ASIG5V.n657 ASIG5V.n656 0.0380882
R47060 ASIG5V.n658 ASIG5V.n657 0.0380882
R47061 ASIG5V.n659 ASIG5V.n658 0.0380882
R47062 ASIG5V.n660 ASIG5V.n659 0.0380882
R47063 ASIG5V.n661 ASIG5V.n660 0.0380882
R47064 ASIG5V.n1314 ASIG5V.n1313 0.0380882
R47065 ASIG5V.n1313 ASIG5V.n1312 0.0380882
R47066 ASIG5V.n1312 ASIG5V.n1311 0.0380882
R47067 ASIG5V.n1311 ASIG5V.n1310 0.0380882
R47068 ASIG5V.n1310 ASIG5V.n1309 0.0380882
R47069 ASIG5V.n1309 ASIG5V.n1308 0.0380882
R47070 ASIG5V.n1308 ASIG5V.n1307 0.0380882
R47071 ASIG5V.n1307 ASIG5V.n1306 0.0380882
R47072 ASIG5V.n1306 ASIG5V.n1305 0.0380882
R47073 ASIG5V.n1305 ASIG5V.n1304 0.0380882
R47074 ASIG5V.n1304 ASIG5V.n1303 0.0380882
R47075 ASIG5V.n1303 ASIG5V.n1302 0.0380882
R47076 ASIG5V.n1302 ASIG5V.n1301 0.0380882
R47077 ASIG5V.n1301 ASIG5V.n1300 0.0380882
R47078 ASIG5V.n1300 ASIG5V.n1299 0.0380882
R47079 ASIG5V.n1299 ASIG5V.n1298 0.0380882
R47080 ASIG5V.n1298 ASIG5V.n1297 0.0380882
R47081 ASIG5V.n1297 ASIG5V.n1296 0.0380882
R47082 ASIG5V.n1296 ASIG5V.n1295 0.0380882
R47083 ASIG5V.n1295 ASIG5V.n1294 0.0380882
R47084 ASIG5V.n1294 ASIG5V.n1293 0.0380882
R47085 ASIG5V.n1293 ASIG5V.n1292 0.0380882
R47086 ASIG5V.n1292 ASIG5V.n1291 0.0380882
R47087 ASIG5V.n1291 ASIG5V.n1290 0.0380882
R47088 ASIG5V.n1290 ASIG5V.n1289 0.0380882
R47089 ASIG5V.n1289 ASIG5V.n1288 0.0380882
R47090 ASIG5V.n1288 ASIG5V.n1287 0.0380882
R47091 ASIG5V.n1287 ASIG5V.n1286 0.0380882
R47092 ASIG5V.n1286 ASIG5V.n1285 0.0380882
R47093 ASIG5V.n1285 ASIG5V.n1284 0.0380882
R47094 ASIG5V.n1284 ASIG5V.n1283 0.0380882
R47095 ASIG5V.n1283 ASIG5V.n1282 0.0380882
R47096 ASIG5V.n1282 ASIG5V.n1281 0.0380882
R47097 ASIG5V.n1281 ASIG5V.n1280 0.0380882
R47098 ASIG5V.n1280 ASIG5V.n1279 0.0380882
R47099 ASIG5V.n1279 ASIG5V.n1278 0.0380882
R47100 ASIG5V.n1278 ASIG5V.n1277 0.0380882
R47101 ASIG5V.n1277 ASIG5V.n1276 0.0380882
R47102 ASIG5V.n1276 ASIG5V.n1275 0.0380882
R47103 ASIG5V.n1275 ASIG5V.n1274 0.0380882
R47104 ASIG5V.n1274 ASIG5V.n1273 0.0380882
R47105 ASIG5V.n1273 ASIG5V.n1272 0.0380882
R47106 ASIG5V.n1272 ASIG5V.n1271 0.0380882
R47107 ASIG5V.n1271 ASIG5V.n1270 0.0380882
R47108 ASIG5V.n1270 ASIG5V.n1269 0.0380882
R47109 ASIG5V.n1269 ASIG5V.n1268 0.0380882
R47110 ASIG5V.n1268 ASIG5V.n1267 0.0380882
R47111 ASIG5V.n1267 ASIG5V.n1266 0.0380882
R47112 ASIG5V.n1266 ASIG5V.n1265 0.0380882
R47113 ASIG5V.n1265 ASIG5V.n1264 0.0380882
R47114 ASIG5V.n1264 ASIG5V.n1263 0.0380882
R47115 ASIG5V.n1263 ASIG5V.n1262 0.0380882
R47116 ASIG5V.n1262 ASIG5V.n1261 0.0380882
R47117 ASIG5V.n1261 ASIG5V.n1260 0.0380882
R47118 ASIG5V.n778 ASIG5V.n777 0.0380882
R47119 ASIG5V.n779 ASIG5V.n778 0.0380882
R47120 ASIG5V.n780 ASIG5V.n779 0.0380882
R47121 ASIG5V.n781 ASIG5V.n780 0.0380882
R47122 ASIG5V.n782 ASIG5V.n781 0.0380882
R47123 ASIG5V.n783 ASIG5V.n782 0.0380882
R47124 ASIG5V.n784 ASIG5V.n783 0.0380882
R47125 ASIG5V.n785 ASIG5V.n784 0.0380882
R47126 ASIG5V.n786 ASIG5V.n785 0.0380882
R47127 ASIG5V.n787 ASIG5V.n786 0.0380882
R47128 ASIG5V.n788 ASIG5V.n787 0.0380882
R47129 ASIG5V.n789 ASIG5V.n788 0.0380882
R47130 ASIG5V.n790 ASIG5V.n789 0.0380882
R47131 ASIG5V.n791 ASIG5V.n790 0.0380882
R47132 ASIG5V.n792 ASIG5V.n791 0.0380882
R47133 ASIG5V.n793 ASIG5V.n792 0.0380882
R47134 ASIG5V.n794 ASIG5V.n793 0.0380882
R47135 ASIG5V.n795 ASIG5V.n794 0.0380882
R47136 ASIG5V.n796 ASIG5V.n795 0.0380882
R47137 ASIG5V.n797 ASIG5V.n796 0.0380882
R47138 ASIG5V.n798 ASIG5V.n797 0.0380882
R47139 ASIG5V.n799 ASIG5V.n798 0.0380882
R47140 ASIG5V.n800 ASIG5V.n799 0.0380882
R47141 ASIG5V.n801 ASIG5V.n800 0.0380882
R47142 ASIG5V.n802 ASIG5V.n801 0.0380882
R47143 ASIG5V.n803 ASIG5V.n802 0.0380882
R47144 ASIG5V.n804 ASIG5V.n803 0.0380882
R47145 ASIG5V.n805 ASIG5V.n804 0.0380882
R47146 ASIG5V.n2730 ASIG5V.n2729 0.0380882
R47147 ASIG5V.n2729 ASIG5V.n2728 0.0380882
R47148 ASIG5V.n2728 ASIG5V.n2727 0.0380882
R47149 ASIG5V.n2727 ASIG5V.n2726 0.0380882
R47150 ASIG5V.n2726 ASIG5V.n2725 0.0380882
R47151 ASIG5V.n2725 ASIG5V.n2724 0.0380882
R47152 ASIG5V.n2724 ASIG5V.n2723 0.0380882
R47153 ASIG5V.n2723 ASIG5V.n2722 0.0380882
R47154 ASIG5V.n2722 ASIG5V.n2721 0.0380882
R47155 ASIG5V.n2721 ASIG5V.n2720 0.0380882
R47156 ASIG5V.n2720 ASIG5V.n2719 0.0380882
R47157 ASIG5V.n2719 ASIG5V.n2718 0.0380882
R47158 ASIG5V.n2718 ASIG5V.n2717 0.0380882
R47159 ASIG5V.n2717 ASIG5V.n2716 0.0380882
R47160 ASIG5V.n2716 ASIG5V.n2715 0.0380882
R47161 ASIG5V.n2715 ASIG5V.n2714 0.0380882
R47162 ASIG5V.n2714 ASIG5V.n2713 0.0380882
R47163 ASIG5V.n2713 ASIG5V.n2712 0.0380882
R47164 ASIG5V.n2712 ASIG5V.n2711 0.0380882
R47165 ASIG5V.n2711 ASIG5V.n2710 0.0380882
R47166 ASIG5V.n2710 ASIG5V.n2709 0.0380882
R47167 ASIG5V.n2709 ASIG5V.n2708 0.0380882
R47168 ASIG5V.n2708 ASIG5V.n2707 0.0380882
R47169 ASIG5V.n2707 ASIG5V.n2706 0.0380882
R47170 ASIG5V.n2706 ASIG5V.n2705 0.0380882
R47171 ASIG5V.n2705 ASIG5V.n2704 0.0380882
R47172 ASIG5V.n2704 ASIG5V.n2703 0.0380882
R47173 ASIG5V.n2703 ASIG5V.n2702 0.0380882
R47174 ASIG5V.n2702 ASIG5V.n2701 0.0380882
R47175 ASIG5V.n2701 ASIG5V.n2700 0.0380882
R47176 ASIG5V.n2700 ASIG5V.n2699 0.0380882
R47177 ASIG5V.n663 ASIG5V.n662 0.0380882
R47178 ASIG5V.n664 ASIG5V.n663 0.0380882
R47179 ASIG5V.n665 ASIG5V.n664 0.0380882
R47180 ASIG5V.n666 ASIG5V.n665 0.0380882
R47181 ASIG5V.n667 ASIG5V.n666 0.0380882
R47182 ASIG5V.n668 ASIG5V.n667 0.0380882
R47183 ASIG5V.n669 ASIG5V.n668 0.0380882
R47184 ASIG5V.n670 ASIG5V.n669 0.0380882
R47185 ASIG5V.n671 ASIG5V.n670 0.0380882
R47186 ASIG5V.n672 ASIG5V.n671 0.0380882
R47187 ASIG5V.n673 ASIG5V.n672 0.0380882
R47188 ASIG5V.n1368 ASIG5V.n1367 0.0380882
R47189 ASIG5V.n1367 ASIG5V.n1366 0.0380882
R47190 ASIG5V.n1366 ASIG5V.n1365 0.0380882
R47191 ASIG5V.n1365 ASIG5V.n1364 0.0380882
R47192 ASIG5V.n1364 ASIG5V.n1363 0.0380882
R47193 ASIG5V.n1363 ASIG5V.n1362 0.0380882
R47194 ASIG5V.n1362 ASIG5V.n1361 0.0380882
R47195 ASIG5V.n1361 ASIG5V.n1360 0.0380882
R47196 ASIG5V.n1360 ASIG5V.n1359 0.0380882
R47197 ASIG5V.n1359 ASIG5V.n1358 0.0380882
R47198 ASIG5V.n1358 ASIG5V.n1357 0.0380882
R47199 ASIG5V.n1357 ASIG5V.n1356 0.0380882
R47200 ASIG5V.n1356 ASIG5V.n1355 0.0380882
R47201 ASIG5V.n1355 ASIG5V.n1354 0.0380882
R47202 ASIG5V.n1354 ASIG5V.n1353 0.0380882
R47203 ASIG5V.n1353 ASIG5V.n1352 0.0380882
R47204 ASIG5V.n1352 ASIG5V.n1351 0.0380882
R47205 ASIG5V.n1351 ASIG5V.n1350 0.0380882
R47206 ASIG5V.n1350 ASIG5V.n1349 0.0380882
R47207 ASIG5V.n1349 ASIG5V.n1348 0.0380882
R47208 ASIG5V.n1348 ASIG5V.n1347 0.0380882
R47209 ASIG5V.n1347 ASIG5V.n1346 0.0380882
R47210 ASIG5V.n1346 ASIG5V.n1345 0.0380882
R47211 ASIG5V.n1345 ASIG5V.n1344 0.0380882
R47212 ASIG5V.n1344 ASIG5V.n1343 0.0380882
R47213 ASIG5V.n1343 ASIG5V.n1342 0.0380882
R47214 ASIG5V.n1342 ASIG5V.n1341 0.0380882
R47215 ASIG5V.n1341 ASIG5V.n1340 0.0380882
R47216 ASIG5V.n1340 ASIG5V.n1339 0.0380882
R47217 ASIG5V.n1339 ASIG5V.n1338 0.0380882
R47218 ASIG5V.n1338 ASIG5V.n1337 0.0380882
R47219 ASIG5V.n1337 ASIG5V.n1336 0.0380882
R47220 ASIG5V.n1336 ASIG5V.n1335 0.0380882
R47221 ASIG5V.n1335 ASIG5V.n1334 0.0380882
R47222 ASIG5V.n1334 ASIG5V.n1333 0.0380882
R47223 ASIG5V.n1333 ASIG5V.n1332 0.0380882
R47224 ASIG5V.n1332 ASIG5V.n1331 0.0380882
R47225 ASIG5V.n1331 ASIG5V.n1330 0.0380882
R47226 ASIG5V.n1330 ASIG5V.n1329 0.0380882
R47227 ASIG5V.n1329 ASIG5V.n1328 0.0380882
R47228 ASIG5V.n1328 ASIG5V.n1327 0.0380882
R47229 ASIG5V.n1327 ASIG5V.n1326 0.0380882
R47230 ASIG5V.n1326 ASIG5V.n1325 0.0380882
R47231 ASIG5V.n1325 ASIG5V.n1324 0.0380882
R47232 ASIG5V.n1324 ASIG5V.n1323 0.0380882
R47233 ASIG5V.n1323 ASIG5V.n1322 0.0380882
R47234 ASIG5V.n1322 ASIG5V.n1321 0.0380882
R47235 ASIG5V.n1321 ASIG5V.n1320 0.0380882
R47236 ASIG5V.n1320 ASIG5V.n1319 0.0380882
R47237 ASIG5V.n1319 ASIG5V.n1318 0.0380882
R47238 ASIG5V.n1318 ASIG5V.n1317 0.0380882
R47239 ASIG5V.n1317 ASIG5V.n1316 0.0380882
R47240 ASIG5V.n1316 ASIG5V.n1315 0.0380882
R47241 ASIG5V.n807 ASIG5V.n806 0.0380882
R47242 ASIG5V.n808 ASIG5V.n807 0.0380882
R47243 ASIG5V.n809 ASIG5V.n808 0.0380882
R47244 ASIG5V.n810 ASIG5V.n809 0.0380882
R47245 ASIG5V.n811 ASIG5V.n810 0.0380882
R47246 ASIG5V.n812 ASIG5V.n811 0.0380882
R47247 ASIG5V.n813 ASIG5V.n812 0.0380882
R47248 ASIG5V.n814 ASIG5V.n813 0.0380882
R47249 ASIG5V.n815 ASIG5V.n814 0.0380882
R47250 ASIG5V.n816 ASIG5V.n815 0.0380882
R47251 ASIG5V.n817 ASIG5V.n816 0.0380882
R47252 ASIG5V.n818 ASIG5V.n817 0.0380882
R47253 ASIG5V.n819 ASIG5V.n818 0.0380882
R47254 ASIG5V.n820 ASIG5V.n819 0.0380882
R47255 ASIG5V.n821 ASIG5V.n820 0.0380882
R47256 ASIG5V.n822 ASIG5V.n821 0.0380882
R47257 ASIG5V.n823 ASIG5V.n822 0.0380882
R47258 ASIG5V.n824 ASIG5V.n823 0.0380882
R47259 ASIG5V.n825 ASIG5V.n824 0.0380882
R47260 ASIG5V.n826 ASIG5V.n825 0.0380882
R47261 ASIG5V.n827 ASIG5V.n826 0.0380882
R47262 ASIG5V.n828 ASIG5V.n827 0.0380882
R47263 ASIG5V.n829 ASIG5V.n828 0.0380882
R47264 ASIG5V.n830 ASIG5V.n829 0.0380882
R47265 ASIG5V.n831 ASIG5V.n830 0.0380882
R47266 ASIG5V.n832 ASIG5V.n831 0.0380882
R47267 ASIG5V.n3619 ASIG5V.n3618 0.0380882
R47268 ASIG5V.n3618 ASIG5V.n3617 0.0380882
R47269 ASIG5V.n3617 ASIG5V.n3616 0.0380882
R47270 ASIG5V.n3616 ASIG5V.n3615 0.0380882
R47271 ASIG5V.n3615 ASIG5V.n3614 0.0380882
R47272 ASIG5V.n3614 ASIG5V.n3613 0.0380882
R47273 ASIG5V.n3613 ASIG5V.n3612 0.0380882
R47274 ASIG5V.n3612 ASIG5V.n3611 0.0380882
R47275 ASIG5V.n3611 ASIG5V.n3610 0.0380882
R47276 ASIG5V.n3610 ASIG5V.n3609 0.0380882
R47277 ASIG5V.n3609 ASIG5V.n3608 0.0380882
R47278 ASIG5V.n3608 ASIG5V.n3607 0.0380882
R47279 ASIG5V.n3607 ASIG5V.n3606 0.0380882
R47280 ASIG5V.n3606 ASIG5V.n3605 0.0380882
R47281 ASIG5V.n3605 ASIG5V.n3604 0.0380882
R47282 ASIG5V.n3604 ASIG5V.n3603 0.0380882
R47283 ASIG5V.n3603 ASIG5V.n3602 0.0380882
R47284 ASIG5V.n3602 ASIG5V.n3601 0.0380882
R47285 ASIG5V.n3601 ASIG5V.n3600 0.0380882
R47286 ASIG5V.n3600 ASIG5V.n3599 0.0380882
R47287 ASIG5V.n3599 ASIG5V.n3598 0.0380882
R47288 ASIG5V.n3598 ASIG5V.n3597 0.0380882
R47289 ASIG5V.n3597 ASIG5V.n3596 0.0380882
R47290 ASIG5V.n3596 ASIG5V.n3595 0.0380882
R47291 ASIG5V.n3595 ASIG5V.n3594 0.0380882
R47292 ASIG5V.n3594 ASIG5V.n3593 0.0380882
R47293 ASIG5V.n3593 ASIG5V.n3592 0.0380882
R47294 ASIG5V.n3592 ASIG5V.n3591 0.0380882
R47295 ASIG5V.n3591 ASIG5V.n3590 0.0380882
R47296 ASIG5V.n3590 ASIG5V.n3589 0.0380882
R47297 ASIG5V.n675 ASIG5V.n674 0.0380882
R47298 ASIG5V.n676 ASIG5V.n675 0.0380882
R47299 ASIG5V.n677 ASIG5V.n676 0.0380882
R47300 ASIG5V.n678 ASIG5V.n677 0.0380882
R47301 ASIG5V.n679 ASIG5V.n678 0.0380882
R47302 ASIG5V.n680 ASIG5V.n679 0.0380882
R47303 ASIG5V.n681 ASIG5V.n680 0.0380882
R47304 ASIG5V.n682 ASIG5V.n681 0.0380882
R47305 ASIG5V.n683 ASIG5V.n682 0.0380882
R47306 ASIG5V.n1728 ASIG5V.n1727 0.0380882
R47307 ASIG5V.n1727 ASIG5V.n1726 0.0380882
R47308 ASIG5V.n1726 ASIG5V.n1725 0.0380882
R47309 ASIG5V.n1725 ASIG5V.n1724 0.0380882
R47310 ASIG5V.n1724 ASIG5V.n1723 0.0380882
R47311 ASIG5V.n1723 ASIG5V.n1722 0.0380882
R47312 ASIG5V.n1722 ASIG5V.n1721 0.0380882
R47313 ASIG5V.n1721 ASIG5V.n1720 0.0380882
R47314 ASIG5V.n1720 ASIG5V.n1719 0.0380882
R47315 ASIG5V.n1719 ASIG5V.n1718 0.0380882
R47316 ASIG5V.n1718 ASIG5V.n1717 0.0380882
R47317 ASIG5V.n1717 ASIG5V.n1716 0.0380882
R47318 ASIG5V.n1716 ASIG5V.n1715 0.0380882
R47319 ASIG5V.n1715 ASIG5V.n1714 0.0380882
R47320 ASIG5V.n1714 ASIG5V.n1713 0.0380882
R47321 ASIG5V.n1713 ASIG5V.n1712 0.0380882
R47322 ASIG5V.n1712 ASIG5V.n1711 0.0380882
R47323 ASIG5V.n1711 ASIG5V.n1710 0.0380882
R47324 ASIG5V.n1710 ASIG5V.n1709 0.0380882
R47325 ASIG5V.n1709 ASIG5V.n1708 0.0380882
R47326 ASIG5V.n1708 ASIG5V.n1707 0.0380882
R47327 ASIG5V.n1707 ASIG5V.n1706 0.0380882
R47328 ASIG5V.n1706 ASIG5V.n1705 0.0380882
R47329 ASIG5V.n1705 ASIG5V.n1704 0.0380882
R47330 ASIG5V.n1704 ASIG5V.n1703 0.0380882
R47331 ASIG5V.n1703 ASIG5V.n1702 0.0380882
R47332 ASIG5V.n1702 ASIG5V.n1701 0.0380882
R47333 ASIG5V.n1701 ASIG5V.n1700 0.0380882
R47334 ASIG5V.n1700 ASIG5V.n1699 0.0380882
R47335 ASIG5V.n1699 ASIG5V.n1698 0.0380882
R47336 ASIG5V.n1698 ASIG5V.n1697 0.0380882
R47337 ASIG5V.n1697 ASIG5V.n1696 0.0380882
R47338 ASIG5V.n1696 ASIG5V.n1695 0.0380882
R47339 ASIG5V.n1695 ASIG5V.n1694 0.0380882
R47340 ASIG5V.n1694 ASIG5V.n1693 0.0380882
R47341 ASIG5V.n1693 ASIG5V.n1692 0.0380882
R47342 ASIG5V.n1692 ASIG5V.n1691 0.0380882
R47343 ASIG5V.n1691 ASIG5V.n1690 0.0380882
R47344 ASIG5V.n1690 ASIG5V.n1689 0.0380882
R47345 ASIG5V.n1689 ASIG5V.n1688 0.0380882
R47346 ASIG5V.n1688 ASIG5V.n1687 0.0380882
R47347 ASIG5V.n1687 ASIG5V.n1686 0.0380882
R47348 ASIG5V.n1686 ASIG5V.n1685 0.0380882
R47349 ASIG5V.n1685 ASIG5V.n1684 0.0380882
R47350 ASIG5V.n1684 ASIG5V.n1683 0.0380882
R47351 ASIG5V.n1683 ASIG5V.n1682 0.0380882
R47352 ASIG5V.n1682 ASIG5V.n1681 0.0380882
R47353 ASIG5V.n1681 ASIG5V.n1680 0.0380882
R47354 ASIG5V.n1680 ASIG5V.n1679 0.0380882
R47355 ASIG5V.n1679 ASIG5V.n1678 0.0380882
R47356 ASIG5V.n1678 ASIG5V.n1677 0.0380882
R47357 ASIG5V.n1677 ASIG5V.n1676 0.0380882
R47358 ASIG5V.n834 ASIG5V.n833 0.0380882
R47359 ASIG5V.n835 ASIG5V.n834 0.0380882
R47360 ASIG5V.n836 ASIG5V.n835 0.0380882
R47361 ASIG5V.n837 ASIG5V.n836 0.0380882
R47362 ASIG5V.n838 ASIG5V.n837 0.0380882
R47363 ASIG5V.n839 ASIG5V.n838 0.0380882
R47364 ASIG5V.n840 ASIG5V.n839 0.0380882
R47365 ASIG5V.n841 ASIG5V.n840 0.0380882
R47366 ASIG5V.n842 ASIG5V.n841 0.0380882
R47367 ASIG5V.n843 ASIG5V.n842 0.0380882
R47368 ASIG5V.n844 ASIG5V.n843 0.0380882
R47369 ASIG5V.n845 ASIG5V.n844 0.0380882
R47370 ASIG5V.n846 ASIG5V.n845 0.0380882
R47371 ASIG5V.n847 ASIG5V.n846 0.0380882
R47372 ASIG5V.n848 ASIG5V.n847 0.0380882
R47373 ASIG5V.n849 ASIG5V.n848 0.0380882
R47374 ASIG5V.n850 ASIG5V.n849 0.0380882
R47375 ASIG5V.n851 ASIG5V.n850 0.0380882
R47376 ASIG5V.n852 ASIG5V.n851 0.0380882
R47377 ASIG5V.n853 ASIG5V.n852 0.0380882
R47378 ASIG5V.n854 ASIG5V.n853 0.0380882
R47379 ASIG5V.n855 ASIG5V.n854 0.0380882
R47380 ASIG5V.n856 ASIG5V.n855 0.0380882
R47381 ASIG5V.n857 ASIG5V.n856 0.0380882
R47382 ASIG5V.n3893 ASIG5V.n3892 0.0380882
R47383 ASIG5V.n3892 ASIG5V.n3891 0.0380882
R47384 ASIG5V.n3891 ASIG5V.n3890 0.0380882
R47385 ASIG5V.n3890 ASIG5V.n3889 0.0380882
R47386 ASIG5V.n3889 ASIG5V.n3888 0.0380882
R47387 ASIG5V.n3888 ASIG5V.n3887 0.0380882
R47388 ASIG5V.n3887 ASIG5V.n3886 0.0380882
R47389 ASIG5V.n3886 ASIG5V.n3885 0.0380882
R47390 ASIG5V.n3885 ASIG5V.n3884 0.0380882
R47391 ASIG5V.n3884 ASIG5V.n3883 0.0380882
R47392 ASIG5V.n3883 ASIG5V.n3882 0.0380882
R47393 ASIG5V.n3882 ASIG5V.n3881 0.0380882
R47394 ASIG5V.n3881 ASIG5V.n3880 0.0380882
R47395 ASIG5V.n3880 ASIG5V.n3879 0.0380882
R47396 ASIG5V.n3879 ASIG5V.n3878 0.0380882
R47397 ASIG5V.n3878 ASIG5V.n3877 0.0380882
R47398 ASIG5V.n3877 ASIG5V.n3876 0.0380882
R47399 ASIG5V.n3876 ASIG5V.n3875 0.0380882
R47400 ASIG5V.n3875 ASIG5V.n3874 0.0380882
R47401 ASIG5V.n3874 ASIG5V.n3873 0.0380882
R47402 ASIG5V.n3873 ASIG5V.n3872 0.0380882
R47403 ASIG5V.n3872 ASIG5V.n3871 0.0380882
R47404 ASIG5V.n3871 ASIG5V.n3870 0.0380882
R47405 ASIG5V.n3870 ASIG5V.n3869 0.0380882
R47406 ASIG5V.n3869 ASIG5V.n3868 0.0380882
R47407 ASIG5V.n3868 ASIG5V.n3867 0.0380882
R47408 ASIG5V.n3867 ASIG5V.n3866 0.0380882
R47409 ASIG5V.n3866 ASIG5V.n3865 0.0380882
R47410 ASIG5V.n3865 ASIG5V.n3864 0.0380882
R47411 ASIG5V.n3864 ASIG5V.n3863 0.0380882
R47412 ASIG5V.n685 ASIG5V.n684 0.0380882
R47413 ASIG5V.n686 ASIG5V.n685 0.0380882
R47414 ASIG5V.n687 ASIG5V.n686 0.0380882
R47415 ASIG5V.n688 ASIG5V.n687 0.0380882
R47416 ASIG5V.n689 ASIG5V.n688 0.0380882
R47417 ASIG5V.n690 ASIG5V.n689 0.0380882
R47418 ASIG5V.n691 ASIG5V.n690 0.0380882
R47419 ASIG5V.n1780 ASIG5V.n1779 0.0380882
R47420 ASIG5V.n1779 ASIG5V.n1778 0.0380882
R47421 ASIG5V.n1778 ASIG5V.n1777 0.0380882
R47422 ASIG5V.n1777 ASIG5V.n1776 0.0380882
R47423 ASIG5V.n1776 ASIG5V.n1775 0.0380882
R47424 ASIG5V.n1775 ASIG5V.n1774 0.0380882
R47425 ASIG5V.n1774 ASIG5V.n1773 0.0380882
R47426 ASIG5V.n1773 ASIG5V.n1772 0.0380882
R47427 ASIG5V.n1772 ASIG5V.n1771 0.0380882
R47428 ASIG5V.n1771 ASIG5V.n1770 0.0380882
R47429 ASIG5V.n1770 ASIG5V.n1769 0.0380882
R47430 ASIG5V.n1769 ASIG5V.n1768 0.0380882
R47431 ASIG5V.n1768 ASIG5V.n1767 0.0380882
R47432 ASIG5V.n1767 ASIG5V.n1766 0.0380882
R47433 ASIG5V.n1766 ASIG5V.n1765 0.0380882
R47434 ASIG5V.n1765 ASIG5V.n1764 0.0380882
R47435 ASIG5V.n1764 ASIG5V.n1763 0.0380882
R47436 ASIG5V.n1763 ASIG5V.n1762 0.0380882
R47437 ASIG5V.n1762 ASIG5V.n1761 0.0380882
R47438 ASIG5V.n1761 ASIG5V.n1760 0.0380882
R47439 ASIG5V.n1760 ASIG5V.n1759 0.0380882
R47440 ASIG5V.n1759 ASIG5V.n1758 0.0380882
R47441 ASIG5V.n1758 ASIG5V.n1757 0.0380882
R47442 ASIG5V.n1757 ASIG5V.n1756 0.0380882
R47443 ASIG5V.n1756 ASIG5V.n1755 0.0380882
R47444 ASIG5V.n1755 ASIG5V.n1754 0.0380882
R47445 ASIG5V.n1754 ASIG5V.n1753 0.0380882
R47446 ASIG5V.n1753 ASIG5V.n1752 0.0380882
R47447 ASIG5V.n1752 ASIG5V.n1751 0.0380882
R47448 ASIG5V.n1751 ASIG5V.n1750 0.0380882
R47449 ASIG5V.n1750 ASIG5V.n1749 0.0380882
R47450 ASIG5V.n1749 ASIG5V.n1748 0.0380882
R47451 ASIG5V.n1748 ASIG5V.n1747 0.0380882
R47452 ASIG5V.n1747 ASIG5V.n1746 0.0380882
R47453 ASIG5V.n1746 ASIG5V.n1745 0.0380882
R47454 ASIG5V.n1745 ASIG5V.n1744 0.0380882
R47455 ASIG5V.n1744 ASIG5V.n1743 0.0380882
R47456 ASIG5V.n1743 ASIG5V.n1742 0.0380882
R47457 ASIG5V.n1742 ASIG5V.n1741 0.0380882
R47458 ASIG5V.n1741 ASIG5V.n1740 0.0380882
R47459 ASIG5V.n1740 ASIG5V.n1739 0.0380882
R47460 ASIG5V.n1739 ASIG5V.n1738 0.0380882
R47461 ASIG5V.n1738 ASIG5V.n1737 0.0380882
R47462 ASIG5V.n1737 ASIG5V.n1736 0.0380882
R47463 ASIG5V.n1736 ASIG5V.n1735 0.0380882
R47464 ASIG5V.n1735 ASIG5V.n1734 0.0380882
R47465 ASIG5V.n1734 ASIG5V.n1733 0.0380882
R47466 ASIG5V.n1733 ASIG5V.n1732 0.0380882
R47467 ASIG5V.n1732 ASIG5V.n1731 0.0380882
R47468 ASIG5V.n1731 ASIG5V.n1730 0.0380882
R47469 ASIG5V.n1730 ASIG5V.n1729 0.0380882
R47470 ASIG5V.n859 ASIG5V.n858 0.0380882
R47471 ASIG5V.n860 ASIG5V.n859 0.0380882
R47472 ASIG5V.n861 ASIG5V.n860 0.0380882
R47473 ASIG5V.n862 ASIG5V.n861 0.0380882
R47474 ASIG5V.n863 ASIG5V.n862 0.0380882
R47475 ASIG5V.n864 ASIG5V.n863 0.0380882
R47476 ASIG5V.n865 ASIG5V.n864 0.0380882
R47477 ASIG5V.n866 ASIG5V.n865 0.0380882
R47478 ASIG5V.n867 ASIG5V.n866 0.0380882
R47479 ASIG5V.n868 ASIG5V.n867 0.0380882
R47480 ASIG5V.n869 ASIG5V.n868 0.0380882
R47481 ASIG5V.n870 ASIG5V.n869 0.0380882
R47482 ASIG5V.n871 ASIG5V.n870 0.0380882
R47483 ASIG5V.n872 ASIG5V.n871 0.0380882
R47484 ASIG5V.n873 ASIG5V.n872 0.0380882
R47485 ASIG5V.n874 ASIG5V.n873 0.0380882
R47486 ASIG5V.n875 ASIG5V.n874 0.0380882
R47487 ASIG5V.n876 ASIG5V.n875 0.0380882
R47488 ASIG5V.n877 ASIG5V.n876 0.0380882
R47489 ASIG5V.n878 ASIG5V.n877 0.0380882
R47490 ASIG5V.n879 ASIG5V.n878 0.0380882
R47491 ASIG5V.n4160 ASIG5V.n4159 0.0380882
R47492 ASIG5V.n4159 ASIG5V.n4158 0.0380882
R47493 ASIG5V.n4158 ASIG5V.n4157 0.0380882
R47494 ASIG5V.n4157 ASIG5V.n4156 0.0380882
R47495 ASIG5V.n4156 ASIG5V.n4155 0.0380882
R47496 ASIG5V.n4155 ASIG5V.n4154 0.0380882
R47497 ASIG5V.n4154 ASIG5V.n4153 0.0380882
R47498 ASIG5V.n4153 ASIG5V.n4152 0.0380882
R47499 ASIG5V.n4152 ASIG5V.n4151 0.0380882
R47500 ASIG5V.n4151 ASIG5V.n4150 0.0380882
R47501 ASIG5V.n4150 ASIG5V.n4149 0.0380882
R47502 ASIG5V.n4149 ASIG5V.n4148 0.0380882
R47503 ASIG5V.n4148 ASIG5V.n4147 0.0380882
R47504 ASIG5V.n4147 ASIG5V.n4146 0.0380882
R47505 ASIG5V.n4146 ASIG5V.n4145 0.0380882
R47506 ASIG5V.n4145 ASIG5V.n4144 0.0380882
R47507 ASIG5V.n4144 ASIG5V.n4143 0.0380882
R47508 ASIG5V.n4143 ASIG5V.n4142 0.0380882
R47509 ASIG5V.n4142 ASIG5V.n4141 0.0380882
R47510 ASIG5V.n4141 ASIG5V.n4140 0.0380882
R47511 ASIG5V.n4140 ASIG5V.n4139 0.0380882
R47512 ASIG5V.n4139 ASIG5V.n4138 0.0380882
R47513 ASIG5V.n4138 ASIG5V.n4137 0.0380882
R47514 ASIG5V.n4137 ASIG5V.n4136 0.0380882
R47515 ASIG5V.n4136 ASIG5V.n4135 0.0380882
R47516 ASIG5V.n4135 ASIG5V.n4134 0.0380882
R47517 ASIG5V.n4134 ASIG5V.n4133 0.0380882
R47518 ASIG5V.n4133 ASIG5V.n4132 0.0380882
R47519 ASIG5V.n4132 ASIG5V.n4131 0.0380882
R47520 ASIG5V.n4131 ASIG5V.n4130 0.0380882
R47521 ASIG5V.n693 ASIG5V.n692 0.0380882
R47522 ASIG5V.n694 ASIG5V.n693 0.0380882
R47523 ASIG5V.n695 ASIG5V.n694 0.0380882
R47524 ASIG5V.n696 ASIG5V.n695 0.0380882
R47525 ASIG5V.n697 ASIG5V.n696 0.0380882
R47526 ASIG5V.n1830 ASIG5V.n1829 0.0380882
R47527 ASIG5V.n1829 ASIG5V.n1828 0.0380882
R47528 ASIG5V.n1828 ASIG5V.n1827 0.0380882
R47529 ASIG5V.n1827 ASIG5V.n1826 0.0380882
R47530 ASIG5V.n1826 ASIG5V.n1825 0.0380882
R47531 ASIG5V.n1825 ASIG5V.n1824 0.0380882
R47532 ASIG5V.n1824 ASIG5V.n1823 0.0380882
R47533 ASIG5V.n1823 ASIG5V.n1822 0.0380882
R47534 ASIG5V.n1822 ASIG5V.n1821 0.0380882
R47535 ASIG5V.n1821 ASIG5V.n1820 0.0380882
R47536 ASIG5V.n1820 ASIG5V.n1819 0.0380882
R47537 ASIG5V.n1819 ASIG5V.n1818 0.0380882
R47538 ASIG5V.n1818 ASIG5V.n1817 0.0380882
R47539 ASIG5V.n1817 ASIG5V.n1816 0.0380882
R47540 ASIG5V.n1816 ASIG5V.n1815 0.0380882
R47541 ASIG5V.n1815 ASIG5V.n1814 0.0380882
R47542 ASIG5V.n1814 ASIG5V.n1813 0.0380882
R47543 ASIG5V.n1813 ASIG5V.n1812 0.0380882
R47544 ASIG5V.n1812 ASIG5V.n1811 0.0380882
R47545 ASIG5V.n1811 ASIG5V.n1810 0.0380882
R47546 ASIG5V.n1810 ASIG5V.n1809 0.0380882
R47547 ASIG5V.n1809 ASIG5V.n1808 0.0380882
R47548 ASIG5V.n1808 ASIG5V.n1807 0.0380882
R47549 ASIG5V.n1807 ASIG5V.n1806 0.0380882
R47550 ASIG5V.n1806 ASIG5V.n1805 0.0380882
R47551 ASIG5V.n1805 ASIG5V.n1804 0.0380882
R47552 ASIG5V.n1804 ASIG5V.n1803 0.0380882
R47553 ASIG5V.n1803 ASIG5V.n1802 0.0380882
R47554 ASIG5V.n1802 ASIG5V.n1801 0.0380882
R47555 ASIG5V.n1801 ASIG5V.n1800 0.0380882
R47556 ASIG5V.n1800 ASIG5V.n1799 0.0380882
R47557 ASIG5V.n1799 ASIG5V.n1798 0.0380882
R47558 ASIG5V.n1798 ASIG5V.n1797 0.0380882
R47559 ASIG5V.n1797 ASIG5V.n1796 0.0380882
R47560 ASIG5V.n1796 ASIG5V.n1795 0.0380882
R47561 ASIG5V.n1795 ASIG5V.n1794 0.0380882
R47562 ASIG5V.n1794 ASIG5V.n1793 0.0380882
R47563 ASIG5V.n1793 ASIG5V.n1792 0.0380882
R47564 ASIG5V.n1792 ASIG5V.n1791 0.0380882
R47565 ASIG5V.n1791 ASIG5V.n1790 0.0380882
R47566 ASIG5V.n1790 ASIG5V.n1789 0.0380882
R47567 ASIG5V.n1789 ASIG5V.n1788 0.0380882
R47568 ASIG5V.n1788 ASIG5V.n1787 0.0380882
R47569 ASIG5V.n1787 ASIG5V.n1786 0.0380882
R47570 ASIG5V.n1786 ASIG5V.n1785 0.0380882
R47571 ASIG5V.n1785 ASIG5V.n1784 0.0380882
R47572 ASIG5V.n1784 ASIG5V.n1783 0.0380882
R47573 ASIG5V.n1783 ASIG5V.n1782 0.0380882
R47574 ASIG5V.n1782 ASIG5V.n1781 0.0380882
R47575 ASIG5V.n881 ASIG5V.n880 0.0380882
R47576 ASIG5V.n882 ASIG5V.n881 0.0380882
R47577 ASIG5V.n883 ASIG5V.n882 0.0380882
R47578 ASIG5V.n884 ASIG5V.n883 0.0380882
R47579 ASIG5V.n885 ASIG5V.n884 0.0380882
R47580 ASIG5V.n886 ASIG5V.n885 0.0380882
R47581 ASIG5V.n887 ASIG5V.n886 0.0380882
R47582 ASIG5V.n888 ASIG5V.n887 0.0380882
R47583 ASIG5V.n889 ASIG5V.n888 0.0380882
R47584 ASIG5V.n890 ASIG5V.n889 0.0380882
R47585 ASIG5V.n891 ASIG5V.n890 0.0380882
R47586 ASIG5V.n892 ASIG5V.n891 0.0380882
R47587 ASIG5V.n893 ASIG5V.n892 0.0380882
R47588 ASIG5V.n894 ASIG5V.n893 0.0380882
R47589 ASIG5V.n895 ASIG5V.n894 0.0380882
R47590 ASIG5V.n896 ASIG5V.n895 0.0380882
R47591 ASIG5V.n897 ASIG5V.n896 0.0380882
R47592 ASIG5V.n898 ASIG5V.n897 0.0380882
R47593 ASIG5V.n899 ASIG5V.n898 0.0380882
R47594 ASIG5V.n4436 ASIG5V.n4435 0.0380882
R47595 ASIG5V.n4435 ASIG5V.n4434 0.0380882
R47596 ASIG5V.n4434 ASIG5V.n4433 0.0380882
R47597 ASIG5V.n4433 ASIG5V.n4432 0.0380882
R47598 ASIG5V.n4432 ASIG5V.n4431 0.0380882
R47599 ASIG5V.n4431 ASIG5V.n4430 0.0380882
R47600 ASIG5V.n4430 ASIG5V.n4429 0.0380882
R47601 ASIG5V.n4429 ASIG5V.n4428 0.0380882
R47602 ASIG5V.n4428 ASIG5V.n4427 0.0380882
R47603 ASIG5V.n4427 ASIG5V.n4426 0.0380882
R47604 ASIG5V.n4426 ASIG5V.n4425 0.0380882
R47605 ASIG5V.n4425 ASIG5V.n4424 0.0380882
R47606 ASIG5V.n4424 ASIG5V.n4423 0.0380882
R47607 ASIG5V.n4423 ASIG5V.n4422 0.0380882
R47608 ASIG5V.n4422 ASIG5V.n4421 0.0380882
R47609 ASIG5V.n4421 ASIG5V.n4420 0.0380882
R47610 ASIG5V.n4420 ASIG5V.n4419 0.0380882
R47611 ASIG5V.n4419 ASIG5V.n4418 0.0380882
R47612 ASIG5V.n4418 ASIG5V.n4417 0.0380882
R47613 ASIG5V.n4417 ASIG5V.n4416 0.0380882
R47614 ASIG5V.n4416 ASIG5V.n4415 0.0380882
R47615 ASIG5V.n4415 ASIG5V.n4414 0.0380882
R47616 ASIG5V.n4414 ASIG5V.n4413 0.0380882
R47617 ASIG5V.n4413 ASIG5V.n4412 0.0380882
R47618 ASIG5V.n4412 ASIG5V.n4411 0.0380882
R47619 ASIG5V.n4411 ASIG5V.n4410 0.0380882
R47620 ASIG5V.n4410 ASIG5V.n4409 0.0380882
R47621 ASIG5V.n4409 ASIG5V.n4408 0.0380882
R47622 ASIG5V.n4408 ASIG5V.n4407 0.0380882
R47623 ASIG5V.n4407 ASIG5V.n4406 0.0380882
R47624 ASIG5V.n699 ASIG5V.n698 0.0380882
R47625 ASIG5V.n700 ASIG5V.n699 0.0380882
R47626 ASIG5V.n701 ASIG5V.n700 0.0380882
R47627 ASIG5V.n1879 ASIG5V.n1878 0.0380882
R47628 ASIG5V.n1878 ASIG5V.n1877 0.0380882
R47629 ASIG5V.n1877 ASIG5V.n1876 0.0380882
R47630 ASIG5V.n1876 ASIG5V.n1875 0.0380882
R47631 ASIG5V.n1875 ASIG5V.n1874 0.0380882
R47632 ASIG5V.n1874 ASIG5V.n1873 0.0380882
R47633 ASIG5V.n1873 ASIG5V.n1872 0.0380882
R47634 ASIG5V.n1872 ASIG5V.n1871 0.0380882
R47635 ASIG5V.n1871 ASIG5V.n1870 0.0380882
R47636 ASIG5V.n1870 ASIG5V.n1869 0.0380882
R47637 ASIG5V.n1869 ASIG5V.n1868 0.0380882
R47638 ASIG5V.n1868 ASIG5V.n1867 0.0380882
R47639 ASIG5V.n1867 ASIG5V.n1866 0.0380882
R47640 ASIG5V.n1866 ASIG5V.n1865 0.0380882
R47641 ASIG5V.n1865 ASIG5V.n1864 0.0380882
R47642 ASIG5V.n1864 ASIG5V.n1863 0.0380882
R47643 ASIG5V.n1863 ASIG5V.n1862 0.0380882
R47644 ASIG5V.n1862 ASIG5V.n1861 0.0380882
R47645 ASIG5V.n1861 ASIG5V.n1860 0.0380882
R47646 ASIG5V.n1860 ASIG5V.n1859 0.0380882
R47647 ASIG5V.n1859 ASIG5V.n1858 0.0380882
R47648 ASIG5V.n1858 ASIG5V.n1857 0.0380882
R47649 ASIG5V.n1857 ASIG5V.n1856 0.0380882
R47650 ASIG5V.n1856 ASIG5V.n1855 0.0380882
R47651 ASIG5V.n1855 ASIG5V.n1854 0.0380882
R47652 ASIG5V.n1854 ASIG5V.n1853 0.0380882
R47653 ASIG5V.n1853 ASIG5V.n1852 0.0380882
R47654 ASIG5V.n1852 ASIG5V.n1851 0.0380882
R47655 ASIG5V.n1851 ASIG5V.n1850 0.0380882
R47656 ASIG5V.n1850 ASIG5V.n1849 0.0380882
R47657 ASIG5V.n1849 ASIG5V.n1848 0.0380882
R47658 ASIG5V.n1848 ASIG5V.n1847 0.0380882
R47659 ASIG5V.n1847 ASIG5V.n1846 0.0380882
R47660 ASIG5V.n1846 ASIG5V.n1845 0.0380882
R47661 ASIG5V.n1845 ASIG5V.n1844 0.0380882
R47662 ASIG5V.n1844 ASIG5V.n1843 0.0380882
R47663 ASIG5V.n1843 ASIG5V.n1842 0.0380882
R47664 ASIG5V.n1842 ASIG5V.n1841 0.0380882
R47665 ASIG5V.n1841 ASIG5V.n1840 0.0380882
R47666 ASIG5V.n1840 ASIG5V.n1839 0.0380882
R47667 ASIG5V.n1839 ASIG5V.n1838 0.0380882
R47668 ASIG5V.n1838 ASIG5V.n1837 0.0380882
R47669 ASIG5V.n1837 ASIG5V.n1836 0.0380882
R47670 ASIG5V.n1836 ASIG5V.n1835 0.0380882
R47671 ASIG5V.n1835 ASIG5V.n1834 0.0380882
R47672 ASIG5V.n1834 ASIG5V.n1833 0.0380882
R47673 ASIG5V.n1833 ASIG5V.n1832 0.0380882
R47674 ASIG5V.n1832 ASIG5V.n1831 0.0380882
R47675 ASIG5V.n901 ASIG5V.n900 0.0380882
R47676 ASIG5V.n902 ASIG5V.n901 0.0380882
R47677 ASIG5V.n903 ASIG5V.n902 0.0380882
R47678 ASIG5V.n904 ASIG5V.n903 0.0380882
R47679 ASIG5V.n905 ASIG5V.n904 0.0380882
R47680 ASIG5V.n906 ASIG5V.n905 0.0380882
R47681 ASIG5V.n907 ASIG5V.n906 0.0380882
R47682 ASIG5V.n908 ASIG5V.n907 0.0380882
R47683 ASIG5V.n909 ASIG5V.n908 0.0380882
R47684 ASIG5V.n910 ASIG5V.n909 0.0380882
R47685 ASIG5V.n911 ASIG5V.n910 0.0380882
R47686 ASIG5V.n912 ASIG5V.n911 0.0380882
R47687 ASIG5V.n913 ASIG5V.n912 0.0380882
R47688 ASIG5V.n914 ASIG5V.n913 0.0380882
R47689 ASIG5V.n915 ASIG5V.n914 0.0380882
R47690 ASIG5V.n916 ASIG5V.n915 0.0380882
R47691 ASIG5V.n917 ASIG5V.n916 0.0380882
R47692 ASIG5V.n4694 ASIG5V.n4693 0.0380882
R47693 ASIG5V.n4693 ASIG5V.n4692 0.0380882
R47694 ASIG5V.n4692 ASIG5V.n4691 0.0380882
R47695 ASIG5V.n4691 ASIG5V.n4690 0.0380882
R47696 ASIG5V.n4690 ASIG5V.n4689 0.0380882
R47697 ASIG5V.n4689 ASIG5V.n4688 0.0380882
R47698 ASIG5V.n4688 ASIG5V.n4687 0.0380882
R47699 ASIG5V.n4687 ASIG5V.n4686 0.0380882
R47700 ASIG5V.n4686 ASIG5V.n4685 0.0380882
R47701 ASIG5V.n4685 ASIG5V.n4684 0.0380882
R47702 ASIG5V.n4684 ASIG5V.n4683 0.0380882
R47703 ASIG5V.n4683 ASIG5V.n4682 0.0380882
R47704 ASIG5V.n4682 ASIG5V.n4681 0.0380882
R47705 ASIG5V.n4681 ASIG5V.n4680 0.0380882
R47706 ASIG5V.n4680 ASIG5V.n4679 0.0380882
R47707 ASIG5V.n4679 ASIG5V.n4678 0.0380882
R47708 ASIG5V.n4678 ASIG5V.n4677 0.0380882
R47709 ASIG5V.n4677 ASIG5V.n4676 0.0380882
R47710 ASIG5V.n4676 ASIG5V.n4675 0.0380882
R47711 ASIG5V.n4675 ASIG5V.n4674 0.0380882
R47712 ASIG5V.n4674 ASIG5V.n4673 0.0380882
R47713 ASIG5V.n4673 ASIG5V.n4672 0.0380882
R47714 ASIG5V.n4672 ASIG5V.n4671 0.0380882
R47715 ASIG5V.n4671 ASIG5V.n4670 0.0380882
R47716 ASIG5V.n4670 ASIG5V.n4669 0.0380882
R47717 ASIG5V.n4669 ASIG5V.n4668 0.0380882
R47718 ASIG5V.n4668 ASIG5V.n4667 0.0380882
R47719 ASIG5V.n4667 ASIG5V.n4666 0.0380882
R47720 ASIG5V.n4666 ASIG5V.n4665 0.0380882
R47721 ASIG5V.n4665 ASIG5V.n4664 0.0380882
R47722 ASIG5V.n703 ASIG5V.n702 0.0380882
R47723 ASIG5V.n1926 ASIG5V.n1925 0.0380882
R47724 ASIG5V.n1925 ASIG5V.n1924 0.0380882
R47725 ASIG5V.n1924 ASIG5V.n1923 0.0380882
R47726 ASIG5V.n1923 ASIG5V.n1922 0.0380882
R47727 ASIG5V.n1922 ASIG5V.n1921 0.0380882
R47728 ASIG5V.n1921 ASIG5V.n1920 0.0380882
R47729 ASIG5V.n1920 ASIG5V.n1919 0.0380882
R47730 ASIG5V.n1919 ASIG5V.n1918 0.0380882
R47731 ASIG5V.n1918 ASIG5V.n1917 0.0380882
R47732 ASIG5V.n1917 ASIG5V.n1916 0.0380882
R47733 ASIG5V.n1916 ASIG5V.n1915 0.0380882
R47734 ASIG5V.n1915 ASIG5V.n1914 0.0380882
R47735 ASIG5V.n1914 ASIG5V.n1913 0.0380882
R47736 ASIG5V.n1913 ASIG5V.n1912 0.0380882
R47737 ASIG5V.n1912 ASIG5V.n1911 0.0380882
R47738 ASIG5V.n1911 ASIG5V.n1910 0.0380882
R47739 ASIG5V.n1910 ASIG5V.n1909 0.0380882
R47740 ASIG5V.n1909 ASIG5V.n1908 0.0380882
R47741 ASIG5V.n1908 ASIG5V.n1907 0.0380882
R47742 ASIG5V.n1907 ASIG5V.n1906 0.0380882
R47743 ASIG5V.n1906 ASIG5V.n1905 0.0380882
R47744 ASIG5V.n1905 ASIG5V.n1904 0.0380882
R47745 ASIG5V.n1904 ASIG5V.n1903 0.0380882
R47746 ASIG5V.n1903 ASIG5V.n1902 0.0380882
R47747 ASIG5V.n1902 ASIG5V.n1901 0.0380882
R47748 ASIG5V.n1901 ASIG5V.n1900 0.0380882
R47749 ASIG5V.n1900 ASIG5V.n1899 0.0380882
R47750 ASIG5V.n1899 ASIG5V.n1898 0.0380882
R47751 ASIG5V.n1898 ASIG5V.n1897 0.0380882
R47752 ASIG5V.n1897 ASIG5V.n1896 0.0380882
R47753 ASIG5V.n1896 ASIG5V.n1895 0.0380882
R47754 ASIG5V.n1895 ASIG5V.n1894 0.0380882
R47755 ASIG5V.n1894 ASIG5V.n1893 0.0380882
R47756 ASIG5V.n1893 ASIG5V.n1892 0.0380882
R47757 ASIG5V.n1892 ASIG5V.n1891 0.0380882
R47758 ASIG5V.n1891 ASIG5V.n1890 0.0380882
R47759 ASIG5V.n1890 ASIG5V.n1889 0.0380882
R47760 ASIG5V.n1889 ASIG5V.n1888 0.0380882
R47761 ASIG5V.n1888 ASIG5V.n1887 0.0380882
R47762 ASIG5V.n1887 ASIG5V.n1886 0.0380882
R47763 ASIG5V.n1886 ASIG5V.n1885 0.0380882
R47764 ASIG5V.n1885 ASIG5V.n1884 0.0380882
R47765 ASIG5V.n1884 ASIG5V.n1883 0.0380882
R47766 ASIG5V.n1883 ASIG5V.n1882 0.0380882
R47767 ASIG5V.n1882 ASIG5V.n1881 0.0380882
R47768 ASIG5V.n1881 ASIG5V.n1880 0.0380882
R47769 ASIG5V.n919 ASIG5V.n918 0.0380882
R47770 ASIG5V.n920 ASIG5V.n919 0.0380882
R47771 ASIG5V.n921 ASIG5V.n920 0.0380882
R47772 ASIG5V.n922 ASIG5V.n921 0.0380882
R47773 ASIG5V.n923 ASIG5V.n922 0.0380882
R47774 ASIG5V.n924 ASIG5V.n923 0.0380882
R47775 ASIG5V.n925 ASIG5V.n924 0.0380882
R47776 ASIG5V.n926 ASIG5V.n925 0.0380882
R47777 ASIG5V.n927 ASIG5V.n926 0.0380882
R47778 ASIG5V.n928 ASIG5V.n927 0.0380882
R47779 ASIG5V.n929 ASIG5V.n928 0.0380882
R47780 ASIG5V.n930 ASIG5V.n929 0.0380882
R47781 ASIG5V.n931 ASIG5V.n930 0.0380882
R47782 ASIG5V.n932 ASIG5V.n931 0.0380882
R47783 ASIG5V.n4962 ASIG5V.n4961 0.0380882
R47784 ASIG5V.n4961 ASIG5V.n4960 0.0380882
R47785 ASIG5V.n4960 ASIG5V.n4959 0.0380882
R47786 ASIG5V.n4959 ASIG5V.n4958 0.0380882
R47787 ASIG5V.n4958 ASIG5V.n4957 0.0380882
R47788 ASIG5V.n4957 ASIG5V.n4956 0.0380882
R47789 ASIG5V.n4956 ASIG5V.n4955 0.0380882
R47790 ASIG5V.n4955 ASIG5V.n4954 0.0380882
R47791 ASIG5V.n4954 ASIG5V.n4953 0.0380882
R47792 ASIG5V.n4953 ASIG5V.n4952 0.0380882
R47793 ASIG5V.n4952 ASIG5V.n4951 0.0380882
R47794 ASIG5V.n4951 ASIG5V.n4950 0.0380882
R47795 ASIG5V.n4950 ASIG5V.n4949 0.0380882
R47796 ASIG5V.n4949 ASIG5V.n4948 0.0380882
R47797 ASIG5V.n4948 ASIG5V.n4947 0.0380882
R47798 ASIG5V.n4947 ASIG5V.n4946 0.0380882
R47799 ASIG5V.n4946 ASIG5V.n4945 0.0380882
R47800 ASIG5V.n4945 ASIG5V.n4944 0.0380882
R47801 ASIG5V.n4944 ASIG5V.n4943 0.0380882
R47802 ASIG5V.n4943 ASIG5V.n4942 0.0380882
R47803 ASIG5V.n4942 ASIG5V.n4941 0.0380882
R47804 ASIG5V.n4941 ASIG5V.n4940 0.0380882
R47805 ASIG5V.n4940 ASIG5V.n4939 0.0380882
R47806 ASIG5V.n4939 ASIG5V.n4938 0.0380882
R47807 ASIG5V.n4938 ASIG5V.n4937 0.0380882
R47808 ASIG5V.n4937 ASIG5V.n4936 0.0380882
R47809 ASIG5V.n4936 ASIG5V.n4935 0.0380882
R47810 ASIG5V.n4935 ASIG5V.n4934 0.0380882
R47811 ASIG5V.n4934 ASIG5V.n4933 0.0380882
R47812 ASIG5V.n4933 ASIG5V.n4932 0.0380882
R47813 ASIG5V.n1972 ASIG5V.n1971 0.0380882
R47814 ASIG5V.n1971 ASIG5V.n1970 0.0380882
R47815 ASIG5V.n1970 ASIG5V.n1969 0.0380882
R47816 ASIG5V.n1969 ASIG5V.n1968 0.0380882
R47817 ASIG5V.n1968 ASIG5V.n1967 0.0380882
R47818 ASIG5V.n1967 ASIG5V.n1966 0.0380882
R47819 ASIG5V.n1966 ASIG5V.n1965 0.0380882
R47820 ASIG5V.n1965 ASIG5V.n1964 0.0380882
R47821 ASIG5V.n1964 ASIG5V.n1963 0.0380882
R47822 ASIG5V.n1963 ASIG5V.n1962 0.0380882
R47823 ASIG5V.n1962 ASIG5V.n1961 0.0380882
R47824 ASIG5V.n1961 ASIG5V.n1960 0.0380882
R47825 ASIG5V.n1960 ASIG5V.n1959 0.0380882
R47826 ASIG5V.n1959 ASIG5V.n1958 0.0380882
R47827 ASIG5V.n1958 ASIG5V.n1957 0.0380882
R47828 ASIG5V.n1957 ASIG5V.n1956 0.0380882
R47829 ASIG5V.n1956 ASIG5V.n1955 0.0380882
R47830 ASIG5V.n1955 ASIG5V.n1954 0.0380882
R47831 ASIG5V.n1954 ASIG5V.n1953 0.0380882
R47832 ASIG5V.n1953 ASIG5V.n1952 0.0380882
R47833 ASIG5V.n1952 ASIG5V.n1951 0.0380882
R47834 ASIG5V.n1951 ASIG5V.n1950 0.0380882
R47835 ASIG5V.n1950 ASIG5V.n1949 0.0380882
R47836 ASIG5V.n1949 ASIG5V.n1948 0.0380882
R47837 ASIG5V.n1948 ASIG5V.n1947 0.0380882
R47838 ASIG5V.n1947 ASIG5V.n1946 0.0380882
R47839 ASIG5V.n1946 ASIG5V.n1945 0.0380882
R47840 ASIG5V.n1945 ASIG5V.n1944 0.0380882
R47841 ASIG5V.n1944 ASIG5V.n1943 0.0380882
R47842 ASIG5V.n1943 ASIG5V.n1942 0.0380882
R47843 ASIG5V.n1942 ASIG5V.n1941 0.0380882
R47844 ASIG5V.n1941 ASIG5V.n1940 0.0380882
R47845 ASIG5V.n1940 ASIG5V.n1939 0.0380882
R47846 ASIG5V.n1939 ASIG5V.n1938 0.0380882
R47847 ASIG5V.n1938 ASIG5V.n1937 0.0380882
R47848 ASIG5V.n1937 ASIG5V.n1936 0.0380882
R47849 ASIG5V.n1936 ASIG5V.n1935 0.0380882
R47850 ASIG5V.n1935 ASIG5V.n1934 0.0380882
R47851 ASIG5V.n1934 ASIG5V.n1933 0.0380882
R47852 ASIG5V.n1933 ASIG5V.n1932 0.0380882
R47853 ASIG5V.n1932 ASIG5V.n1931 0.0380882
R47854 ASIG5V.n1931 ASIG5V.n1930 0.0380882
R47855 ASIG5V.n1930 ASIG5V.n1929 0.0380882
R47856 ASIG5V.n1929 ASIG5V.n1928 0.0380882
R47857 ASIG5V.n1928 ASIG5V.n1927 0.0380882
R47858 ASIG5V.n934 ASIG5V.n933 0.0380882
R47859 ASIG5V.n935 ASIG5V.n934 0.0380882
R47860 ASIG5V.n936 ASIG5V.n935 0.0380882
R47861 ASIG5V.n937 ASIG5V.n936 0.0380882
R47862 ASIG5V.n938 ASIG5V.n937 0.0380882
R47863 ASIG5V.n939 ASIG5V.n938 0.0380882
R47864 ASIG5V.n940 ASIG5V.n939 0.0380882
R47865 ASIG5V.n941 ASIG5V.n940 0.0380882
R47866 ASIG5V.n942 ASIG5V.n941 0.0380882
R47867 ASIG5V.n943 ASIG5V.n942 0.0380882
R47868 ASIG5V.n944 ASIG5V.n943 0.0380882
R47869 ASIG5V.n945 ASIG5V.n944 0.0380882
R47870 ASIG5V.n5389 ASIG5V.n5388 0.0380882
R47871 ASIG5V.n5388 ASIG5V.n5387 0.0380882
R47872 ASIG5V.n5387 ASIG5V.n5386 0.0380882
R47873 ASIG5V.n5386 ASIG5V.n5385 0.0380882
R47874 ASIG5V.n5385 ASIG5V.n5384 0.0380882
R47875 ASIG5V.n5384 ASIG5V.n5383 0.0380882
R47876 ASIG5V.n5383 ASIG5V.n5382 0.0380882
R47877 ASIG5V.n5382 ASIG5V.n5381 0.0380882
R47878 ASIG5V.n5381 ASIG5V.n5380 0.0380882
R47879 ASIG5V.n5380 ASIG5V.n5379 0.0380882
R47880 ASIG5V.n5379 ASIG5V.n5378 0.0380882
R47881 ASIG5V.n5378 ASIG5V.n5377 0.0380882
R47882 ASIG5V.n5377 ASIG5V.n5376 0.0380882
R47883 ASIG5V.n5376 ASIG5V.n5375 0.0380882
R47884 ASIG5V.n5375 ASIG5V.n5374 0.0380882
R47885 ASIG5V.n5374 ASIG5V.n5373 0.0380882
R47886 ASIG5V.n5373 ASIG5V.n5372 0.0380882
R47887 ASIG5V.n5372 ASIG5V.n5371 0.0380882
R47888 ASIG5V.n5371 ASIG5V.n5370 0.0380882
R47889 ASIG5V.n5370 ASIG5V.n5369 0.0380882
R47890 ASIG5V.n5369 ASIG5V.n5368 0.0380882
R47891 ASIG5V.n5368 ASIG5V.n5367 0.0380882
R47892 ASIG5V.n5367 ASIG5V.n5366 0.0380882
R47893 ASIG5V.n5366 ASIG5V.n5365 0.0380882
R47894 ASIG5V.n5365 ASIG5V.n5364 0.0380882
R47895 ASIG5V.n5364 ASIG5V.n5363 0.0380882
R47896 ASIG5V.n5363 ASIG5V.n5362 0.0380882
R47897 ASIG5V.n5362 ASIG5V.n5361 0.0380882
R47898 ASIG5V.n5361 ASIG5V.n5360 0.0380882
R47899 ASIG5V.n5360 ASIG5V.n5359 0.0380882
R47900 ASIG5V.n5666 ASIG5V.n5665 0.0380882
R47901 ASIG5V.n5665 ASIG5V.n5664 0.0380882
R47902 ASIG5V.n5664 ASIG5V.n5663 0.0380882
R47903 ASIG5V.n5663 ASIG5V.n5662 0.0380882
R47904 ASIG5V.n5662 ASIG5V.n5661 0.0380882
R47905 ASIG5V.n5661 ASIG5V.n5660 0.0380882
R47906 ASIG5V.n5660 ASIG5V.n5659 0.0380882
R47907 ASIG5V.n5659 ASIG5V.n5658 0.0380882
R47908 ASIG5V.n5658 ASIG5V.n5657 0.0380882
R47909 ASIG5V.n5657 ASIG5V.n5656 0.0380882
R47910 ASIG5V.n5656 ASIG5V.n5655 0.0380882
R47911 ASIG5V.n5655 ASIG5V.n5654 0.0380882
R47912 ASIG5V.n5654 ASIG5V.n5653 0.0380882
R47913 ASIG5V.n5653 ASIG5V.n5652 0.0380882
R47914 ASIG5V.n5652 ASIG5V.n5651 0.0380882
R47915 ASIG5V.n5651 ASIG5V.n5650 0.0380882
R47916 ASIG5V.n5650 ASIG5V.n5649 0.0380882
R47917 ASIG5V.n5649 ASIG5V.n5648 0.0380882
R47918 ASIG5V.n5648 ASIG5V.n5647 0.0380882
R47919 ASIG5V.n5647 ASIG5V.n5646 0.0380882
R47920 ASIG5V.n5646 ASIG5V.n5645 0.0380882
R47921 ASIG5V.n5645 ASIG5V.n5644 0.0380882
R47922 ASIG5V.n5644 ASIG5V.n5643 0.0380882
R47923 ASIG5V.n5643 ASIG5V.n5642 0.0380882
R47924 ASIG5V.n5642 ASIG5V.n5641 0.0380882
R47925 ASIG5V.n5641 ASIG5V.n5640 0.0380882
R47926 ASIG5V.n5640 ASIG5V.n5639 0.0380882
R47927 ASIG5V.n5639 ASIG5V.n5638 0.0380882
R47928 ASIG5V.n5638 ASIG5V.n5637 0.0380882
R47929 ASIG5V.n5637 ASIG5V.n5636 0.0380882
R47930 ASIG5V.n5636 ASIG5V.n5635 0.0380882
R47931 ASIG5V.n5635 ASIG5V.n5634 0.0380882
R47932 ASIG5V.n5634 ASIG5V.n5633 0.0380882
R47933 ASIG5V.n5633 ASIG5V.n5632 0.0380882
R47934 ASIG5V.n5632 ASIG5V.n5631 0.0380882
R47935 ASIG5V.n5631 ASIG5V.n5630 0.0380882
R47936 ASIG5V.n5630 ASIG5V.n5629 0.0380882
R47937 ASIG5V.n5629 ASIG5V.n5628 0.0380882
R47938 ASIG5V.n5628 ASIG5V.n5627 0.0380882
R47939 ASIG5V.n5627 ASIG5V.n5626 0.0380882
R47940 ASIG5V.n5626 ASIG5V.n5625 0.0380882
R47941 ASIG5V.n5625 ASIG5V.n5624 0.0380882
R47942 ASIG5V.n5624 ASIG5V.n5623 0.0380882
R47943 ASIG5V.n5623 ASIG5V.n5622 0.0380882
R47944 ASIG5V.n947 ASIG5V.n946 0.0380882
R47945 ASIG5V.n948 ASIG5V.n947 0.0380882
R47946 ASIG5V.n949 ASIG5V.n948 0.0380882
R47947 ASIG5V.n950 ASIG5V.n949 0.0380882
R47948 ASIG5V.n951 ASIG5V.n950 0.0380882
R47949 ASIG5V.n952 ASIG5V.n951 0.0380882
R47950 ASIG5V.n953 ASIG5V.n952 0.0380882
R47951 ASIG5V.n954 ASIG5V.n953 0.0380882
R47952 ASIG5V.n955 ASIG5V.n954 0.0380882
R47953 ASIG5V.n956 ASIG5V.n955 0.0380882
R47954 ASIG5V.n5620 ASIG5V.n5619 0.0380882
R47955 ASIG5V.n5619 ASIG5V.n5618 0.0380882
R47956 ASIG5V.n5618 ASIG5V.n5617 0.0380882
R47957 ASIG5V.n5617 ASIG5V.n5616 0.0380882
R47958 ASIG5V.n5616 ASIG5V.n5615 0.0380882
R47959 ASIG5V.n5615 ASIG5V.n5614 0.0380882
R47960 ASIG5V.n5614 ASIG5V.n5613 0.0380882
R47961 ASIG5V.n5613 ASIG5V.n5612 0.0380882
R47962 ASIG5V.n5612 ASIG5V.n5611 0.0380882
R47963 ASIG5V.n5611 ASIG5V.n5610 0.0380882
R47964 ASIG5V.n5610 ASIG5V.n5609 0.0380882
R47965 ASIG5V.n5609 ASIG5V.n5608 0.0380882
R47966 ASIG5V.n5608 ASIG5V.n5607 0.0380882
R47967 ASIG5V.n5607 ASIG5V.n5606 0.0380882
R47968 ASIG5V.n5606 ASIG5V.n5605 0.0380882
R47969 ASIG5V.n5605 ASIG5V.n5604 0.0380882
R47970 ASIG5V.n5604 ASIG5V.n5603 0.0380882
R47971 ASIG5V.n5603 ASIG5V.n5602 0.0380882
R47972 ASIG5V.n5602 ASIG5V.n5601 0.0380882
R47973 ASIG5V.n5601 ASIG5V.n5600 0.0380882
R47974 ASIG5V.n5600 ASIG5V.n5599 0.0380882
R47975 ASIG5V.n5599 ASIG5V.n5598 0.0380882
R47976 ASIG5V.n5598 ASIG5V.n5597 0.0380882
R47977 ASIG5V.n5597 ASIG5V.n5596 0.0380882
R47978 ASIG5V.n5596 ASIG5V.n5595 0.0380882
R47979 ASIG5V.n5595 ASIG5V.n5594 0.0380882
R47980 ASIG5V.n5594 ASIG5V.n5593 0.0380882
R47981 ASIG5V.n5593 ASIG5V.n5592 0.0380882
R47982 ASIG5V.n5592 ASIG5V.n5591 0.0380882
R47983 ASIG5V.n5591 ASIG5V.n5590 0.0380882
R47984 ASIG5V.n5967 ASIG5V.n5966 0.0380882
R47985 ASIG5V.n5966 ASIG5V.n5965 0.0380882
R47986 ASIG5V.n5965 ASIG5V.n5964 0.0380882
R47987 ASIG5V.n5964 ASIG5V.n5963 0.0380882
R47988 ASIG5V.n5963 ASIG5V.n5962 0.0380882
R47989 ASIG5V.n5962 ASIG5V.n5961 0.0380882
R47990 ASIG5V.n5961 ASIG5V.n5960 0.0380882
R47991 ASIG5V.n5960 ASIG5V.n5959 0.0380882
R47992 ASIG5V.n5959 ASIG5V.n5958 0.0380882
R47993 ASIG5V.n5958 ASIG5V.n5957 0.0380882
R47994 ASIG5V.n5957 ASIG5V.n5956 0.0380882
R47995 ASIG5V.n5956 ASIG5V.n5955 0.0380882
R47996 ASIG5V.n5955 ASIG5V.n5954 0.0380882
R47997 ASIG5V.n5954 ASIG5V.n5953 0.0380882
R47998 ASIG5V.n5953 ASIG5V.n5952 0.0380882
R47999 ASIG5V.n5952 ASIG5V.n5951 0.0380882
R48000 ASIG5V.n5951 ASIG5V.n5950 0.0380882
R48001 ASIG5V.n5950 ASIG5V.n5949 0.0380882
R48002 ASIG5V.n5949 ASIG5V.n5948 0.0380882
R48003 ASIG5V.n5948 ASIG5V.n5947 0.0380882
R48004 ASIG5V.n5947 ASIG5V.n5946 0.0380882
R48005 ASIG5V.n5946 ASIG5V.n5945 0.0380882
R48006 ASIG5V.n5945 ASIG5V.n5944 0.0380882
R48007 ASIG5V.n5944 ASIG5V.n5943 0.0380882
R48008 ASIG5V.n5943 ASIG5V.n5942 0.0380882
R48009 ASIG5V.n5942 ASIG5V.n5941 0.0380882
R48010 ASIG5V.n5941 ASIG5V.n5940 0.0380882
R48011 ASIG5V.n5940 ASIG5V.n5939 0.0380882
R48012 ASIG5V.n5939 ASIG5V.n5938 0.0380882
R48013 ASIG5V.n5938 ASIG5V.n5937 0.0380882
R48014 ASIG5V.n5937 ASIG5V.n5936 0.0380882
R48015 ASIG5V.n5936 ASIG5V.n5935 0.0380882
R48016 ASIG5V.n5935 ASIG5V.n5934 0.0380882
R48017 ASIG5V.n5934 ASIG5V.n5933 0.0380882
R48018 ASIG5V.n5933 ASIG5V.n5932 0.0380882
R48019 ASIG5V.n5932 ASIG5V.n5931 0.0380882
R48020 ASIG5V.n5931 ASIG5V.n5930 0.0380882
R48021 ASIG5V.n5930 ASIG5V.n5929 0.0380882
R48022 ASIG5V.n5929 ASIG5V.n5928 0.0380882
R48023 ASIG5V.n5928 ASIG5V.n5927 0.0380882
R48024 ASIG5V.n5927 ASIG5V.n5926 0.0380882
R48025 ASIG5V.n5926 ASIG5V.n5925 0.0380882
R48026 ASIG5V.n5925 ASIG5V.n5924 0.0380882
R48027 ASIG5V.n5924 ASIG5V.n5923 0.0380882
R48028 ASIG5V.n958 ASIG5V.n957 0.0380882
R48029 ASIG5V.n959 ASIG5V.n958 0.0380882
R48030 ASIG5V.n960 ASIG5V.n959 0.0380882
R48031 ASIG5V.n961 ASIG5V.n960 0.0380882
R48032 ASIG5V.n962 ASIG5V.n961 0.0380882
R48033 ASIG5V.n963 ASIG5V.n962 0.0380882
R48034 ASIG5V.n964 ASIG5V.n963 0.0380882
R48035 ASIG5V.n5921 ASIG5V.n5920 0.0380882
R48036 ASIG5V.n5920 ASIG5V.n5919 0.0380882
R48037 ASIG5V.n5919 ASIG5V.n5918 0.0380882
R48038 ASIG5V.n5918 ASIG5V.n5917 0.0380882
R48039 ASIG5V.n5917 ASIG5V.n5916 0.0380882
R48040 ASIG5V.n5916 ASIG5V.n5915 0.0380882
R48041 ASIG5V.n5915 ASIG5V.n5914 0.0380882
R48042 ASIG5V.n5914 ASIG5V.n5913 0.0380882
R48043 ASIG5V.n5913 ASIG5V.n5912 0.0380882
R48044 ASIG5V.n5912 ASIG5V.n5911 0.0380882
R48045 ASIG5V.n5911 ASIG5V.n5910 0.0380882
R48046 ASIG5V.n5910 ASIG5V.n5909 0.0380882
R48047 ASIG5V.n5909 ASIG5V.n5908 0.0380882
R48048 ASIG5V.n5908 ASIG5V.n5907 0.0380882
R48049 ASIG5V.n5907 ASIG5V.n5906 0.0380882
R48050 ASIG5V.n5906 ASIG5V.n5905 0.0380882
R48051 ASIG5V.n5905 ASIG5V.n5904 0.0380882
R48052 ASIG5V.n5904 ASIG5V.n5903 0.0380882
R48053 ASIG5V.n5903 ASIG5V.n5902 0.0380882
R48054 ASIG5V.n5902 ASIG5V.n5901 0.0380882
R48055 ASIG5V.n5901 ASIG5V.n5900 0.0380882
R48056 ASIG5V.n5900 ASIG5V.n5899 0.0380882
R48057 ASIG5V.n5899 ASIG5V.n5898 0.0380882
R48058 ASIG5V.n5898 ASIG5V.n5897 0.0380882
R48059 ASIG5V.n5897 ASIG5V.n5896 0.0380882
R48060 ASIG5V.n5896 ASIG5V.n5895 0.0380882
R48061 ASIG5V.n5895 ASIG5V.n5894 0.0380882
R48062 ASIG5V.n5894 ASIG5V.n5893 0.0380882
R48063 ASIG5V.n5893 ASIG5V.n5892 0.0380882
R48064 ASIG5V.n5892 ASIG5V.n5891 0.0380882
R48065 ASIG5V.n449 ASIG5V.n448 0.0380882
R48066 ASIG5V.n448 ASIG5V.n447 0.0380882
R48067 ASIG5V.n447 ASIG5V.n446 0.0380882
R48068 ASIG5V.n446 ASIG5V.n445 0.0380882
R48069 ASIG5V.n445 ASIG5V.n444 0.0380882
R48070 ASIG5V.n444 ASIG5V.n443 0.0380882
R48071 ASIG5V.n443 ASIG5V.n442 0.0380882
R48072 ASIG5V.n442 ASIG5V.n441 0.0380882
R48073 ASIG5V.n441 ASIG5V.n440 0.0380882
R48074 ASIG5V.n440 ASIG5V.n439 0.0380882
R48075 ASIG5V.n439 ASIG5V.n438 0.0380882
R48076 ASIG5V.n438 ASIG5V.n437 0.0380882
R48077 ASIG5V.n437 ASIG5V.n436 0.0380882
R48078 ASIG5V.n436 ASIG5V.n435 0.0380882
R48079 ASIG5V.n435 ASIG5V.n434 0.0380882
R48080 ASIG5V.n434 ASIG5V.n433 0.0380882
R48081 ASIG5V.n433 ASIG5V.n432 0.0380882
R48082 ASIG5V.n432 ASIG5V.n431 0.0380882
R48083 ASIG5V.n431 ASIG5V.n430 0.0380882
R48084 ASIG5V.n430 ASIG5V.n429 0.0380882
R48085 ASIG5V.n429 ASIG5V.n428 0.0380882
R48086 ASIG5V.n428 ASIG5V.n427 0.0380882
R48087 ASIG5V.n427 ASIG5V.n426 0.0380882
R48088 ASIG5V.n426 ASIG5V.n425 0.0380882
R48089 ASIG5V.n425 ASIG5V.n424 0.0380882
R48090 ASIG5V.n424 ASIG5V.n423 0.0380882
R48091 ASIG5V.n423 ASIG5V.n422 0.0380882
R48092 ASIG5V.n422 ASIG5V.n421 0.0380882
R48093 ASIG5V.n421 ASIG5V.n420 0.0380882
R48094 ASIG5V.n420 ASIG5V.n419 0.0380882
R48095 ASIG5V.n419 ASIG5V.n418 0.0380882
R48096 ASIG5V.n418 ASIG5V.n417 0.0380882
R48097 ASIG5V.n417 ASIG5V.n416 0.0380882
R48098 ASIG5V.n416 ASIG5V.n415 0.0380882
R48099 ASIG5V.n415 ASIG5V.n414 0.0380882
R48100 ASIG5V.n414 ASIG5V.n413 0.0380882
R48101 ASIG5V.n413 ASIG5V.n412 0.0380882
R48102 ASIG5V.n412 ASIG5V.n411 0.0380882
R48103 ASIG5V.n411 ASIG5V.n410 0.0380882
R48104 ASIG5V.n410 ASIG5V.n409 0.0380882
R48105 ASIG5V.n409 ASIG5V.n408 0.0380882
R48106 ASIG5V.n408 ASIG5V.n407 0.0380882
R48107 ASIG5V.n407 ASIG5V.n406 0.0380882
R48108 ASIG5V.n406 ASIG5V.n405 0.0380882
R48109 ASIG5V.n966 ASIG5V.n965 0.0380882
R48110 ASIG5V.n967 ASIG5V.n966 0.0380882
R48111 ASIG5V.n968 ASIG5V.n967 0.0380882
R48112 ASIG5V.n969 ASIG5V.n968 0.0380882
R48113 ASIG5V.n970 ASIG5V.n969 0.0380882
R48114 ASIG5V.n481 ASIG5V.n480 0.0380882
R48115 ASIG5V.n480 ASIG5V.n479 0.0380882
R48116 ASIG5V.n479 ASIG5V.n478 0.0380882
R48117 ASIG5V.n478 ASIG5V.n477 0.0380882
R48118 ASIG5V.n477 ASIG5V.n476 0.0380882
R48119 ASIG5V.n476 ASIG5V.n475 0.0380882
R48120 ASIG5V.n475 ASIG5V.n474 0.0380882
R48121 ASIG5V.n474 ASIG5V.n473 0.0380882
R48122 ASIG5V.n473 ASIG5V.n472 0.0380882
R48123 ASIG5V.n472 ASIG5V.n471 0.0380882
R48124 ASIG5V.n471 ASIG5V.n470 0.0380882
R48125 ASIG5V.n470 ASIG5V.n469 0.0380882
R48126 ASIG5V.n469 ASIG5V.n468 0.0380882
R48127 ASIG5V.n468 ASIG5V.n467 0.0380882
R48128 ASIG5V.n467 ASIG5V.n466 0.0380882
R48129 ASIG5V.n466 ASIG5V.n465 0.0380882
R48130 ASIG5V.n465 ASIG5V.n464 0.0380882
R48131 ASIG5V.n464 ASIG5V.n463 0.0380882
R48132 ASIG5V.n463 ASIG5V.n462 0.0380882
R48133 ASIG5V.n462 ASIG5V.n461 0.0380882
R48134 ASIG5V.n461 ASIG5V.n460 0.0380882
R48135 ASIG5V.n460 ASIG5V.n459 0.0380882
R48136 ASIG5V.n459 ASIG5V.n458 0.0380882
R48137 ASIG5V.n458 ASIG5V.n457 0.0380882
R48138 ASIG5V.n457 ASIG5V.n456 0.0380882
R48139 ASIG5V.n456 ASIG5V.n455 0.0380882
R48140 ASIG5V.n455 ASIG5V.n454 0.0380882
R48141 ASIG5V.n454 ASIG5V.n453 0.0380882
R48142 ASIG5V.n453 ASIG5V.n452 0.0380882
R48143 ASIG5V.n452 ASIG5V.n451 0.0380882
R48144 ASIG5V.n7043 ASIG5V.n7042 0.0380882
R48145 ASIG5V.n7042 ASIG5V.n7041 0.0380882
R48146 ASIG5V.n7041 ASIG5V.n7040 0.0380882
R48147 ASIG5V.n7040 ASIG5V.n7039 0.0380882
R48148 ASIG5V.n7039 ASIG5V.n7038 0.0380882
R48149 ASIG5V.n7038 ASIG5V.n7037 0.0380882
R48150 ASIG5V.n7037 ASIG5V.n7036 0.0380882
R48151 ASIG5V.n7036 ASIG5V.n7035 0.0380882
R48152 ASIG5V.n7035 ASIG5V.n7034 0.0380882
R48153 ASIG5V.n7034 ASIG5V.n7033 0.0380882
R48154 ASIG5V.n7033 ASIG5V.n7032 0.0380882
R48155 ASIG5V.n7032 ASIG5V.n7031 0.0380882
R48156 ASIG5V.n7031 ASIG5V.n7030 0.0380882
R48157 ASIG5V.n7030 ASIG5V.n7029 0.0380882
R48158 ASIG5V.n7029 ASIG5V.n7028 0.0380882
R48159 ASIG5V.n7028 ASIG5V.n7027 0.0380882
R48160 ASIG5V.n7027 ASIG5V.n7026 0.0380882
R48161 ASIG5V.n7026 ASIG5V.n7025 0.0380882
R48162 ASIG5V.n7025 ASIG5V.n7024 0.0380882
R48163 ASIG5V.n7024 ASIG5V.n7023 0.0380882
R48164 ASIG5V.n7023 ASIG5V.n7022 0.0380882
R48165 ASIG5V.n7022 ASIG5V.n7021 0.0380882
R48166 ASIG5V.n7021 ASIG5V.n7020 0.0380882
R48167 ASIG5V.n7020 ASIG5V.n7019 0.0380882
R48168 ASIG5V.n7019 ASIG5V.n7018 0.0380882
R48169 ASIG5V.n7018 ASIG5V.n7017 0.0380882
R48170 ASIG5V.n7017 ASIG5V.n7016 0.0380882
R48171 ASIG5V.n7016 ASIG5V.n7015 0.0380882
R48172 ASIG5V.n7015 ASIG5V.n7014 0.0380882
R48173 ASIG5V.n7014 ASIG5V.n7013 0.0380882
R48174 ASIG5V.n7013 ASIG5V.n7012 0.0380882
R48175 ASIG5V.n7012 ASIG5V.n7011 0.0380882
R48176 ASIG5V.n7011 ASIG5V.n7010 0.0380882
R48177 ASIG5V.n7010 ASIG5V.n7009 0.0380882
R48178 ASIG5V.n7009 ASIG5V.n7008 0.0380882
R48179 ASIG5V.n7008 ASIG5V.n7007 0.0380882
R48180 ASIG5V.n7007 ASIG5V.n7006 0.0380882
R48181 ASIG5V.n7006 ASIG5V.n7005 0.0380882
R48182 ASIG5V.n7005 ASIG5V.n7004 0.0380882
R48183 ASIG5V.n7004 ASIG5V.n7003 0.0380882
R48184 ASIG5V.n7003 ASIG5V.n7002 0.0380882
R48185 ASIG5V.n7002 ASIG5V.n7001 0.0380882
R48186 ASIG5V.n7001 ASIG5V.n7000 0.0380882
R48187 ASIG5V.n7000 ASIG5V.n6999 0.0380882
R48188 ASIG5V.n6999 ASIG5V.n6998 0.0380882
R48189 ASIG5V.n972 ASIG5V.n971 0.0380882
R48190 ASIG5V.n973 ASIG5V.n972 0.0380882
R48191 ASIG5V.n6996 ASIG5V.n6995 0.0380882
R48192 ASIG5V.n6995 ASIG5V.n6994 0.0380882
R48193 ASIG5V.n6994 ASIG5V.n6993 0.0380882
R48194 ASIG5V.n6993 ASIG5V.n6992 0.0380882
R48195 ASIG5V.n6992 ASIG5V.n6991 0.0380882
R48196 ASIG5V.n6991 ASIG5V.n6990 0.0380882
R48197 ASIG5V.n6990 ASIG5V.n6989 0.0380882
R48198 ASIG5V.n6989 ASIG5V.n6988 0.0380882
R48199 ASIG5V.n6988 ASIG5V.n6987 0.0380882
R48200 ASIG5V.n6987 ASIG5V.n6986 0.0380882
R48201 ASIG5V.n6986 ASIG5V.n6985 0.0380882
R48202 ASIG5V.n6985 ASIG5V.n6984 0.0380882
R48203 ASIG5V.n6984 ASIG5V.n6983 0.0380882
R48204 ASIG5V.n6983 ASIG5V.n6982 0.0380882
R48205 ASIG5V.n6982 ASIG5V.n6981 0.0380882
R48206 ASIG5V.n6981 ASIG5V.n6980 0.0380882
R48207 ASIG5V.n6980 ASIG5V.n6979 0.0380882
R48208 ASIG5V.n6979 ASIG5V.n6978 0.0380882
R48209 ASIG5V.n6978 ASIG5V.n6977 0.0380882
R48210 ASIG5V.n6977 ASIG5V.n6976 0.0380882
R48211 ASIG5V.n6976 ASIG5V.n6975 0.0380882
R48212 ASIG5V.n6975 ASIG5V.n6974 0.0380882
R48213 ASIG5V.n6974 ASIG5V.n6973 0.0380882
R48214 ASIG5V.n6973 ASIG5V.n6972 0.0380882
R48215 ASIG5V.n6972 ASIG5V.n6971 0.0380882
R48216 ASIG5V.n6971 ASIG5V.n6970 0.0380882
R48217 ASIG5V.n6970 ASIG5V.n6969 0.0380882
R48218 ASIG5V.n6969 ASIG5V.n6968 0.0380882
R48219 ASIG5V.n6968 ASIG5V.n6967 0.0380882
R48220 ASIG5V.n6967 ASIG5V.n6966 0.0380882
R48221 ASIG5V.n6764 ASIG5V.n6763 0.0380882
R48222 ASIG5V.n6763 ASIG5V.n6762 0.0380882
R48223 ASIG5V.n6762 ASIG5V.n6761 0.0380882
R48224 ASIG5V.n6761 ASIG5V.n6760 0.0380882
R48225 ASIG5V.n6760 ASIG5V.n6759 0.0380882
R48226 ASIG5V.n6759 ASIG5V.n6758 0.0380882
R48227 ASIG5V.n6758 ASIG5V.n6757 0.0380882
R48228 ASIG5V.n6757 ASIG5V.n6756 0.0380882
R48229 ASIG5V.n6756 ASIG5V.n6755 0.0380882
R48230 ASIG5V.n6755 ASIG5V.n6754 0.0380882
R48231 ASIG5V.n6754 ASIG5V.n6753 0.0380882
R48232 ASIG5V.n6753 ASIG5V.n6752 0.0380882
R48233 ASIG5V.n6752 ASIG5V.n6751 0.0380882
R48234 ASIG5V.n6751 ASIG5V.n6750 0.0380882
R48235 ASIG5V.n6750 ASIG5V.n6749 0.0380882
R48236 ASIG5V.n6749 ASIG5V.n6748 0.0380882
R48237 ASIG5V.n6748 ASIG5V.n6747 0.0380882
R48238 ASIG5V.n6747 ASIG5V.n6746 0.0380882
R48239 ASIG5V.n6746 ASIG5V.n6745 0.0380882
R48240 ASIG5V.n6745 ASIG5V.n6744 0.0380882
R48241 ASIG5V.n6744 ASIG5V.n6743 0.0380882
R48242 ASIG5V.n6743 ASIG5V.n6742 0.0380882
R48243 ASIG5V.n6742 ASIG5V.n6741 0.0380882
R48244 ASIG5V.n6741 ASIG5V.n6740 0.0380882
R48245 ASIG5V.n6740 ASIG5V.n6739 0.0380882
R48246 ASIG5V.n6739 ASIG5V.n6738 0.0380882
R48247 ASIG5V.n6738 ASIG5V.n6737 0.0380882
R48248 ASIG5V.n6737 ASIG5V.n6736 0.0380882
R48249 ASIG5V.n6736 ASIG5V.n6735 0.0380882
R48250 ASIG5V.n6735 ASIG5V.n6734 0.0380882
R48251 ASIG5V.n6734 ASIG5V.n6733 0.0380882
R48252 ASIG5V.n6733 ASIG5V.n6732 0.0380882
R48253 ASIG5V.n6732 ASIG5V.n6731 0.0380882
R48254 ASIG5V.n6731 ASIG5V.n6730 0.0380882
R48255 ASIG5V.n6730 ASIG5V.n6729 0.0380882
R48256 ASIG5V.n6729 ASIG5V.n6728 0.0380882
R48257 ASIG5V.n6728 ASIG5V.n6727 0.0380882
R48258 ASIG5V.n6727 ASIG5V.n6726 0.0380882
R48259 ASIG5V.n6726 ASIG5V.n6725 0.0380882
R48260 ASIG5V.n6725 ASIG5V.n6724 0.0380882
R48261 ASIG5V.n6724 ASIG5V.n6723 0.0380882
R48262 ASIG5V.n6723 ASIG5V.n6722 0.0380882
R48263 ASIG5V.n6722 ASIG5V.n6721 0.0380882
R48264 ASIG5V.n6721 ASIG5V.n6720 0.0380882
R48265 ASIG5V.n6718 ASIG5V.n6717 0.0380882
R48266 ASIG5V.n6717 ASIG5V.n6716 0.0380882
R48267 ASIG5V.n6716 ASIG5V.n6715 0.0380882
R48268 ASIG5V.n6715 ASIG5V.n6714 0.0380882
R48269 ASIG5V.n6714 ASIG5V.n6713 0.0380882
R48270 ASIG5V.n6713 ASIG5V.n6712 0.0380882
R48271 ASIG5V.n6712 ASIG5V.n6711 0.0380882
R48272 ASIG5V.n6711 ASIG5V.n6710 0.0380882
R48273 ASIG5V.n6710 ASIG5V.n6709 0.0380882
R48274 ASIG5V.n6709 ASIG5V.n6708 0.0380882
R48275 ASIG5V.n6708 ASIG5V.n6707 0.0380882
R48276 ASIG5V.n6707 ASIG5V.n6706 0.0380882
R48277 ASIG5V.n6706 ASIG5V.n6705 0.0380882
R48278 ASIG5V.n6705 ASIG5V.n6704 0.0380882
R48279 ASIG5V.n6704 ASIG5V.n6703 0.0380882
R48280 ASIG5V.n6703 ASIG5V.n6702 0.0380882
R48281 ASIG5V.n6702 ASIG5V.n6701 0.0380882
R48282 ASIG5V.n6701 ASIG5V.n6700 0.0380882
R48283 ASIG5V.n6700 ASIG5V.n6699 0.0380882
R48284 ASIG5V.n6699 ASIG5V.n6698 0.0380882
R48285 ASIG5V.n6698 ASIG5V.n6697 0.0380882
R48286 ASIG5V.n6697 ASIG5V.n6696 0.0380882
R48287 ASIG5V.n6696 ASIG5V.n6695 0.0380882
R48288 ASIG5V.n6695 ASIG5V.n6694 0.0380882
R48289 ASIG5V.n6694 ASIG5V.n6693 0.0380882
R48290 ASIG5V.n6693 ASIG5V.n6692 0.0380882
R48291 ASIG5V.n6692 ASIG5V.n6691 0.0380882
R48292 ASIG5V.n6691 ASIG5V.n6690 0.0380882
R48293 ASIG5V.n6690 ASIG5V.n6689 0.0380882
R48294 ASIG5V.n6689 ASIG5V.n6688 0.0380882
R48295 ASIG5V.n13602 ASIG5V.n13601 0.0380882
R48296 ASIG5V.n13601 ASIG5V.n13600 0.0380882
R48297 ASIG5V.n13600 ASIG5V.n13599 0.0380882
R48298 ASIG5V.n13599 ASIG5V.n13598 0.0380882
R48299 ASIG5V.n13598 ASIG5V.n13597 0.0380882
R48300 ASIG5V.n13597 ASIG5V.n13596 0.0380882
R48301 ASIG5V.n13596 ASIG5V.n13595 0.0380882
R48302 ASIG5V.n13595 ASIG5V.n13594 0.0380882
R48303 ASIG5V.n13594 ASIG5V.n13593 0.0380882
R48304 ASIG5V.n13593 ASIG5V.n13592 0.0380882
R48305 ASIG5V.n13592 ASIG5V.n13591 0.0380882
R48306 ASIG5V.n13591 ASIG5V.n13590 0.0380882
R48307 ASIG5V.n13590 ASIG5V.n13589 0.0380882
R48308 ASIG5V.n13589 ASIG5V.n13588 0.0380882
R48309 ASIG5V.n13588 ASIG5V.n13587 0.0380882
R48310 ASIG5V.n13587 ASIG5V.n13586 0.0380882
R48311 ASIG5V.n13586 ASIG5V.n13585 0.0380882
R48312 ASIG5V.n13585 ASIG5V.n13584 0.0380882
R48313 ASIG5V.n13584 ASIG5V.n13583 0.0380882
R48314 ASIG5V.n13583 ASIG5V.n13582 0.0380882
R48315 ASIG5V.n13582 ASIG5V.n13581 0.0380882
R48316 ASIG5V.n13581 ASIG5V.n13580 0.0380882
R48317 ASIG5V.n13580 ASIG5V.n13579 0.0380882
R48318 ASIG5V.n13579 ASIG5V.n13578 0.0380882
R48319 ASIG5V.n13578 ASIG5V.n13577 0.0380882
R48320 ASIG5V.n13577 ASIG5V.n13576 0.0380882
R48321 ASIG5V.n13576 ASIG5V.n13575 0.0380882
R48322 ASIG5V.n13575 ASIG5V.n13574 0.0380882
R48323 ASIG5V.n13574 ASIG5V.n13573 0.0380882
R48324 ASIG5V.n13573 ASIG5V.n13572 0.0380882
R48325 ASIG5V.n13572 ASIG5V.n13571 0.0380882
R48326 ASIG5V.n13571 ASIG5V.n13570 0.0380882
R48327 ASIG5V.n13570 ASIG5V.n13569 0.0380882
R48328 ASIG5V.n13569 ASIG5V.n13568 0.0380882
R48329 ASIG5V.n13568 ASIG5V.n13567 0.0380882
R48330 ASIG5V.n13567 ASIG5V.n13566 0.0380882
R48331 ASIG5V.n13566 ASIG5V.n13565 0.0380882
R48332 ASIG5V.n13565 ASIG5V.n13564 0.0380882
R48333 ASIG5V.n13564 ASIG5V.n13563 0.0380882
R48334 ASIG5V.n13563 ASIG5V.n13562 0.0380882
R48335 ASIG5V.n13562 ASIG5V.n13561 0.0380882
R48336 ASIG5V.n13561 ASIG5V.n13560 0.0380882
R48337 ASIG5V.n13560 ASIG5V.n13559 0.0380882
R48338 ASIG5V.n13559 ASIG5V.n13558 0.0380882
R48339 ASIG5V.n9370 ASIG5V.n9369 0.0380882
R48340 ASIG5V.n9371 ASIG5V.n9370 0.0380882
R48341 ASIG5V.n13556 ASIG5V.n13555 0.0380882
R48342 ASIG5V.n13555 ASIG5V.n13554 0.0380882
R48343 ASIG5V.n13554 ASIG5V.n13553 0.0380882
R48344 ASIG5V.n13553 ASIG5V.n13552 0.0380882
R48345 ASIG5V.n13552 ASIG5V.n13551 0.0380882
R48346 ASIG5V.n13551 ASIG5V.n13550 0.0380882
R48347 ASIG5V.n13550 ASIG5V.n13549 0.0380882
R48348 ASIG5V.n13549 ASIG5V.n13548 0.0380882
R48349 ASIG5V.n13548 ASIG5V.n13547 0.0380882
R48350 ASIG5V.n13547 ASIG5V.n13546 0.0380882
R48351 ASIG5V.n13546 ASIG5V.n13545 0.0380882
R48352 ASIG5V.n13545 ASIG5V.n13544 0.0380882
R48353 ASIG5V.n13544 ASIG5V.n13543 0.0380882
R48354 ASIG5V.n13543 ASIG5V.n13542 0.0380882
R48355 ASIG5V.n13542 ASIG5V.n13541 0.0380882
R48356 ASIG5V.n13541 ASIG5V.n13540 0.0380882
R48357 ASIG5V.n13540 ASIG5V.n13539 0.0380882
R48358 ASIG5V.n13539 ASIG5V.n13538 0.0380882
R48359 ASIG5V.n13538 ASIG5V.n13537 0.0380882
R48360 ASIG5V.n13537 ASIG5V.n13536 0.0380882
R48361 ASIG5V.n13536 ASIG5V.n13535 0.0380882
R48362 ASIG5V.n13535 ASIG5V.n13534 0.0380882
R48363 ASIG5V.n13534 ASIG5V.n13533 0.0380882
R48364 ASIG5V.n13533 ASIG5V.n13532 0.0380882
R48365 ASIG5V.n13532 ASIG5V.n13531 0.0380882
R48366 ASIG5V.n13531 ASIG5V.n13530 0.0380882
R48367 ASIG5V.n13530 ASIG5V.n13529 0.0380882
R48368 ASIG5V.n13529 ASIG5V.n13528 0.0380882
R48369 ASIG5V.n13528 ASIG5V.n13527 0.0380882
R48370 ASIG5V.n13527 ASIG5V.n13526 0.0380882
R48371 ASIG5V.n13347 ASIG5V.n13346 0.0380882
R48372 ASIG5V.n13346 ASIG5V.n13345 0.0380882
R48373 ASIG5V.n13345 ASIG5V.n13344 0.0380882
R48374 ASIG5V.n13344 ASIG5V.n13343 0.0380882
R48375 ASIG5V.n13343 ASIG5V.n13342 0.0380882
R48376 ASIG5V.n13342 ASIG5V.n13341 0.0380882
R48377 ASIG5V.n13341 ASIG5V.n13340 0.0380882
R48378 ASIG5V.n13340 ASIG5V.n13339 0.0380882
R48379 ASIG5V.n13339 ASIG5V.n13338 0.0380882
R48380 ASIG5V.n13338 ASIG5V.n13337 0.0380882
R48381 ASIG5V.n13337 ASIG5V.n13336 0.0380882
R48382 ASIG5V.n13336 ASIG5V.n13335 0.0380882
R48383 ASIG5V.n13335 ASIG5V.n13334 0.0380882
R48384 ASIG5V.n13334 ASIG5V.n13333 0.0380882
R48385 ASIG5V.n13333 ASIG5V.n13332 0.0380882
R48386 ASIG5V.n13332 ASIG5V.n13331 0.0380882
R48387 ASIG5V.n13331 ASIG5V.n13330 0.0380882
R48388 ASIG5V.n13330 ASIG5V.n13329 0.0380882
R48389 ASIG5V.n13329 ASIG5V.n13328 0.0380882
R48390 ASIG5V.n13328 ASIG5V.n13327 0.0380882
R48391 ASIG5V.n13327 ASIG5V.n13326 0.0380882
R48392 ASIG5V.n13326 ASIG5V.n13325 0.0380882
R48393 ASIG5V.n13325 ASIG5V.n13324 0.0380882
R48394 ASIG5V.n13324 ASIG5V.n13323 0.0380882
R48395 ASIG5V.n13323 ASIG5V.n13322 0.0380882
R48396 ASIG5V.n13322 ASIG5V.n13321 0.0380882
R48397 ASIG5V.n13321 ASIG5V.n13320 0.0380882
R48398 ASIG5V.n13320 ASIG5V.n13319 0.0380882
R48399 ASIG5V.n13319 ASIG5V.n13318 0.0380882
R48400 ASIG5V.n13318 ASIG5V.n13317 0.0380882
R48401 ASIG5V.n13317 ASIG5V.n13316 0.0380882
R48402 ASIG5V.n13316 ASIG5V.n13315 0.0380882
R48403 ASIG5V.n13315 ASIG5V.n13314 0.0380882
R48404 ASIG5V.n13314 ASIG5V.n13313 0.0380882
R48405 ASIG5V.n13313 ASIG5V.n13312 0.0380882
R48406 ASIG5V.n13312 ASIG5V.n13311 0.0380882
R48407 ASIG5V.n13311 ASIG5V.n13310 0.0380882
R48408 ASIG5V.n13310 ASIG5V.n13309 0.0380882
R48409 ASIG5V.n13309 ASIG5V.n13308 0.0380882
R48410 ASIG5V.n13308 ASIG5V.n13307 0.0380882
R48411 ASIG5V.n13307 ASIG5V.n13306 0.0380882
R48412 ASIG5V.n13306 ASIG5V.n13305 0.0380882
R48413 ASIG5V.n13305 ASIG5V.n13304 0.0380882
R48414 ASIG5V.n13304 ASIG5V.n13303 0.0380882
R48415 ASIG5V.n9365 ASIG5V.n9364 0.0380882
R48416 ASIG5V.n9366 ASIG5V.n9365 0.0380882
R48417 ASIG5V.n9367 ASIG5V.n9366 0.0380882
R48418 ASIG5V.n9368 ASIG5V.n9367 0.0380882
R48419 ASIG5V.n392 ASIG5V.n391 0.0380882
R48420 ASIG5V.n391 ASIG5V.n390 0.0380882
R48421 ASIG5V.n390 ASIG5V.n389 0.0380882
R48422 ASIG5V.n389 ASIG5V.n388 0.0380882
R48423 ASIG5V.n388 ASIG5V.n387 0.0380882
R48424 ASIG5V.n387 ASIG5V.n386 0.0380882
R48425 ASIG5V.n386 ASIG5V.n385 0.0380882
R48426 ASIG5V.n385 ASIG5V.n384 0.0380882
R48427 ASIG5V.n384 ASIG5V.n383 0.0380882
R48428 ASIG5V.n383 ASIG5V.n382 0.0380882
R48429 ASIG5V.n382 ASIG5V.n381 0.0380882
R48430 ASIG5V.n381 ASIG5V.n380 0.0380882
R48431 ASIG5V.n380 ASIG5V.n379 0.0380882
R48432 ASIG5V.n379 ASIG5V.n378 0.0380882
R48433 ASIG5V.n378 ASIG5V.n377 0.0380882
R48434 ASIG5V.n377 ASIG5V.n376 0.0380882
R48435 ASIG5V.n376 ASIG5V.n375 0.0380882
R48436 ASIG5V.n375 ASIG5V.n374 0.0380882
R48437 ASIG5V.n374 ASIG5V.n373 0.0380882
R48438 ASIG5V.n373 ASIG5V.n372 0.0380882
R48439 ASIG5V.n372 ASIG5V.n371 0.0380882
R48440 ASIG5V.n371 ASIG5V.n370 0.0380882
R48441 ASIG5V.n370 ASIG5V.n369 0.0380882
R48442 ASIG5V.n369 ASIG5V.n368 0.0380882
R48443 ASIG5V.n368 ASIG5V.n367 0.0380882
R48444 ASIG5V.n367 ASIG5V.n366 0.0380882
R48445 ASIG5V.n366 ASIG5V.n365 0.0380882
R48446 ASIG5V.n365 ASIG5V.n364 0.0380882
R48447 ASIG5V.n364 ASIG5V.n363 0.0380882
R48448 ASIG5V.n363 ASIG5V.n362 0.0380882
R48449 ASIG5V.n7514 ASIG5V.n7513 0.0380882
R48450 ASIG5V.n7513 ASIG5V.n7512 0.0380882
R48451 ASIG5V.n7512 ASIG5V.n7511 0.0380882
R48452 ASIG5V.n7511 ASIG5V.n7510 0.0380882
R48453 ASIG5V.n7510 ASIG5V.n7509 0.0380882
R48454 ASIG5V.n7509 ASIG5V.n7508 0.0380882
R48455 ASIG5V.n7508 ASIG5V.n7507 0.0380882
R48456 ASIG5V.n7507 ASIG5V.n7506 0.0380882
R48457 ASIG5V.n7506 ASIG5V.n7505 0.0380882
R48458 ASIG5V.n7505 ASIG5V.n7504 0.0380882
R48459 ASIG5V.n7504 ASIG5V.n7503 0.0380882
R48460 ASIG5V.n7503 ASIG5V.n7502 0.0380882
R48461 ASIG5V.n7502 ASIG5V.n7501 0.0380882
R48462 ASIG5V.n7501 ASIG5V.n7500 0.0380882
R48463 ASIG5V.n7500 ASIG5V.n7499 0.0380882
R48464 ASIG5V.n7499 ASIG5V.n7498 0.0380882
R48465 ASIG5V.n7498 ASIG5V.n7497 0.0380882
R48466 ASIG5V.n7497 ASIG5V.n7496 0.0380882
R48467 ASIG5V.n7496 ASIG5V.n7495 0.0380882
R48468 ASIG5V.n7495 ASIG5V.n7494 0.0380882
R48469 ASIG5V.n7494 ASIG5V.n7493 0.0380882
R48470 ASIG5V.n7493 ASIG5V.n7492 0.0380882
R48471 ASIG5V.n7492 ASIG5V.n7491 0.0380882
R48472 ASIG5V.n7491 ASIG5V.n7490 0.0380882
R48473 ASIG5V.n7490 ASIG5V.n7489 0.0380882
R48474 ASIG5V.n7489 ASIG5V.n7488 0.0380882
R48475 ASIG5V.n7488 ASIG5V.n7487 0.0380882
R48476 ASIG5V.n7487 ASIG5V.n7486 0.0380882
R48477 ASIG5V.n7486 ASIG5V.n7485 0.0380882
R48478 ASIG5V.n7485 ASIG5V.n7484 0.0380882
R48479 ASIG5V.n7484 ASIG5V.n7483 0.0380882
R48480 ASIG5V.n7483 ASIG5V.n7482 0.0380882
R48481 ASIG5V.n7482 ASIG5V.n7481 0.0380882
R48482 ASIG5V.n7481 ASIG5V.n7480 0.0380882
R48483 ASIG5V.n7480 ASIG5V.n7479 0.0380882
R48484 ASIG5V.n7479 ASIG5V.n7478 0.0380882
R48485 ASIG5V.n7478 ASIG5V.n7477 0.0380882
R48486 ASIG5V.n7477 ASIG5V.n7476 0.0380882
R48487 ASIG5V.n7476 ASIG5V.n7475 0.0380882
R48488 ASIG5V.n7475 ASIG5V.n7474 0.0380882
R48489 ASIG5V.n7474 ASIG5V.n7473 0.0380882
R48490 ASIG5V.n7473 ASIG5V.n7472 0.0380882
R48491 ASIG5V.n7472 ASIG5V.n7471 0.0380882
R48492 ASIG5V.n7471 ASIG5V.n7470 0.0380882
R48493 ASIG5V.n7470 ASIG5V.n7469 0.0380882
R48494 ASIG5V.n9357 ASIG5V.n9356 0.0380882
R48495 ASIG5V.n9358 ASIG5V.n9357 0.0380882
R48496 ASIG5V.n9359 ASIG5V.n9358 0.0380882
R48497 ASIG5V.n9360 ASIG5V.n9359 0.0380882
R48498 ASIG5V.n9361 ASIG5V.n9360 0.0380882
R48499 ASIG5V.n9362 ASIG5V.n9361 0.0380882
R48500 ASIG5V.n9363 ASIG5V.n9362 0.0380882
R48501 ASIG5V.n7467 ASIG5V.n7466 0.0380882
R48502 ASIG5V.n7466 ASIG5V.n7465 0.0380882
R48503 ASIG5V.n7465 ASIG5V.n7464 0.0380882
R48504 ASIG5V.n7464 ASIG5V.n7463 0.0380882
R48505 ASIG5V.n7463 ASIG5V.n7462 0.0380882
R48506 ASIG5V.n7462 ASIG5V.n7461 0.0380882
R48507 ASIG5V.n7461 ASIG5V.n7460 0.0380882
R48508 ASIG5V.n7460 ASIG5V.n7459 0.0380882
R48509 ASIG5V.n7459 ASIG5V.n7458 0.0380882
R48510 ASIG5V.n7458 ASIG5V.n7457 0.0380882
R48511 ASIG5V.n7457 ASIG5V.n7456 0.0380882
R48512 ASIG5V.n7456 ASIG5V.n7455 0.0380882
R48513 ASIG5V.n7455 ASIG5V.n7454 0.0380882
R48514 ASIG5V.n7454 ASIG5V.n7453 0.0380882
R48515 ASIG5V.n7453 ASIG5V.n7452 0.0380882
R48516 ASIG5V.n7452 ASIG5V.n7451 0.0380882
R48517 ASIG5V.n7451 ASIG5V.n7450 0.0380882
R48518 ASIG5V.n7450 ASIG5V.n7449 0.0380882
R48519 ASIG5V.n7449 ASIG5V.n7448 0.0380882
R48520 ASIG5V.n7448 ASIG5V.n7447 0.0380882
R48521 ASIG5V.n7447 ASIG5V.n7446 0.0380882
R48522 ASIG5V.n7446 ASIG5V.n7445 0.0380882
R48523 ASIG5V.n7445 ASIG5V.n7444 0.0380882
R48524 ASIG5V.n7444 ASIG5V.n7443 0.0380882
R48525 ASIG5V.n7443 ASIG5V.n7442 0.0380882
R48526 ASIG5V.n7442 ASIG5V.n7441 0.0380882
R48527 ASIG5V.n7441 ASIG5V.n7440 0.0380882
R48528 ASIG5V.n7440 ASIG5V.n7439 0.0380882
R48529 ASIG5V.n7439 ASIG5V.n7438 0.0380882
R48530 ASIG5V.n7438 ASIG5V.n7437 0.0380882
R48531 ASIG5V.n7931 ASIG5V.n7930 0.0380882
R48532 ASIG5V.n7930 ASIG5V.n7929 0.0380882
R48533 ASIG5V.n7929 ASIG5V.n7928 0.0380882
R48534 ASIG5V.n7928 ASIG5V.n7927 0.0380882
R48535 ASIG5V.n7927 ASIG5V.n7926 0.0380882
R48536 ASIG5V.n7926 ASIG5V.n7925 0.0380882
R48537 ASIG5V.n7925 ASIG5V.n7924 0.0380882
R48538 ASIG5V.n7924 ASIG5V.n7923 0.0380882
R48539 ASIG5V.n7923 ASIG5V.n7922 0.0380882
R48540 ASIG5V.n7922 ASIG5V.n7921 0.0380882
R48541 ASIG5V.n7921 ASIG5V.n7920 0.0380882
R48542 ASIG5V.n7920 ASIG5V.n7919 0.0380882
R48543 ASIG5V.n7919 ASIG5V.n7918 0.0380882
R48544 ASIG5V.n7918 ASIG5V.n7917 0.0380882
R48545 ASIG5V.n7917 ASIG5V.n7916 0.0380882
R48546 ASIG5V.n7916 ASIG5V.n7915 0.0380882
R48547 ASIG5V.n7915 ASIG5V.n7914 0.0380882
R48548 ASIG5V.n7914 ASIG5V.n7913 0.0380882
R48549 ASIG5V.n7913 ASIG5V.n7912 0.0380882
R48550 ASIG5V.n7912 ASIG5V.n7911 0.0380882
R48551 ASIG5V.n7911 ASIG5V.n7910 0.0380882
R48552 ASIG5V.n7910 ASIG5V.n7909 0.0380882
R48553 ASIG5V.n7909 ASIG5V.n7908 0.0380882
R48554 ASIG5V.n7908 ASIG5V.n7907 0.0380882
R48555 ASIG5V.n7907 ASIG5V.n7906 0.0380882
R48556 ASIG5V.n7906 ASIG5V.n7905 0.0380882
R48557 ASIG5V.n7905 ASIG5V.n7904 0.0380882
R48558 ASIG5V.n7904 ASIG5V.n7903 0.0380882
R48559 ASIG5V.n7903 ASIG5V.n7902 0.0380882
R48560 ASIG5V.n7902 ASIG5V.n7901 0.0380882
R48561 ASIG5V.n7901 ASIG5V.n7900 0.0380882
R48562 ASIG5V.n7900 ASIG5V.n7899 0.0380882
R48563 ASIG5V.n7899 ASIG5V.n7898 0.0380882
R48564 ASIG5V.n7898 ASIG5V.n7897 0.0380882
R48565 ASIG5V.n7897 ASIG5V.n7896 0.0380882
R48566 ASIG5V.n7896 ASIG5V.n7895 0.0380882
R48567 ASIG5V.n7895 ASIG5V.n7894 0.0380882
R48568 ASIG5V.n7894 ASIG5V.n7893 0.0380882
R48569 ASIG5V.n7893 ASIG5V.n7892 0.0380882
R48570 ASIG5V.n7892 ASIG5V.n7891 0.0380882
R48571 ASIG5V.n7891 ASIG5V.n7890 0.0380882
R48572 ASIG5V.n7890 ASIG5V.n7889 0.0380882
R48573 ASIG5V.n7889 ASIG5V.n7888 0.0380882
R48574 ASIG5V.n7888 ASIG5V.n7887 0.0380882
R48575 ASIG5V.n7887 ASIG5V.n7886 0.0380882
R48576 ASIG5V.n9347 ASIG5V.n9346 0.0380882
R48577 ASIG5V.n9348 ASIG5V.n9347 0.0380882
R48578 ASIG5V.n9349 ASIG5V.n9348 0.0380882
R48579 ASIG5V.n9350 ASIG5V.n9349 0.0380882
R48580 ASIG5V.n9351 ASIG5V.n9350 0.0380882
R48581 ASIG5V.n9352 ASIG5V.n9351 0.0380882
R48582 ASIG5V.n9353 ASIG5V.n9352 0.0380882
R48583 ASIG5V.n9354 ASIG5V.n9353 0.0380882
R48584 ASIG5V.n9355 ASIG5V.n9354 0.0380882
R48585 ASIG5V.n7884 ASIG5V.n7883 0.0380882
R48586 ASIG5V.n7883 ASIG5V.n7882 0.0380882
R48587 ASIG5V.n7882 ASIG5V.n7881 0.0380882
R48588 ASIG5V.n7881 ASIG5V.n7880 0.0380882
R48589 ASIG5V.n7880 ASIG5V.n7879 0.0380882
R48590 ASIG5V.n7879 ASIG5V.n7878 0.0380882
R48591 ASIG5V.n7878 ASIG5V.n7877 0.0380882
R48592 ASIG5V.n7877 ASIG5V.n7876 0.0380882
R48593 ASIG5V.n7876 ASIG5V.n7875 0.0380882
R48594 ASIG5V.n7875 ASIG5V.n7874 0.0380882
R48595 ASIG5V.n7874 ASIG5V.n7873 0.0380882
R48596 ASIG5V.n7873 ASIG5V.n7872 0.0380882
R48597 ASIG5V.n7872 ASIG5V.n7871 0.0380882
R48598 ASIG5V.n7871 ASIG5V.n7870 0.0380882
R48599 ASIG5V.n7870 ASIG5V.n7869 0.0380882
R48600 ASIG5V.n7869 ASIG5V.n7868 0.0380882
R48601 ASIG5V.n7868 ASIG5V.n7867 0.0380882
R48602 ASIG5V.n7867 ASIG5V.n7866 0.0380882
R48603 ASIG5V.n7866 ASIG5V.n7865 0.0380882
R48604 ASIG5V.n7865 ASIG5V.n7864 0.0380882
R48605 ASIG5V.n7864 ASIG5V.n7863 0.0380882
R48606 ASIG5V.n7863 ASIG5V.n7862 0.0380882
R48607 ASIG5V.n7862 ASIG5V.n7861 0.0380882
R48608 ASIG5V.n7861 ASIG5V.n7860 0.0380882
R48609 ASIG5V.n7860 ASIG5V.n7859 0.0380882
R48610 ASIG5V.n7859 ASIG5V.n7858 0.0380882
R48611 ASIG5V.n7858 ASIG5V.n7857 0.0380882
R48612 ASIG5V.n7857 ASIG5V.n7856 0.0380882
R48613 ASIG5V.n7856 ASIG5V.n7855 0.0380882
R48614 ASIG5V.n7855 ASIG5V.n7854 0.0380882
R48615 ASIG5V.n10713 ASIG5V.n10712 0.0380882
R48616 ASIG5V.n10712 ASIG5V.n10711 0.0380882
R48617 ASIG5V.n10711 ASIG5V.n10710 0.0380882
R48618 ASIG5V.n10710 ASIG5V.n10709 0.0380882
R48619 ASIG5V.n10709 ASIG5V.n10708 0.0380882
R48620 ASIG5V.n10708 ASIG5V.n10707 0.0380882
R48621 ASIG5V.n10707 ASIG5V.n10706 0.0380882
R48622 ASIG5V.n10706 ASIG5V.n10705 0.0380882
R48623 ASIG5V.n10705 ASIG5V.n10704 0.0380882
R48624 ASIG5V.n10704 ASIG5V.n10703 0.0380882
R48625 ASIG5V.n10703 ASIG5V.n10702 0.0380882
R48626 ASIG5V.n10702 ASIG5V.n10701 0.0380882
R48627 ASIG5V.n10701 ASIG5V.n10700 0.0380882
R48628 ASIG5V.n10700 ASIG5V.n10699 0.0380882
R48629 ASIG5V.n10699 ASIG5V.n10698 0.0380882
R48630 ASIG5V.n10698 ASIG5V.n10697 0.0380882
R48631 ASIG5V.n10697 ASIG5V.n10696 0.0380882
R48632 ASIG5V.n10696 ASIG5V.n10695 0.0380882
R48633 ASIG5V.n10695 ASIG5V.n10694 0.0380882
R48634 ASIG5V.n10694 ASIG5V.n10693 0.0380882
R48635 ASIG5V.n10693 ASIG5V.n10692 0.0380882
R48636 ASIG5V.n10692 ASIG5V.n10691 0.0380882
R48637 ASIG5V.n10691 ASIG5V.n10690 0.0380882
R48638 ASIG5V.n10690 ASIG5V.n10689 0.0380882
R48639 ASIG5V.n10689 ASIG5V.n10688 0.0380882
R48640 ASIG5V.n10688 ASIG5V.n10687 0.0380882
R48641 ASIG5V.n10687 ASIG5V.n10686 0.0380882
R48642 ASIG5V.n10686 ASIG5V.n10685 0.0380882
R48643 ASIG5V.n10685 ASIG5V.n10684 0.0380882
R48644 ASIG5V.n10684 ASIG5V.n10683 0.0380882
R48645 ASIG5V.n10683 ASIG5V.n10682 0.0380882
R48646 ASIG5V.n10682 ASIG5V.n10681 0.0380882
R48647 ASIG5V.n10681 ASIG5V.n10680 0.0380882
R48648 ASIG5V.n10680 ASIG5V.n10679 0.0380882
R48649 ASIG5V.n10679 ASIG5V.n10678 0.0380882
R48650 ASIG5V.n10678 ASIG5V.n10677 0.0380882
R48651 ASIG5V.n10677 ASIG5V.n10676 0.0380882
R48652 ASIG5V.n10676 ASIG5V.n10675 0.0380882
R48653 ASIG5V.n10675 ASIG5V.n10674 0.0380882
R48654 ASIG5V.n10674 ASIG5V.n10673 0.0380882
R48655 ASIG5V.n10673 ASIG5V.n10672 0.0380882
R48656 ASIG5V.n10672 ASIG5V.n10671 0.0380882
R48657 ASIG5V.n10671 ASIG5V.n10670 0.0380882
R48658 ASIG5V.n10670 ASIG5V.n10669 0.0380882
R48659 ASIG5V.n10669 ASIG5V.n10668 0.0380882
R48660 ASIG5V.n9335 ASIG5V.n9334 0.0380882
R48661 ASIG5V.n9336 ASIG5V.n9335 0.0380882
R48662 ASIG5V.n9337 ASIG5V.n9336 0.0380882
R48663 ASIG5V.n9338 ASIG5V.n9337 0.0380882
R48664 ASIG5V.n9339 ASIG5V.n9338 0.0380882
R48665 ASIG5V.n9340 ASIG5V.n9339 0.0380882
R48666 ASIG5V.n9341 ASIG5V.n9340 0.0380882
R48667 ASIG5V.n9342 ASIG5V.n9341 0.0380882
R48668 ASIG5V.n9343 ASIG5V.n9342 0.0380882
R48669 ASIG5V.n9344 ASIG5V.n9343 0.0380882
R48670 ASIG5V.n9345 ASIG5V.n9344 0.0380882
R48671 ASIG5V.n7240 ASIG5V.n7239 0.0380882
R48672 ASIG5V.n7239 ASIG5V.n7238 0.0380882
R48673 ASIG5V.n7238 ASIG5V.n7237 0.0380882
R48674 ASIG5V.n7237 ASIG5V.n7236 0.0380882
R48675 ASIG5V.n7236 ASIG5V.n7235 0.0380882
R48676 ASIG5V.n7235 ASIG5V.n7234 0.0380882
R48677 ASIG5V.n7234 ASIG5V.n7233 0.0380882
R48678 ASIG5V.n7233 ASIG5V.n7232 0.0380882
R48679 ASIG5V.n7232 ASIG5V.n7231 0.0380882
R48680 ASIG5V.n7231 ASIG5V.n7230 0.0380882
R48681 ASIG5V.n7230 ASIG5V.n7229 0.0380882
R48682 ASIG5V.n7229 ASIG5V.n7228 0.0380882
R48683 ASIG5V.n7228 ASIG5V.n7227 0.0380882
R48684 ASIG5V.n7227 ASIG5V.n7226 0.0380882
R48685 ASIG5V.n7226 ASIG5V.n7225 0.0380882
R48686 ASIG5V.n7225 ASIG5V.n7224 0.0380882
R48687 ASIG5V.n7224 ASIG5V.n7223 0.0380882
R48688 ASIG5V.n7223 ASIG5V.n7222 0.0380882
R48689 ASIG5V.n7222 ASIG5V.n7221 0.0380882
R48690 ASIG5V.n7221 ASIG5V.n7220 0.0380882
R48691 ASIG5V.n7220 ASIG5V.n7219 0.0380882
R48692 ASIG5V.n7219 ASIG5V.n7218 0.0380882
R48693 ASIG5V.n7218 ASIG5V.n7217 0.0380882
R48694 ASIG5V.n7217 ASIG5V.n7216 0.0380882
R48695 ASIG5V.n7216 ASIG5V.n7215 0.0380882
R48696 ASIG5V.n7215 ASIG5V.n7214 0.0380882
R48697 ASIG5V.n7214 ASIG5V.n7213 0.0380882
R48698 ASIG5V.n7213 ASIG5V.n7212 0.0380882
R48699 ASIG5V.n7212 ASIG5V.n7211 0.0380882
R48700 ASIG5V.n7211 ASIG5V.n7210 0.0380882
R48701 ASIG5V.n10667 ASIG5V.n10666 0.0380882
R48702 ASIG5V.n10666 ASIG5V.n10665 0.0380882
R48703 ASIG5V.n10665 ASIG5V.n10664 0.0380882
R48704 ASIG5V.n10664 ASIG5V.n10663 0.0380882
R48705 ASIG5V.n10663 ASIG5V.n10662 0.0380882
R48706 ASIG5V.n10662 ASIG5V.n10661 0.0380882
R48707 ASIG5V.n10661 ASIG5V.n10660 0.0380882
R48708 ASIG5V.n10660 ASIG5V.n10659 0.0380882
R48709 ASIG5V.n10659 ASIG5V.n10658 0.0380882
R48710 ASIG5V.n10658 ASIG5V.n10657 0.0380882
R48711 ASIG5V.n10657 ASIG5V.n10656 0.0380882
R48712 ASIG5V.n10656 ASIG5V.n10655 0.0380882
R48713 ASIG5V.n10655 ASIG5V.n10654 0.0380882
R48714 ASIG5V.n10654 ASIG5V.n10653 0.0380882
R48715 ASIG5V.n10653 ASIG5V.n10652 0.0380882
R48716 ASIG5V.n10652 ASIG5V.n10651 0.0380882
R48717 ASIG5V.n10651 ASIG5V.n10650 0.0380882
R48718 ASIG5V.n10650 ASIG5V.n10649 0.0380882
R48719 ASIG5V.n10649 ASIG5V.n10648 0.0380882
R48720 ASIG5V.n10648 ASIG5V.n10647 0.0380882
R48721 ASIG5V.n10647 ASIG5V.n10646 0.0380882
R48722 ASIG5V.n10646 ASIG5V.n10645 0.0380882
R48723 ASIG5V.n10645 ASIG5V.n10644 0.0380882
R48724 ASIG5V.n10644 ASIG5V.n10643 0.0380882
R48725 ASIG5V.n10643 ASIG5V.n10642 0.0380882
R48726 ASIG5V.n10642 ASIG5V.n10641 0.0380882
R48727 ASIG5V.n10641 ASIG5V.n10640 0.0380882
R48728 ASIG5V.n10640 ASIG5V.n10639 0.0380882
R48729 ASIG5V.n10639 ASIG5V.n10638 0.0380882
R48730 ASIG5V.n10638 ASIG5V.n10637 0.0380882
R48731 ASIG5V.n10637 ASIG5V.n10636 0.0380882
R48732 ASIG5V.n10636 ASIG5V.n10635 0.0380882
R48733 ASIG5V.n10635 ASIG5V.n10634 0.0380882
R48734 ASIG5V.n10634 ASIG5V.n10633 0.0380882
R48735 ASIG5V.n10633 ASIG5V.n10632 0.0380882
R48736 ASIG5V.n10632 ASIG5V.n10631 0.0380882
R48737 ASIG5V.n10631 ASIG5V.n10630 0.0380882
R48738 ASIG5V.n10630 ASIG5V.n10629 0.0380882
R48739 ASIG5V.n10629 ASIG5V.n10628 0.0380882
R48740 ASIG5V.n10628 ASIG5V.n10627 0.0380882
R48741 ASIG5V.n10627 ASIG5V.n10626 0.0380882
R48742 ASIG5V.n10626 ASIG5V.n10625 0.0380882
R48743 ASIG5V.n10625 ASIG5V.n10624 0.0380882
R48744 ASIG5V.n10624 ASIG5V.n10623 0.0380882
R48745 ASIG5V.n10623 ASIG5V.n10622 0.0380882
R48746 ASIG5V.n10622 ASIG5V.n10621 0.0380882
R48747 ASIG5V.n9320 ASIG5V.n9319 0.0380882
R48748 ASIG5V.n9321 ASIG5V.n9320 0.0380882
R48749 ASIG5V.n9322 ASIG5V.n9321 0.0380882
R48750 ASIG5V.n9323 ASIG5V.n9322 0.0380882
R48751 ASIG5V.n9324 ASIG5V.n9323 0.0380882
R48752 ASIG5V.n9325 ASIG5V.n9324 0.0380882
R48753 ASIG5V.n9326 ASIG5V.n9325 0.0380882
R48754 ASIG5V.n9327 ASIG5V.n9326 0.0380882
R48755 ASIG5V.n9328 ASIG5V.n9327 0.0380882
R48756 ASIG5V.n9329 ASIG5V.n9328 0.0380882
R48757 ASIG5V.n9330 ASIG5V.n9329 0.0380882
R48758 ASIG5V.n9331 ASIG5V.n9330 0.0380882
R48759 ASIG5V.n9332 ASIG5V.n9331 0.0380882
R48760 ASIG5V.n9333 ASIG5V.n9332 0.0380882
R48761 ASIG5V.n12642 ASIG5V.n12641 0.0380882
R48762 ASIG5V.n12641 ASIG5V.n12640 0.0380882
R48763 ASIG5V.n12640 ASIG5V.n12639 0.0380882
R48764 ASIG5V.n12639 ASIG5V.n12638 0.0380882
R48765 ASIG5V.n12638 ASIG5V.n12637 0.0380882
R48766 ASIG5V.n12637 ASIG5V.n12636 0.0380882
R48767 ASIG5V.n12636 ASIG5V.n12635 0.0380882
R48768 ASIG5V.n12635 ASIG5V.n12634 0.0380882
R48769 ASIG5V.n12634 ASIG5V.n12633 0.0380882
R48770 ASIG5V.n12633 ASIG5V.n12632 0.0380882
R48771 ASIG5V.n12632 ASIG5V.n12631 0.0380882
R48772 ASIG5V.n12631 ASIG5V.n12630 0.0380882
R48773 ASIG5V.n12630 ASIG5V.n12629 0.0380882
R48774 ASIG5V.n12629 ASIG5V.n12628 0.0380882
R48775 ASIG5V.n12628 ASIG5V.n12627 0.0380882
R48776 ASIG5V.n12627 ASIG5V.n12626 0.0380882
R48777 ASIG5V.n12626 ASIG5V.n12625 0.0380882
R48778 ASIG5V.n12625 ASIG5V.n12624 0.0380882
R48779 ASIG5V.n12624 ASIG5V.n12623 0.0380882
R48780 ASIG5V.n12623 ASIG5V.n12622 0.0380882
R48781 ASIG5V.n12622 ASIG5V.n12621 0.0380882
R48782 ASIG5V.n12621 ASIG5V.n12620 0.0380882
R48783 ASIG5V.n12620 ASIG5V.n12619 0.0380882
R48784 ASIG5V.n12619 ASIG5V.n12618 0.0380882
R48785 ASIG5V.n12618 ASIG5V.n12617 0.0380882
R48786 ASIG5V.n12617 ASIG5V.n12616 0.0380882
R48787 ASIG5V.n12616 ASIG5V.n12615 0.0380882
R48788 ASIG5V.n12615 ASIG5V.n12614 0.0380882
R48789 ASIG5V.n12614 ASIG5V.n12613 0.0380882
R48790 ASIG5V.n12613 ASIG5V.n12612 0.0380882
R48791 ASIG5V.n10620 ASIG5V.n10619 0.0380882
R48792 ASIG5V.n10619 ASIG5V.n10618 0.0380882
R48793 ASIG5V.n10618 ASIG5V.n10617 0.0380882
R48794 ASIG5V.n10617 ASIG5V.n10616 0.0380882
R48795 ASIG5V.n10616 ASIG5V.n10615 0.0380882
R48796 ASIG5V.n10615 ASIG5V.n10614 0.0380882
R48797 ASIG5V.n10614 ASIG5V.n10613 0.0380882
R48798 ASIG5V.n10613 ASIG5V.n10612 0.0380882
R48799 ASIG5V.n10612 ASIG5V.n10611 0.0380882
R48800 ASIG5V.n10611 ASIG5V.n10610 0.0380882
R48801 ASIG5V.n10610 ASIG5V.n10609 0.0380882
R48802 ASIG5V.n10609 ASIG5V.n10608 0.0380882
R48803 ASIG5V.n10608 ASIG5V.n10607 0.0380882
R48804 ASIG5V.n10607 ASIG5V.n10606 0.0380882
R48805 ASIG5V.n10606 ASIG5V.n10605 0.0380882
R48806 ASIG5V.n10605 ASIG5V.n10604 0.0380882
R48807 ASIG5V.n10604 ASIG5V.n10603 0.0380882
R48808 ASIG5V.n10603 ASIG5V.n10602 0.0380882
R48809 ASIG5V.n10602 ASIG5V.n10601 0.0380882
R48810 ASIG5V.n10601 ASIG5V.n10600 0.0380882
R48811 ASIG5V.n10600 ASIG5V.n10599 0.0380882
R48812 ASIG5V.n10599 ASIG5V.n10598 0.0380882
R48813 ASIG5V.n10598 ASIG5V.n10597 0.0380882
R48814 ASIG5V.n10597 ASIG5V.n10596 0.0380882
R48815 ASIG5V.n10596 ASIG5V.n10595 0.0380882
R48816 ASIG5V.n10595 ASIG5V.n10594 0.0380882
R48817 ASIG5V.n10594 ASIG5V.n10593 0.0380882
R48818 ASIG5V.n10593 ASIG5V.n10592 0.0380882
R48819 ASIG5V.n10592 ASIG5V.n10591 0.0380882
R48820 ASIG5V.n10591 ASIG5V.n10590 0.0380882
R48821 ASIG5V.n10590 ASIG5V.n10589 0.0380882
R48822 ASIG5V.n10589 ASIG5V.n10588 0.0380882
R48823 ASIG5V.n10588 ASIG5V.n10587 0.0380882
R48824 ASIG5V.n10587 ASIG5V.n10586 0.0380882
R48825 ASIG5V.n10586 ASIG5V.n10585 0.0380882
R48826 ASIG5V.n10585 ASIG5V.n10584 0.0380882
R48827 ASIG5V.n10584 ASIG5V.n10583 0.0380882
R48828 ASIG5V.n10583 ASIG5V.n10582 0.0380882
R48829 ASIG5V.n10582 ASIG5V.n10581 0.0380882
R48830 ASIG5V.n10581 ASIG5V.n10580 0.0380882
R48831 ASIG5V.n10580 ASIG5V.n10579 0.0380882
R48832 ASIG5V.n10579 ASIG5V.n10578 0.0380882
R48833 ASIG5V.n10578 ASIG5V.n10577 0.0380882
R48834 ASIG5V.n10577 ASIG5V.n10576 0.0380882
R48835 ASIG5V.n10576 ASIG5V.n10575 0.0380882
R48836 ASIG5V.n10575 ASIG5V.n10574 0.0380882
R48837 ASIG5V.n10574 ASIG5V.n10573 0.0380882
R48838 ASIG5V.n9303 ASIG5V.n9302 0.0380882
R48839 ASIG5V.n9304 ASIG5V.n9303 0.0380882
R48840 ASIG5V.n9305 ASIG5V.n9304 0.0380882
R48841 ASIG5V.n9306 ASIG5V.n9305 0.0380882
R48842 ASIG5V.n9307 ASIG5V.n9306 0.0380882
R48843 ASIG5V.n9308 ASIG5V.n9307 0.0380882
R48844 ASIG5V.n9309 ASIG5V.n9308 0.0380882
R48845 ASIG5V.n9310 ASIG5V.n9309 0.0380882
R48846 ASIG5V.n9311 ASIG5V.n9310 0.0380882
R48847 ASIG5V.n9312 ASIG5V.n9311 0.0380882
R48848 ASIG5V.n9313 ASIG5V.n9312 0.0380882
R48849 ASIG5V.n9314 ASIG5V.n9313 0.0380882
R48850 ASIG5V.n9315 ASIG5V.n9314 0.0380882
R48851 ASIG5V.n9316 ASIG5V.n9315 0.0380882
R48852 ASIG5V.n9317 ASIG5V.n9316 0.0380882
R48853 ASIG5V.n9318 ASIG5V.n9317 0.0380882
R48854 ASIG5V.n12416 ASIG5V.n12415 0.0380882
R48855 ASIG5V.n12415 ASIG5V.n12414 0.0380882
R48856 ASIG5V.n12414 ASIG5V.n12413 0.0380882
R48857 ASIG5V.n12413 ASIG5V.n12412 0.0380882
R48858 ASIG5V.n12412 ASIG5V.n12411 0.0380882
R48859 ASIG5V.n12411 ASIG5V.n12410 0.0380882
R48860 ASIG5V.n12410 ASIG5V.n12409 0.0380882
R48861 ASIG5V.n12409 ASIG5V.n12408 0.0380882
R48862 ASIG5V.n12408 ASIG5V.n12407 0.0380882
R48863 ASIG5V.n12407 ASIG5V.n12406 0.0380882
R48864 ASIG5V.n12406 ASIG5V.n12405 0.0380882
R48865 ASIG5V.n12405 ASIG5V.n12404 0.0380882
R48866 ASIG5V.n12404 ASIG5V.n12403 0.0380882
R48867 ASIG5V.n12403 ASIG5V.n12402 0.0380882
R48868 ASIG5V.n12402 ASIG5V.n12401 0.0380882
R48869 ASIG5V.n12401 ASIG5V.n12400 0.0380882
R48870 ASIG5V.n12400 ASIG5V.n12399 0.0380882
R48871 ASIG5V.n12399 ASIG5V.n12398 0.0380882
R48872 ASIG5V.n12398 ASIG5V.n12397 0.0380882
R48873 ASIG5V.n12397 ASIG5V.n12396 0.0380882
R48874 ASIG5V.n12396 ASIG5V.n12395 0.0380882
R48875 ASIG5V.n12395 ASIG5V.n12394 0.0380882
R48876 ASIG5V.n12394 ASIG5V.n12393 0.0380882
R48877 ASIG5V.n12393 ASIG5V.n12392 0.0380882
R48878 ASIG5V.n12392 ASIG5V.n12391 0.0380882
R48879 ASIG5V.n12391 ASIG5V.n12390 0.0380882
R48880 ASIG5V.n12390 ASIG5V.n12389 0.0380882
R48881 ASIG5V.n12389 ASIG5V.n12388 0.0380882
R48882 ASIG5V.n12388 ASIG5V.n12387 0.0380882
R48883 ASIG5V.n12387 ASIG5V.n12386 0.0380882
R48884 ASIG5V.n9061 ASIG5V.n9060 0.0380882
R48885 ASIG5V.n10292 ASIG5V.n10291 0.0380882
R48886 ASIG5V.n10291 ASIG5V.n10290 0.0380882
R48887 ASIG5V.n10290 ASIG5V.n10289 0.0380882
R48888 ASIG5V.n10289 ASIG5V.n10288 0.0380882
R48889 ASIG5V.n10288 ASIG5V.n10287 0.0380882
R48890 ASIG5V.n10287 ASIG5V.n10286 0.0380882
R48891 ASIG5V.n10286 ASIG5V.n10285 0.0380882
R48892 ASIG5V.n10285 ASIG5V.n10284 0.0380882
R48893 ASIG5V.n10284 ASIG5V.n10283 0.0380882
R48894 ASIG5V.n10283 ASIG5V.n10282 0.0380882
R48895 ASIG5V.n10282 ASIG5V.n10281 0.0380882
R48896 ASIG5V.n10281 ASIG5V.n10280 0.0380882
R48897 ASIG5V.n10280 ASIG5V.n10279 0.0380882
R48898 ASIG5V.n10279 ASIG5V.n10278 0.0380882
R48899 ASIG5V.n10278 ASIG5V.n10277 0.0380882
R48900 ASIG5V.n10277 ASIG5V.n10276 0.0380882
R48901 ASIG5V.n10276 ASIG5V.n10275 0.0380882
R48902 ASIG5V.n10275 ASIG5V.n10274 0.0380882
R48903 ASIG5V.n10274 ASIG5V.n10273 0.0380882
R48904 ASIG5V.n10273 ASIG5V.n10272 0.0380882
R48905 ASIG5V.n10272 ASIG5V.n10271 0.0380882
R48906 ASIG5V.n10271 ASIG5V.n10270 0.0380882
R48907 ASIG5V.n10270 ASIG5V.n10269 0.0380882
R48908 ASIG5V.n10269 ASIG5V.n10268 0.0380882
R48909 ASIG5V.n10268 ASIG5V.n10267 0.0380882
R48910 ASIG5V.n10267 ASIG5V.n10266 0.0380882
R48911 ASIG5V.n10266 ASIG5V.n10265 0.0380882
R48912 ASIG5V.n10265 ASIG5V.n10264 0.0380882
R48913 ASIG5V.n10264 ASIG5V.n10263 0.0380882
R48914 ASIG5V.n10263 ASIG5V.n10262 0.0380882
R48915 ASIG5V.n10262 ASIG5V.n10261 0.0380882
R48916 ASIG5V.n10261 ASIG5V.n10260 0.0380882
R48917 ASIG5V.n10260 ASIG5V.n10259 0.0380882
R48918 ASIG5V.n10259 ASIG5V.n10258 0.0380882
R48919 ASIG5V.n10258 ASIG5V.n10257 0.0380882
R48920 ASIG5V.n10257 ASIG5V.n10256 0.0380882
R48921 ASIG5V.n10256 ASIG5V.n10255 0.0380882
R48922 ASIG5V.n10255 ASIG5V.n10254 0.0380882
R48923 ASIG5V.n10254 ASIG5V.n10253 0.0380882
R48924 ASIG5V.n10253 ASIG5V.n10252 0.0380882
R48925 ASIG5V.n10252 ASIG5V.n10251 0.0380882
R48926 ASIG5V.n10251 ASIG5V.n10250 0.0380882
R48927 ASIG5V.n10250 ASIG5V.n10249 0.0380882
R48928 ASIG5V.n10249 ASIG5V.n10248 0.0380882
R48929 ASIG5V.n10248 ASIG5V.n10247 0.0380882
R48930 ASIG5V.n10247 ASIG5V.n10246 0.0380882
R48931 ASIG5V.n10246 ASIG5V.n10245 0.0380882
R48932 ASIG5V.n10245 ASIG5V.n10244 0.0380882
R48933 ASIG5V.n10244 ASIG5V.n10243 0.0380882
R48934 ASIG5V.n9284 ASIG5V.n9283 0.0380882
R48935 ASIG5V.n9285 ASIG5V.n9284 0.0380882
R48936 ASIG5V.n9286 ASIG5V.n9285 0.0380882
R48937 ASIG5V.n9287 ASIG5V.n9286 0.0380882
R48938 ASIG5V.n9288 ASIG5V.n9287 0.0380882
R48939 ASIG5V.n9289 ASIG5V.n9288 0.0380882
R48940 ASIG5V.n9290 ASIG5V.n9289 0.0380882
R48941 ASIG5V.n9291 ASIG5V.n9290 0.0380882
R48942 ASIG5V.n9292 ASIG5V.n9291 0.0380882
R48943 ASIG5V.n9293 ASIG5V.n9292 0.0380882
R48944 ASIG5V.n9294 ASIG5V.n9293 0.0380882
R48945 ASIG5V.n9295 ASIG5V.n9294 0.0380882
R48946 ASIG5V.n9296 ASIG5V.n9295 0.0380882
R48947 ASIG5V.n9297 ASIG5V.n9296 0.0380882
R48948 ASIG5V.n9298 ASIG5V.n9297 0.0380882
R48949 ASIG5V.n9299 ASIG5V.n9298 0.0380882
R48950 ASIG5V.n9300 ASIG5V.n9299 0.0380882
R48951 ASIG5V.n9301 ASIG5V.n9300 0.0380882
R48952 ASIG5V.n12299 ASIG5V.n12298 0.0380882
R48953 ASIG5V.n12298 ASIG5V.n12297 0.0380882
R48954 ASIG5V.n12297 ASIG5V.n12296 0.0380882
R48955 ASIG5V.n12296 ASIG5V.n12295 0.0380882
R48956 ASIG5V.n12295 ASIG5V.n12294 0.0380882
R48957 ASIG5V.n12294 ASIG5V.n12293 0.0380882
R48958 ASIG5V.n12293 ASIG5V.n12292 0.0380882
R48959 ASIG5V.n12292 ASIG5V.n12291 0.0380882
R48960 ASIG5V.n12291 ASIG5V.n12290 0.0380882
R48961 ASIG5V.n12290 ASIG5V.n12289 0.0380882
R48962 ASIG5V.n12289 ASIG5V.n12288 0.0380882
R48963 ASIG5V.n12288 ASIG5V.n12287 0.0380882
R48964 ASIG5V.n12287 ASIG5V.n12286 0.0380882
R48965 ASIG5V.n12286 ASIG5V.n12285 0.0380882
R48966 ASIG5V.n12285 ASIG5V.n12284 0.0380882
R48967 ASIG5V.n12284 ASIG5V.n12283 0.0380882
R48968 ASIG5V.n12283 ASIG5V.n12282 0.0380882
R48969 ASIG5V.n12282 ASIG5V.n12281 0.0380882
R48970 ASIG5V.n12281 ASIG5V.n12280 0.0380882
R48971 ASIG5V.n12280 ASIG5V.n12279 0.0380882
R48972 ASIG5V.n12279 ASIG5V.n12278 0.0380882
R48973 ASIG5V.n12278 ASIG5V.n12277 0.0380882
R48974 ASIG5V.n12277 ASIG5V.n12276 0.0380882
R48975 ASIG5V.n12276 ASIG5V.n12275 0.0380882
R48976 ASIG5V.n12275 ASIG5V.n12274 0.0380882
R48977 ASIG5V.n12274 ASIG5V.n12273 0.0380882
R48978 ASIG5V.n12273 ASIG5V.n12272 0.0380882
R48979 ASIG5V.n12272 ASIG5V.n12271 0.0380882
R48980 ASIG5V.n12271 ASIG5V.n12270 0.0380882
R48981 ASIG5V.n12270 ASIG5V.n12269 0.0380882
R48982 ASIG5V.n9057 ASIG5V.n9056 0.0380882
R48983 ASIG5V.n9058 ASIG5V.n9057 0.0380882
R48984 ASIG5V.n9059 ASIG5V.n9058 0.0380882
R48985 ASIG5V.n10242 ASIG5V.n10241 0.0380882
R48986 ASIG5V.n10241 ASIG5V.n10240 0.0380882
R48987 ASIG5V.n10240 ASIG5V.n10239 0.0380882
R48988 ASIG5V.n10239 ASIG5V.n10238 0.0380882
R48989 ASIG5V.n10238 ASIG5V.n10237 0.0380882
R48990 ASIG5V.n10237 ASIG5V.n10236 0.0380882
R48991 ASIG5V.n10236 ASIG5V.n10235 0.0380882
R48992 ASIG5V.n10235 ASIG5V.n10234 0.0380882
R48993 ASIG5V.n10234 ASIG5V.n10233 0.0380882
R48994 ASIG5V.n10233 ASIG5V.n10232 0.0380882
R48995 ASIG5V.n10232 ASIG5V.n10231 0.0380882
R48996 ASIG5V.n10231 ASIG5V.n10230 0.0380882
R48997 ASIG5V.n10230 ASIG5V.n10229 0.0380882
R48998 ASIG5V.n10229 ASIG5V.n10228 0.0380882
R48999 ASIG5V.n10228 ASIG5V.n10227 0.0380882
R49000 ASIG5V.n10227 ASIG5V.n10226 0.0380882
R49001 ASIG5V.n10226 ASIG5V.n10225 0.0380882
R49002 ASIG5V.n10225 ASIG5V.n10224 0.0380882
R49003 ASIG5V.n10224 ASIG5V.n10223 0.0380882
R49004 ASIG5V.n10223 ASIG5V.n10222 0.0380882
R49005 ASIG5V.n10222 ASIG5V.n10221 0.0380882
R49006 ASIG5V.n10221 ASIG5V.n10220 0.0380882
R49007 ASIG5V.n10220 ASIG5V.n10219 0.0380882
R49008 ASIG5V.n10219 ASIG5V.n10218 0.0380882
R49009 ASIG5V.n10218 ASIG5V.n10217 0.0380882
R49010 ASIG5V.n10217 ASIG5V.n10216 0.0380882
R49011 ASIG5V.n10216 ASIG5V.n10215 0.0380882
R49012 ASIG5V.n10215 ASIG5V.n10214 0.0380882
R49013 ASIG5V.n10214 ASIG5V.n10213 0.0380882
R49014 ASIG5V.n10213 ASIG5V.n10212 0.0380882
R49015 ASIG5V.n10212 ASIG5V.n10211 0.0380882
R49016 ASIG5V.n10211 ASIG5V.n10210 0.0380882
R49017 ASIG5V.n10210 ASIG5V.n10209 0.0380882
R49018 ASIG5V.n10209 ASIG5V.n10208 0.0380882
R49019 ASIG5V.n10208 ASIG5V.n10207 0.0380882
R49020 ASIG5V.n10207 ASIG5V.n10206 0.0380882
R49021 ASIG5V.n10206 ASIG5V.n10205 0.0380882
R49022 ASIG5V.n10205 ASIG5V.n10204 0.0380882
R49023 ASIG5V.n10204 ASIG5V.n10203 0.0380882
R49024 ASIG5V.n10203 ASIG5V.n10202 0.0380882
R49025 ASIG5V.n10202 ASIG5V.n10201 0.0380882
R49026 ASIG5V.n10201 ASIG5V.n10200 0.0380882
R49027 ASIG5V.n10200 ASIG5V.n10199 0.0380882
R49028 ASIG5V.n10199 ASIG5V.n10198 0.0380882
R49029 ASIG5V.n10198 ASIG5V.n10197 0.0380882
R49030 ASIG5V.n10197 ASIG5V.n10196 0.0380882
R49031 ASIG5V.n10196 ASIG5V.n10195 0.0380882
R49032 ASIG5V.n10195 ASIG5V.n10194 0.0380882
R49033 ASIG5V.n10194 ASIG5V.n10193 0.0380882
R49034 ASIG5V.n10193 ASIG5V.n10192 0.0380882
R49035 ASIG5V.n9262 ASIG5V.n9261 0.0380882
R49036 ASIG5V.n9263 ASIG5V.n9262 0.0380882
R49037 ASIG5V.n9264 ASIG5V.n9263 0.0380882
R49038 ASIG5V.n9265 ASIG5V.n9264 0.0380882
R49039 ASIG5V.n9266 ASIG5V.n9265 0.0380882
R49040 ASIG5V.n9267 ASIG5V.n9266 0.0380882
R49041 ASIG5V.n9268 ASIG5V.n9267 0.0380882
R49042 ASIG5V.n9269 ASIG5V.n9268 0.0380882
R49043 ASIG5V.n9270 ASIG5V.n9269 0.0380882
R49044 ASIG5V.n9271 ASIG5V.n9270 0.0380882
R49045 ASIG5V.n9272 ASIG5V.n9271 0.0380882
R49046 ASIG5V.n9273 ASIG5V.n9272 0.0380882
R49047 ASIG5V.n9274 ASIG5V.n9273 0.0380882
R49048 ASIG5V.n9275 ASIG5V.n9274 0.0380882
R49049 ASIG5V.n9276 ASIG5V.n9275 0.0380882
R49050 ASIG5V.n9277 ASIG5V.n9276 0.0380882
R49051 ASIG5V.n9278 ASIG5V.n9277 0.0380882
R49052 ASIG5V.n9279 ASIG5V.n9278 0.0380882
R49053 ASIG5V.n9280 ASIG5V.n9279 0.0380882
R49054 ASIG5V.n9281 ASIG5V.n9280 0.0380882
R49055 ASIG5V.n9282 ASIG5V.n9281 0.0380882
R49056 ASIG5V.n12146 ASIG5V.n12145 0.0380882
R49057 ASIG5V.n12145 ASIG5V.n12144 0.0380882
R49058 ASIG5V.n12144 ASIG5V.n12143 0.0380882
R49059 ASIG5V.n12143 ASIG5V.n12142 0.0380882
R49060 ASIG5V.n12142 ASIG5V.n12141 0.0380882
R49061 ASIG5V.n12141 ASIG5V.n12140 0.0380882
R49062 ASIG5V.n12140 ASIG5V.n12139 0.0380882
R49063 ASIG5V.n12139 ASIG5V.n12138 0.0380882
R49064 ASIG5V.n12138 ASIG5V.n12137 0.0380882
R49065 ASIG5V.n12137 ASIG5V.n12136 0.0380882
R49066 ASIG5V.n12136 ASIG5V.n12135 0.0380882
R49067 ASIG5V.n12135 ASIG5V.n12134 0.0380882
R49068 ASIG5V.n12134 ASIG5V.n12133 0.0380882
R49069 ASIG5V.n12133 ASIG5V.n12132 0.0380882
R49070 ASIG5V.n12132 ASIG5V.n12131 0.0380882
R49071 ASIG5V.n12131 ASIG5V.n12130 0.0380882
R49072 ASIG5V.n12130 ASIG5V.n12129 0.0380882
R49073 ASIG5V.n12129 ASIG5V.n12128 0.0380882
R49074 ASIG5V.n12128 ASIG5V.n12127 0.0380882
R49075 ASIG5V.n12127 ASIG5V.n12126 0.0380882
R49076 ASIG5V.n12126 ASIG5V.n12125 0.0380882
R49077 ASIG5V.n12125 ASIG5V.n12124 0.0380882
R49078 ASIG5V.n12124 ASIG5V.n12123 0.0380882
R49079 ASIG5V.n12123 ASIG5V.n12122 0.0380882
R49080 ASIG5V.n12122 ASIG5V.n12121 0.0380882
R49081 ASIG5V.n12121 ASIG5V.n12120 0.0380882
R49082 ASIG5V.n12120 ASIG5V.n12119 0.0380882
R49083 ASIG5V.n12119 ASIG5V.n12118 0.0380882
R49084 ASIG5V.n12118 ASIG5V.n12117 0.0380882
R49085 ASIG5V.n12117 ASIG5V.n12116 0.0380882
R49086 ASIG5V.n9051 ASIG5V.n9050 0.0380882
R49087 ASIG5V.n9052 ASIG5V.n9051 0.0380882
R49088 ASIG5V.n9053 ASIG5V.n9052 0.0380882
R49089 ASIG5V.n9054 ASIG5V.n9053 0.0380882
R49090 ASIG5V.n9055 ASIG5V.n9054 0.0380882
R49091 ASIG5V.n10191 ASIG5V.n10190 0.0380882
R49092 ASIG5V.n10190 ASIG5V.n10189 0.0380882
R49093 ASIG5V.n10189 ASIG5V.n10188 0.0380882
R49094 ASIG5V.n10188 ASIG5V.n10187 0.0380882
R49095 ASIG5V.n10187 ASIG5V.n10186 0.0380882
R49096 ASIG5V.n10186 ASIG5V.n10185 0.0380882
R49097 ASIG5V.n10185 ASIG5V.n10184 0.0380882
R49098 ASIG5V.n10184 ASIG5V.n10183 0.0380882
R49099 ASIG5V.n10183 ASIG5V.n10182 0.0380882
R49100 ASIG5V.n10182 ASIG5V.n10181 0.0380882
R49101 ASIG5V.n10181 ASIG5V.n10180 0.0380882
R49102 ASIG5V.n10180 ASIG5V.n10179 0.0380882
R49103 ASIG5V.n10179 ASIG5V.n10178 0.0380882
R49104 ASIG5V.n10178 ASIG5V.n10177 0.0380882
R49105 ASIG5V.n10177 ASIG5V.n10176 0.0380882
R49106 ASIG5V.n10176 ASIG5V.n10175 0.0380882
R49107 ASIG5V.n10175 ASIG5V.n10174 0.0380882
R49108 ASIG5V.n10174 ASIG5V.n10173 0.0380882
R49109 ASIG5V.n10173 ASIG5V.n10172 0.0380882
R49110 ASIG5V.n10172 ASIG5V.n10171 0.0380882
R49111 ASIG5V.n10171 ASIG5V.n10170 0.0380882
R49112 ASIG5V.n10170 ASIG5V.n10169 0.0380882
R49113 ASIG5V.n10169 ASIG5V.n10168 0.0380882
R49114 ASIG5V.n10168 ASIG5V.n10167 0.0380882
R49115 ASIG5V.n10167 ASIG5V.n10166 0.0380882
R49116 ASIG5V.n10166 ASIG5V.n10165 0.0380882
R49117 ASIG5V.n10165 ASIG5V.n10164 0.0380882
R49118 ASIG5V.n10164 ASIG5V.n10163 0.0380882
R49119 ASIG5V.n10163 ASIG5V.n10162 0.0380882
R49120 ASIG5V.n10162 ASIG5V.n10161 0.0380882
R49121 ASIG5V.n10161 ASIG5V.n10160 0.0380882
R49122 ASIG5V.n10160 ASIG5V.n10159 0.0380882
R49123 ASIG5V.n10159 ASIG5V.n10158 0.0380882
R49124 ASIG5V.n10158 ASIG5V.n10157 0.0380882
R49125 ASIG5V.n10157 ASIG5V.n10156 0.0380882
R49126 ASIG5V.n10156 ASIG5V.n10155 0.0380882
R49127 ASIG5V.n10155 ASIG5V.n10154 0.0380882
R49128 ASIG5V.n10154 ASIG5V.n10153 0.0380882
R49129 ASIG5V.n10153 ASIG5V.n10152 0.0380882
R49130 ASIG5V.n10152 ASIG5V.n10151 0.0380882
R49131 ASIG5V.n10151 ASIG5V.n10150 0.0380882
R49132 ASIG5V.n10150 ASIG5V.n10149 0.0380882
R49133 ASIG5V.n10149 ASIG5V.n10148 0.0380882
R49134 ASIG5V.n10148 ASIG5V.n10147 0.0380882
R49135 ASIG5V.n10147 ASIG5V.n10146 0.0380882
R49136 ASIG5V.n10146 ASIG5V.n10145 0.0380882
R49137 ASIG5V.n10145 ASIG5V.n10144 0.0380882
R49138 ASIG5V.n10144 ASIG5V.n10143 0.0380882
R49139 ASIG5V.n10143 ASIG5V.n10142 0.0380882
R49140 ASIG5V.n10142 ASIG5V.n10141 0.0380882
R49141 ASIG5V.n10141 ASIG5V.n10140 0.0380882
R49142 ASIG5V.n10140 ASIG5V.n10139 0.0380882
R49143 ASIG5V.n9238 ASIG5V.n9237 0.0380882
R49144 ASIG5V.n9239 ASIG5V.n9238 0.0380882
R49145 ASIG5V.n9240 ASIG5V.n9239 0.0380882
R49146 ASIG5V.n9241 ASIG5V.n9240 0.0380882
R49147 ASIG5V.n9242 ASIG5V.n9241 0.0380882
R49148 ASIG5V.n9243 ASIG5V.n9242 0.0380882
R49149 ASIG5V.n9244 ASIG5V.n9243 0.0380882
R49150 ASIG5V.n9245 ASIG5V.n9244 0.0380882
R49151 ASIG5V.n9246 ASIG5V.n9245 0.0380882
R49152 ASIG5V.n9247 ASIG5V.n9246 0.0380882
R49153 ASIG5V.n9248 ASIG5V.n9247 0.0380882
R49154 ASIG5V.n9249 ASIG5V.n9248 0.0380882
R49155 ASIG5V.n9250 ASIG5V.n9249 0.0380882
R49156 ASIG5V.n9251 ASIG5V.n9250 0.0380882
R49157 ASIG5V.n9252 ASIG5V.n9251 0.0380882
R49158 ASIG5V.n9253 ASIG5V.n9252 0.0380882
R49159 ASIG5V.n9254 ASIG5V.n9253 0.0380882
R49160 ASIG5V.n9255 ASIG5V.n9254 0.0380882
R49161 ASIG5V.n9256 ASIG5V.n9255 0.0380882
R49162 ASIG5V.n9257 ASIG5V.n9256 0.0380882
R49163 ASIG5V.n9258 ASIG5V.n9257 0.0380882
R49164 ASIG5V.n9259 ASIG5V.n9258 0.0380882
R49165 ASIG5V.n9260 ASIG5V.n9259 0.0380882
R49166 ASIG5V.n11993 ASIG5V.n11992 0.0380882
R49167 ASIG5V.n11992 ASIG5V.n11991 0.0380882
R49168 ASIG5V.n11991 ASIG5V.n11990 0.0380882
R49169 ASIG5V.n11990 ASIG5V.n11989 0.0380882
R49170 ASIG5V.n11989 ASIG5V.n11988 0.0380882
R49171 ASIG5V.n11988 ASIG5V.n11987 0.0380882
R49172 ASIG5V.n11987 ASIG5V.n11986 0.0380882
R49173 ASIG5V.n11986 ASIG5V.n11985 0.0380882
R49174 ASIG5V.n11985 ASIG5V.n11984 0.0380882
R49175 ASIG5V.n11984 ASIG5V.n11983 0.0380882
R49176 ASIG5V.n11983 ASIG5V.n11982 0.0380882
R49177 ASIG5V.n11982 ASIG5V.n11981 0.0380882
R49178 ASIG5V.n11981 ASIG5V.n11980 0.0380882
R49179 ASIG5V.n11980 ASIG5V.n11979 0.0380882
R49180 ASIG5V.n11979 ASIG5V.n11978 0.0380882
R49181 ASIG5V.n11978 ASIG5V.n11977 0.0380882
R49182 ASIG5V.n11977 ASIG5V.n11976 0.0380882
R49183 ASIG5V.n11976 ASIG5V.n11975 0.0380882
R49184 ASIG5V.n11975 ASIG5V.n11974 0.0380882
R49185 ASIG5V.n11974 ASIG5V.n11973 0.0380882
R49186 ASIG5V.n11973 ASIG5V.n11972 0.0380882
R49187 ASIG5V.n11972 ASIG5V.n11971 0.0380882
R49188 ASIG5V.n11971 ASIG5V.n11970 0.0380882
R49189 ASIG5V.n11970 ASIG5V.n11969 0.0380882
R49190 ASIG5V.n11969 ASIG5V.n11968 0.0380882
R49191 ASIG5V.n11968 ASIG5V.n11967 0.0380882
R49192 ASIG5V.n11967 ASIG5V.n11966 0.0380882
R49193 ASIG5V.n11966 ASIG5V.n11965 0.0380882
R49194 ASIG5V.n11965 ASIG5V.n11964 0.0380882
R49195 ASIG5V.n11964 ASIG5V.n11963 0.0380882
R49196 ASIG5V.n9043 ASIG5V.n9042 0.0380882
R49197 ASIG5V.n9044 ASIG5V.n9043 0.0380882
R49198 ASIG5V.n9045 ASIG5V.n9044 0.0380882
R49199 ASIG5V.n9046 ASIG5V.n9045 0.0380882
R49200 ASIG5V.n9047 ASIG5V.n9046 0.0380882
R49201 ASIG5V.n9048 ASIG5V.n9047 0.0380882
R49202 ASIG5V.n9049 ASIG5V.n9048 0.0380882
R49203 ASIG5V.n9733 ASIG5V.n9732 0.0380882
R49204 ASIG5V.n9732 ASIG5V.n9731 0.0380882
R49205 ASIG5V.n9731 ASIG5V.n9730 0.0380882
R49206 ASIG5V.n9730 ASIG5V.n9729 0.0380882
R49207 ASIG5V.n9729 ASIG5V.n9728 0.0380882
R49208 ASIG5V.n9728 ASIG5V.n9727 0.0380882
R49209 ASIG5V.n9727 ASIG5V.n9726 0.0380882
R49210 ASIG5V.n9726 ASIG5V.n9725 0.0380882
R49211 ASIG5V.n9725 ASIG5V.n9724 0.0380882
R49212 ASIG5V.n9724 ASIG5V.n9723 0.0380882
R49213 ASIG5V.n9723 ASIG5V.n9722 0.0380882
R49214 ASIG5V.n9722 ASIG5V.n9721 0.0380882
R49215 ASIG5V.n9721 ASIG5V.n9720 0.0380882
R49216 ASIG5V.n9720 ASIG5V.n9719 0.0380882
R49217 ASIG5V.n9719 ASIG5V.n9718 0.0380882
R49218 ASIG5V.n9718 ASIG5V.n9717 0.0380882
R49219 ASIG5V.n9717 ASIG5V.n9716 0.0380882
R49220 ASIG5V.n9716 ASIG5V.n9715 0.0380882
R49221 ASIG5V.n9715 ASIG5V.n9714 0.0380882
R49222 ASIG5V.n9714 ASIG5V.n9713 0.0380882
R49223 ASIG5V.n9713 ASIG5V.n9712 0.0380882
R49224 ASIG5V.n9712 ASIG5V.n9711 0.0380882
R49225 ASIG5V.n9711 ASIG5V.n9710 0.0380882
R49226 ASIG5V.n9710 ASIG5V.n9709 0.0380882
R49227 ASIG5V.n9709 ASIG5V.n9708 0.0380882
R49228 ASIG5V.n9708 ASIG5V.n9707 0.0380882
R49229 ASIG5V.n9707 ASIG5V.n9706 0.0380882
R49230 ASIG5V.n9706 ASIG5V.n9705 0.0380882
R49231 ASIG5V.n9705 ASIG5V.n9704 0.0380882
R49232 ASIG5V.n9704 ASIG5V.n9703 0.0380882
R49233 ASIG5V.n9703 ASIG5V.n9702 0.0380882
R49234 ASIG5V.n9702 ASIG5V.n9701 0.0380882
R49235 ASIG5V.n9701 ASIG5V.n9700 0.0380882
R49236 ASIG5V.n9700 ASIG5V.n9699 0.0380882
R49237 ASIG5V.n9699 ASIG5V.n9698 0.0380882
R49238 ASIG5V.n9698 ASIG5V.n9697 0.0380882
R49239 ASIG5V.n9697 ASIG5V.n9696 0.0380882
R49240 ASIG5V.n9696 ASIG5V.n9695 0.0380882
R49241 ASIG5V.n9695 ASIG5V.n9694 0.0380882
R49242 ASIG5V.n9694 ASIG5V.n9693 0.0380882
R49243 ASIG5V.n9693 ASIG5V.n9692 0.0380882
R49244 ASIG5V.n9692 ASIG5V.n9691 0.0380882
R49245 ASIG5V.n9691 ASIG5V.n9690 0.0380882
R49246 ASIG5V.n9690 ASIG5V.n9689 0.0380882
R49247 ASIG5V.n9689 ASIG5V.n9688 0.0380882
R49248 ASIG5V.n9688 ASIG5V.n9687 0.0380882
R49249 ASIG5V.n9687 ASIG5V.n9686 0.0380882
R49250 ASIG5V.n9686 ASIG5V.n9685 0.0380882
R49251 ASIG5V.n9685 ASIG5V.n9684 0.0380882
R49252 ASIG5V.n9684 ASIG5V.n9683 0.0380882
R49253 ASIG5V.n9683 ASIG5V.n9682 0.0380882
R49254 ASIG5V.n9682 ASIG5V.n9681 0.0380882
R49255 ASIG5V.n9681 ASIG5V.n9680 0.0380882
R49256 ASIG5V.n9211 ASIG5V.n9210 0.0380882
R49257 ASIG5V.n9212 ASIG5V.n9211 0.0380882
R49258 ASIG5V.n9213 ASIG5V.n9212 0.0380882
R49259 ASIG5V.n9214 ASIG5V.n9213 0.0380882
R49260 ASIG5V.n9215 ASIG5V.n9214 0.0380882
R49261 ASIG5V.n9216 ASIG5V.n9215 0.0380882
R49262 ASIG5V.n9217 ASIG5V.n9216 0.0380882
R49263 ASIG5V.n9218 ASIG5V.n9217 0.0380882
R49264 ASIG5V.n9219 ASIG5V.n9218 0.0380882
R49265 ASIG5V.n9220 ASIG5V.n9219 0.0380882
R49266 ASIG5V.n9221 ASIG5V.n9220 0.0380882
R49267 ASIG5V.n9222 ASIG5V.n9221 0.0380882
R49268 ASIG5V.n9223 ASIG5V.n9222 0.0380882
R49269 ASIG5V.n9224 ASIG5V.n9223 0.0380882
R49270 ASIG5V.n9225 ASIG5V.n9224 0.0380882
R49271 ASIG5V.n9226 ASIG5V.n9225 0.0380882
R49272 ASIG5V.n9227 ASIG5V.n9226 0.0380882
R49273 ASIG5V.n9228 ASIG5V.n9227 0.0380882
R49274 ASIG5V.n9229 ASIG5V.n9228 0.0380882
R49275 ASIG5V.n9230 ASIG5V.n9229 0.0380882
R49276 ASIG5V.n9231 ASIG5V.n9230 0.0380882
R49277 ASIG5V.n9232 ASIG5V.n9231 0.0380882
R49278 ASIG5V.n9233 ASIG5V.n9232 0.0380882
R49279 ASIG5V.n9234 ASIG5V.n9233 0.0380882
R49280 ASIG5V.n9235 ASIG5V.n9234 0.0380882
R49281 ASIG5V.n9236 ASIG5V.n9235 0.0380882
R49282 ASIG5V.n11824 ASIG5V.n11823 0.0380882
R49283 ASIG5V.n11823 ASIG5V.n11822 0.0380882
R49284 ASIG5V.n11822 ASIG5V.n11821 0.0380882
R49285 ASIG5V.n11821 ASIG5V.n11820 0.0380882
R49286 ASIG5V.n11820 ASIG5V.n11819 0.0380882
R49287 ASIG5V.n11819 ASIG5V.n11818 0.0380882
R49288 ASIG5V.n11818 ASIG5V.n11817 0.0380882
R49289 ASIG5V.n11817 ASIG5V.n11816 0.0380882
R49290 ASIG5V.n11816 ASIG5V.n11815 0.0380882
R49291 ASIG5V.n11815 ASIG5V.n11814 0.0380882
R49292 ASIG5V.n11814 ASIG5V.n11813 0.0380882
R49293 ASIG5V.n11813 ASIG5V.n11812 0.0380882
R49294 ASIG5V.n11812 ASIG5V.n11811 0.0380882
R49295 ASIG5V.n11811 ASIG5V.n11810 0.0380882
R49296 ASIG5V.n11810 ASIG5V.n11809 0.0380882
R49297 ASIG5V.n11809 ASIG5V.n11808 0.0380882
R49298 ASIG5V.n11808 ASIG5V.n11807 0.0380882
R49299 ASIG5V.n11807 ASIG5V.n11806 0.0380882
R49300 ASIG5V.n11806 ASIG5V.n11805 0.0380882
R49301 ASIG5V.n11805 ASIG5V.n11804 0.0380882
R49302 ASIG5V.n11804 ASIG5V.n11803 0.0380882
R49303 ASIG5V.n11803 ASIG5V.n11802 0.0380882
R49304 ASIG5V.n11802 ASIG5V.n11801 0.0380882
R49305 ASIG5V.n11801 ASIG5V.n11800 0.0380882
R49306 ASIG5V.n11800 ASIG5V.n11799 0.0380882
R49307 ASIG5V.n11799 ASIG5V.n11798 0.0380882
R49308 ASIG5V.n11798 ASIG5V.n11797 0.0380882
R49309 ASIG5V.n11797 ASIG5V.n11796 0.0380882
R49310 ASIG5V.n11796 ASIG5V.n11795 0.0380882
R49311 ASIG5V.n11795 ASIG5V.n11794 0.0380882
R49312 ASIG5V.n9033 ASIG5V.n9032 0.0380882
R49313 ASIG5V.n9034 ASIG5V.n9033 0.0380882
R49314 ASIG5V.n9035 ASIG5V.n9034 0.0380882
R49315 ASIG5V.n9036 ASIG5V.n9035 0.0380882
R49316 ASIG5V.n9037 ASIG5V.n9036 0.0380882
R49317 ASIG5V.n9038 ASIG5V.n9037 0.0380882
R49318 ASIG5V.n9039 ASIG5V.n9038 0.0380882
R49319 ASIG5V.n9040 ASIG5V.n9039 0.0380882
R49320 ASIG5V.n9041 ASIG5V.n9040 0.0380882
R49321 ASIG5V.n9679 ASIG5V.n9678 0.0380882
R49322 ASIG5V.n9678 ASIG5V.n9677 0.0380882
R49323 ASIG5V.n9677 ASIG5V.n9676 0.0380882
R49324 ASIG5V.n9676 ASIG5V.n9675 0.0380882
R49325 ASIG5V.n9675 ASIG5V.n9674 0.0380882
R49326 ASIG5V.n9674 ASIG5V.n9673 0.0380882
R49327 ASIG5V.n9673 ASIG5V.n9672 0.0380882
R49328 ASIG5V.n9672 ASIG5V.n9671 0.0380882
R49329 ASIG5V.n9671 ASIG5V.n9670 0.0380882
R49330 ASIG5V.n9670 ASIG5V.n9669 0.0380882
R49331 ASIG5V.n9669 ASIG5V.n9668 0.0380882
R49332 ASIG5V.n9668 ASIG5V.n9667 0.0380882
R49333 ASIG5V.n9667 ASIG5V.n9666 0.0380882
R49334 ASIG5V.n9666 ASIG5V.n9665 0.0380882
R49335 ASIG5V.n9665 ASIG5V.n9664 0.0380882
R49336 ASIG5V.n9664 ASIG5V.n9663 0.0380882
R49337 ASIG5V.n9663 ASIG5V.n9662 0.0380882
R49338 ASIG5V.n9662 ASIG5V.n9661 0.0380882
R49339 ASIG5V.n9661 ASIG5V.n9660 0.0380882
R49340 ASIG5V.n9660 ASIG5V.n9659 0.0380882
R49341 ASIG5V.n9659 ASIG5V.n9658 0.0380882
R49342 ASIG5V.n9658 ASIG5V.n9657 0.0380882
R49343 ASIG5V.n9657 ASIG5V.n9656 0.0380882
R49344 ASIG5V.n9656 ASIG5V.n9655 0.0380882
R49345 ASIG5V.n9655 ASIG5V.n9654 0.0380882
R49346 ASIG5V.n9654 ASIG5V.n9653 0.0380882
R49347 ASIG5V.n9653 ASIG5V.n9652 0.0380882
R49348 ASIG5V.n9652 ASIG5V.n9651 0.0380882
R49349 ASIG5V.n9651 ASIG5V.n9650 0.0380882
R49350 ASIG5V.n9650 ASIG5V.n9649 0.0380882
R49351 ASIG5V.n9649 ASIG5V.n9648 0.0380882
R49352 ASIG5V.n9648 ASIG5V.n9647 0.0380882
R49353 ASIG5V.n9647 ASIG5V.n9646 0.0380882
R49354 ASIG5V.n9646 ASIG5V.n9645 0.0380882
R49355 ASIG5V.n9645 ASIG5V.n9644 0.0380882
R49356 ASIG5V.n9644 ASIG5V.n9643 0.0380882
R49357 ASIG5V.n9643 ASIG5V.n9642 0.0380882
R49358 ASIG5V.n9642 ASIG5V.n9641 0.0380882
R49359 ASIG5V.n9641 ASIG5V.n9640 0.0380882
R49360 ASIG5V.n9640 ASIG5V.n9639 0.0380882
R49361 ASIG5V.n9639 ASIG5V.n9638 0.0380882
R49362 ASIG5V.n9638 ASIG5V.n9637 0.0380882
R49363 ASIG5V.n9637 ASIG5V.n9636 0.0380882
R49364 ASIG5V.n9636 ASIG5V.n9635 0.0380882
R49365 ASIG5V.n9635 ASIG5V.n9634 0.0380882
R49366 ASIG5V.n9634 ASIG5V.n9633 0.0380882
R49367 ASIG5V.n9633 ASIG5V.n9632 0.0380882
R49368 ASIG5V.n9632 ASIG5V.n9631 0.0380882
R49369 ASIG5V.n9631 ASIG5V.n9630 0.0380882
R49370 ASIG5V.n9630 ASIG5V.n9629 0.0380882
R49371 ASIG5V.n9629 ASIG5V.n9628 0.0380882
R49372 ASIG5V.n9628 ASIG5V.n9627 0.0380882
R49373 ASIG5V.n9627 ASIG5V.n9626 0.0380882
R49374 ASIG5V.n9626 ASIG5V.n9625 0.0380882
R49375 ASIG5V.n9182 ASIG5V.n9181 0.0380882
R49376 ASIG5V.n9183 ASIG5V.n9182 0.0380882
R49377 ASIG5V.n9184 ASIG5V.n9183 0.0380882
R49378 ASIG5V.n9185 ASIG5V.n9184 0.0380882
R49379 ASIG5V.n9186 ASIG5V.n9185 0.0380882
R49380 ASIG5V.n9187 ASIG5V.n9186 0.0380882
R49381 ASIG5V.n9188 ASIG5V.n9187 0.0380882
R49382 ASIG5V.n9189 ASIG5V.n9188 0.0380882
R49383 ASIG5V.n9190 ASIG5V.n9189 0.0380882
R49384 ASIG5V.n9191 ASIG5V.n9190 0.0380882
R49385 ASIG5V.n9192 ASIG5V.n9191 0.0380882
R49386 ASIG5V.n9193 ASIG5V.n9192 0.0380882
R49387 ASIG5V.n9194 ASIG5V.n9193 0.0380882
R49388 ASIG5V.n9195 ASIG5V.n9194 0.0380882
R49389 ASIG5V.n9196 ASIG5V.n9195 0.0380882
R49390 ASIG5V.n9197 ASIG5V.n9196 0.0380882
R49391 ASIG5V.n9198 ASIG5V.n9197 0.0380882
R49392 ASIG5V.n9199 ASIG5V.n9198 0.0380882
R49393 ASIG5V.n9200 ASIG5V.n9199 0.0380882
R49394 ASIG5V.n9201 ASIG5V.n9200 0.0380882
R49395 ASIG5V.n9202 ASIG5V.n9201 0.0380882
R49396 ASIG5V.n9203 ASIG5V.n9202 0.0380882
R49397 ASIG5V.n9204 ASIG5V.n9203 0.0380882
R49398 ASIG5V.n9205 ASIG5V.n9204 0.0380882
R49399 ASIG5V.n9206 ASIG5V.n9205 0.0380882
R49400 ASIG5V.n9207 ASIG5V.n9206 0.0380882
R49401 ASIG5V.n9208 ASIG5V.n9207 0.0380882
R49402 ASIG5V.n9209 ASIG5V.n9208 0.0380882
R49403 ASIG5V.n10922 ASIG5V.n10921 0.0380882
R49404 ASIG5V.n10921 ASIG5V.n10920 0.0380882
R49405 ASIG5V.n10920 ASIG5V.n10919 0.0380882
R49406 ASIG5V.n10919 ASIG5V.n10918 0.0380882
R49407 ASIG5V.n10918 ASIG5V.n10917 0.0380882
R49408 ASIG5V.n10917 ASIG5V.n10916 0.0380882
R49409 ASIG5V.n10916 ASIG5V.n10915 0.0380882
R49410 ASIG5V.n10915 ASIG5V.n10914 0.0380882
R49411 ASIG5V.n10914 ASIG5V.n10913 0.0380882
R49412 ASIG5V.n10913 ASIG5V.n10912 0.0380882
R49413 ASIG5V.n10912 ASIG5V.n10911 0.0380882
R49414 ASIG5V.n10911 ASIG5V.n10910 0.0380882
R49415 ASIG5V.n10910 ASIG5V.n10909 0.0380882
R49416 ASIG5V.n10909 ASIG5V.n10908 0.0380882
R49417 ASIG5V.n10908 ASIG5V.n10907 0.0380882
R49418 ASIG5V.n10907 ASIG5V.n10906 0.0380882
R49419 ASIG5V.n10906 ASIG5V.n10905 0.0380882
R49420 ASIG5V.n10905 ASIG5V.n10904 0.0380882
R49421 ASIG5V.n10904 ASIG5V.n10903 0.0380882
R49422 ASIG5V.n10903 ASIG5V.n10902 0.0380882
R49423 ASIG5V.n10902 ASIG5V.n10901 0.0380882
R49424 ASIG5V.n10901 ASIG5V.n10900 0.0380882
R49425 ASIG5V.n10900 ASIG5V.n10899 0.0380882
R49426 ASIG5V.n10899 ASIG5V.n10898 0.0380882
R49427 ASIG5V.n10898 ASIG5V.n10897 0.0380882
R49428 ASIG5V.n10897 ASIG5V.n10896 0.0380882
R49429 ASIG5V.n10896 ASIG5V.n10895 0.0380882
R49430 ASIG5V.n10895 ASIG5V.n10894 0.0380882
R49431 ASIG5V.n10894 ASIG5V.n10893 0.0380882
R49432 ASIG5V.n10893 ASIG5V.n10892 0.0380882
R49433 ASIG5V.n10892 ASIG5V.n10891 0.0380882
R49434 ASIG5V.n9021 ASIG5V.n9020 0.0380882
R49435 ASIG5V.n9022 ASIG5V.n9021 0.0380882
R49436 ASIG5V.n9023 ASIG5V.n9022 0.0380882
R49437 ASIG5V.n9024 ASIG5V.n9023 0.0380882
R49438 ASIG5V.n9025 ASIG5V.n9024 0.0380882
R49439 ASIG5V.n9026 ASIG5V.n9025 0.0380882
R49440 ASIG5V.n9027 ASIG5V.n9026 0.0380882
R49441 ASIG5V.n9028 ASIG5V.n9027 0.0380882
R49442 ASIG5V.n9029 ASIG5V.n9028 0.0380882
R49443 ASIG5V.n9030 ASIG5V.n9029 0.0380882
R49444 ASIG5V.n9031 ASIG5V.n9030 0.0380882
R49445 ASIG5V.n2665 ASIG5V.n2664 0.0380882
R49446 ASIG5V.n2664 ASIG5V.n2663 0.0380882
R49447 ASIG5V.n2663 ASIG5V.n2662 0.0380882
R49448 ASIG5V.n2662 ASIG5V.n2661 0.0380882
R49449 ASIG5V.n2661 ASIG5V.n2660 0.0380882
R49450 ASIG5V.n2660 ASIG5V.n2659 0.0380882
R49451 ASIG5V.n2659 ASIG5V.n2658 0.0380882
R49452 ASIG5V.n2658 ASIG5V.n2657 0.0380882
R49453 ASIG5V.n2657 ASIG5V.n2656 0.0380882
R49454 ASIG5V.n2656 ASIG5V.n2655 0.0380882
R49455 ASIG5V.n2655 ASIG5V.n2654 0.0380882
R49456 ASIG5V.n2654 ASIG5V.n2653 0.0380882
R49457 ASIG5V.n2653 ASIG5V.n2652 0.0380882
R49458 ASIG5V.n2652 ASIG5V.n2651 0.0380882
R49459 ASIG5V.n2651 ASIG5V.n2650 0.0380882
R49460 ASIG5V.n2650 ASIG5V.n2649 0.0380882
R49461 ASIG5V.n2649 ASIG5V.n2648 0.0380882
R49462 ASIG5V.n2648 ASIG5V.n2647 0.0380882
R49463 ASIG5V.n2647 ASIG5V.n2646 0.0380882
R49464 ASIG5V.n2646 ASIG5V.n2645 0.0380882
R49465 ASIG5V.n2645 ASIG5V.n2644 0.0380882
R49466 ASIG5V.n2644 ASIG5V.n2643 0.0380882
R49467 ASIG5V.n2643 ASIG5V.n2642 0.0380882
R49468 ASIG5V.n2642 ASIG5V.n2641 0.0380882
R49469 ASIG5V.n2641 ASIG5V.n2640 0.0380882
R49470 ASIG5V.n2640 ASIG5V.n2639 0.0380882
R49471 ASIG5V.n2639 ASIG5V.n2638 0.0380882
R49472 ASIG5V.n2638 ASIG5V.n2637 0.0380882
R49473 ASIG5V.n2637 ASIG5V.n2636 0.0380882
R49474 ASIG5V.n2636 ASIG5V.n2635 0.0380882
R49475 ASIG5V.n2635 ASIG5V.n2634 0.0380882
R49476 ASIG5V.n2634 ASIG5V.n2633 0.0380882
R49477 ASIG5V.n2633 ASIG5V.n2632 0.0380882
R49478 ASIG5V.n631 ASIG5V.n630 0.0380882
R49479 ASIG5V.n632 ASIG5V.n631 0.0380882
R49480 ASIG5V.n633 ASIG5V.n632 0.0380882
R49481 ASIG5V.n634 ASIG5V.n633 0.0380882
R49482 ASIG5V.n635 ASIG5V.n634 0.0380882
R49483 ASIG5V.n636 ASIG5V.n635 0.0380882
R49484 ASIG5V.n637 ASIG5V.n636 0.0380882
R49485 ASIG5V.n638 ASIG5V.n637 0.0380882
R49486 ASIG5V.n639 ASIG5V.n638 0.0380882
R49487 ASIG5V.n640 ASIG5V.n639 0.0380882
R49488 ASIG5V.n641 ASIG5V.n640 0.0380882
R49489 ASIG5V.n642 ASIG5V.n641 0.0380882
R49490 ASIG5V.n643 ASIG5V.n642 0.0380882
R49491 ASIG5V.n644 ASIG5V.n643 0.0380882
R49492 ASIG5V.n645 ASIG5V.n644 0.0380882
R49493 ASIG5V.n646 ASIG5V.n645 0.0380882
R49494 ASIG5V.n10980 ASIG5V.n10979 0.0380882
R49495 ASIG5V.n10979 ASIG5V.n10978 0.0380882
R49496 ASIG5V.n10978 ASIG5V.n10977 0.0380882
R49497 ASIG5V.n10977 ASIG5V.n10976 0.0380882
R49498 ASIG5V.n10976 ASIG5V.n10975 0.0380882
R49499 ASIG5V.n10975 ASIG5V.n10974 0.0380882
R49500 ASIG5V.n10974 ASIG5V.n10973 0.0380882
R49501 ASIG5V.n10973 ASIG5V.n10972 0.0380882
R49502 ASIG5V.n10972 ASIG5V.n10971 0.0380882
R49503 ASIG5V.n10971 ASIG5V.n10970 0.0380882
R49504 ASIG5V.n10970 ASIG5V.n10969 0.0380882
R49505 ASIG5V.n10969 ASIG5V.n10968 0.0380882
R49506 ASIG5V.n10968 ASIG5V.n10967 0.0380882
R49507 ASIG5V.n10967 ASIG5V.n10966 0.0380882
R49508 ASIG5V.n10966 ASIG5V.n10965 0.0380882
R49509 ASIG5V.n10965 ASIG5V.n10964 0.0380882
R49510 ASIG5V.n10964 ASIG5V.n10963 0.0380882
R49511 ASIG5V.n10963 ASIG5V.n10962 0.0380882
R49512 ASIG5V.n10962 ASIG5V.n10961 0.0380882
R49513 ASIG5V.n10961 ASIG5V.n10960 0.0380882
R49514 ASIG5V.n10960 ASIG5V.n10959 0.0380882
R49515 ASIG5V.n10959 ASIG5V.n10958 0.0380882
R49516 ASIG5V.n10958 ASIG5V.n10957 0.0380882
R49517 ASIG5V.n10957 ASIG5V.n10956 0.0380882
R49518 ASIG5V.n10956 ASIG5V.n10955 0.0380882
R49519 ASIG5V.n10955 ASIG5V.n10954 0.0380882
R49520 ASIG5V.n10954 ASIG5V.n10953 0.0380882
R49521 ASIG5V.n10953 ASIG5V.n10952 0.0380882
R49522 ASIG5V.n10952 ASIG5V.n10951 0.0380882
R49523 ASIG5V.n10951 ASIG5V.n10950 0.0380882
R49524 ASIG5V.n10950 ASIG5V.n10949 0.0380882
R49525 ASIG5V.n10949 ASIG5V.n10948 0.0380882
R49526 ASIG5V.n10948 ASIG5V.n10947 0.0380882
R49527 ASIG5V.n10947 ASIG5V.n10946 0.0380882
R49528 ASIG5V.n10946 ASIG5V.n10945 0.0380882
R49529 ASIG5V.n10945 ASIG5V.n10944 0.0380882
R49530 ASIG5V.n10944 ASIG5V.n10943 0.0380882
R49531 ASIG5V.n10943 ASIG5V.n10942 0.0380882
R49532 ASIG5V.n10942 ASIG5V.n10941 0.0380882
R49533 ASIG5V.n10941 ASIG5V.n10940 0.0380882
R49534 ASIG5V.n10940 ASIG5V.n10939 0.0380882
R49535 ASIG5V.n10939 ASIG5V.n10938 0.0380882
R49536 ASIG5V.n10938 ASIG5V.n10937 0.0380882
R49537 ASIG5V.n10937 ASIG5V.n10936 0.0380882
R49538 ASIG5V.n10936 ASIG5V.n10935 0.0380882
R49539 ASIG5V.n10935 ASIG5V.n10934 0.0380882
R49540 ASIG5V.n10934 ASIG5V.n10933 0.0380882
R49541 ASIG5V.n10933 ASIG5V.n10932 0.0380882
R49542 ASIG5V.n10932 ASIG5V.n10931 0.0380882
R49543 ASIG5V.n10931 ASIG5V.n10930 0.0380882
R49544 ASIG5V.n8988 ASIG5V.n8987 0.0380882
R49545 ASIG5V.n8989 ASIG5V.n8988 0.0380882
R49546 ASIG5V.n8990 ASIG5V.n8989 0.0380882
R49547 ASIG5V.n8991 ASIG5V.n8990 0.0380882
R49548 ASIG5V.n8992 ASIG5V.n8991 0.0380882
R49549 ASIG5V.n8993 ASIG5V.n8992 0.0380882
R49550 ASIG5V.n8994 ASIG5V.n8993 0.0380882
R49551 ASIG5V.n8995 ASIG5V.n8994 0.0380882
R49552 ASIG5V.n8996 ASIG5V.n8995 0.0380882
R49553 ASIG5V.n8997 ASIG5V.n8996 0.0380882
R49554 ASIG5V.n8998 ASIG5V.n8997 0.0380882
R49555 ASIG5V.n8999 ASIG5V.n8998 0.0380882
R49556 ASIG5V.n9000 ASIG5V.n8999 0.0380882
R49557 ASIG5V.n9001 ASIG5V.n9000 0.0380882
R49558 ASIG5V.n9002 ASIG5V.n9001 0.0380882
R49559 ASIG5V.n9003 ASIG5V.n9002 0.0380882
R49560 ASIG5V.n9004 ASIG5V.n9003 0.0380882
R49561 ASIG5V.n9005 ASIG5V.n9004 0.0380882
R49562 ASIG5V.n9006 ASIG5V.n9005 0.0380882
R49563 ASIG5V.n9007 ASIG5V.n9006 0.0380882
R49564 ASIG5V.n9008 ASIG5V.n9007 0.0380882
R49565 ASIG5V.n9009 ASIG5V.n9008 0.0380882
R49566 ASIG5V.n9010 ASIG5V.n9009 0.0380882
R49567 ASIG5V.n9011 ASIG5V.n9010 0.0380882
R49568 ASIG5V.n9012 ASIG5V.n9011 0.0380882
R49569 ASIG5V.n9013 ASIG5V.n9012 0.0380882
R49570 ASIG5V.n9014 ASIG5V.n9013 0.0380882
R49571 ASIG5V.n9015 ASIG5V.n9014 0.0380882
R49572 ASIG5V.n9016 ASIG5V.n9015 0.0380882
R49573 ASIG5V.n9017 ASIG5V.n9016 0.0380882
R49574 ASIG5V.n9018 ASIG5V.n9017 0.0380882
R49575 ASIG5V.n9019 ASIG5V.n9018 0.0380882
R49576 ASIG5V.n11018 ASIG5V.n11017 0.0380882
R49577 ASIG5V.n11017 ASIG5V.n11016 0.0380882
R49578 ASIG5V.n11016 ASIG5V.n11015 0.0380882
R49579 ASIG5V.n11015 ASIG5V.n11014 0.0380882
R49580 ASIG5V.n11014 ASIG5V.n11013 0.0380882
R49581 ASIG5V.n11013 ASIG5V.n11012 0.0380882
R49582 ASIG5V.n11012 ASIG5V.n11011 0.0380882
R49583 ASIG5V.n11011 ASIG5V.n11010 0.0380882
R49584 ASIG5V.n11010 ASIG5V.n11009 0.0380882
R49585 ASIG5V.n11009 ASIG5V.n11008 0.0380882
R49586 ASIG5V.n11008 ASIG5V.n11007 0.0380882
R49587 ASIG5V.n11007 ASIG5V.n11006 0.0380882
R49588 ASIG5V.n11006 ASIG5V.n11005 0.0380882
R49589 ASIG5V.n11005 ASIG5V.n11004 0.0380882
R49590 ASIG5V.n11004 ASIG5V.n11003 0.0380882
R49591 ASIG5V.n11003 ASIG5V.n11002 0.0380882
R49592 ASIG5V.n11002 ASIG5V.n11001 0.0380882
R49593 ASIG5V.n11001 ASIG5V.n11000 0.0380882
R49594 ASIG5V.n11000 ASIG5V.n10999 0.0380882
R49595 ASIG5V.n10999 ASIG5V.n10998 0.0380882
R49596 ASIG5V.n10998 ASIG5V.n10997 0.0380882
R49597 ASIG5V.n10997 ASIG5V.n10996 0.0380882
R49598 ASIG5V.n10996 ASIG5V.n10995 0.0380882
R49599 ASIG5V.n10995 ASIG5V.n10994 0.0380882
R49600 ASIG5V.n10994 ASIG5V.n10993 0.0380882
R49601 ASIG5V.n10993 ASIG5V.n10992 0.0380882
R49602 ASIG5V.n10992 ASIG5V.n10991 0.0380882
R49603 ASIG5V.n10991 ASIG5V.n10990 0.0380882
R49604 ASIG5V.n10990 ASIG5V.n10989 0.0380882
R49605 ASIG5V.n10989 ASIG5V.n10988 0.0380882
R49606 ASIG5V.n10988 ASIG5V.n10987 0.0380882
R49607 ASIG5V.n10987 ASIG5V.n10986 0.0380882
R49608 ASIG5V.n10986 ASIG5V.n10985 0.0380882
R49609 ASIG5V.n9092 ASIG5V.n9091 0.0380882
R49610 ASIG5V.n9093 ASIG5V.n9092 0.0380882
R49611 ASIG5V.n9094 ASIG5V.n9093 0.0380882
R49612 ASIG5V.n9095 ASIG5V.n9094 0.0380882
R49613 ASIG5V.n9096 ASIG5V.n9095 0.0380882
R49614 ASIG5V.n9097 ASIG5V.n9096 0.0380882
R49615 ASIG5V.n9098 ASIG5V.n9097 0.0380882
R49616 ASIG5V.n9099 ASIG5V.n9098 0.0380882
R49617 ASIG5V.n9100 ASIG5V.n9099 0.0380882
R49618 ASIG5V.n9101 ASIG5V.n9100 0.0380882
R49619 ASIG5V.n9102 ASIG5V.n9101 0.0380882
R49620 ASIG5V.n9103 ASIG5V.n9102 0.0380882
R49621 ASIG5V.n9104 ASIG5V.n9103 0.0380882
R49622 ASIG5V.n9105 ASIG5V.n9104 0.0380882
R49623 ASIG5V.n9106 ASIG5V.n9105 0.0380882
R49624 ASIG5V.n9569 ASIG5V.n9568 0.0380882
R49625 ASIG5V.n9568 ASIG5V.n9567 0.0380882
R49626 ASIG5V.n9567 ASIG5V.n9566 0.0380882
R49627 ASIG5V.n9566 ASIG5V.n9565 0.0380882
R49628 ASIG5V.n9565 ASIG5V.n9564 0.0380882
R49629 ASIG5V.n9564 ASIG5V.n9563 0.0380882
R49630 ASIG5V.n9563 ASIG5V.n9562 0.0380882
R49631 ASIG5V.n9562 ASIG5V.n9561 0.0380882
R49632 ASIG5V.n9561 ASIG5V.n9560 0.0380882
R49633 ASIG5V.n9560 ASIG5V.n9559 0.0380882
R49634 ASIG5V.n9559 ASIG5V.n9558 0.0380882
R49635 ASIG5V.n9558 ASIG5V.n9557 0.0380882
R49636 ASIG5V.n9557 ASIG5V.n9556 0.0380882
R49637 ASIG5V.n9556 ASIG5V.n9555 0.0380882
R49638 ASIG5V.n9555 ASIG5V.n9554 0.0380882
R49639 ASIG5V.n9554 ASIG5V.n9553 0.0380882
R49640 ASIG5V.n9553 ASIG5V.n9552 0.0380882
R49641 ASIG5V.n9552 ASIG5V.n9551 0.0380882
R49642 ASIG5V.n9551 ASIG5V.n9550 0.0380882
R49643 ASIG5V.n9550 ASIG5V.n9549 0.0380882
R49644 ASIG5V.n9549 ASIG5V.n9548 0.0380882
R49645 ASIG5V.n9548 ASIG5V.n9547 0.0380882
R49646 ASIG5V.n9547 ASIG5V.n9546 0.0380882
R49647 ASIG5V.n9546 ASIG5V.n9545 0.0380882
R49648 ASIG5V.n9545 ASIG5V.n9544 0.0380882
R49649 ASIG5V.n9544 ASIG5V.n9543 0.0380882
R49650 ASIG5V.n9543 ASIG5V.n9542 0.0380882
R49651 ASIG5V.n9542 ASIG5V.n9541 0.0380882
R49652 ASIG5V.n9541 ASIG5V.n9540 0.0380882
R49653 ASIG5V.n9540 ASIG5V.n9539 0.0380882
R49654 ASIG5V.n9539 ASIG5V.n9538 0.0380882
R49655 ASIG5V.n9538 ASIG5V.n9537 0.0380882
R49656 ASIG5V.n9537 ASIG5V.n9536 0.0380882
R49657 ASIG5V.n9536 ASIG5V.n9535 0.0380882
R49658 ASIG5V.n9535 ASIG5V.n9534 0.0380882
R49659 ASIG5V.n9534 ASIG5V.n9533 0.0380882
R49660 ASIG5V.n9533 ASIG5V.n9532 0.0380882
R49661 ASIG5V.n9532 ASIG5V.n9531 0.0380882
R49662 ASIG5V.n9531 ASIG5V.n9530 0.0380882
R49663 ASIG5V.n9530 ASIG5V.n9529 0.0380882
R49664 ASIG5V.n9529 ASIG5V.n9528 0.0380882
R49665 ASIG5V.n9528 ASIG5V.n9527 0.0380882
R49666 ASIG5V.n9527 ASIG5V.n9526 0.0380882
R49667 ASIG5V.n9526 ASIG5V.n9525 0.0380882
R49668 ASIG5V.n9525 ASIG5V.n9524 0.0380882
R49669 ASIG5V.n9524 ASIG5V.n9523 0.0380882
R49670 ASIG5V.n9523 ASIG5V.n9522 0.0380882
R49671 ASIG5V.n9522 ASIG5V.n9521 0.0380882
R49672 ASIG5V.n9521 ASIG5V.n9520 0.0380882
R49673 ASIG5V.n9520 ASIG5V.n9519 0.0380882
R49674 ASIG5V.n9519 ASIG5V.n9518 0.0380882
R49675 ASIG5V.n9518 ASIG5V.n9517 0.0380882
R49676 ASIG5V.n9517 ASIG5V.n9516 0.0380882
R49677 ASIG5V.n9123 ASIG5V.n9122 0.0380882
R49678 ASIG5V.n9124 ASIG5V.n9123 0.0380882
R49679 ASIG5V.n9125 ASIG5V.n9124 0.0380882
R49680 ASIG5V.n9126 ASIG5V.n9125 0.0380882
R49681 ASIG5V.n9127 ASIG5V.n9126 0.0380882
R49682 ASIG5V.n9128 ASIG5V.n9127 0.0380882
R49683 ASIG5V.n9129 ASIG5V.n9128 0.0380882
R49684 ASIG5V.n9130 ASIG5V.n9129 0.0380882
R49685 ASIG5V.n9131 ASIG5V.n9130 0.0380882
R49686 ASIG5V.n9132 ASIG5V.n9131 0.0380882
R49687 ASIG5V.n9133 ASIG5V.n9132 0.0380882
R49688 ASIG5V.n9134 ASIG5V.n9133 0.0380882
R49689 ASIG5V.n9135 ASIG5V.n9134 0.0380882
R49690 ASIG5V.n9136 ASIG5V.n9135 0.0380882
R49691 ASIG5V.n9137 ASIG5V.n9136 0.0380882
R49692 ASIG5V.n9138 ASIG5V.n9137 0.0380882
R49693 ASIG5V.n9139 ASIG5V.n9138 0.0380882
R49694 ASIG5V.n9140 ASIG5V.n9139 0.0380882
R49695 ASIG5V.n9141 ASIG5V.n9140 0.0380882
R49696 ASIG5V.n9142 ASIG5V.n9141 0.0380882
R49697 ASIG5V.n9143 ASIG5V.n9142 0.0380882
R49698 ASIG5V.n9144 ASIG5V.n9143 0.0380882
R49699 ASIG5V.n9145 ASIG5V.n9144 0.0380882
R49700 ASIG5V.n9146 ASIG5V.n9145 0.0380882
R49701 ASIG5V.n9147 ASIG5V.n9146 0.0380882
R49702 ASIG5V.n9148 ASIG5V.n9147 0.0380882
R49703 ASIG5V.n9149 ASIG5V.n9148 0.0380882
R49704 ASIG5V.n9150 ASIG5V.n9149 0.0380882
R49705 ASIG5V.n9151 ASIG5V.n9150 0.0380882
R49706 ASIG5V.n1204 ASIG5V.n1203 0.0380882
R49707 ASIG5V.n1203 ASIG5V.n1202 0.0380882
R49708 ASIG5V.n1202 ASIG5V.n1201 0.0380882
R49709 ASIG5V.n1201 ASIG5V.n1200 0.0380882
R49710 ASIG5V.n1200 ASIG5V.n1199 0.0380882
R49711 ASIG5V.n1199 ASIG5V.n1198 0.0380882
R49712 ASIG5V.n1198 ASIG5V.n1197 0.0380882
R49713 ASIG5V.n1197 ASIG5V.n1196 0.0380882
R49714 ASIG5V.n1196 ASIG5V.n1195 0.0380882
R49715 ASIG5V.n1195 ASIG5V.n1194 0.0380882
R49716 ASIG5V.n1194 ASIG5V.n1193 0.0380882
R49717 ASIG5V.n1193 ASIG5V.n1192 0.0380882
R49718 ASIG5V.n1192 ASIG5V.n1191 0.0380882
R49719 ASIG5V.n1191 ASIG5V.n1190 0.0380882
R49720 ASIG5V.n1190 ASIG5V.n1189 0.0380882
R49721 ASIG5V.n1189 ASIG5V.n1188 0.0380882
R49722 ASIG5V.n1188 ASIG5V.n1187 0.0380882
R49723 ASIG5V.n1187 ASIG5V.n1186 0.0380882
R49724 ASIG5V.n1186 ASIG5V.n1185 0.0380882
R49725 ASIG5V.n1185 ASIG5V.n1184 0.0380882
R49726 ASIG5V.n1184 ASIG5V.n1183 0.0380882
R49727 ASIG5V.n1183 ASIG5V.n1182 0.0380882
R49728 ASIG5V.n1182 ASIG5V.n1181 0.0380882
R49729 ASIG5V.n1181 ASIG5V.n1180 0.0380882
R49730 ASIG5V.n1180 ASIG5V.n1179 0.0380882
R49731 ASIG5V.n1179 ASIG5V.n1178 0.0380882
R49732 ASIG5V.n1178 ASIG5V.n1177 0.0380882
R49733 ASIG5V.n1177 ASIG5V.n1176 0.0380882
R49734 ASIG5V.n1176 ASIG5V.n1175 0.0380882
R49735 ASIG5V.n1175 ASIG5V.n1174 0.0380882
R49736 ASIG5V.n1174 ASIG5V.n1173 0.0380882
R49737 ASIG5V.n1173 ASIG5V.n1172 0.0380882
R49738 ASIG5V.n1172 ASIG5V.n1171 0.0380882
R49739 ASIG5V.n1171 ASIG5V.n1170 0.0380882
R49740 ASIG5V.n1170 ASIG5V.n1169 0.0380882
R49741 ASIG5V.n1169 ASIG5V.n1168 0.0380882
R49742 ASIG5V.n1168 ASIG5V.n1167 0.0380882
R49743 ASIG5V.n1167 ASIG5V.n1166 0.0380882
R49744 ASIG5V.n1166 ASIG5V.n1165 0.0380882
R49745 ASIG5V.n1165 ASIG5V.n1164 0.0380882
R49746 ASIG5V.n1164 ASIG5V.n1163 0.0380882
R49747 ASIG5V.n1163 ASIG5V.n1162 0.0380882
R49748 ASIG5V.n1162 ASIG5V.n1161 0.0380882
R49749 ASIG5V.n1161 ASIG5V.n1160 0.0380882
R49750 ASIG5V.n1160 ASIG5V.n1159 0.0380882
R49751 ASIG5V.n1159 ASIG5V.n1158 0.0380882
R49752 ASIG5V.n1158 ASIG5V.n1157 0.0380882
R49753 ASIG5V.n1157 ASIG5V.n1156 0.0380882
R49754 ASIG5V.n1156 ASIG5V.n1155 0.0380882
R49755 ASIG5V.n1155 ASIG5V.n1154 0.0380882
R49756 ASIG5V.n1154 ASIG5V.n1153 0.0380882
R49757 ASIG5V.n1153 ASIG5V.n1152 0.0380882
R49758 ASIG5V.n1152 ASIG5V.n1151 0.0380882
R49759 ASIG5V.n1030 ASIG5V.n1029 0.0380882
R49760 ASIG5V.n1031 ASIG5V.n1030 0.0380882
R49761 ASIG5V.n1032 ASIG5V.n1031 0.0380882
R49762 ASIG5V.n1033 ASIG5V.n1032 0.0380882
R49763 ASIG5V.n1034 ASIG5V.n1033 0.0380882
R49764 ASIG5V.n1035 ASIG5V.n1034 0.0380882
R49765 ASIG5V.n1036 ASIG5V.n1035 0.0380882
R49766 ASIG5V.n1037 ASIG5V.n1036 0.0380882
R49767 ASIG5V.n1038 ASIG5V.n1037 0.0380882
R49768 ASIG5V.n1039 ASIG5V.n1038 0.0380882
R49769 ASIG5V.n1040 ASIG5V.n1039 0.0380882
R49770 ASIG5V.n1041 ASIG5V.n1040 0.0380882
R49771 ASIG5V.n1042 ASIG5V.n1041 0.0380882
R49772 ASIG5V.n1043 ASIG5V.n1042 0.0380882
R49773 ASIG5V.n1044 ASIG5V.n1043 0.0380882
R49774 ASIG5V.n1045 ASIG5V.n1044 0.0380882
R49775 ASIG5V.n1046 ASIG5V.n1045 0.0380882
R49776 ASIG5V.n1047 ASIG5V.n1046 0.0380882
R49777 ASIG5V.n1048 ASIG5V.n1047 0.0380882
R49778 ASIG5V.n1049 ASIG5V.n1048 0.0380882
R49779 ASIG5V.n1050 ASIG5V.n1049 0.0380882
R49780 ASIG5V.n1051 ASIG5V.n1050 0.0380882
R49781 ASIG5V.n1052 ASIG5V.n1051 0.0380882
R49782 ASIG5V.n1053 ASIG5V.n1052 0.0380882
R49783 ASIG5V.n1054 ASIG5V.n1053 0.0380882
R49784 ASIG5V.n1055 ASIG5V.n1054 0.0380882
R49785 ASIG5V.n1056 ASIG5V.n1055 0.0380882
R49786 ASIG5V.n1057 ASIG5V.n1056 0.0380882
R49787 ASIG5V.n1058 ASIG5V.n1057 0.0380882
R49788 ASIG5V.n1062 ASIG5V.n1061 0.03245
R49789 ASIG5V.n1061 ASIG5V.n1060 0.03245
R49790 ASIG5V.n1028 ASIG5V.n1027 0.03245
R49791 ASIG5V.n1027 ASIG5V.n1026 0.03245
R49792 ASIG5V.n1024 ASIG5V.n1023 0.03245
R49793 ASIG5V.n1021 ASIG5V.n1020 0.03245
R49794 ASIG5V.n1020 ASIG5V.n1019 0.03245
R49795 ASIG5V.n1017 ASIG5V.n1016 0.03245
R49796 ASIG5V.n1016 ASIG5V.n1015 0.03245
R49797 ASIG5V.n1013 ASIG5V.n1012 0.03245
R49798 ASIG5V.n1012 ASIG5V.n1011 0.03245
R49799 ASIG5V.n1009 ASIG5V.n1008 0.03245
R49800 ASIG5V.n1008 ASIG5V.n1007 0.03245
R49801 ASIG5V.n1005 ASIG5V.n1004 0.03245
R49802 ASIG5V.n1004 ASIG5V.n1003 0.03245
R49803 ASIG5V.n1001 ASIG5V.n1000 0.03245
R49804 ASIG5V.n998 ASIG5V.n997 0.03245
R49805 ASIG5V.n997 ASIG5V.n996 0.03245
R49806 ASIG5V.n994 ASIG5V.n993 0.03245
R49807 ASIG5V.n993 ASIG5V.n992 0.03245
R49808 ASIG5V.n990 ASIG5V.n989 0.03245
R49809 ASIG5V.n989 ASIG5V.n988 0.03245
R49810 ASIG5V.n986 ASIG5V.n985 0.03245
R49811 ASIG5V.n985 ASIG5V.n984 0.03245
R49812 ASIG5V.n982 ASIG5V.n981 0.03245
R49813 ASIG5V.n979 ASIG5V.n978 0.03245
R49814 ASIG5V.n978 ASIG5V.n977 0.03245
R49815 ASIG5V.n9373 ASIG5V.n9372 0.03245
R49816 ASIG5V.n9376 ASIG5V.n9375 0.03245
R49817 ASIG5V.n9377 ASIG5V.n9376 0.03245
R49818 ASIG5V.n9380 ASIG5V.n9379 0.03245
R49819 ASIG5V.n9381 ASIG5V.n9380 0.03245
R49820 ASIG5V.n9384 ASIG5V.n9383 0.03245
R49821 ASIG5V.n9385 ASIG5V.n9384 0.03245
R49822 ASIG5V.n9388 ASIG5V.n9387 0.03245
R49823 ASIG5V.n9391 ASIG5V.n9390 0.03245
R49824 ASIG5V.n9392 ASIG5V.n9391 0.03245
R49825 ASIG5V.n9395 ASIG5V.n9394 0.03245
R49826 ASIG5V.n9396 ASIG5V.n9395 0.03245
R49827 ASIG5V.n9399 ASIG5V.n9398 0.03245
R49828 ASIG5V.n9400 ASIG5V.n9399 0.03245
R49829 ASIG5V.n9403 ASIG5V.n9402 0.03245
R49830 ASIG5V.n9404 ASIG5V.n9403 0.03245
R49831 ASIG5V.n9407 ASIG5V.n9406 0.03245
R49832 ASIG5V.n9410 ASIG5V.n9409 0.03245
R49833 ASIG5V.n9411 ASIG5V.n9410 0.03245
R49834 ASIG5V.n9414 ASIG5V.n9413 0.03245
R49835 ASIG5V.n9415 ASIG5V.n9414 0.03245
R49836 ASIG5V.n9418 ASIG5V.n9417 0.03245
R49837 ASIG5V.n9419 ASIG5V.n9418 0.03245
R49838 ASIG5V.n9422 ASIG5V.n9421 0.03245
R49839 ASIG5V.n9423 ASIG5V.n9422 0.03245
R49840 ASIG5V.n9426 ASIG5V.n9425 0.03245
R49841 ASIG5V.n9427 ASIG5V.n9426 0.03245
R49842 ASIG5V.n1023 ASIG5V.n1022 0.031775
R49843 ASIG5V.n10750 ASIG5V.n9624 0.0317353
R49844 ASIG5V.n2489 ASIG5V.n1259 0.0317353
R49845 ASIG5V.n2485 ASIG5V.n1314 0.0317353
R49846 ASIG5V.n2481 ASIG5V.n1368 0.0317353
R49847 ASIG5V.n2476 ASIG5V.n1728 0.0317353
R49848 ASIG5V.n2472 ASIG5V.n1780 0.0317353
R49849 ASIG5V.n2468 ASIG5V.n1830 0.0317353
R49850 ASIG5V.n2186 ASIG5V.n1879 0.0317353
R49851 ASIG5V.n2182 ASIG5V.n1926 0.0317353
R49852 ASIG5V.n2177 ASIG5V.n1972 0.0317353
R49853 ASIG5V.n5667 ASIG5V.n5666 0.0317353
R49854 ASIG5V.n5968 ASIG5V.n5967 0.0317353
R49855 ASIG5V.n450 ASIG5V.n449 0.0317353
R49856 ASIG5V.n7044 ASIG5V.n7043 0.0317353
R49857 ASIG5V.n6765 ASIG5V.n6764 0.0317353
R49858 ASIG5V.n13603 ASIG5V.n13602 0.0317353
R49859 ASIG5V.n13348 ASIG5V.n13347 0.0317353
R49860 ASIG5V.n7515 ASIG5V.n7514 0.0317353
R49861 ASIG5V.n7932 ASIG5V.n7931 0.0317353
R49862 ASIG5V.n10714 ASIG5V.n10713 0.0317353
R49863 ASIG5V.n10718 ASIG5V.n10667 0.0317353
R49864 ASIG5V.n10722 ASIG5V.n10620 0.0317353
R49865 ASIG5V.n10728 ASIG5V.n10292 0.0317353
R49866 ASIG5V.n10732 ASIG5V.n10242 0.0317353
R49867 ASIG5V.n10736 ASIG5V.n10191 0.0317353
R49868 ASIG5V.n10741 ASIG5V.n9733 0.0317353
R49869 ASIG5V.n10745 ASIG5V.n9679 0.0317353
R49870 ASIG5V.n10754 ASIG5V.n9569 0.0317353
R49871 ASIG5V.n2493 ASIG5V.n1204 0.0317353
R49872 ASIG5V.n981 ASIG5V.n980 0.031325
R49873 ASIG5V.n9387 ASIG5V.n9386 0.030875
R49874 ASIG5V.n9408 ASIG5V.n9407 0.030875
R49875 ASIG5V.n1002 ASIG5V.n1001 0.030425
R49876 ASIG5V.n1000 ASIG5V.n999 0.028625
R49877 ASIG5V.n736 ASIG5V.n735 0.0284039
R49878 ASIG5V.n735 ASIG5V.n734 0.0284039
R49879 ASIG5V.n732 ASIG5V.n731 0.0284039
R49880 ASIG5V.n731 ASIG5V.n730 0.0284039
R49881 ASIG5V.n728 ASIG5V.n727 0.0284039
R49882 ASIG5V.n725 ASIG5V.n724 0.0284039
R49883 ASIG5V.n724 ASIG5V.n723 0.0284039
R49884 ASIG5V.n721 ASIG5V.n720 0.0284039
R49885 ASIG5V.n720 ASIG5V.n719 0.0284039
R49886 ASIG5V.n717 ASIG5V.n716 0.0284039
R49887 ASIG5V.n716 ASIG5V.n715 0.0284039
R49888 ASIG5V.n713 ASIG5V.n712 0.0284039
R49889 ASIG5V.n712 ASIG5V.n711 0.0284039
R49890 ASIG5V.n709 ASIG5V.n708 0.0284039
R49891 ASIG5V.n708 ASIG5V.n707 0.0284039
R49892 ASIG5V.n705 ASIG5V.n704 0.0284039
R49893 ASIG5V.n9063 ASIG5V.n9062 0.0284039
R49894 ASIG5V.n9066 ASIG5V.n9065 0.0284039
R49895 ASIG5V.n9067 ASIG5V.n9066 0.0284039
R49896 ASIG5V.n9070 ASIG5V.n9069 0.0284039
R49897 ASIG5V.n9071 ASIG5V.n9070 0.0284039
R49898 ASIG5V.n9074 ASIG5V.n9073 0.0284039
R49899 ASIG5V.n9077 ASIG5V.n9076 0.0284039
R49900 ASIG5V.n9078 ASIG5V.n9077 0.0284039
R49901 ASIG5V.n9081 ASIG5V.n9080 0.0284039
R49902 ASIG5V.n9082 ASIG5V.n9081 0.0284039
R49903 ASIG5V.n9085 ASIG5V.n9084 0.0284039
R49904 ASIG5V.n9086 ASIG5V.n9085 0.0284039
R49905 ASIG5V.n9089 ASIG5V.n9088 0.0284039
R49906 ASIG5V.n9090 ASIG5V.n9089 0.0284039
R49907 ASIG5V.n9109 ASIG5V.n9108 0.0284039
R49908 ASIG5V.n9110 ASIG5V.n9109 0.0284039
R49909 ASIG5V.n9389 ASIG5V.n9388 0.028175
R49910 ASIG5V.n9406 ASIG5V.n9405 0.028175
R49911 ASIG5V.n727 ASIG5V.n726 0.0278144
R49912 ASIG5V.n983 ASIG5V.n982 0.027725
R49913 ASIG5V.n1025 ASIG5V.n1024 0.027275
R49914 ASIG5V.n2194 ASIG5V.n2193 0.0272535
R49915 ASIG5V.n9075 ASIG5V.n9074 0.0270284
R49916 ASIG5V.n2215 ASIG5V.n2214 0.0269689
R49917 ASIG5V.n2205 ASIG5V.n2204 0.0269689
R49918 ASIG5V.n1393 ASIG5V.n1392 0.0269689
R49919 ASIG5V.n1384 ASIG5V.n1383 0.0269689
R49920 ASIG5V.n13185 ASIG5V.n13184 0.0269689
R49921 ASIG5V.n12859 ASIG5V.n12858 0.0269689
R49922 ASIG5V.n10484 ASIG5V.n10483 0.0269689
R49923 ASIG5V.n12805 ASIG5V.n12804 0.0269689
R49924 ASIG5V.n10515 ASIG5V.n10514 0.0269689
R49925 ASIG5V.n7141 ASIG5V.n7140 0.0269689
R49926 ASIG5V.n12775 ASIG5V.n12774 0.0269689
R49927 ASIG5V.n10544 ASIG5V.n10543 0.0269689
R49928 ASIG5V.n10560 ASIG5V.n10559 0.0269689
R49929 ASIG5V.n706 ASIG5V.n705 0.0266354
R49930 ASIG5V.n11412 ASIG5V.n11411 0.0265863
R49931 ASIG5V.n1019 ASIG5V.n1018 0.025925
R49932 ASIG5V.n11482 ASIG5V.n11481 0.0259201
R49933 ASIG5V.n9420 ASIG5V.n9180 0.0259118
R49934 ASIG5V.n1025 ASIG5V.n776 0.0259118
R49935 ASIG5V.n1022 ASIG5V.n805 0.0259118
R49936 ASIG5V.n1018 ASIG5V.n832 0.0259118
R49937 ASIG5V.n1014 ASIG5V.n857 0.0259118
R49938 ASIG5V.n1010 ASIG5V.n879 0.0259118
R49939 ASIG5V.n1006 ASIG5V.n899 0.0259118
R49940 ASIG5V.n1002 ASIG5V.n917 0.0259118
R49941 ASIG5V.n999 ASIG5V.n932 0.0259118
R49942 ASIG5V.n995 ASIG5V.n945 0.0259118
R49943 ASIG5V.n991 ASIG5V.n956 0.0259118
R49944 ASIG5V.n987 ASIG5V.n964 0.0259118
R49945 ASIG5V.n983 ASIG5V.n970 0.0259118
R49946 ASIG5V.n980 ASIG5V.n973 0.0259118
R49947 ASIG5V.n976 ASIG5V.n974 0.0259118
R49948 ASIG5V.n9374 ASIG5V.n9371 0.0259118
R49949 ASIG5V.n9378 ASIG5V.n9368 0.0259118
R49950 ASIG5V.n9382 ASIG5V.n9363 0.0259118
R49951 ASIG5V.n9386 ASIG5V.n9355 0.0259118
R49952 ASIG5V.n9389 ASIG5V.n9345 0.0259118
R49953 ASIG5V.n9393 ASIG5V.n9333 0.0259118
R49954 ASIG5V.n9397 ASIG5V.n9318 0.0259118
R49955 ASIG5V.n9401 ASIG5V.n9301 0.0259118
R49956 ASIG5V.n9405 ASIG5V.n9282 0.0259118
R49957 ASIG5V.n9408 ASIG5V.n9260 0.0259118
R49958 ASIG5V.n9412 ASIG5V.n9236 0.0259118
R49959 ASIG5V.n9416 ASIG5V.n9209 0.0259118
R49960 ASIG5V.n9424 ASIG5V.n9151 0.0259118
R49961 ASIG5V.n1059 ASIG5V.n1058 0.0259118
R49962 ASIG5V.n977 ASIG5V.n976 0.025475
R49963 ASIG5V.n9425 ASIG5V.n9424 0.025475
R49964 ASIG5V.n1149 ASIG5V.n1148 0.0251375
R49965 ASIG5V.n2816 ASIG5V.n2815 0.0251375
R49966 ASIG5V.n9514 ASIG5V.n9513 0.0251375
R49967 ASIG5V.n11093 ASIG5V.n11092 0.0251375
R49968 ASIG5V.n10889 ASIG5V.n10888 0.0251375
R49969 ASIG5V.n2630 ASIG5V.n2629 0.0251375
R49970 ASIG5V.n9383 ASIG5V.n9382 0.025025
R49971 ASIG5V.n9412 ASIG5V.n9411 0.025025
R49972 ASIG5V.n9073 ASIG5V.n9072 0.0246703
R49973 ASIG5V.n1006 ASIG5V.n1005 0.024575
R49974 ASIG5V.n13154 ASIG5V.n13153 0.0243788
R49975 ASIG5V.n12888 ASIG5V.n12887 0.0243788
R49976 ASIG5V.n7177 ASIG5V.n7176 0.0243788
R49977 ASIG5V.n10315 ASIG5V.n10314 0.0243788
R49978 ASIG5V.n10323 ASIG5V.n10322 0.0243788
R49979 ASIG5V.n13038 ASIG5V.n13037 0.0243788
R49980 ASIG5V.n10328 ASIG5V.n10327 0.0243788
R49981 ASIG5V.n10336 ASIG5V.n10335 0.0243788
R49982 ASIG5V.n1481 ASIG5V.n1480 0.0243788
R49983 ASIG5V.n2261 ASIG5V.n2260 0.0243788
R49984 ASIG5V.n13011 ASIG5V.n13010 0.0243788
R49985 ASIG5V.n12985 ASIG5V.n12984 0.0243788
R49986 ASIG5V.n9796 ASIG5V.n9795 0.0243788
R49987 ASIG5V.n9804 ASIG5V.n9803 0.0243788
R49988 ASIG5V.n1432 ASIG5V.n1431 0.0243788
R49989 ASIG5V.n729 ASIG5V.n728 0.0238843
R49990 ASIG5V.n996 ASIG5V.n995 0.022775
R49991 ASIG5V.n723 ASIG5V.n722 0.0227052
R49992 ASIG5V.n9974 ASIG5V 0.0226037
R49993 ASIG5V ASIG5V.n13126 0.0226037
R49994 ASIG5V.n13047 ASIG5V 0.0226037
R49995 ASIG5V ASIG5V.n12993 0.0226037
R49996 ASIG5V.n9393 ASIG5V.n9392 0.022325
R49997 ASIG5V.n9402 ASIG5V.n9401 0.022325
R49998 ASIG5V.n9108 ASIG5V.n9107 0.0223122
R49999 ASIG5V.n9079 ASIG5V.n9078 0.0219192
R50000 ASIG5V.n987 ASIG5V.n986 0.021875
R50001 ASIG5V.n710 ASIG5V.n709 0.0215262
R50002 ASIG5V.n1059 ASIG5V.n1028 0.021425
R50003 ASIG5V.n3145 ASIG5V.n3143 0.0202635
R50004 ASIG5V.n3337 ASIG5V.n3335 0.0202635
R50005 ASIG5V.n4169 ASIG5V.n4167 0.0202635
R50006 ASIG5V.n4452 ASIG5V.n4450 0.0202635
R50007 ASIG5V.n4706 ASIG5V.n4703 0.0202635
R50008 ASIG5V.n4981 ASIG5V.n4978 0.0202635
R50009 ASIG5V.n5404 ASIG5V.n5403 0.0202635
R50010 ASIG5V.n5686 ASIG5V.n5683 0.0202635
R50011 ASIG5V.n5982 ASIG5V.n5979 0.0202635
R50012 ASIG5V.n6337 ASIG5V.n6336 0.0202635
R50013 ASIG5V.n6422 ASIG5V.n6421 0.0202635
R50014 ASIG5V.n149 ASIG5V.n146 0.0202635
R50015 ASIG5V.n7525 ASIG5V.n7524 0.0202635
R50016 ASIG5V.n8128 ASIG5V.n8127 0.0202635
R50017 ASIG5V.n8195 ASIG5V.n8192 0.0202635
R50018 ASIG5V.n8613 ASIG5V.n8612 0.0202635
R50019 ASIG5V.n8718 ASIG5V.n8716 0.0202635
R50020 ASIG5V.n8856 ASIG5V.n8854 0.0202635
R50021 ASIG5V.n11662 ASIG5V.n11661 0.0202635
R50022 ASIG5V.n11791 ASIG5V.n11790 0.0202635
R50023 ASIG5V.n11954 ASIG5V.n11953 0.0202635
R50024 ASIG5V.n12113 ASIG5V.n12112 0.0202635
R50025 ASIG5V.n12266 ASIG5V.n12265 0.0202635
R50026 ASIG5V.n12383 ASIG5V.n12382 0.0202635
R50027 ASIG5V.n12609 ASIG5V.n12608 0.0202635
R50028 ASIG5V.n7269 ASIG5V.n7268 0.0202635
R50029 ASIG5V.n7851 ASIG5V.n7850 0.0202635
R50030 ASIG5V.n7434 ASIG5V.n7433 0.0202635
R50031 ASIG5V.n359 ASIG5V.n358 0.0202635
R50032 ASIG5V.n13523 ASIG5V.n13522 0.0202635
R50033 ASIG5V.n6685 ASIG5V.n6684 0.0202635
R50034 ASIG5V.n6963 ASIG5V.n6962 0.0202635
R50035 ASIG5V.n510 ASIG5V.n509 0.0202635
R50036 ASIG5V.n5888 ASIG5V.n5887 0.0202635
R50037 ASIG5V.n5587 ASIG5V.n5586 0.0202635
R50038 ASIG5V.n5356 ASIG5V.n5355 0.0202635
R50039 ASIG5V.n4929 ASIG5V.n4928 0.0202635
R50040 ASIG5V.n4661 ASIG5V.n4660 0.0202635
R50041 ASIG5V.n4403 ASIG5V.n4402 0.0202635
R50042 ASIG5V.n4127 ASIG5V.n4126 0.0202635
R50043 ASIG5V.n3861 ASIG5V.n3860 0.0202635
R50044 ASIG5V.n3586 ASIG5V.n3585 0.0202635
R50045 ASIG5V.n3327 ASIG5V.n3326 0.0202635
R50046 ASIG5V.n3132 ASIG5V.n3131 0.0202635
R50047 ASIG5V.n11659 ASIG5V.n11658 0.0202635
R50048 ASIG5V.n11788 ASIG5V.n11787 0.0202635
R50049 ASIG5V.n11951 ASIG5V.n11950 0.0202635
R50050 ASIG5V.n12110 ASIG5V.n12109 0.0202635
R50051 ASIG5V.n12263 ASIG5V.n12262 0.0202635
R50052 ASIG5V.n12380 ASIG5V.n12379 0.0202635
R50053 ASIG5V.n12606 ASIG5V.n12605 0.0202635
R50054 ASIG5V.n7266 ASIG5V.n7265 0.0202635
R50055 ASIG5V.n7848 ASIG5V.n7847 0.0202635
R50056 ASIG5V.n7431 ASIG5V.n7430 0.0202635
R50057 ASIG5V.n356 ASIG5V.n355 0.0202635
R50058 ASIG5V.n13520 ASIG5V.n13519 0.0202635
R50059 ASIG5V.n6682 ASIG5V.n6681 0.0202635
R50060 ASIG5V.n6960 ASIG5V.n6959 0.0202635
R50061 ASIG5V.n507 ASIG5V.n506 0.0202635
R50062 ASIG5V.n5885 ASIG5V.n5884 0.0202635
R50063 ASIG5V.n5584 ASIG5V.n5583 0.0202635
R50064 ASIG5V.n5353 ASIG5V.n5352 0.0202635
R50065 ASIG5V.n4926 ASIG5V.n4925 0.0202635
R50066 ASIG5V.n4658 ASIG5V.n4657 0.0202635
R50067 ASIG5V.n4400 ASIG5V.n4399 0.0202635
R50068 ASIG5V.n4124 ASIG5V.n4123 0.0202635
R50069 ASIG5V.n3858 ASIG5V.n3857 0.0202635
R50070 ASIG5V.n3583 ASIG5V.n3582 0.0202635
R50071 ASIG5V.n3324 ASIG5V.n3323 0.0202635
R50072 ASIG5V.n3129 ASIG5V.n3128 0.0202635
R50073 ASIG5V.n3125 ASIG5V.n3124 0.0202635
R50074 ASIG5V.n3320 ASIG5V.n3319 0.0202635
R50075 ASIG5V.n3579 ASIG5V.n3578 0.0202635
R50076 ASIG5V.n3854 ASIG5V.n3853 0.0202635
R50077 ASIG5V.n4120 ASIG5V.n4119 0.0202635
R50078 ASIG5V.n4396 ASIG5V.n4395 0.0202635
R50079 ASIG5V.n4654 ASIG5V.n4653 0.0202635
R50080 ASIG5V.n4922 ASIG5V.n4921 0.0202635
R50081 ASIG5V.n5349 ASIG5V.n5348 0.0202635
R50082 ASIG5V.n5580 ASIG5V.n5579 0.0202635
R50083 ASIG5V.n5881 ASIG5V.n5880 0.0202635
R50084 ASIG5V.n503 ASIG5V.n502 0.0202635
R50085 ASIG5V.n6956 ASIG5V.n6955 0.0202635
R50086 ASIG5V.n6678 ASIG5V.n6677 0.0202635
R50087 ASIG5V.n13516 ASIG5V.n13515 0.0202635
R50088 ASIG5V.n352 ASIG5V.n351 0.0202635
R50089 ASIG5V.n7427 ASIG5V.n7426 0.0202635
R50090 ASIG5V.n7844 ASIG5V.n7843 0.0202635
R50091 ASIG5V.n7262 ASIG5V.n7261 0.0202635
R50092 ASIG5V.n12602 ASIG5V.n12601 0.0202635
R50093 ASIG5V.n12376 ASIG5V.n12375 0.0202635
R50094 ASIG5V.n12259 ASIG5V.n12258 0.0202635
R50095 ASIG5V.n12106 ASIG5V.n12105 0.0202635
R50096 ASIG5V.n11947 ASIG5V.n11946 0.0202635
R50097 ASIG5V.n11784 ASIG5V.n11783 0.0202635
R50098 ASIG5V.n11655 ASIG5V.n11654 0.0202635
R50099 ASIG5V.n3121 ASIG5V.n3120 0.0202635
R50100 ASIG5V.n3316 ASIG5V.n3315 0.0202635
R50101 ASIG5V.n3575 ASIG5V.n3574 0.0202635
R50102 ASIG5V.n3850 ASIG5V.n3849 0.0202635
R50103 ASIG5V.n4116 ASIG5V.n4115 0.0202635
R50104 ASIG5V.n4392 ASIG5V.n4391 0.0202635
R50105 ASIG5V.n4650 ASIG5V.n4649 0.0202635
R50106 ASIG5V.n4918 ASIG5V.n4917 0.0202635
R50107 ASIG5V.n5345 ASIG5V.n5344 0.0202635
R50108 ASIG5V.n5576 ASIG5V.n5575 0.0202635
R50109 ASIG5V.n5877 ASIG5V.n5876 0.0202635
R50110 ASIG5V.n499 ASIG5V.n498 0.0202635
R50111 ASIG5V.n6952 ASIG5V.n6951 0.0202635
R50112 ASIG5V.n6674 ASIG5V.n6673 0.0202635
R50113 ASIG5V.n13512 ASIG5V.n13511 0.0202635
R50114 ASIG5V.n348 ASIG5V.n347 0.0202635
R50115 ASIG5V.n7423 ASIG5V.n7422 0.0202635
R50116 ASIG5V.n7840 ASIG5V.n7839 0.0202635
R50117 ASIG5V.n7258 ASIG5V.n7257 0.0202635
R50118 ASIG5V.n12598 ASIG5V.n12597 0.0202635
R50119 ASIG5V.n12372 ASIG5V.n12371 0.0202635
R50120 ASIG5V.n12255 ASIG5V.n12254 0.0202635
R50121 ASIG5V.n12102 ASIG5V.n12101 0.0202635
R50122 ASIG5V.n11943 ASIG5V.n11942 0.0202635
R50123 ASIG5V.n11780 ASIG5V.n11779 0.0202635
R50124 ASIG5V.n11651 ASIG5V.n11650 0.0202635
R50125 ASIG5V.n11647 ASIG5V.n11646 0.0202635
R50126 ASIG5V.n11776 ASIG5V.n11775 0.0202635
R50127 ASIG5V.n11939 ASIG5V.n11938 0.0202635
R50128 ASIG5V.n12098 ASIG5V.n12097 0.0202635
R50129 ASIG5V.n12251 ASIG5V.n12250 0.0202635
R50130 ASIG5V.n12368 ASIG5V.n12367 0.0202635
R50131 ASIG5V.n12594 ASIG5V.n12593 0.0202635
R50132 ASIG5V.n7254 ASIG5V.n7253 0.0202635
R50133 ASIG5V.n7836 ASIG5V.n7835 0.0202635
R50134 ASIG5V.n7419 ASIG5V.n7418 0.0202635
R50135 ASIG5V.n344 ASIG5V.n343 0.0202635
R50136 ASIG5V.n13508 ASIG5V.n13507 0.0202635
R50137 ASIG5V.n6670 ASIG5V.n6669 0.0202635
R50138 ASIG5V.n6948 ASIG5V.n6947 0.0202635
R50139 ASIG5V.n495 ASIG5V.n494 0.0202635
R50140 ASIG5V.n5873 ASIG5V.n5872 0.0202635
R50141 ASIG5V.n5572 ASIG5V.n5571 0.0202635
R50142 ASIG5V.n5341 ASIG5V.n5340 0.0202635
R50143 ASIG5V.n4914 ASIG5V.n4913 0.0202635
R50144 ASIG5V.n4646 ASIG5V.n4645 0.0202635
R50145 ASIG5V.n4388 ASIG5V.n4387 0.0202635
R50146 ASIG5V.n4112 ASIG5V.n4111 0.0202635
R50147 ASIG5V.n3846 ASIG5V.n3845 0.0202635
R50148 ASIG5V.n3571 ASIG5V.n3570 0.0202635
R50149 ASIG5V.n3312 ASIG5V.n3311 0.0202635
R50150 ASIG5V.n3117 ASIG5V.n3116 0.0202635
R50151 ASIG5V.n11643 ASIG5V.n11642 0.0202635
R50152 ASIG5V.n11772 ASIG5V.n11771 0.0202635
R50153 ASIG5V.n11935 ASIG5V.n11934 0.0202635
R50154 ASIG5V.n12094 ASIG5V.n12093 0.0202635
R50155 ASIG5V.n12247 ASIG5V.n12246 0.0202635
R50156 ASIG5V.n12364 ASIG5V.n12363 0.0202635
R50157 ASIG5V.n12590 ASIG5V.n12589 0.0202635
R50158 ASIG5V.n7250 ASIG5V.n7249 0.0202635
R50159 ASIG5V.n7832 ASIG5V.n7831 0.0202635
R50160 ASIG5V.n7415 ASIG5V.n7414 0.0202635
R50161 ASIG5V.n340 ASIG5V.n339 0.0202635
R50162 ASIG5V.n13504 ASIG5V.n13503 0.0202635
R50163 ASIG5V.n6666 ASIG5V.n6665 0.0202635
R50164 ASIG5V.n6944 ASIG5V.n6943 0.0202635
R50165 ASIG5V.n491 ASIG5V.n490 0.0202635
R50166 ASIG5V.n5869 ASIG5V.n5868 0.0202635
R50167 ASIG5V.n5568 ASIG5V.n5567 0.0202635
R50168 ASIG5V.n5337 ASIG5V.n5336 0.0202635
R50169 ASIG5V.n4910 ASIG5V.n4909 0.0202635
R50170 ASIG5V.n4642 ASIG5V.n4641 0.0202635
R50171 ASIG5V.n4384 ASIG5V.n4383 0.0202635
R50172 ASIG5V.n4108 ASIG5V.n4107 0.0202635
R50173 ASIG5V.n3842 ASIG5V.n3841 0.0202635
R50174 ASIG5V.n3567 ASIG5V.n3566 0.0202635
R50175 ASIG5V.n3308 ASIG5V.n3307 0.0202635
R50176 ASIG5V.n3113 ASIG5V.n3112 0.0202635
R50177 ASIG5V.n3109 ASIG5V.n3108 0.0202635
R50178 ASIG5V.n3304 ASIG5V.n3303 0.0202635
R50179 ASIG5V.n3563 ASIG5V.n3562 0.0202635
R50180 ASIG5V.n3838 ASIG5V.n3837 0.0202635
R50181 ASIG5V.n4104 ASIG5V.n4103 0.0202635
R50182 ASIG5V.n4380 ASIG5V.n4379 0.0202635
R50183 ASIG5V.n4638 ASIG5V.n4637 0.0202635
R50184 ASIG5V.n4906 ASIG5V.n4905 0.0202635
R50185 ASIG5V.n5333 ASIG5V.n5332 0.0202635
R50186 ASIG5V.n5564 ASIG5V.n5563 0.0202635
R50187 ASIG5V.n5865 ASIG5V.n5864 0.0202635
R50188 ASIG5V.n487 ASIG5V.n486 0.0202635
R50189 ASIG5V.n6940 ASIG5V.n6939 0.0202635
R50190 ASIG5V.n6662 ASIG5V.n6661 0.0202635
R50191 ASIG5V.n13500 ASIG5V.n13499 0.0202635
R50192 ASIG5V.n336 ASIG5V.n335 0.0202635
R50193 ASIG5V.n7411 ASIG5V.n7410 0.0202635
R50194 ASIG5V.n7828 ASIG5V.n7827 0.0202635
R50195 ASIG5V.n7246 ASIG5V.n7245 0.0202635
R50196 ASIG5V.n12586 ASIG5V.n12585 0.0202635
R50197 ASIG5V.n12360 ASIG5V.n12359 0.0202635
R50198 ASIG5V.n12243 ASIG5V.n12242 0.0202635
R50199 ASIG5V.n12090 ASIG5V.n12089 0.0202635
R50200 ASIG5V.n11931 ASIG5V.n11930 0.0202635
R50201 ASIG5V.n11768 ASIG5V.n11767 0.0202635
R50202 ASIG5V.n11639 ASIG5V.n11638 0.0202635
R50203 ASIG5V.n11557 ASIG5V.n11555 0.0202635
R50204 ASIG5V.n11714 ASIG5V.n11713 0.0202635
R50205 ASIG5V.n12195 ASIG5V.n12194 0.0202635
R50206 ASIG5V.n12490 ASIG5V.n12488 0.0202635
R50207 ASIG5V.n7567 ASIG5V.n7565 0.0202635
R50208 ASIG5V.n234 ASIG5V.n232 0.0202635
R50209 ASIG5V.n6618 ASIG5V.n6616 0.0202635
R50210 ASIG5V.n6831 ASIG5V.n6829 0.0202635
R50211 ASIG5V.n6065 ASIG5V.n6063 0.0202635
R50212 ASIG5V.n5737 ASIG5V.n5736 0.0202635
R50213 ASIG5V.n5060 ASIG5V.n5058 0.0202635
R50214 ASIG5V.n4770 ASIG5V.n4768 0.0202635
R50215 ASIG5V.n4503 ASIG5V.n4501 0.0202635
R50216 ASIG5V.n4220 ASIG5V.n4218 0.0202635
R50217 ASIG5V.n3950 ASIG5V.n3949 0.0202635
R50218 ASIG5V.n3682 ASIG5V.n3680 0.0202635
R50219 ASIG5V.n3402 ASIG5V.n3400 0.0202635
R50220 ASIG5V.n3197 ASIG5V.n3195 0.0202635
R50221 ASIG5V.n3200 ASIG5V.n3198 0.0202635
R50222 ASIG5V.n3405 ASIG5V.n3403 0.0202635
R50223 ASIG5V.n3684 ASIG5V.n3683 0.0202635
R50224 ASIG5V.n3953 ASIG5V.n3951 0.0202635
R50225 ASIG5V.n4223 ASIG5V.n4221 0.0202635
R50226 ASIG5V.n4506 ASIG5V.n4504 0.0202635
R50227 ASIG5V.n4773 ASIG5V.n4771 0.0202635
R50228 ASIG5V.n5063 ASIG5V.n5061 0.0202635
R50229 ASIG5V.n5739 ASIG5V.n5738 0.0202635
R50230 ASIG5V.n6068 ASIG5V.n6066 0.0202635
R50231 ASIG5V.n6834 ASIG5V.n6832 0.0202635
R50232 ASIG5V.n6621 ASIG5V.n6619 0.0202635
R50233 ASIG5V.n237 ASIG5V.n235 0.0202635
R50234 ASIG5V.n7569 ASIG5V.n7568 0.0202635
R50235 ASIG5V.n12493 ASIG5V.n12491 0.0202635
R50236 ASIG5V.n12197 ASIG5V.n12196 0.0202635
R50237 ASIG5V.n12043 ASIG5V.n12042 0.0202635
R50238 ASIG5V.n11716 ASIG5V.n11715 0.0202635
R50239 ASIG5V.n11560 ASIG5V.n11558 0.0202635
R50240 ASIG5V.n3150 ASIG5V.n3148 0.0202635
R50241 ASIG5V.n3342 ASIG5V.n3340 0.0202635
R50242 ASIG5V.n3906 ASIG5V.n3905 0.0202635
R50243 ASIG5V.n4174 ASIG5V.n4172 0.0202635
R50244 ASIG5V.n4456 ASIG5V.n4455 0.0202635
R50245 ASIG5V.n4711 ASIG5V.n4709 0.0202635
R50246 ASIG5V.n4986 ASIG5V.n4984 0.0202635
R50247 ASIG5V.n5690 ASIG5V.n5688 0.0202635
R50248 ASIG5V.n5987 ASIG5V.n5985 0.0202635
R50249 ASIG5V.n154 ASIG5V.n152 0.0202635
R50250 ASIG5V.n12671 ASIG5V.n12670 0.0202635
R50251 ASIG5V.n12438 ASIG5V.n12437 0.0202635
R50252 ASIG5V.n12012 ASIG5V.n12011 0.0202635
R50253 ASIG5V.n11844 ASIG5V.n11843 0.0202635
R50254 ASIG5V.n11679 ASIG5V.n11678 0.0202635
R50255 ASIG5V.n11497 ASIG5V.n11495 0.0202635
R50256 ASIG5V.n11563 ASIG5V.n11561 0.0202635
R50257 ASIG5V.n11718 ASIG5V.n11717 0.0202635
R50258 ASIG5V.n11882 ASIG5V.n11881 0.0202635
R50259 ASIG5V.n12045 ASIG5V.n12044 0.0202635
R50260 ASIG5V.n12199 ASIG5V.n12198 0.0202635
R50261 ASIG5V.n12496 ASIG5V.n12494 0.0202635
R50262 ASIG5V.n12707 ASIG5V.n12706 0.0202635
R50263 ASIG5V.n240 ASIG5V.n238 0.0202635
R50264 ASIG5V.n6624 ASIG5V.n6622 0.0202635
R50265 ASIG5V.n6837 ASIG5V.n6835 0.0202635
R50266 ASIG5V.n6071 ASIG5V.n6069 0.0202635
R50267 ASIG5V.n5741 ASIG5V.n5740 0.0202635
R50268 ASIG5V.n5066 ASIG5V.n5064 0.0202635
R50269 ASIG5V.n4776 ASIG5V.n4774 0.0202635
R50270 ASIG5V.n4508 ASIG5V.n4507 0.0202635
R50271 ASIG5V.n4226 ASIG5V.n4224 0.0202635
R50272 ASIG5V.n3955 ASIG5V.n3954 0.0202635
R50273 ASIG5V.n3408 ASIG5V.n3406 0.0202635
R50274 ASIG5V.n3202 ASIG5V.n3201 0.0202635
R50275 ASIG5V.n3204 ASIG5V.n3203 0.0202635
R50276 ASIG5V.n3411 ASIG5V.n3409 0.0202635
R50277 ASIG5V.n3957 ASIG5V.n3956 0.0202635
R50278 ASIG5V.n4229 ASIG5V.n4227 0.0202635
R50279 ASIG5V.n4510 ASIG5V.n4509 0.0202635
R50280 ASIG5V.n4779 ASIG5V.n4777 0.0202635
R50281 ASIG5V.n5069 ASIG5V.n5067 0.0202635
R50282 ASIG5V.n5743 ASIG5V.n5742 0.0202635
R50283 ASIG5V.n6074 ASIG5V.n6072 0.0202635
R50284 ASIG5V.n6840 ASIG5V.n6838 0.0202635
R50285 ASIG5V.n6627 ASIG5V.n6625 0.0202635
R50286 ASIG5V.n243 ASIG5V.n241 0.0202635
R50287 ASIG5V.n7572 ASIG5V.n7571 0.0202635
R50288 ASIG5V.n12709 ASIG5V.n12708 0.0202635
R50289 ASIG5V.n12499 ASIG5V.n12497 0.0202635
R50290 ASIG5V.n12047 ASIG5V.n12046 0.0202635
R50291 ASIG5V.n11884 ASIG5V.n11883 0.0202635
R50292 ASIG5V.n11720 ASIG5V.n11719 0.0202635
R50293 ASIG5V.n11566 ASIG5V.n11564 0.0202635
R50294 ASIG5V.n3153 ASIG5V.n3151 0.0202635
R50295 ASIG5V.n3345 ASIG5V.n3343 0.0202635
R50296 ASIG5V.n3635 ASIG5V.n3633 0.0202635
R50297 ASIG5V.n3908 ASIG5V.n3907 0.0202635
R50298 ASIG5V.n4177 ASIG5V.n4175 0.0202635
R50299 ASIG5V.n4458 ASIG5V.n4457 0.0202635
R50300 ASIG5V.n4714 ASIG5V.n4712 0.0202635
R50301 ASIG5V.n4989 ASIG5V.n4987 0.0202635
R50302 ASIG5V.n5990 ASIG5V.n5988 0.0202635
R50303 ASIG5V.n6795 ASIG5V.n6794 0.0202635
R50304 ASIG5V.n6560 ASIG5V.n6559 0.0202635
R50305 ASIG5V.n157 ASIG5V.n155 0.0202635
R50306 ASIG5V.n12673 ASIG5V.n12672 0.0202635
R50307 ASIG5V.n12440 ASIG5V.n12439 0.0202635
R50308 ASIG5V.n11846 ASIG5V.n11845 0.0202635
R50309 ASIG5V.n11681 ASIG5V.n11680 0.0202635
R50310 ASIG5V.n11500 ASIG5V.n11498 0.0202635
R50311 ASIG5V.n3155 ASIG5V.n3154 0.0202635
R50312 ASIG5V.n3348 ASIG5V.n3346 0.0202635
R50313 ASIG5V.n3638 ASIG5V.n3636 0.0202635
R50314 ASIG5V.n3910 ASIG5V.n3909 0.0202635
R50315 ASIG5V.n4180 ASIG5V.n4178 0.0202635
R50316 ASIG5V.n4460 ASIG5V.n4459 0.0202635
R50317 ASIG5V.n4717 ASIG5V.n4715 0.0202635
R50318 ASIG5V.n4992 ASIG5V.n4990 0.0202635
R50319 ASIG5V.n5993 ASIG5V.n5991 0.0202635
R50320 ASIG5V.n6797 ASIG5V.n6796 0.0202635
R50321 ASIG5V.n13376 ASIG5V.n13375 0.0202635
R50322 ASIG5V.n160 ASIG5V.n158 0.0202635
R50323 ASIG5V.n12675 ASIG5V.n12674 0.0202635
R50324 ASIG5V.n12443 ASIG5V.n12441 0.0202635
R50325 ASIG5V.n12169 ASIG5V.n12168 0.0202635
R50326 ASIG5V.n12015 ASIG5V.n12014 0.0202635
R50327 ASIG5V.n11848 ASIG5V.n11847 0.0202635
R50328 ASIG5V.n11503 ASIG5V.n11501 0.0202635
R50329 ASIG5V.n11569 ASIG5V.n11567 0.0202635
R50330 ASIG5V.n11722 ASIG5V.n11721 0.0202635
R50331 ASIG5V.n12049 ASIG5V.n12048 0.0202635
R50332 ASIG5V.n12202 ASIG5V.n12201 0.0202635
R50333 ASIG5V.n12503 ASIG5V.n12500 0.0202635
R50334 ASIG5V.n12711 ASIG5V.n12710 0.0202635
R50335 ASIG5V.n7574 ASIG5V.n7573 0.0202635
R50336 ASIG5V.n247 ASIG5V.n244 0.0202635
R50337 ASIG5V.n13416 ASIG5V.n13413 0.0202635
R50338 ASIG5V.n6629 ASIG5V.n6628 0.0202635
R50339 ASIG5V.n6844 ASIG5V.n6841 0.0202635
R50340 ASIG5V.n6078 ASIG5V.n6075 0.0202635
R50341 ASIG5V.n5745 ASIG5V.n5744 0.0202635
R50342 ASIG5V.n5073 ASIG5V.n5070 0.0202635
R50343 ASIG5V.n4783 ASIG5V.n4780 0.0202635
R50344 ASIG5V.n4512 ASIG5V.n4511 0.0202635
R50345 ASIG5V.n4231 ASIG5V.n4230 0.0202635
R50346 ASIG5V.n3961 ASIG5V.n3958 0.0202635
R50347 ASIG5V.n3414 ASIG5V.n3412 0.0202635
R50348 ASIG5V.n3206 ASIG5V.n3205 0.0202635
R50349 ASIG5V.n3157 ASIG5V.n3156 0.0202635
R50350 ASIG5V.n3353 ASIG5V.n3350 0.0202635
R50351 ASIG5V.n3643 ASIG5V.n3640 0.0202635
R50352 ASIG5V.n3915 ASIG5V.n3912 0.0202635
R50353 ASIG5V.n4183 ASIG5V.n4182 0.0202635
R50354 ASIG5V.n4463 ASIG5V.n4462 0.0202635
R50355 ASIG5V.n4722 ASIG5V.n4719 0.0202635
R50356 ASIG5V.n4997 ASIG5V.n4994 0.0202635
R50357 ASIG5V.n5695 ASIG5V.n5694 0.0202635
R50358 ASIG5V.n5998 ASIG5V.n5995 0.0202635
R50359 ASIG5V.n6564 ASIG5V.n6563 0.0202635
R50360 ASIG5V.n13379 ASIG5V.n13378 0.0202635
R50361 ASIG5V.n165 ASIG5V.n162 0.0202635
R50362 ASIG5V.n7533 ASIG5V.n7532 0.0202635
R50363 ASIG5V.n12678 ASIG5V.n12677 0.0202635
R50364 ASIG5V.n12446 ASIG5V.n12445 0.0202635
R50365 ASIG5V.n12018 ASIG5V.n12017 0.0202635
R50366 ASIG5V.n11851 ASIG5V.n11850 0.0202635
R50367 ASIG5V.n11685 ASIG5V.n11684 0.0202635
R50368 ASIG5V.n11508 ASIG5V.n11505 0.0202635
R50369 ASIG5V.n3162 ASIG5V.n3159 0.0202635
R50370 ASIG5V.n3358 ASIG5V.n3355 0.0202635
R50371 ASIG5V.n3648 ASIG5V.n3645 0.0202635
R50372 ASIG5V.n3918 ASIG5V.n3917 0.0202635
R50373 ASIG5V.n4188 ASIG5V.n4185 0.0202635
R50374 ASIG5V.n4468 ASIG5V.n4465 0.0202635
R50375 ASIG5V.n4727 ASIG5V.n4724 0.0202635
R50376 ASIG5V.n5002 ASIG5V.n4999 0.0202635
R50377 ASIG5V.n5698 ASIG5V.n5697 0.0202635
R50378 ASIG5V.n6003 ASIG5V.n6000 0.0202635
R50379 ASIG5V.n6801 ASIG5V.n6800 0.0202635
R50380 ASIG5V.n13382 ASIG5V.n13381 0.0202635
R50381 ASIG5V.n170 ASIG5V.n167 0.0202635
R50382 ASIG5V.n7536 ASIG5V.n7535 0.0202635
R50383 ASIG5V.n12683 ASIG5V.n12680 0.0202635
R50384 ASIG5V.n12449 ASIG5V.n12448 0.0202635
R50385 ASIG5V.n12173 ASIG5V.n12172 0.0202635
R50386 ASIG5V.n12021 ASIG5V.n12020 0.0202635
R50387 ASIG5V.n11854 ASIG5V.n11853 0.0202635
R50388 ASIG5V.n11513 ASIG5V.n11510 0.0202635
R50389 ASIG5V.n11574 ASIG5V.n11571 0.0202635
R50390 ASIG5V.n11725 ASIG5V.n11724 0.0202635
R50391 ASIG5V.n11888 ASIG5V.n11887 0.0202635
R50392 ASIG5V.n12052 ASIG5V.n12051 0.0202635
R50393 ASIG5V.n12205 ASIG5V.n12204 0.0202635
R50394 ASIG5V.n12508 ASIG5V.n12505 0.0202635
R50395 ASIG5V.n12714 ASIG5V.n12713 0.0202635
R50396 ASIG5V.n7577 ASIG5V.n7576 0.0202635
R50397 ASIG5V.n252 ASIG5V.n249 0.0202635
R50398 ASIG5V.n13419 ASIG5V.n13418 0.0202635
R50399 ASIG5V.n6632 ASIG5V.n6631 0.0202635
R50400 ASIG5V.n6849 ASIG5V.n6846 0.0202635
R50401 ASIG5V.n6083 ASIG5V.n6080 0.0202635
R50402 ASIG5V.n5748 ASIG5V.n5747 0.0202635
R50403 ASIG5V.n5427 ASIG5V.n5426 0.0202635
R50404 ASIG5V.n5078 ASIG5V.n5075 0.0202635
R50405 ASIG5V.n4788 ASIG5V.n4785 0.0202635
R50406 ASIG5V.n4515 ASIG5V.n4514 0.0202635
R50407 ASIG5V.n4234 ASIG5V.n4233 0.0202635
R50408 ASIG5V.n3966 ASIG5V.n3963 0.0202635
R50409 ASIG5V.n3693 ASIG5V.n3692 0.0202635
R50410 ASIG5V.n3419 ASIG5V.n3416 0.0202635
R50411 ASIG5V.n3209 ASIG5V.n3208 0.0202635
R50412 ASIG5V.n3214 ASIG5V.n3211 0.0202635
R50413 ASIG5V.n3424 ASIG5V.n3421 0.0202635
R50414 ASIG5V.n3969 ASIG5V.n3968 0.0202635
R50415 ASIG5V.n4239 ASIG5V.n4236 0.0202635
R50416 ASIG5V.n4518 ASIG5V.n4517 0.0202635
R50417 ASIG5V.n4793 ASIG5V.n4790 0.0202635
R50418 ASIG5V.n5083 ASIG5V.n5080 0.0202635
R50419 ASIG5V.n5751 ASIG5V.n5750 0.0202635
R50420 ASIG5V.n6088 ASIG5V.n6085 0.0202635
R50421 ASIG5V.n6854 ASIG5V.n6851 0.0202635
R50422 ASIG5V.n6635 ASIG5V.n6634 0.0202635
R50423 ASIG5V.n13422 ASIG5V.n13421 0.0202635
R50424 ASIG5V.n257 ASIG5V.n254 0.0202635
R50425 ASIG5V.n7582 ASIG5V.n7579 0.0202635
R50426 ASIG5V.n12717 ASIG5V.n12716 0.0202635
R50427 ASIG5V.n12513 ASIG5V.n12510 0.0202635
R50428 ASIG5V.n11891 ASIG5V.n11890 0.0202635
R50429 ASIG5V.n11728 ASIG5V.n11727 0.0202635
R50430 ASIG5V.n11579 ASIG5V.n11576 0.0202635
R50431 ASIG5V.n3167 ASIG5V.n3164 0.0202635
R50432 ASIG5V.n3363 ASIG5V.n3360 0.0202635
R50433 ASIG5V.n4191 ASIG5V.n4190 0.0202635
R50434 ASIG5V.n4471 ASIG5V.n4470 0.0202635
R50435 ASIG5V.n4732 ASIG5V.n4729 0.0202635
R50436 ASIG5V.n5007 ASIG5V.n5004 0.0202635
R50437 ASIG5V.n5701 ASIG5V.n5700 0.0202635
R50438 ASIG5V.n6008 ASIG5V.n6005 0.0202635
R50439 ASIG5V.n6568 ASIG5V.n6567 0.0202635
R50440 ASIG5V.n13385 ASIG5V.n13384 0.0202635
R50441 ASIG5V.n175 ASIG5V.n172 0.0202635
R50442 ASIG5V.n7539 ASIG5V.n7538 0.0202635
R50443 ASIG5V.n12686 ASIG5V.n12685 0.0202635
R50444 ASIG5V.n12452 ASIG5V.n12451 0.0202635
R50445 ASIG5V.n12176 ASIG5V.n12175 0.0202635
R50446 ASIG5V.n11857 ASIG5V.n11856 0.0202635
R50447 ASIG5V.n11689 ASIG5V.n11688 0.0202635
R50448 ASIG5V.n11518 ASIG5V.n11515 0.0202635
R50449 ASIG5V.n11584 ASIG5V.n11581 0.0202635
R50450 ASIG5V.n11731 ASIG5V.n11730 0.0202635
R50451 ASIG5V.n11894 ASIG5V.n11893 0.0202635
R50452 ASIG5V.n12056 ASIG5V.n12055 0.0202635
R50453 ASIG5V.n12518 ASIG5V.n12515 0.0202635
R50454 ASIG5V.n12720 ASIG5V.n12719 0.0202635
R50455 ASIG5V.n7585 ASIG5V.n7584 0.0202635
R50456 ASIG5V.n262 ASIG5V.n259 0.0202635
R50457 ASIG5V.n13425 ASIG5V.n13424 0.0202635
R50458 ASIG5V.n6638 ASIG5V.n6637 0.0202635
R50459 ASIG5V.n6859 ASIG5V.n6856 0.0202635
R50460 ASIG5V.n6093 ASIG5V.n6090 0.0202635
R50461 ASIG5V.n5754 ASIG5V.n5753 0.0202635
R50462 ASIG5V.n5088 ASIG5V.n5085 0.0202635
R50463 ASIG5V.n4796 ASIG5V.n4795 0.0202635
R50464 ASIG5V.n4521 ASIG5V.n4520 0.0202635
R50465 ASIG5V.n4242 ASIG5V.n4241 0.0202635
R50466 ASIG5V.n3972 ASIG5V.n3971 0.0202635
R50467 ASIG5V.n3701 ASIG5V.n3698 0.0202635
R50468 ASIG5V.n3429 ASIG5V.n3426 0.0202635
R50469 ASIG5V.n3219 ASIG5V.n3216 0.0202635
R50470 ASIG5V.n11589 ASIG5V.n11586 0.0202635
R50471 ASIG5V.n11734 ASIG5V.n11733 0.0202635
R50472 ASIG5V.n11897 ASIG5V.n11896 0.0202635
R50473 ASIG5V.n12210 ASIG5V.n12209 0.0202635
R50474 ASIG5V.n12523 ASIG5V.n12520 0.0202635
R50475 ASIG5V.n12723 ASIG5V.n12722 0.0202635
R50476 ASIG5V.n7590 ASIG5V.n7587 0.0202635
R50477 ASIG5V.n268 ASIG5V.n264 0.0202635
R50478 ASIG5V.n13431 ASIG5V.n13427 0.0202635
R50479 ASIG5V.n6864 ASIG5V.n6861 0.0202635
R50480 ASIG5V.n6099 ASIG5V.n6095 0.0202635
R50481 ASIG5V.n5757 ASIG5V.n5756 0.0202635
R50482 ASIG5V.n5093 ASIG5V.n5090 0.0202635
R50483 ASIG5V.n4801 ASIG5V.n4798 0.0202635
R50484 ASIG5V.n4524 ASIG5V.n4523 0.0202635
R50485 ASIG5V.n4245 ASIG5V.n4244 0.0202635
R50486 ASIG5V.n3975 ASIG5V.n3974 0.0202635
R50487 ASIG5V.n3434 ASIG5V.n3431 0.0202635
R50488 ASIG5V.n3222 ASIG5V.n3221 0.0202635
R50489 ASIG5V.n3170 ASIG5V.n3169 0.0202635
R50490 ASIG5V.n3368 ASIG5V.n3365 0.0202635
R50491 ASIG5V.n3656 ASIG5V.n3653 0.0202635
R50492 ASIG5V.n3922 ASIG5V.n3921 0.0202635
R50493 ASIG5V.n4194 ASIG5V.n4193 0.0202635
R50494 ASIG5V.n4474 ASIG5V.n4473 0.0202635
R50495 ASIG5V.n4737 ASIG5V.n4734 0.0202635
R50496 ASIG5V.n5013 ASIG5V.n5009 0.0202635
R50497 ASIG5V.n5705 ASIG5V.n5704 0.0202635
R50498 ASIG5V.n6015 ASIG5V.n6011 0.0202635
R50499 ASIG5V.n6806 ASIG5V.n6805 0.0202635
R50500 ASIG5V.n6572 ASIG5V.n6571 0.0202635
R50501 ASIG5V.n182 ASIG5V.n178 0.0202635
R50502 ASIG5V.n7543 ASIG5V.n7542 0.0202635
R50503 ASIG5V.n12690 ASIG5V.n12689 0.0202635
R50504 ASIG5V.n12458 ASIG5V.n12454 0.0202635
R50505 ASIG5V.n12179 ASIG5V.n12178 0.0202635
R50506 ASIG5V.n12025 ASIG5V.n12024 0.0202635
R50507 ASIG5V.n11860 ASIG5V.n11859 0.0202635
R50508 ASIG5V.n11692 ASIG5V.n11691 0.0202635
R50509 ASIG5V.n11523 ASIG5V.n11520 0.0202635
R50510 ASIG5V.n3175 ASIG5V.n3172 0.0202635
R50511 ASIG5V.n3373 ASIG5V.n3370 0.0202635
R50512 ASIG5V.n3661 ASIG5V.n3658 0.0202635
R50513 ASIG5V.n3925 ASIG5V.n3924 0.0202635
R50514 ASIG5V.n4197 ASIG5V.n4196 0.0202635
R50515 ASIG5V.n4477 ASIG5V.n4476 0.0202635
R50516 ASIG5V.n4740 ASIG5V.n4739 0.0202635
R50517 ASIG5V.n5020 ASIG5V.n5016 0.0202635
R50518 ASIG5V.n5709 ASIG5V.n5708 0.0202635
R50519 ASIG5V.n6022 ASIG5V.n6018 0.0202635
R50520 ASIG5V.n6810 ASIG5V.n6809 0.0202635
R50521 ASIG5V.n6576 ASIG5V.n6575 0.0202635
R50522 ASIG5V.n13390 ASIG5V.n13389 0.0202635
R50523 ASIG5V.n189 ASIG5V.n185 0.0202635
R50524 ASIG5V.n7547 ASIG5V.n7546 0.0202635
R50525 ASIG5V.n12694 ASIG5V.n12693 0.0202635
R50526 ASIG5V.n12462 ASIG5V.n12461 0.0202635
R50527 ASIG5V.n12182 ASIG5V.n12181 0.0202635
R50528 ASIG5V.n12028 ASIG5V.n12027 0.0202635
R50529 ASIG5V.n11695 ASIG5V.n11694 0.0202635
R50530 ASIG5V.n11528 ASIG5V.n11525 0.0202635
R50531 ASIG5V.n11594 ASIG5V.n11591 0.0202635
R50532 ASIG5V.n11737 ASIG5V.n11736 0.0202635
R50533 ASIG5V.n12060 ASIG5V.n12059 0.0202635
R50534 ASIG5V.n12214 ASIG5V.n12213 0.0202635
R50535 ASIG5V.n12530 ASIG5V.n12526 0.0202635
R50536 ASIG5V.n7594 ASIG5V.n7593 0.0202635
R50537 ASIG5V.n275 ASIG5V.n271 0.0202635
R50538 ASIG5V.n13438 ASIG5V.n13434 0.0202635
R50539 ASIG5V.n6871 ASIG5V.n6867 0.0202635
R50540 ASIG5V.n6106 ASIG5V.n6102 0.0202635
R50541 ASIG5V.n5761 ASIG5V.n5760 0.0202635
R50542 ASIG5V.n5100 ASIG5V.n5096 0.0202635
R50543 ASIG5V.n4808 ASIG5V.n4804 0.0202635
R50544 ASIG5V.n4531 ASIG5V.n4527 0.0202635
R50545 ASIG5V.n4248 ASIG5V.n4247 0.0202635
R50546 ASIG5V.n3978 ASIG5V.n3977 0.0202635
R50547 ASIG5V.n3439 ASIG5V.n3436 0.0202635
R50548 ASIG5V.n3225 ASIG5V.n3224 0.0202635
R50549 ASIG5V.n3228 ASIG5V.n3227 0.0202635
R50550 ASIG5V.n3444 ASIG5V.n3441 0.0202635
R50551 ASIG5V.n3712 ASIG5V.n3709 0.0202635
R50552 ASIG5V.n3981 ASIG5V.n3980 0.0202635
R50553 ASIG5V.n4252 ASIG5V.n4251 0.0202635
R50554 ASIG5V.n4535 ASIG5V.n4534 0.0202635
R50555 ASIG5V.n4812 ASIG5V.n4811 0.0202635
R50556 ASIG5V.n5107 ASIG5V.n5103 0.0202635
R50557 ASIG5V.n5765 ASIG5V.n5764 0.0202635
R50558 ASIG5V.n6113 ASIG5V.n6109 0.0202635
R50559 ASIG5V.n6878 ASIG5V.n6874 0.0202635
R50560 ASIG5V.n13445 ASIG5V.n13441 0.0202635
R50561 ASIG5V.n282 ASIG5V.n278 0.0202635
R50562 ASIG5V.n7601 ASIG5V.n7597 0.0202635
R50563 ASIG5V.n12537 ASIG5V.n12533 0.0202635
R50564 ASIG5V.n12064 ASIG5V.n12063 0.0202635
R50565 ASIG5V.n11901 ASIG5V.n11900 0.0202635
R50566 ASIG5V.n11599 ASIG5V.n11596 0.0202635
R50567 ASIG5V.n3178 ASIG5V.n3177 0.0202635
R50568 ASIG5V.n3378 ASIG5V.n3375 0.0202635
R50569 ASIG5V.n3929 ASIG5V.n3928 0.0202635
R50570 ASIG5V.n4201 ASIG5V.n4200 0.0202635
R50571 ASIG5V.n4481 ASIG5V.n4480 0.0202635
R50572 ASIG5V.n5027 ASIG5V.n5023 0.0202635
R50573 ASIG5V.n5713 ASIG5V.n5712 0.0202635
R50574 ASIG5V.n6029 ASIG5V.n6025 0.0202635
R50575 ASIG5V.n6814 ASIG5V.n6813 0.0202635
R50576 ASIG5V.n6583 ASIG5V.n6579 0.0202635
R50577 ASIG5V.n196 ASIG5V.n192 0.0202635
R50578 ASIG5V.n12698 ASIG5V.n12697 0.0202635
R50579 ASIG5V.n12466 ASIG5V.n12465 0.0202635
R50580 ASIG5V.n11865 ASIG5V.n11864 0.0202635
R50581 ASIG5V.n11699 ASIG5V.n11698 0.0202635
R50582 ASIG5V.n11533 ASIG5V.n11530 0.0202635
R50583 ASIG5V.n11604 ASIG5V.n11601 0.0202635
R50584 ASIG5V.n11742 ASIG5V.n11741 0.0202635
R50585 ASIG5V.n11905 ASIG5V.n11904 0.0202635
R50586 ASIG5V.n12068 ASIG5V.n12067 0.0202635
R50587 ASIG5V.n12219 ASIG5V.n12218 0.0202635
R50588 ASIG5V.n12544 ASIG5V.n12540 0.0202635
R50589 ASIG5V.n12729 ASIG5V.n12728 0.0202635
R50590 ASIG5V.n7605 ASIG5V.n7604 0.0202635
R50591 ASIG5V.n289 ASIG5V.n285 0.0202635
R50592 ASIG5V.n13452 ASIG5V.n13448 0.0202635
R50593 ASIG5V.n6645 ASIG5V.n6644 0.0202635
R50594 ASIG5V.n6885 ASIG5V.n6881 0.0202635
R50595 ASIG5V.n6120 ASIG5V.n6116 0.0202635
R50596 ASIG5V.n5772 ASIG5V.n5768 0.0202635
R50597 ASIG5V.n5114 ASIG5V.n5110 0.0202635
R50598 ASIG5V.n4819 ASIG5V.n4815 0.0202635
R50599 ASIG5V.n4539 ASIG5V.n4538 0.0202635
R50600 ASIG5V.n4256 ASIG5V.n4255 0.0202635
R50601 ASIG5V.n3985 ASIG5V.n3984 0.0202635
R50602 ASIG5V.n3449 ASIG5V.n3446 0.0202635
R50603 ASIG5V.n3231 ASIG5V.n3230 0.0202635
R50604 ASIG5V.n11609 ASIG5V.n11606 0.0202635
R50605 ASIG5V.n11745 ASIG5V.n11744 0.0202635
R50606 ASIG5V.n11909 ASIG5V.n11908 0.0202635
R50607 ASIG5V.n12072 ASIG5V.n12071 0.0202635
R50608 ASIG5V.n12223 ASIG5V.n12222 0.0202635
R50609 ASIG5V.n12551 ASIG5V.n12547 0.0202635
R50610 ASIG5V.n12733 ASIG5V.n12732 0.0202635
R50611 ASIG5V.n7609 ASIG5V.n7608 0.0202635
R50612 ASIG5V.n296 ASIG5V.n292 0.0202635
R50613 ASIG5V.n13459 ASIG5V.n13455 0.0202635
R50614 ASIG5V.n6892 ASIG5V.n6888 0.0202635
R50615 ASIG5V.n6127 ASIG5V.n6123 0.0202635
R50616 ASIG5V.n5779 ASIG5V.n5775 0.0202635
R50617 ASIG5V.n5121 ASIG5V.n5117 0.0202635
R50618 ASIG5V.n4826 ASIG5V.n4822 0.0202635
R50619 ASIG5V.n4543 ASIG5V.n4542 0.0202635
R50620 ASIG5V.n4260 ASIG5V.n4259 0.0202635
R50621 ASIG5V.n3989 ASIG5V.n3988 0.0202635
R50622 ASIG5V.n3720 ASIG5V.n3717 0.0202635
R50623 ASIG5V.n3454 ASIG5V.n3451 0.0202635
R50624 ASIG5V.n3236 ASIG5V.n3233 0.0202635
R50625 ASIG5V.n3181 ASIG5V.n3180 0.0202635
R50626 ASIG5V.n3383 ASIG5V.n3380 0.0202635
R50627 ASIG5V.n3670 ASIG5V.n3667 0.0202635
R50628 ASIG5V.n3932 ASIG5V.n3931 0.0202635
R50629 ASIG5V.n4205 ASIG5V.n4204 0.0202635
R50630 ASIG5V.n4485 ASIG5V.n4484 0.0202635
R50631 ASIG5V.n4748 ASIG5V.n4744 0.0202635
R50632 ASIG5V.n5034 ASIG5V.n5030 0.0202635
R50633 ASIG5V.n5717 ASIG5V.n5716 0.0202635
R50634 ASIG5V.n6036 ASIG5V.n6032 0.0202635
R50635 ASIG5V.n6818 ASIG5V.n6817 0.0202635
R50636 ASIG5V.n6590 ASIG5V.n6586 0.0202635
R50637 ASIG5V.n13398 ASIG5V.n13394 0.0202635
R50638 ASIG5V.n203 ASIG5V.n199 0.0202635
R50639 ASIG5V.n12187 ASIG5V.n12186 0.0202635
R50640 ASIG5V.n11868 ASIG5V.n11867 0.0202635
R50641 ASIG5V.n11702 ASIG5V.n11701 0.0202635
R50642 ASIG5V.n11538 ASIG5V.n11535 0.0202635
R50643 ASIG5V.n3186 ASIG5V.n3183 0.0202635
R50644 ASIG5V.n3388 ASIG5V.n3385 0.0202635
R50645 ASIG5V.n3937 ASIG5V.n3934 0.0202635
R50646 ASIG5V.n4208 ASIG5V.n4207 0.0202635
R50647 ASIG5V.n4489 ASIG5V.n4488 0.0202635
R50648 ASIG5V.n4752 ASIG5V.n4751 0.0202635
R50649 ASIG5V.n5041 ASIG5V.n5037 0.0202635
R50650 ASIG5V.n5721 ASIG5V.n5720 0.0202635
R50651 ASIG5V.n6043 ASIG5V.n6039 0.0202635
R50652 ASIG5V.n6597 ASIG5V.n6593 0.0202635
R50653 ASIG5V.n13402 ASIG5V.n13401 0.0202635
R50654 ASIG5V.n210 ASIG5V.n206 0.0202635
R50655 ASIG5V.n7553 ASIG5V.n7552 0.0202635
R50656 ASIG5V.n12471 ASIG5V.n12470 0.0202635
R50657 ASIG5V.n12033 ASIG5V.n12032 0.0202635
R50658 ASIG5V.n11871 ASIG5V.n11870 0.0202635
R50659 ASIG5V.n11705 ASIG5V.n11704 0.0202635
R50660 ASIG5V.n11543 ASIG5V.n11540 0.0202635
R50661 ASIG5V.n11614 ASIG5V.n11611 0.0202635
R50662 ASIG5V.n11748 ASIG5V.n11747 0.0202635
R50663 ASIG5V.n11912 ASIG5V.n11911 0.0202635
R50664 ASIG5V.n12075 ASIG5V.n12074 0.0202635
R50665 ASIG5V.n12227 ASIG5V.n12226 0.0202635
R50666 ASIG5V.n12558 ASIG5V.n12554 0.0202635
R50667 ASIG5V.n12737 ASIG5V.n12736 0.0202635
R50668 ASIG5V.n7613 ASIG5V.n7612 0.0202635
R50669 ASIG5V.n303 ASIG5V.n299 0.0202635
R50670 ASIG5V.n13466 ASIG5V.n13462 0.0202635
R50671 ASIG5V.n6899 ASIG5V.n6895 0.0202635
R50672 ASIG5V.n7113 ASIG5V.n7112 0.0202635
R50673 ASIG5V.n6134 ASIG5V.n6130 0.0202635
R50674 ASIG5V.n5128 ASIG5V.n5124 0.0202635
R50675 ASIG5V.n4830 ASIG5V.n4829 0.0202635
R50676 ASIG5V.n4546 ASIG5V.n4545 0.0202635
R50677 ASIG5V.n4263 ASIG5V.n4262 0.0202635
R50678 ASIG5V.n3725 ASIG5V.n3722 0.0202635
R50679 ASIG5V.n3459 ASIG5V.n3456 0.0202635
R50680 ASIG5V.n3239 ASIG5V.n3238 0.0202635
R50681 ASIG5V.n3244 ASIG5V.n3241 0.0202635
R50682 ASIG5V.n3464 ASIG5V.n3461 0.0202635
R50683 ASIG5V.n3995 ASIG5V.n3994 0.0202635
R50684 ASIG5V.n4266 ASIG5V.n4265 0.0202635
R50685 ASIG5V.n4549 ASIG5V.n4548 0.0202635
R50686 ASIG5V.n4835 ASIG5V.n4832 0.0202635
R50687 ASIG5V.n5132 ASIG5V.n5131 0.0202635
R50688 ASIG5V.n5784 ASIG5V.n5783 0.0202635
R50689 ASIG5V.n7117 ASIG5V.n7116 0.0202635
R50690 ASIG5V.n6906 ASIG5V.n6902 0.0202635
R50691 ASIG5V.n13473 ASIG5V.n13469 0.0202635
R50692 ASIG5V.n310 ASIG5V.n306 0.0202635
R50693 ASIG5V.n7617 ASIG5V.n7616 0.0202635
R50694 ASIG5V.n12741 ASIG5V.n12740 0.0202635
R50695 ASIG5V.n12565 ASIG5V.n12561 0.0202635
R50696 ASIG5V.n12230 ASIG5V.n12229 0.0202635
R50697 ASIG5V.n11917 ASIG5V.n11914 0.0202635
R50698 ASIG5V.n11751 ASIG5V.n11750 0.0202635
R50699 ASIG5V.n11619 ASIG5V.n11616 0.0202635
R50700 ASIG5V.n3189 ASIG5V.n3188 0.0202635
R50701 ASIG5V.n3393 ASIG5V.n3390 0.0202635
R50702 ASIG5V.n3942 ASIG5V.n3939 0.0202635
R50703 ASIG5V.n4211 ASIG5V.n4210 0.0202635
R50704 ASIG5V.n4492 ASIG5V.n4491 0.0202635
R50705 ASIG5V.n4757 ASIG5V.n4754 0.0202635
R50706 ASIG5V.n5047 ASIG5V.n5044 0.0202635
R50707 ASIG5V.n5725 ASIG5V.n5724 0.0202635
R50708 ASIG5V.n6050 ASIG5V.n6046 0.0202635
R50709 ASIG5V.n7088 ASIG5V.n7084 0.0202635
R50710 ASIG5V.n6604 ASIG5V.n6600 0.0202635
R50711 ASIG5V.n217 ASIG5V.n213 0.0202635
R50712 ASIG5V.n7557 ASIG5V.n7556 0.0202635
R50713 ASIG5V.n12477 ASIG5V.n12474 0.0202635
R50714 ASIG5V.n12191 ASIG5V.n12190 0.0202635
R50715 ASIG5V.n12036 ASIG5V.n12035 0.0202635
R50716 ASIG5V.n11874 ASIG5V.n11873 0.0202635
R50717 ASIG5V.n11708 ASIG5V.n11707 0.0202635
R50718 ASIG5V.n11548 ASIG5V.n11545 0.0202635
R50719 ASIG5V.n11624 ASIG5V.n11621 0.0202635
R50720 ASIG5V.n11754 ASIG5V.n11753 0.0202635
R50721 ASIG5V.n11920 ASIG5V.n11919 0.0202635
R50722 ASIG5V.n12079 ASIG5V.n12078 0.0202635
R50723 ASIG5V.n12570 ASIG5V.n12567 0.0202635
R50724 ASIG5V.n12745 ASIG5V.n12744 0.0202635
R50725 ASIG5V.n7621 ASIG5V.n7620 0.0202635
R50726 ASIG5V.n317 ASIG5V.n313 0.0202635
R50727 ASIG5V.n13480 ASIG5V.n13476 0.0202635
R50728 ASIG5V.n6913 ASIG5V.n6909 0.0202635
R50729 ASIG5V.n6142 ASIG5V.n6138 0.0202635
R50730 ASIG5V.n5788 ASIG5V.n5787 0.0202635
R50731 ASIG5V.n5135 ASIG5V.n5134 0.0202635
R50732 ASIG5V.n4840 ASIG5V.n4837 0.0202635
R50733 ASIG5V.n4552 ASIG5V.n4551 0.0202635
R50734 ASIG5V.n4271 ASIG5V.n4268 0.0202635
R50735 ASIG5V.n3469 ASIG5V.n3466 0.0202635
R50736 ASIG5V.n3246 ASIG5V.n3245 0.0202635
R50737 ASIG5V.n11627 ASIG5V.n11625 0.0202635
R50738 ASIG5V.n11757 ASIG5V.n11756 0.0202635
R50739 ASIG5V.n11923 ASIG5V.n11922 0.0202635
R50740 ASIG5V.n12234 ASIG5V.n12233 0.0202635
R50741 ASIG5V.n12575 ASIG5V.n12572 0.0202635
R50742 ASIG5V.n12748 ASIG5V.n12747 0.0202635
R50743 ASIG5V.n324 ASIG5V.n320 0.0202635
R50744 ASIG5V.n13487 ASIG5V.n13483 0.0202635
R50745 ASIG5V.n6920 ASIG5V.n6916 0.0202635
R50746 ASIG5V.n5138 ASIG5V.n5137 0.0202635
R50747 ASIG5V.n4843 ASIG5V.n4842 0.0202635
R50748 ASIG5V.n4555 ASIG5V.n4554 0.0202635
R50749 ASIG5V.n4274 ASIG5V.n4273 0.0202635
R50750 ASIG5V.n4001 ASIG5V.n3998 0.0202635
R50751 ASIG5V.n3472 ASIG5V.n3470 0.0202635
R50752 ASIG5V.n3248 ASIG5V.n3247 0.0202635
R50753 ASIG5V.n3192 ASIG5V.n3190 0.0202635
R50754 ASIG5V.n3396 ASIG5V.n3394 0.0202635
R50755 ASIG5V.n3677 ASIG5V.n3675 0.0202635
R50756 ASIG5V.n3945 ASIG5V.n3944 0.0202635
R50757 ASIG5V.n4214 ASIG5V.n4213 0.0202635
R50758 ASIG5V.n4497 ASIG5V.n4494 0.0202635
R50759 ASIG5V.n4762 ASIG5V.n4759 0.0202635
R50760 ASIG5V.n5052 ASIG5V.n5049 0.0202635
R50761 ASIG5V.n5730 ASIG5V.n5727 0.0202635
R50762 ASIG5V.n6057 ASIG5V.n6053 0.0202635
R50763 ASIG5V.n7092 ASIG5V.n7091 0.0202635
R50764 ASIG5V.n6824 ASIG5V.n6823 0.0202635
R50765 ASIG5V.n6611 ASIG5V.n6607 0.0202635
R50766 ASIG5V.n224 ASIG5V.n220 0.0202635
R50767 ASIG5V.n7561 ASIG5V.n7560 0.0202635
R50768 ASIG5V.n12482 ASIG5V.n12479 0.0202635
R50769 ASIG5V.n12039 ASIG5V.n12038 0.0202635
R50770 ASIG5V.n11877 ASIG5V.n11876 0.0202635
R50771 ASIG5V.n11710 ASIG5V.n11709 0.0202635
R50772 ASIG5V.n11551 ASIG5V.n11549 0.0202635
R50773 ASIG5V.n3194 ASIG5V.n3193 0.0202635
R50774 ASIG5V.n3399 ASIG5V.n3397 0.0202635
R50775 ASIG5V.n3948 ASIG5V.n3946 0.0202635
R50776 ASIG5V.n4217 ASIG5V.n4216 0.0202635
R50777 ASIG5V.n4500 ASIG5V.n4499 0.0202635
R50778 ASIG5V.n4767 ASIG5V.n4764 0.0202635
R50779 ASIG5V.n5057 ASIG5V.n5054 0.0202635
R50780 ASIG5V.n5735 ASIG5V.n5732 0.0202635
R50781 ASIG5V.n6062 ASIG5V.n6059 0.0202635
R50782 ASIG5V.n7096 ASIG5V.n7095 0.0202635
R50783 ASIG5V.n6828 ASIG5V.n6827 0.0202635
R50784 ASIG5V.n13408 ASIG5V.n13407 0.0202635
R50785 ASIG5V.n231 ASIG5V.n227 0.0202635
R50786 ASIG5V.n7564 ASIG5V.n7563 0.0202635
R50787 ASIG5V.n12487 ASIG5V.n12484 0.0202635
R50788 ASIG5V.n11712 ASIG5V.n11711 0.0202635
R50789 ASIG5V.n11554 ASIG5V.n11552 0.0202635
R50790 ASIG5V.n11630 ASIG5V.n11628 0.0202635
R50791 ASIG5V.n11925 ASIG5V.n11924 0.0202635
R50792 ASIG5V.n12237 ASIG5V.n12236 0.0202635
R50793 ASIG5V.n12580 ASIG5V.n12577 0.0202635
R50794 ASIG5V.n12751 ASIG5V.n12750 0.0202635
R50795 ASIG5V.n7625 ASIG5V.n7624 0.0202635
R50796 ASIG5V.n330 ASIG5V.n327 0.0202635
R50797 ASIG5V.n13494 ASIG5V.n13490 0.0202635
R50798 ASIG5V.n6927 ASIG5V.n6923 0.0202635
R50799 ASIG5V.n7122 ASIG5V.n7121 0.0202635
R50800 ASIG5V.n6148 ASIG5V.n6145 0.0202635
R50801 ASIG5V.n5792 ASIG5V.n5791 0.0202635
R50802 ASIG5V.n5141 ASIG5V.n5140 0.0202635
R50803 ASIG5V.n4846 ASIG5V.n4845 0.0202635
R50804 ASIG5V.n4560 ASIG5V.n4557 0.0202635
R50805 ASIG5V.n4276 ASIG5V.n4275 0.0202635
R50806 ASIG5V.n4003 ASIG5V.n4002 0.0202635
R50807 ASIG5V.n3474 ASIG5V.n3473 0.0202635
R50808 ASIG5V.n3250 ASIG5V.n3249 0.0202635
R50809 ASIG5V.n3131 ASIG5V.n3130 0.0202635
R50810 ASIG5V.n3127 ASIG5V.n3126 0.0202635
R50811 ASIG5V.n3123 ASIG5V.n3122 0.0202635
R50812 ASIG5V.n3119 ASIG5V.n3118 0.0202635
R50813 ASIG5V.n3115 ASIG5V.n3114 0.0202635
R50814 ASIG5V.n3111 ASIG5V.n3110 0.0202635
R50815 ASIG5V.n3107 ASIG5V.n3106 0.0202635
R50816 ASIG5V.n3098 ASIG5V.n3097 0.0202635
R50817 ASIG5V.n3096 ASIG5V.n3095 0.0202635
R50818 ASIG5V.n3093 ASIG5V.n3092 0.0202635
R50819 ASIG5V.n3091 ASIG5V.n3090 0.0202635
R50820 ASIG5V.n3089 ASIG5V.n3088 0.0202635
R50821 ASIG5V.n3085 ASIG5V.n3084 0.0202635
R50822 ASIG5V.n3079 ASIG5V.n3078 0.0202635
R50823 ASIG5V.n3076 ASIG5V.n3075 0.0202635
R50824 ASIG5V.n3072 ASIG5V.n3071 0.0202635
R50825 ASIG5V.n3069 ASIG5V.n3068 0.0202635
R50826 ASIG5V.n3066 ASIG5V.n3065 0.0202635
R50827 ASIG5V.n3063 ASIG5V.n3062 0.0202635
R50828 ASIG5V.n3059 ASIG5V.n3058 0.0202635
R50829 ASIG5V.n3055 ASIG5V.n3054 0.0202635
R50830 ASIG5V.n3051 ASIG5V.n3050 0.0202635
R50831 ASIG5V.n3049 ASIG5V.n3048 0.0202635
R50832 ASIG5V.n3047 ASIG5V.n3046 0.0202635
R50833 ASIG5V.n3044 ASIG5V.n3043 0.0202635
R50834 ASIG5V.n3042 ASIG5V.n3041 0.0202635
R50835 ASIG5V.n3326 ASIG5V.n3325 0.0202635
R50836 ASIG5V.n3322 ASIG5V.n3321 0.0202635
R50837 ASIG5V.n3318 ASIG5V.n3317 0.0202635
R50838 ASIG5V.n3314 ASIG5V.n3313 0.0202635
R50839 ASIG5V.n3310 ASIG5V.n3309 0.0202635
R50840 ASIG5V.n3306 ASIG5V.n3305 0.0202635
R50841 ASIG5V.n3302 ASIG5V.n3301 0.0202635
R50842 ASIG5V.n3261 ASIG5V.n3260 0.0202635
R50843 ASIG5V.n3585 ASIG5V.n3584 0.0202635
R50844 ASIG5V.n3581 ASIG5V.n3580 0.0202635
R50845 ASIG5V.n3577 ASIG5V.n3576 0.0202635
R50846 ASIG5V.n3573 ASIG5V.n3572 0.0202635
R50847 ASIG5V.n3569 ASIG5V.n3568 0.0202635
R50848 ASIG5V.n3565 ASIG5V.n3564 0.0202635
R50849 ASIG5V.n3561 ASIG5V.n3560 0.0202635
R50850 ASIG5V.n3552 ASIG5V.n3550 0.0202635
R50851 ASIG5V.n3549 ASIG5V.n3547 0.0202635
R50852 ASIG5V.n3546 ASIG5V.n3544 0.0202635
R50853 ASIG5V.n3536 ASIG5V.n3533 0.0202635
R50854 ASIG5V.n3505 ASIG5V.n3504 0.0202635
R50855 ASIG5V.n3860 ASIG5V.n3859 0.0202635
R50856 ASIG5V.n3856 ASIG5V.n3855 0.0202635
R50857 ASIG5V.n3852 ASIG5V.n3851 0.0202635
R50858 ASIG5V.n3848 ASIG5V.n3847 0.0202635
R50859 ASIG5V.n3844 ASIG5V.n3843 0.0202635
R50860 ASIG5V.n3840 ASIG5V.n3839 0.0202635
R50861 ASIG5V.n3836 ASIG5V.n3835 0.0202635
R50862 ASIG5V.n3830 ASIG5V.n3829 0.0202635
R50863 ASIG5V.n3828 ASIG5V.n3827 0.0202635
R50864 ASIG5V.n3825 ASIG5V.n3824 0.0202635
R50865 ASIG5V.n3823 ASIG5V.n3822 0.0202635
R50866 ASIG5V.n3821 ASIG5V.n3820 0.0202635
R50867 ASIG5V.n3819 ASIG5V.n3818 0.0202635
R50868 ASIG5V.n3817 ASIG5V.n3816 0.0202635
R50869 ASIG5V.n3813 ASIG5V.n3812 0.0202635
R50870 ASIG5V.n3809 ASIG5V.n3806 0.0202635
R50871 ASIG5V.n3804 ASIG5V.n3803 0.0202635
R50872 ASIG5V.n3801 ASIG5V.n3800 0.0202635
R50873 ASIG5V.n3798 ASIG5V.n3797 0.0202635
R50874 ASIG5V.n3795 ASIG5V.n3794 0.0202635
R50875 ASIG5V.n3792 ASIG5V.n3791 0.0202635
R50876 ASIG5V.n3789 ASIG5V.n3788 0.0202635
R50877 ASIG5V.n3786 ASIG5V.n3785 0.0202635
R50878 ASIG5V.n3782 ASIG5V.n3781 0.0202635
R50879 ASIG5V.n3778 ASIG5V.n3777 0.0202635
R50880 ASIG5V.n3774 ASIG5V.n3773 0.0202635
R50881 ASIG5V.n3771 ASIG5V.n3770 0.0202635
R50882 ASIG5V.n3764 ASIG5V.n3763 0.0202635
R50883 ASIG5V.n3758 ASIG5V.n3757 0.0202635
R50884 ASIG5V.n3754 ASIG5V.n3753 0.0202635
R50885 ASIG5V.n3750 ASIG5V.n3748 0.0202635
R50886 ASIG5V.n4126 ASIG5V.n4125 0.0202635
R50887 ASIG5V.n4122 ASIG5V.n4121 0.0202635
R50888 ASIG5V.n4118 ASIG5V.n4117 0.0202635
R50889 ASIG5V.n4114 ASIG5V.n4113 0.0202635
R50890 ASIG5V.n4110 ASIG5V.n4109 0.0202635
R50891 ASIG5V.n4106 ASIG5V.n4105 0.0202635
R50892 ASIG5V.n4102 ASIG5V.n4101 0.0202635
R50893 ASIG5V.n4085 ASIG5V.n4084 0.0202635
R50894 ASIG5V.n4082 ASIG5V.n4081 0.0202635
R50895 ASIG5V.n4078 ASIG5V.n4077 0.0202635
R50896 ASIG5V.n4074 ASIG5V.n4073 0.0202635
R50897 ASIG5V.n4071 ASIG5V.n4070 0.0202635
R50898 ASIG5V.n4068 ASIG5V.n4067 0.0202635
R50899 ASIG5V.n4065 ASIG5V.n4064 0.0202635
R50900 ASIG5V.n4062 ASIG5V.n4061 0.0202635
R50901 ASIG5V.n4059 ASIG5V.n4058 0.0202635
R50902 ASIG5V.n4056 ASIG5V.n4055 0.0202635
R50903 ASIG5V.n4052 ASIG5V.n4051 0.0202635
R50904 ASIG5V.n4048 ASIG5V.n4047 0.0202635
R50905 ASIG5V.n4044 ASIG5V.n4043 0.0202635
R50906 ASIG5V.n4040 ASIG5V.n4039 0.0202635
R50907 ASIG5V.n4036 ASIG5V.n4035 0.0202635
R50908 ASIG5V.n4033 ASIG5V.n4032 0.0202635
R50909 ASIG5V.n4030 ASIG5V.n4029 0.0202635
R50910 ASIG5V.n4027 ASIG5V.n4026 0.0202635
R50911 ASIG5V.n4023 ASIG5V.n4022 0.0202635
R50912 ASIG5V.n4020 ASIG5V.n4019 0.0202635
R50913 ASIG5V.n4017 ASIG5V.n4016 0.0202635
R50914 ASIG5V.n4014 ASIG5V.n4013 0.0202635
R50915 ASIG5V.n4402 ASIG5V.n4401 0.0202635
R50916 ASIG5V.n4398 ASIG5V.n4397 0.0202635
R50917 ASIG5V.n4394 ASIG5V.n4393 0.0202635
R50918 ASIG5V.n4390 ASIG5V.n4389 0.0202635
R50919 ASIG5V.n4386 ASIG5V.n4385 0.0202635
R50920 ASIG5V.n4382 ASIG5V.n4381 0.0202635
R50921 ASIG5V.n4378 ASIG5V.n4377 0.0202635
R50922 ASIG5V.n4370 ASIG5V.n4369 0.0202635
R50923 ASIG5V.n4368 ASIG5V.n4367 0.0202635
R50924 ASIG5V.n4366 ASIG5V.n4365 0.0202635
R50925 ASIG5V.n4364 ASIG5V.n4363 0.0202635
R50926 ASIG5V.n4362 ASIG5V.n4361 0.0202635
R50927 ASIG5V.n4360 ASIG5V.n4359 0.0202635
R50928 ASIG5V.n4357 ASIG5V.n4356 0.0202635
R50929 ASIG5V.n4353 ASIG5V.n4352 0.0202635
R50930 ASIG5V.n4350 ASIG5V.n4349 0.0202635
R50931 ASIG5V.n4347 ASIG5V.n4346 0.0202635
R50932 ASIG5V.n4344 ASIG5V.n4343 0.0202635
R50933 ASIG5V.n4341 ASIG5V.n4340 0.0202635
R50934 ASIG5V.n4338 ASIG5V.n4337 0.0202635
R50935 ASIG5V.n4335 ASIG5V.n4334 0.0202635
R50936 ASIG5V.n4331 ASIG5V.n4330 0.0202635
R50937 ASIG5V.n4327 ASIG5V.n4326 0.0202635
R50938 ASIG5V.n4323 ASIG5V.n4322 0.0202635
R50939 ASIG5V.n4319 ASIG5V.n4318 0.0202635
R50940 ASIG5V.n4315 ASIG5V.n4314 0.0202635
R50941 ASIG5V.n4311 ASIG5V.n4310 0.0202635
R50942 ASIG5V.n4307 ASIG5V.n4306 0.0202635
R50943 ASIG5V.n4304 ASIG5V.n4303 0.0202635
R50944 ASIG5V.n4301 ASIG5V.n4300 0.0202635
R50945 ASIG5V.n4298 ASIG5V.n4297 0.0202635
R50946 ASIG5V.n4295 ASIG5V.n4294 0.0202635
R50947 ASIG5V.n4291 ASIG5V.n4290 0.0202635
R50948 ASIG5V.n4660 ASIG5V.n4659 0.0202635
R50949 ASIG5V.n4656 ASIG5V.n4655 0.0202635
R50950 ASIG5V.n4652 ASIG5V.n4651 0.0202635
R50951 ASIG5V.n4648 ASIG5V.n4647 0.0202635
R50952 ASIG5V.n4644 ASIG5V.n4643 0.0202635
R50953 ASIG5V.n4640 ASIG5V.n4639 0.0202635
R50954 ASIG5V.n4636 ASIG5V.n4635 0.0202635
R50955 ASIG5V.n4614 ASIG5V.n4613 0.0202635
R50956 ASIG5V.n4609 ASIG5V.n4608 0.0202635
R50957 ASIG5V.n4604 ASIG5V.n4600 0.0202635
R50958 ASIG5V.n4597 ASIG5V.n4596 0.0202635
R50959 ASIG5V.n4590 ASIG5V.n4589 0.0202635
R50960 ASIG5V.n4586 ASIG5V.n4585 0.0202635
R50961 ASIG5V.n4579 ASIG5V.n4578 0.0202635
R50962 ASIG5V.n4574 ASIG5V.n4573 0.0202635
R50963 ASIG5V.n4928 ASIG5V.n4927 0.0202635
R50964 ASIG5V.n4924 ASIG5V.n4923 0.0202635
R50965 ASIG5V.n4920 ASIG5V.n4919 0.0202635
R50966 ASIG5V.n4916 ASIG5V.n4915 0.0202635
R50967 ASIG5V.n4912 ASIG5V.n4911 0.0202635
R50968 ASIG5V.n4908 ASIG5V.n4907 0.0202635
R50969 ASIG5V.n4904 ASIG5V.n4903 0.0202635
R50970 ASIG5V.n4873 ASIG5V.n4872 0.0202635
R50971 ASIG5V.n4868 ASIG5V.n4867 0.0202635
R50972 ASIG5V.n4865 ASIG5V.n4864 0.0202635
R50973 ASIG5V.n4860 ASIG5V.n4859 0.0202635
R50974 ASIG5V.n5355 ASIG5V.n5354 0.0202635
R50975 ASIG5V.n5351 ASIG5V.n5350 0.0202635
R50976 ASIG5V.n5347 ASIG5V.n5346 0.0202635
R50977 ASIG5V.n5343 ASIG5V.n5342 0.0202635
R50978 ASIG5V.n5339 ASIG5V.n5338 0.0202635
R50979 ASIG5V.n5335 ASIG5V.n5334 0.0202635
R50980 ASIG5V.n5331 ASIG5V.n5330 0.0202635
R50981 ASIG5V.n5322 ASIG5V.n5320 0.0202635
R50982 ASIG5V.n5319 ASIG5V.n5317 0.0202635
R50983 ASIG5V.n5316 ASIG5V.n5314 0.0202635
R50984 ASIG5V.n5313 ASIG5V.n5311 0.0202635
R50985 ASIG5V.n5310 ASIG5V.n5308 0.0202635
R50986 ASIG5V.n5307 ASIG5V.n5305 0.0202635
R50987 ASIG5V.n5304 ASIG5V.n5302 0.0202635
R50988 ASIG5V.n5301 ASIG5V.n5299 0.0202635
R50989 ASIG5V.n5298 ASIG5V.n5295 0.0202635
R50990 ASIG5V.n5293 ASIG5V.n5290 0.0202635
R50991 ASIG5V.n5288 ASIG5V.n5287 0.0202635
R50992 ASIG5V.n5285 ASIG5V.n5282 0.0202635
R50993 ASIG5V.n5280 ASIG5V.n5277 0.0202635
R50994 ASIG5V.n5275 ASIG5V.n5272 0.0202635
R50995 ASIG5V.n5270 ASIG5V.n5267 0.0202635
R50996 ASIG5V.n5265 ASIG5V.n5261 0.0202635
R50997 ASIG5V.n5259 ASIG5V.n5255 0.0202635
R50998 ASIG5V.n5252 ASIG5V.n5248 0.0202635
R50999 ASIG5V.n5245 ASIG5V.n5241 0.0202635
R51000 ASIG5V.n5238 ASIG5V.n5234 0.0202635
R51001 ASIG5V.n5231 ASIG5V.n5227 0.0202635
R51002 ASIG5V.n5224 ASIG5V.n5220 0.0202635
R51003 ASIG5V.n5217 ASIG5V.n5213 0.0202635
R51004 ASIG5V.n5210 ASIG5V.n5206 0.0202635
R51005 ASIG5V.n5203 ASIG5V.n5199 0.0202635
R51006 ASIG5V.n5196 ASIG5V.n5192 0.0202635
R51007 ASIG5V.n5189 ASIG5V.n5185 0.0202635
R51008 ASIG5V.n5182 ASIG5V.n5178 0.0202635
R51009 ASIG5V.n5175 ASIG5V.n5172 0.0202635
R51010 ASIG5V.n5170 ASIG5V.n5167 0.0202635
R51011 ASIG5V.n5165 ASIG5V.n5162 0.0202635
R51012 ASIG5V.n5160 ASIG5V.n5157 0.0202635
R51013 ASIG5V.n5586 ASIG5V.n5585 0.0202635
R51014 ASIG5V.n5582 ASIG5V.n5581 0.0202635
R51015 ASIG5V.n5578 ASIG5V.n5577 0.0202635
R51016 ASIG5V.n5574 ASIG5V.n5573 0.0202635
R51017 ASIG5V.n5570 ASIG5V.n5569 0.0202635
R51018 ASIG5V.n5566 ASIG5V.n5565 0.0202635
R51019 ASIG5V.n5562 ASIG5V.n5561 0.0202635
R51020 ASIG5V.n5557 ASIG5V.n5556 0.0202635
R51021 ASIG5V.n5555 ASIG5V.n5554 0.0202635
R51022 ASIG5V.n5553 ASIG5V.n5552 0.0202635
R51023 ASIG5V.n5550 ASIG5V.n5549 0.0202635
R51024 ASIG5V.n5548 ASIG5V.n5546 0.0202635
R51025 ASIG5V.n5545 ASIG5V.n5543 0.0202635
R51026 ASIG5V.n5542 ASIG5V.n5541 0.0202635
R51027 ASIG5V.n5540 ASIG5V.n5539 0.0202635
R51028 ASIG5V.n5537 ASIG5V.n5536 0.0202635
R51029 ASIG5V.n5534 ASIG5V.n5533 0.0202635
R51030 ASIG5V.n5531 ASIG5V.n5530 0.0202635
R51031 ASIG5V.n5528 ASIG5V.n5527 0.0202635
R51032 ASIG5V.n5525 ASIG5V.n5524 0.0202635
R51033 ASIG5V.n5522 ASIG5V.n5521 0.0202635
R51034 ASIG5V.n5519 ASIG5V.n5518 0.0202635
R51035 ASIG5V.n5515 ASIG5V.n5514 0.0202635
R51036 ASIG5V.n5511 ASIG5V.n5510 0.0202635
R51037 ASIG5V.n5507 ASIG5V.n5506 0.0202635
R51038 ASIG5V.n5503 ASIG5V.n5502 0.0202635
R51039 ASIG5V.n5499 ASIG5V.n5498 0.0202635
R51040 ASIG5V.n5493 ASIG5V.n5492 0.0202635
R51041 ASIG5V.n5489 ASIG5V.n5485 0.0202635
R51042 ASIG5V.n5482 ASIG5V.n5481 0.0202635
R51043 ASIG5V.n5478 ASIG5V.n5477 0.0202635
R51044 ASIG5V.n5474 ASIG5V.n5473 0.0202635
R51045 ASIG5V.n5470 ASIG5V.n5466 0.0202635
R51046 ASIG5V.n5463 ASIG5V.n5462 0.0202635
R51047 ASIG5V.n5458 ASIG5V.n5457 0.0202635
R51048 ASIG5V.n5887 ASIG5V.n5886 0.0202635
R51049 ASIG5V.n5883 ASIG5V.n5882 0.0202635
R51050 ASIG5V.n5879 ASIG5V.n5878 0.0202635
R51051 ASIG5V.n5875 ASIG5V.n5874 0.0202635
R51052 ASIG5V.n5871 ASIG5V.n5870 0.0202635
R51053 ASIG5V.n5867 ASIG5V.n5866 0.0202635
R51054 ASIG5V.n5863 ASIG5V.n5862 0.0202635
R51055 ASIG5V.n5824 ASIG5V.n5823 0.0202635
R51056 ASIG5V.n5815 ASIG5V.n5814 0.0202635
R51057 ASIG5V.n509 ASIG5V.n508 0.0202635
R51058 ASIG5V.n505 ASIG5V.n504 0.0202635
R51059 ASIG5V.n501 ASIG5V.n500 0.0202635
R51060 ASIG5V.n497 ASIG5V.n496 0.0202635
R51061 ASIG5V.n493 ASIG5V.n492 0.0202635
R51062 ASIG5V.n489 ASIG5V.n488 0.0202635
R51063 ASIG5V.n485 ASIG5V.n484 0.0202635
R51064 ASIG5V.n6320 ASIG5V.n6318 0.0202635
R51065 ASIG5V.n6317 ASIG5V.n6315 0.0202635
R51066 ASIG5V.n6314 ASIG5V.n6312 0.0202635
R51067 ASIG5V.n6311 ASIG5V.n6309 0.0202635
R51068 ASIG5V.n6308 ASIG5V.n6306 0.0202635
R51069 ASIG5V.n6305 ASIG5V.n6303 0.0202635
R51070 ASIG5V.n6302 ASIG5V.n6300 0.0202635
R51071 ASIG5V.n6299 ASIG5V.n6297 0.0202635
R51072 ASIG5V.n6296 ASIG5V.n6293 0.0202635
R51073 ASIG5V.n6291 ASIG5V.n6288 0.0202635
R51074 ASIG5V.n6286 ASIG5V.n6283 0.0202635
R51075 ASIG5V.n6281 ASIG5V.n6278 0.0202635
R51076 ASIG5V.n6276 ASIG5V.n6273 0.0202635
R51077 ASIG5V.n6271 ASIG5V.n6268 0.0202635
R51078 ASIG5V.n6266 ASIG5V.n6263 0.0202635
R51079 ASIG5V.n6261 ASIG5V.n6257 0.0202635
R51080 ASIG5V.n6254 ASIG5V.n6250 0.0202635
R51081 ASIG5V.n6247 ASIG5V.n6243 0.0202635
R51082 ASIG5V.n6240 ASIG5V.n6236 0.0202635
R51083 ASIG5V.n6233 ASIG5V.n6229 0.0202635
R51084 ASIG5V.n6226 ASIG5V.n6222 0.0202635
R51085 ASIG5V.n6219 ASIG5V.n6215 0.0202635
R51086 ASIG5V.n6212 ASIG5V.n6208 0.0202635
R51087 ASIG5V.n6205 ASIG5V.n6201 0.0202635
R51088 ASIG5V.n6197 ASIG5V.n6196 0.0202635
R51089 ASIG5V.n6193 ASIG5V.n6192 0.0202635
R51090 ASIG5V.n6185 ASIG5V.n6181 0.0202635
R51091 ASIG5V.n6178 ASIG5V.n6177 0.0202635
R51092 ASIG5V.n6174 ASIG5V.n6173 0.0202635
R51093 ASIG5V.n6170 ASIG5V.n6169 0.0202635
R51094 ASIG5V.n6166 ASIG5V.n6165 0.0202635
R51095 ASIG5V.n6962 ASIG5V.n6961 0.0202635
R51096 ASIG5V.n6958 ASIG5V.n6957 0.0202635
R51097 ASIG5V.n6954 ASIG5V.n6953 0.0202635
R51098 ASIG5V.n6950 ASIG5V.n6949 0.0202635
R51099 ASIG5V.n6946 ASIG5V.n6945 0.0202635
R51100 ASIG5V.n6942 ASIG5V.n6941 0.0202635
R51101 ASIG5V.n6938 ASIG5V.n6937 0.0202635
R51102 ASIG5V.n6415 ASIG5V.n6414 0.0202635
R51103 ASIG5V.n6410 ASIG5V.n6409 0.0202635
R51104 ASIG5V.n6406 ASIG5V.n6405 0.0202635
R51105 ASIG5V.n6404 ASIG5V.n6403 0.0202635
R51106 ASIG5V.n6399 ASIG5V.n6398 0.0202635
R51107 ASIG5V.n6396 ASIG5V.n6395 0.0202635
R51108 ASIG5V.n6389 ASIG5V.n6388 0.0202635
R51109 ASIG5V.n6384 ASIG5V.n6383 0.0202635
R51110 ASIG5V.n6380 ASIG5V.n6379 0.0202635
R51111 ASIG5V.n6374 ASIG5V.n6373 0.0202635
R51112 ASIG5V.n6368 ASIG5V.n6364 0.0202635
R51113 ASIG5V.n6361 ASIG5V.n6360 0.0202635
R51114 ASIG5V.n6352 ASIG5V.n6351 0.0202635
R51115 ASIG5V.n6346 ASIG5V.n6345 0.0202635
R51116 ASIG5V.n6342 ASIG5V.n6341 0.0202635
R51117 ASIG5V.n6684 ASIG5V.n6683 0.0202635
R51118 ASIG5V.n6680 ASIG5V.n6679 0.0202635
R51119 ASIG5V.n6676 ASIG5V.n6675 0.0202635
R51120 ASIG5V.n6672 ASIG5V.n6671 0.0202635
R51121 ASIG5V.n6668 ASIG5V.n6667 0.0202635
R51122 ASIG5V.n6664 ASIG5V.n6663 0.0202635
R51123 ASIG5V.n6660 ASIG5V.n6659 0.0202635
R51124 ASIG5V.n6545 ASIG5V.n6544 0.0202635
R51125 ASIG5V.n6540 ASIG5V.n6539 0.0202635
R51126 ASIG5V.n6536 ASIG5V.n6534 0.0202635
R51127 ASIG5V.n6533 ASIG5V.n6532 0.0202635
R51128 ASIG5V.n6531 ASIG5V.n6530 0.0202635
R51129 ASIG5V.n6528 ASIG5V.n6525 0.0202635
R51130 ASIG5V.n6523 ASIG5V.n6522 0.0202635
R51131 ASIG5V.n6520 ASIG5V.n6519 0.0202635
R51132 ASIG5V.n6517 ASIG5V.n6516 0.0202635
R51133 ASIG5V.n6514 ASIG5V.n6513 0.0202635
R51134 ASIG5V.n6511 ASIG5V.n6508 0.0202635
R51135 ASIG5V.n6506 ASIG5V.n6505 0.0202635
R51136 ASIG5V.n6502 ASIG5V.n6501 0.0202635
R51137 ASIG5V.n6498 ASIG5V.n6494 0.0202635
R51138 ASIG5V.n6491 ASIG5V.n6487 0.0202635
R51139 ASIG5V.n6484 ASIG5V.n6483 0.0202635
R51140 ASIG5V.n6479 ASIG5V.n6475 0.0202635
R51141 ASIG5V.n6472 ASIG5V.n6471 0.0202635
R51142 ASIG5V.n6463 ASIG5V.n6459 0.0202635
R51143 ASIG5V.n6456 ASIG5V.n6455 0.0202635
R51144 ASIG5V.n6448 ASIG5V.n6444 0.0202635
R51145 ASIG5V.n6441 ASIG5V.n6440 0.0202635
R51146 ASIG5V.n6429 ASIG5V.n6425 0.0202635
R51147 ASIG5V.n13522 ASIG5V.n13521 0.0202635
R51148 ASIG5V.n13518 ASIG5V.n13517 0.0202635
R51149 ASIG5V.n13514 ASIG5V.n13513 0.0202635
R51150 ASIG5V.n13510 ASIG5V.n13509 0.0202635
R51151 ASIG5V.n13506 ASIG5V.n13505 0.0202635
R51152 ASIG5V.n13502 ASIG5V.n13501 0.0202635
R51153 ASIG5V.n13498 ASIG5V.n13497 0.0202635
R51154 ASIG5V.n98 ASIG5V.n96 0.0202635
R51155 ASIG5V.n95 ASIG5V.n93 0.0202635
R51156 ASIG5V.n92 ASIG5V.n90 0.0202635
R51157 ASIG5V.n89 ASIG5V.n87 0.0202635
R51158 ASIG5V.n86 ASIG5V.n84 0.0202635
R51159 ASIG5V.n83 ASIG5V.n81 0.0202635
R51160 ASIG5V.n80 ASIG5V.n79 0.0202635
R51161 ASIG5V.n78 ASIG5V.n77 0.0202635
R51162 ASIG5V.n75 ASIG5V.n74 0.0202635
R51163 ASIG5V.n72 ASIG5V.n71 0.0202635
R51164 ASIG5V.n69 ASIG5V.n68 0.0202635
R51165 ASIG5V.n66 ASIG5V.n65 0.0202635
R51166 ASIG5V.n63 ASIG5V.n62 0.0202635
R51167 ASIG5V.n60 ASIG5V.n59 0.0202635
R51168 ASIG5V.n53 ASIG5V.n52 0.0202635
R51169 ASIG5V.n49 ASIG5V.n48 0.0202635
R51170 ASIG5V.n40 ASIG5V.n39 0.0202635
R51171 ASIG5V.n33 ASIG5V.n32 0.0202635
R51172 ASIG5V.n24 ASIG5V.n23 0.0202635
R51173 ASIG5V.n15 ASIG5V.n14 0.0202635
R51174 ASIG5V.n11 ASIG5V.n10 0.0202635
R51175 ASIG5V.n358 ASIG5V.n357 0.0202635
R51176 ASIG5V.n354 ASIG5V.n353 0.0202635
R51177 ASIG5V.n350 ASIG5V.n349 0.0202635
R51178 ASIG5V.n346 ASIG5V.n345 0.0202635
R51179 ASIG5V.n342 ASIG5V.n341 0.0202635
R51180 ASIG5V.n338 ASIG5V.n337 0.0202635
R51181 ASIG5V.n334 ASIG5V.n333 0.0202635
R51182 ASIG5V.n7433 ASIG5V.n7432 0.0202635
R51183 ASIG5V.n7429 ASIG5V.n7428 0.0202635
R51184 ASIG5V.n7425 ASIG5V.n7424 0.0202635
R51185 ASIG5V.n7421 ASIG5V.n7420 0.0202635
R51186 ASIG5V.n7417 ASIG5V.n7416 0.0202635
R51187 ASIG5V.n7413 ASIG5V.n7412 0.0202635
R51188 ASIG5V.n7409 ASIG5V.n7408 0.0202635
R51189 ASIG5V.n7395 ASIG5V.n7394 0.0202635
R51190 ASIG5V.n7392 ASIG5V.n7390 0.0202635
R51191 ASIG5V.n7387 ASIG5V.n7386 0.0202635
R51192 ASIG5V.n7385 ASIG5V.n7383 0.0202635
R51193 ASIG5V.n7382 ASIG5V.n7380 0.0202635
R51194 ASIG5V.n7379 ASIG5V.n7378 0.0202635
R51195 ASIG5V.n7377 ASIG5V.n7376 0.0202635
R51196 ASIG5V.n7374 ASIG5V.n7373 0.0202635
R51197 ASIG5V.n7371 ASIG5V.n7370 0.0202635
R51198 ASIG5V.n7368 ASIG5V.n7367 0.0202635
R51199 ASIG5V.n7364 ASIG5V.n7363 0.0202635
R51200 ASIG5V.n7361 ASIG5V.n7360 0.0202635
R51201 ASIG5V.n7357 ASIG5V.n7356 0.0202635
R51202 ASIG5V.n7353 ASIG5V.n7352 0.0202635
R51203 ASIG5V.n7349 ASIG5V.n7348 0.0202635
R51204 ASIG5V.n7341 ASIG5V.n7340 0.0202635
R51205 ASIG5V.n7337 ASIG5V.n7336 0.0202635
R51206 ASIG5V.n7333 ASIG5V.n7329 0.0202635
R51207 ASIG5V.n7326 ASIG5V.n7325 0.0202635
R51208 ASIG5V.n7322 ASIG5V.n7321 0.0202635
R51209 ASIG5V.n7318 ASIG5V.n7317 0.0202635
R51210 ASIG5V.n7314 ASIG5V.n7313 0.0202635
R51211 ASIG5V.n7310 ASIG5V.n7309 0.0202635
R51212 ASIG5V.n7306 ASIG5V.n7302 0.0202635
R51213 ASIG5V.n7299 ASIG5V.n7298 0.0202635
R51214 ASIG5V.n7295 ASIG5V.n7294 0.0202635
R51215 ASIG5V.n7291 ASIG5V.n7290 0.0202635
R51216 ASIG5V.n7288 ASIG5V.n7287 0.0202635
R51217 ASIG5V.n7850 ASIG5V.n7849 0.0202635
R51218 ASIG5V.n7846 ASIG5V.n7845 0.0202635
R51219 ASIG5V.n7842 ASIG5V.n7841 0.0202635
R51220 ASIG5V.n7838 ASIG5V.n7837 0.0202635
R51221 ASIG5V.n7834 ASIG5V.n7833 0.0202635
R51222 ASIG5V.n7830 ASIG5V.n7829 0.0202635
R51223 ASIG5V.n7826 ASIG5V.n7825 0.0202635
R51224 ASIG5V.n7817 ASIG5V.n7815 0.0202635
R51225 ASIG5V.n7814 ASIG5V.n7812 0.0202635
R51226 ASIG5V.n7811 ASIG5V.n7809 0.0202635
R51227 ASIG5V.n7808 ASIG5V.n7806 0.0202635
R51228 ASIG5V.n7805 ASIG5V.n7803 0.0202635
R51229 ASIG5V.n7802 ASIG5V.n7800 0.0202635
R51230 ASIG5V.n7799 ASIG5V.n7797 0.0202635
R51231 ASIG5V.n7796 ASIG5V.n7794 0.0202635
R51232 ASIG5V.n7793 ASIG5V.n7790 0.0202635
R51233 ASIG5V.n7788 ASIG5V.n7785 0.0202635
R51234 ASIG5V.n7783 ASIG5V.n7780 0.0202635
R51235 ASIG5V.n7778 ASIG5V.n7775 0.0202635
R51236 ASIG5V.n7773 ASIG5V.n7770 0.0202635
R51237 ASIG5V.n7768 ASIG5V.n7765 0.0202635
R51238 ASIG5V.n7763 ASIG5V.n7760 0.0202635
R51239 ASIG5V.n7758 ASIG5V.n7754 0.0202635
R51240 ASIG5V.n7752 ASIG5V.n7748 0.0202635
R51241 ASIG5V.n7745 ASIG5V.n7741 0.0202635
R51242 ASIG5V.n7738 ASIG5V.n7734 0.0202635
R51243 ASIG5V.n7731 ASIG5V.n7727 0.0202635
R51244 ASIG5V.n7724 ASIG5V.n7720 0.0202635
R51245 ASIG5V.n7717 ASIG5V.n7713 0.0202635
R51246 ASIG5V.n7710 ASIG5V.n7706 0.0202635
R51247 ASIG5V.n7703 ASIG5V.n7699 0.0202635
R51248 ASIG5V.n7696 ASIG5V.n7692 0.0202635
R51249 ASIG5V.n7689 ASIG5V.n7685 0.0202635
R51250 ASIG5V.n7682 ASIG5V.n7678 0.0202635
R51251 ASIG5V.n7675 ASIG5V.n7671 0.0202635
R51252 ASIG5V.n7668 ASIG5V.n7664 0.0202635
R51253 ASIG5V.n7661 ASIG5V.n7658 0.0202635
R51254 ASIG5V.n7655 ASIG5V.n7652 0.0202635
R51255 ASIG5V.n7650 ASIG5V.n7647 0.0202635
R51256 ASIG5V.n7645 ASIG5V.n7642 0.0202635
R51257 ASIG5V.n7268 ASIG5V.n7267 0.0202635
R51258 ASIG5V.n7264 ASIG5V.n7263 0.0202635
R51259 ASIG5V.n7260 ASIG5V.n7259 0.0202635
R51260 ASIG5V.n7256 ASIG5V.n7255 0.0202635
R51261 ASIG5V.n7252 ASIG5V.n7251 0.0202635
R51262 ASIG5V.n7248 ASIG5V.n7247 0.0202635
R51263 ASIG5V.n7244 ASIG5V.n7243 0.0202635
R51264 ASIG5V.n8116 ASIG5V.n8114 0.0202635
R51265 ASIG5V.n8113 ASIG5V.n8111 0.0202635
R51266 ASIG5V.n8110 ASIG5V.n8109 0.0202635
R51267 ASIG5V.n8108 ASIG5V.n8107 0.0202635
R51268 ASIG5V.n8106 ASIG5V.n8105 0.0202635
R51269 ASIG5V.n8104 ASIG5V.n8103 0.0202635
R51270 ASIG5V.n8102 ASIG5V.n8101 0.0202635
R51271 ASIG5V.n8100 ASIG5V.n8099 0.0202635
R51272 ASIG5V.n8098 ASIG5V.n8097 0.0202635
R51273 ASIG5V.n8095 ASIG5V.n8094 0.0202635
R51274 ASIG5V.n8091 ASIG5V.n8090 0.0202635
R51275 ASIG5V.n8088 ASIG5V.n8087 0.0202635
R51276 ASIG5V.n8085 ASIG5V.n8084 0.0202635
R51277 ASIG5V.n8082 ASIG5V.n8081 0.0202635
R51278 ASIG5V.n8079 ASIG5V.n8078 0.0202635
R51279 ASIG5V.n8076 ASIG5V.n8075 0.0202635
R51280 ASIG5V.n8072 ASIG5V.n8068 0.0202635
R51281 ASIG5V.n8065 ASIG5V.n8061 0.0202635
R51282 ASIG5V.n8058 ASIG5V.n8057 0.0202635
R51283 ASIG5V.n8054 ASIG5V.n8053 0.0202635
R51284 ASIG5V.n8050 ASIG5V.n8049 0.0202635
R51285 ASIG5V.n8046 ASIG5V.n8042 0.0202635
R51286 ASIG5V.n8039 ASIG5V.n8035 0.0202635
R51287 ASIG5V.n8032 ASIG5V.n8031 0.0202635
R51288 ASIG5V.n8028 ASIG5V.n8027 0.0202635
R51289 ASIG5V.n8024 ASIG5V.n8020 0.0202635
R51290 ASIG5V.n8017 ASIG5V.n8016 0.0202635
R51291 ASIG5V.n8013 ASIG5V.n8012 0.0202635
R51292 ASIG5V.n8009 ASIG5V.n8006 0.0202635
R51293 ASIG5V.n8004 ASIG5V.n8001 0.0202635
R51294 ASIG5V.n7999 ASIG5V.n7998 0.0202635
R51295 ASIG5V.n7996 ASIG5V.n7995 0.0202635
R51296 ASIG5V.n12608 ASIG5V.n12607 0.0202635
R51297 ASIG5V.n12604 ASIG5V.n12603 0.0202635
R51298 ASIG5V.n12600 ASIG5V.n12599 0.0202635
R51299 ASIG5V.n12596 ASIG5V.n12595 0.0202635
R51300 ASIG5V.n12592 ASIG5V.n12591 0.0202635
R51301 ASIG5V.n12588 ASIG5V.n12587 0.0202635
R51302 ASIG5V.n12584 ASIG5V.n12583 0.0202635
R51303 ASIG5V.n8185 ASIG5V.n8184 0.0202635
R51304 ASIG5V.n8181 ASIG5V.n8180 0.0202635
R51305 ASIG5V.n8177 ASIG5V.n8176 0.0202635
R51306 ASIG5V.n8173 ASIG5V.n8172 0.0202635
R51307 ASIG5V.n8170 ASIG5V.n8169 0.0202635
R51308 ASIG5V.n8165 ASIG5V.n8164 0.0202635
R51309 ASIG5V.n8159 ASIG5V.n8158 0.0202635
R51310 ASIG5V.n8153 ASIG5V.n8152 0.0202635
R51311 ASIG5V.n8144 ASIG5V.n8143 0.0202635
R51312 ASIG5V.n8140 ASIG5V.n8139 0.0202635
R51313 ASIG5V.n12382 ASIG5V.n12381 0.0202635
R51314 ASIG5V.n12378 ASIG5V.n12377 0.0202635
R51315 ASIG5V.n12374 ASIG5V.n12373 0.0202635
R51316 ASIG5V.n12370 ASIG5V.n12369 0.0202635
R51317 ASIG5V.n12366 ASIG5V.n12365 0.0202635
R51318 ASIG5V.n12362 ASIG5V.n12361 0.0202635
R51319 ASIG5V.n12358 ASIG5V.n12357 0.0202635
R51320 ASIG5V.n8363 ASIG5V.n8361 0.0202635
R51321 ASIG5V.n8360 ASIG5V.n8358 0.0202635
R51322 ASIG5V.n8357 ASIG5V.n8355 0.0202635
R51323 ASIG5V.n8354 ASIG5V.n8352 0.0202635
R51324 ASIG5V.n8351 ASIG5V.n8349 0.0202635
R51325 ASIG5V.n8348 ASIG5V.n8346 0.0202635
R51326 ASIG5V.n8345 ASIG5V.n8343 0.0202635
R51327 ASIG5V.n8342 ASIG5V.n8340 0.0202635
R51328 ASIG5V.n8339 ASIG5V.n8336 0.0202635
R51329 ASIG5V.n8334 ASIG5V.n8331 0.0202635
R51330 ASIG5V.n8329 ASIG5V.n8326 0.0202635
R51331 ASIG5V.n8324 ASIG5V.n8321 0.0202635
R51332 ASIG5V.n8319 ASIG5V.n8316 0.0202635
R51333 ASIG5V.n8314 ASIG5V.n8311 0.0202635
R51334 ASIG5V.n8309 ASIG5V.n8306 0.0202635
R51335 ASIG5V.n8304 ASIG5V.n8301 0.0202635
R51336 ASIG5V.n8299 ASIG5V.n8295 0.0202635
R51337 ASIG5V.n8293 ASIG5V.n8289 0.0202635
R51338 ASIG5V.n8286 ASIG5V.n8282 0.0202635
R51339 ASIG5V.n8279 ASIG5V.n8275 0.0202635
R51340 ASIG5V.n8272 ASIG5V.n8268 0.0202635
R51341 ASIG5V.n8265 ASIG5V.n8261 0.0202635
R51342 ASIG5V.n8258 ASIG5V.n8254 0.0202635
R51343 ASIG5V.n8251 ASIG5V.n8247 0.0202635
R51344 ASIG5V.n8244 ASIG5V.n8240 0.0202635
R51345 ASIG5V.n8237 ASIG5V.n8233 0.0202635
R51346 ASIG5V.n8230 ASIG5V.n8227 0.0202635
R51347 ASIG5V.n8225 ASIG5V.n8222 0.0202635
R51348 ASIG5V.n8220 ASIG5V.n8217 0.0202635
R51349 ASIG5V.n8215 ASIG5V.n8212 0.0202635
R51350 ASIG5V.n8210 ASIG5V.n8207 0.0202635
R51351 ASIG5V.n8205 ASIG5V.n8202 0.0202635
R51352 ASIG5V.n8200 ASIG5V.n8197 0.0202635
R51353 ASIG5V.n12265 ASIG5V.n12264 0.0202635
R51354 ASIG5V.n12261 ASIG5V.n12260 0.0202635
R51355 ASIG5V.n12257 ASIG5V.n12256 0.0202635
R51356 ASIG5V.n12253 ASIG5V.n12252 0.0202635
R51357 ASIG5V.n12249 ASIG5V.n12248 0.0202635
R51358 ASIG5V.n12245 ASIG5V.n12244 0.0202635
R51359 ASIG5V.n12241 ASIG5V.n12240 0.0202635
R51360 ASIG5V.n8489 ASIG5V.n8488 0.0202635
R51361 ASIG5V.n8487 ASIG5V.n8486 0.0202635
R51362 ASIG5V.n8485 ASIG5V.n8483 0.0202635
R51363 ASIG5V.n8482 ASIG5V.n8481 0.0202635
R51364 ASIG5V.n8480 ASIG5V.n8478 0.0202635
R51365 ASIG5V.n8477 ASIG5V.n8475 0.0202635
R51366 ASIG5V.n8474 ASIG5V.n8473 0.0202635
R51367 ASIG5V.n8472 ASIG5V.n8471 0.0202635
R51368 ASIG5V.n8470 ASIG5V.n8467 0.0202635
R51369 ASIG5V.n8465 ASIG5V.n8464 0.0202635
R51370 ASIG5V.n8462 ASIG5V.n8461 0.0202635
R51371 ASIG5V.n8459 ASIG5V.n8456 0.0202635
R51372 ASIG5V.n8454 ASIG5V.n8453 0.0202635
R51373 ASIG5V.n8451 ASIG5V.n8448 0.0202635
R51374 ASIG5V.n8446 ASIG5V.n8445 0.0202635
R51375 ASIG5V.n8443 ASIG5V.n8442 0.0202635
R51376 ASIG5V.n8440 ASIG5V.n8439 0.0202635
R51377 ASIG5V.n8437 ASIG5V.n8436 0.0202635
R51378 ASIG5V.n8434 ASIG5V.n8430 0.0202635
R51379 ASIG5V.n8427 ASIG5V.n8423 0.0202635
R51380 ASIG5V.n8420 ASIG5V.n8419 0.0202635
R51381 ASIG5V.n8416 ASIG5V.n8415 0.0202635
R51382 ASIG5V.n8412 ASIG5V.n8411 0.0202635
R51383 ASIG5V.n8408 ASIG5V.n8404 0.0202635
R51384 ASIG5V.n8401 ASIG5V.n8400 0.0202635
R51385 ASIG5V.n8397 ASIG5V.n8396 0.0202635
R51386 ASIG5V.n8394 ASIG5V.n8393 0.0202635
R51387 ASIG5V.n8391 ASIG5V.n8388 0.0202635
R51388 ASIG5V.n8386 ASIG5V.n8385 0.0202635
R51389 ASIG5V.n8383 ASIG5V.n8380 0.0202635
R51390 ASIG5V.n8378 ASIG5V.n8375 0.0202635
R51391 ASIG5V.n8373 ASIG5V.n8372 0.0202635
R51392 ASIG5V.n8370 ASIG5V.n8368 0.0202635
R51393 ASIG5V.n12112 ASIG5V.n12111 0.0202635
R51394 ASIG5V.n12108 ASIG5V.n12107 0.0202635
R51395 ASIG5V.n12104 ASIG5V.n12103 0.0202635
R51396 ASIG5V.n12100 ASIG5V.n12099 0.0202635
R51397 ASIG5V.n12096 ASIG5V.n12095 0.0202635
R51398 ASIG5V.n12092 ASIG5V.n12091 0.0202635
R51399 ASIG5V.n12088 ASIG5V.n12087 0.0202635
R51400 ASIG5V.n8609 ASIG5V.n8607 0.0202635
R51401 ASIG5V.n8606 ASIG5V.n8605 0.0202635
R51402 ASIG5V.n8604 ASIG5V.n8603 0.0202635
R51403 ASIG5V.n8602 ASIG5V.n8601 0.0202635
R51404 ASIG5V.n8600 ASIG5V.n8599 0.0202635
R51405 ASIG5V.n8598 ASIG5V.n8596 0.0202635
R51406 ASIG5V.n8595 ASIG5V.n8594 0.0202635
R51407 ASIG5V.n8593 ASIG5V.n8592 0.0202635
R51408 ASIG5V.n8591 ASIG5V.n8590 0.0202635
R51409 ASIG5V.n8588 ASIG5V.n8587 0.0202635
R51410 ASIG5V.n8585 ASIG5V.n8584 0.0202635
R51411 ASIG5V.n8582 ASIG5V.n8579 0.0202635
R51412 ASIG5V.n8577 ASIG5V.n8574 0.0202635
R51413 ASIG5V.n8572 ASIG5V.n8571 0.0202635
R51414 ASIG5V.n8569 ASIG5V.n8566 0.0202635
R51415 ASIG5V.n8564 ASIG5V.n8563 0.0202635
R51416 ASIG5V.n8561 ASIG5V.n8560 0.0202635
R51417 ASIG5V.n8558 ASIG5V.n8557 0.0202635
R51418 ASIG5V.n8555 ASIG5V.n8554 0.0202635
R51419 ASIG5V.n8551 ASIG5V.n8547 0.0202635
R51420 ASIG5V.n8544 ASIG5V.n8543 0.0202635
R51421 ASIG5V.n8540 ASIG5V.n8539 0.0202635
R51422 ASIG5V.n8536 ASIG5V.n8532 0.0202635
R51423 ASIG5V.n8529 ASIG5V.n8528 0.0202635
R51424 ASIG5V.n8525 ASIG5V.n8524 0.0202635
R51425 ASIG5V.n8522 ASIG5V.n8519 0.0202635
R51426 ASIG5V.n8517 ASIG5V.n8516 0.0202635
R51427 ASIG5V.n8514 ASIG5V.n8513 0.0202635
R51428 ASIG5V.n8511 ASIG5V.n8508 0.0202635
R51429 ASIG5V.n8506 ASIG5V.n8505 0.0202635
R51430 ASIG5V.n8503 ASIG5V.n8500 0.0202635
R51431 ASIG5V.n8498 ASIG5V.n8496 0.0202635
R51432 ASIG5V.n8494 ASIG5V.n8493 0.0202635
R51433 ASIG5V.n11953 ASIG5V.n11952 0.0202635
R51434 ASIG5V.n11949 ASIG5V.n11948 0.0202635
R51435 ASIG5V.n11945 ASIG5V.n11944 0.0202635
R51436 ASIG5V.n11941 ASIG5V.n11940 0.0202635
R51437 ASIG5V.n11937 ASIG5V.n11936 0.0202635
R51438 ASIG5V.n11933 ASIG5V.n11932 0.0202635
R51439 ASIG5V.n11929 ASIG5V.n11928 0.0202635
R51440 ASIG5V.n8712 ASIG5V.n8710 0.0202635
R51441 ASIG5V.n8709 ASIG5V.n8707 0.0202635
R51442 ASIG5V.n8706 ASIG5V.n8705 0.0202635
R51443 ASIG5V.n8704 ASIG5V.n8703 0.0202635
R51444 ASIG5V.n8702 ASIG5V.n8701 0.0202635
R51445 ASIG5V.n8700 ASIG5V.n8699 0.0202635
R51446 ASIG5V.n8698 ASIG5V.n8697 0.0202635
R51447 ASIG5V.n8696 ASIG5V.n8694 0.0202635
R51448 ASIG5V.n8693 ASIG5V.n8692 0.0202635
R51449 ASIG5V.n8690 ASIG5V.n8689 0.0202635
R51450 ASIG5V.n8687 ASIG5V.n8686 0.0202635
R51451 ASIG5V.n8684 ASIG5V.n8683 0.0202635
R51452 ASIG5V.n8681 ASIG5V.n8680 0.0202635
R51453 ASIG5V.n8678 ASIG5V.n8677 0.0202635
R51454 ASIG5V.n8675 ASIG5V.n8674 0.0202635
R51455 ASIG5V.n8672 ASIG5V.n8671 0.0202635
R51456 ASIG5V.n8669 ASIG5V.n8666 0.0202635
R51457 ASIG5V.n8664 ASIG5V.n8661 0.0202635
R51458 ASIG5V.n8659 ASIG5V.n8658 0.0202635
R51459 ASIG5V.n8656 ASIG5V.n8655 0.0202635
R51460 ASIG5V.n8652 ASIG5V.n8651 0.0202635
R51461 ASIG5V.n8648 ASIG5V.n8647 0.0202635
R51462 ASIG5V.n8644 ASIG5V.n8643 0.0202635
R51463 ASIG5V.n8640 ASIG5V.n8639 0.0202635
R51464 ASIG5V.n8637 ASIG5V.n8636 0.0202635
R51465 ASIG5V.n8634 ASIG5V.n8633 0.0202635
R51466 ASIG5V.n8630 ASIG5V.n8629 0.0202635
R51467 ASIG5V.n8627 ASIG5V.n8626 0.0202635
R51468 ASIG5V.n8624 ASIG5V.n8623 0.0202635
R51469 ASIG5V.n8621 ASIG5V.n8619 0.0202635
R51470 ASIG5V.n8617 ASIG5V.n8616 0.0202635
R51471 ASIG5V.n8615 ASIG5V.n8614 0.0202635
R51472 ASIG5V.n11790 ASIG5V.n11789 0.0202635
R51473 ASIG5V.n11786 ASIG5V.n11785 0.0202635
R51474 ASIG5V.n11782 ASIG5V.n11781 0.0202635
R51475 ASIG5V.n11778 ASIG5V.n11777 0.0202635
R51476 ASIG5V.n11774 ASIG5V.n11773 0.0202635
R51477 ASIG5V.n11770 ASIG5V.n11769 0.0202635
R51478 ASIG5V.n11766 ASIG5V.n11765 0.0202635
R51479 ASIG5V.n8813 ASIG5V.n8812 0.0202635
R51480 ASIG5V.n8811 ASIG5V.n8810 0.0202635
R51481 ASIG5V.n8809 ASIG5V.n8808 0.0202635
R51482 ASIG5V.n8807 ASIG5V.n8806 0.0202635
R51483 ASIG5V.n8805 ASIG5V.n8804 0.0202635
R51484 ASIG5V.n8803 ASIG5V.n8802 0.0202635
R51485 ASIG5V.n8801 ASIG5V.n8799 0.0202635
R51486 ASIG5V.n8798 ASIG5V.n8797 0.0202635
R51487 ASIG5V.n8796 ASIG5V.n8795 0.0202635
R51488 ASIG5V.n8793 ASIG5V.n8790 0.0202635
R51489 ASIG5V.n8788 ASIG5V.n8787 0.0202635
R51490 ASIG5V.n8785 ASIG5V.n8784 0.0202635
R51491 ASIG5V.n8782 ASIG5V.n8781 0.0202635
R51492 ASIG5V.n8779 ASIG5V.n8778 0.0202635
R51493 ASIG5V.n8776 ASIG5V.n8775 0.0202635
R51494 ASIG5V.n8773 ASIG5V.n8772 0.0202635
R51495 ASIG5V.n8770 ASIG5V.n8769 0.0202635
R51496 ASIG5V.n8767 ASIG5V.n8766 0.0202635
R51497 ASIG5V.n8764 ASIG5V.n8761 0.0202635
R51498 ASIG5V.n8759 ASIG5V.n8758 0.0202635
R51499 ASIG5V.n8756 ASIG5V.n8755 0.0202635
R51500 ASIG5V.n8752 ASIG5V.n8751 0.0202635
R51501 ASIG5V.n8749 ASIG5V.n8748 0.0202635
R51502 ASIG5V.n8746 ASIG5V.n8745 0.0202635
R51503 ASIG5V.n8743 ASIG5V.n8742 0.0202635
R51504 ASIG5V.n8740 ASIG5V.n8739 0.0202635
R51505 ASIG5V.n8737 ASIG5V.n8736 0.0202635
R51506 ASIG5V.n8734 ASIG5V.n8733 0.0202635
R51507 ASIG5V.n8731 ASIG5V.n8730 0.0202635
R51508 ASIG5V.n8728 ASIG5V.n8727 0.0202635
R51509 ASIG5V.n8725 ASIG5V.n8724 0.0202635
R51510 ASIG5V.n8723 ASIG5V.n8721 0.0202635
R51511 ASIG5V.n11661 ASIG5V.n11660 0.0202635
R51512 ASIG5V.n11657 ASIG5V.n11656 0.0202635
R51513 ASIG5V.n11653 ASIG5V.n11652 0.0202635
R51514 ASIG5V.n11649 ASIG5V.n11648 0.0202635
R51515 ASIG5V.n11645 ASIG5V.n11644 0.0202635
R51516 ASIG5V.n11641 ASIG5V.n11640 0.0202635
R51517 ASIG5V.n11637 ASIG5V.n11636 0.0202635
R51518 ASIG5V.n11422 ASIG5V.n11420 0.0202635
R51519 ASIG5V.n8853 ASIG5V.n8851 0.0202635
R51520 ASIG5V.n8816 ASIG5V.n8814 0.0202635
R51521 ASIG5V.n8715 ASIG5V.n8713 0.0202635
R51522 ASIG5V.n12153 ASIG5V.n12151 0.0202635
R51523 ASIG5V.n12309 ASIG5V.n12307 0.0202635
R51524 ASIG5V.n12424 ASIG5V.n12421 0.0202635
R51525 ASIG5V.n8190 ASIG5V.n8187 0.0202635
R51526 ASIG5V.n8125 ASIG5V.n8122 0.0202635
R51527 ASIG5V.n7822 ASIG5V.n7819 0.0202635
R51528 ASIG5V.n7400 ASIG5V.n7397 0.0202635
R51529 ASIG5V.n144 ASIG5V.n141 0.0202635
R51530 ASIG5V.n103 ASIG5V.n100 0.0202635
R51531 ASIG5V.n6776 ASIG5V.n6772 0.0202635
R51532 ASIG5V.n6418 ASIG5V.n6417 0.0202635
R51533 ASIG5V.n6325 ASIG5V.n6322 0.0202635
R51534 ASIG5V.n5977 ASIG5V.n5974 0.0202635
R51535 ASIG5V.n5681 ASIG5V.n5678 0.0202635
R51536 ASIG5V.n5327 ASIG5V.n5324 0.0202635
R51537 ASIG5V.n4976 ASIG5V.n4973 0.0202635
R51538 ASIG5V.n4701 ASIG5V.n4699 0.0202635
R51539 ASIG5V.n4449 ASIG5V.n4447 0.0202635
R51540 ASIG5V.n4095 ASIG5V.n4094 0.0202635
R51541 ASIG5V.n3832 ASIG5V.n3831 0.0202635
R51542 ASIG5V.n3557 ASIG5V.n3555 0.0202635
R51543 ASIG5V.n3334 ASIG5V.n3332 0.0202635
R51544 ASIG5V.n3142 ASIG5V.n3140 0.0202635
R51545 ASIG5V.n11485 ASIG5V.n11483 0.0202635
R51546 ASIG5V.n1015 ASIG5V.n1014 0.020075
R51547 ASIG5V.n3128 ASIG5V.n3127 0.0200092
R51548 ASIG5V.n3124 ASIG5V.n3123 0.0200092
R51549 ASIG5V.n3116 ASIG5V.n3115 0.0200092
R51550 ASIG5V.n3112 ASIG5V.n3111 0.0200092
R51551 ASIG5V.n3197 ASIG5V.n3196 0.0200092
R51552 ASIG5V.n3200 ASIG5V.n3199 0.0200092
R51553 ASIG5V.n3214 ASIG5V.n3213 0.0200092
R51554 ASIG5V.n3219 ASIG5V.n3218 0.0200092
R51555 ASIG5V.n3236 ASIG5V.n3235 0.0200092
R51556 ASIG5V.n3244 ASIG5V.n3243 0.0200092
R51557 ASIG5V.n3323 ASIG5V.n3322 0.0200092
R51558 ASIG5V.n3319 ASIG5V.n3318 0.0200092
R51559 ASIG5V.n3311 ASIG5V.n3310 0.0200092
R51560 ASIG5V.n3307 ASIG5V.n3306 0.0200092
R51561 ASIG5V.n3402 ASIG5V.n3401 0.0200092
R51562 ASIG5V.n3405 ASIG5V.n3404 0.0200092
R51563 ASIG5V.n3408 ASIG5V.n3407 0.0200092
R51564 ASIG5V.n3411 ASIG5V.n3410 0.0200092
R51565 ASIG5V.n3414 ASIG5V.n3413 0.0200092
R51566 ASIG5V.n3419 ASIG5V.n3418 0.0200092
R51567 ASIG5V.n3424 ASIG5V.n3423 0.0200092
R51568 ASIG5V.n3429 ASIG5V.n3428 0.0200092
R51569 ASIG5V.n3434 ASIG5V.n3433 0.0200092
R51570 ASIG5V.n3439 ASIG5V.n3438 0.0200092
R51571 ASIG5V.n3444 ASIG5V.n3443 0.0200092
R51572 ASIG5V.n3449 ASIG5V.n3448 0.0200092
R51573 ASIG5V.n3454 ASIG5V.n3453 0.0200092
R51574 ASIG5V.n3459 ASIG5V.n3458 0.0200092
R51575 ASIG5V.n3464 ASIG5V.n3463 0.0200092
R51576 ASIG5V.n3469 ASIG5V.n3468 0.0200092
R51577 ASIG5V.n3472 ASIG5V.n3471 0.0200092
R51578 ASIG5V.n3582 ASIG5V.n3581 0.0200092
R51579 ASIG5V.n3578 ASIG5V.n3577 0.0200092
R51580 ASIG5V.n3570 ASIG5V.n3569 0.0200092
R51581 ASIG5V.n3566 ASIG5V.n3565 0.0200092
R51582 ASIG5V.n3682 ASIG5V.n3681 0.0200092
R51583 ASIG5V.n3687 ASIG5V.n3686 0.0200092
R51584 ASIG5V.n3690 ASIG5V.n3689 0.0200092
R51585 ASIG5V.n3696 ASIG5V.n3695 0.0200092
R51586 ASIG5V.n3701 ASIG5V.n3700 0.0200092
R51587 ASIG5V.n3704 ASIG5V.n3703 0.0200092
R51588 ASIG5V.n3707 ASIG5V.n3706 0.0200092
R51589 ASIG5V.n3712 ASIG5V.n3711 0.0200092
R51590 ASIG5V.n3715 ASIG5V.n3714 0.0200092
R51591 ASIG5V.n3720 ASIG5V.n3719 0.0200092
R51592 ASIG5V.n3725 ASIG5V.n3724 0.0200092
R51593 ASIG5V.n3728 ASIG5V.n3727 0.0200092
R51594 ASIG5V.n3731 ASIG5V.n3730 0.0200092
R51595 ASIG5V.n3734 ASIG5V.n3733 0.0200092
R51596 ASIG5V.n3736 ASIG5V.n3735 0.0200092
R51597 ASIG5V.n3857 ASIG5V.n3856 0.0200092
R51598 ASIG5V.n3853 ASIG5V.n3852 0.0200092
R51599 ASIG5V.n3845 ASIG5V.n3844 0.0200092
R51600 ASIG5V.n3841 ASIG5V.n3840 0.0200092
R51601 ASIG5V.n3953 ASIG5V.n3952 0.0200092
R51602 ASIG5V.n3961 ASIG5V.n3960 0.0200092
R51603 ASIG5V.n3966 ASIG5V.n3965 0.0200092
R51604 ASIG5V.n3992 ASIG5V.n3991 0.0200092
R51605 ASIG5V.n4001 ASIG5V.n4000 0.0200092
R51606 ASIG5V.n4123 ASIG5V.n4122 0.0200092
R51607 ASIG5V.n4119 ASIG5V.n4118 0.0200092
R51608 ASIG5V.n4111 ASIG5V.n4110 0.0200092
R51609 ASIG5V.n4107 ASIG5V.n4106 0.0200092
R51610 ASIG5V.n4220 ASIG5V.n4219 0.0200092
R51611 ASIG5V.n4223 ASIG5V.n4222 0.0200092
R51612 ASIG5V.n4226 ASIG5V.n4225 0.0200092
R51613 ASIG5V.n4229 ASIG5V.n4228 0.0200092
R51614 ASIG5V.n4239 ASIG5V.n4238 0.0200092
R51615 ASIG5V.n4271 ASIG5V.n4270 0.0200092
R51616 ASIG5V.n4399 ASIG5V.n4398 0.0200092
R51617 ASIG5V.n4395 ASIG5V.n4394 0.0200092
R51618 ASIG5V.n4387 ASIG5V.n4386 0.0200092
R51619 ASIG5V.n4383 ASIG5V.n4382 0.0200092
R51620 ASIG5V.n4503 ASIG5V.n4502 0.0200092
R51621 ASIG5V.n4506 ASIG5V.n4505 0.0200092
R51622 ASIG5V.n4531 ASIG5V.n4530 0.0200092
R51623 ASIG5V.n4560 ASIG5V.n4559 0.0200092
R51624 ASIG5V.n4657 ASIG5V.n4656 0.0200092
R51625 ASIG5V.n4653 ASIG5V.n4652 0.0200092
R51626 ASIG5V.n4645 ASIG5V.n4644 0.0200092
R51627 ASIG5V.n4641 ASIG5V.n4640 0.0200092
R51628 ASIG5V.n4770 ASIG5V.n4769 0.0200092
R51629 ASIG5V.n4773 ASIG5V.n4772 0.0200092
R51630 ASIG5V.n4776 ASIG5V.n4775 0.0200092
R51631 ASIG5V.n4779 ASIG5V.n4778 0.0200092
R51632 ASIG5V.n4783 ASIG5V.n4782 0.0200092
R51633 ASIG5V.n4788 ASIG5V.n4787 0.0200092
R51634 ASIG5V.n4793 ASIG5V.n4792 0.0200092
R51635 ASIG5V.n4801 ASIG5V.n4800 0.0200092
R51636 ASIG5V.n4808 ASIG5V.n4807 0.0200092
R51637 ASIG5V.n4819 ASIG5V.n4818 0.0200092
R51638 ASIG5V.n4826 ASIG5V.n4825 0.0200092
R51639 ASIG5V.n4835 ASIG5V.n4834 0.0200092
R51640 ASIG5V.n4840 ASIG5V.n4839 0.0200092
R51641 ASIG5V.n4925 ASIG5V.n4924 0.0200092
R51642 ASIG5V.n4921 ASIG5V.n4920 0.0200092
R51643 ASIG5V.n4913 ASIG5V.n4912 0.0200092
R51644 ASIG5V.n4909 ASIG5V.n4908 0.0200092
R51645 ASIG5V.n5060 ASIG5V.n5059 0.0200092
R51646 ASIG5V.n5063 ASIG5V.n5062 0.0200092
R51647 ASIG5V.n5066 ASIG5V.n5065 0.0200092
R51648 ASIG5V.n5069 ASIG5V.n5068 0.0200092
R51649 ASIG5V.n5073 ASIG5V.n5072 0.0200092
R51650 ASIG5V.n5078 ASIG5V.n5077 0.0200092
R51651 ASIG5V.n5083 ASIG5V.n5082 0.0200092
R51652 ASIG5V.n5088 ASIG5V.n5087 0.0200092
R51653 ASIG5V.n5093 ASIG5V.n5092 0.0200092
R51654 ASIG5V.n5100 ASIG5V.n5099 0.0200092
R51655 ASIG5V.n5107 ASIG5V.n5106 0.0200092
R51656 ASIG5V.n5114 ASIG5V.n5113 0.0200092
R51657 ASIG5V.n5121 ASIG5V.n5120 0.0200092
R51658 ASIG5V.n5128 ASIG5V.n5127 0.0200092
R51659 ASIG5V.n5352 ASIG5V.n5351 0.0200092
R51660 ASIG5V.n5348 ASIG5V.n5347 0.0200092
R51661 ASIG5V.n5340 ASIG5V.n5339 0.0200092
R51662 ASIG5V.n5336 ASIG5V.n5335 0.0200092
R51663 ASIG5V.n5441 ASIG5V.n5440 0.0200092
R51664 ASIG5V.n5583 ASIG5V.n5582 0.0200092
R51665 ASIG5V.n5579 ASIG5V.n5578 0.0200092
R51666 ASIG5V.n5571 ASIG5V.n5570 0.0200092
R51667 ASIG5V.n5567 ASIG5V.n5566 0.0200092
R51668 ASIG5V.n5772 ASIG5V.n5771 0.0200092
R51669 ASIG5V.n5779 ASIG5V.n5778 0.0200092
R51670 ASIG5V.n5884 ASIG5V.n5883 0.0200092
R51671 ASIG5V.n5880 ASIG5V.n5879 0.0200092
R51672 ASIG5V.n5872 ASIG5V.n5871 0.0200092
R51673 ASIG5V.n5868 ASIG5V.n5867 0.0200092
R51674 ASIG5V.n6065 ASIG5V.n6064 0.0200092
R51675 ASIG5V.n6068 ASIG5V.n6067 0.0200092
R51676 ASIG5V.n6071 ASIG5V.n6070 0.0200092
R51677 ASIG5V.n6074 ASIG5V.n6073 0.0200092
R51678 ASIG5V.n6078 ASIG5V.n6077 0.0200092
R51679 ASIG5V.n6083 ASIG5V.n6082 0.0200092
R51680 ASIG5V.n6088 ASIG5V.n6087 0.0200092
R51681 ASIG5V.n6093 ASIG5V.n6092 0.0200092
R51682 ASIG5V.n6099 ASIG5V.n6098 0.0200092
R51683 ASIG5V.n6106 ASIG5V.n6105 0.0200092
R51684 ASIG5V.n6113 ASIG5V.n6112 0.0200092
R51685 ASIG5V.n6120 ASIG5V.n6119 0.0200092
R51686 ASIG5V.n6127 ASIG5V.n6126 0.0200092
R51687 ASIG5V.n6134 ASIG5V.n6133 0.0200092
R51688 ASIG5V.n6142 ASIG5V.n6141 0.0200092
R51689 ASIG5V.n6148 ASIG5V.n6147 0.0200092
R51690 ASIG5V.n506 ASIG5V.n505 0.0200092
R51691 ASIG5V.n502 ASIG5V.n501 0.0200092
R51692 ASIG5V.n494 ASIG5V.n493 0.0200092
R51693 ASIG5V.n490 ASIG5V.n489 0.0200092
R51694 ASIG5V.n6959 ASIG5V.n6958 0.0200092
R51695 ASIG5V.n6955 ASIG5V.n6954 0.0200092
R51696 ASIG5V.n6947 ASIG5V.n6946 0.0200092
R51697 ASIG5V.n6943 ASIG5V.n6942 0.0200092
R51698 ASIG5V.n6831 ASIG5V.n6830 0.0200092
R51699 ASIG5V.n6834 ASIG5V.n6833 0.0200092
R51700 ASIG5V.n6837 ASIG5V.n6836 0.0200092
R51701 ASIG5V.n6840 ASIG5V.n6839 0.0200092
R51702 ASIG5V.n6844 ASIG5V.n6843 0.0200092
R51703 ASIG5V.n6849 ASIG5V.n6848 0.0200092
R51704 ASIG5V.n6854 ASIG5V.n6853 0.0200092
R51705 ASIG5V.n6859 ASIG5V.n6858 0.0200092
R51706 ASIG5V.n6864 ASIG5V.n6863 0.0200092
R51707 ASIG5V.n6871 ASIG5V.n6870 0.0200092
R51708 ASIG5V.n6878 ASIG5V.n6877 0.0200092
R51709 ASIG5V.n6885 ASIG5V.n6884 0.0200092
R51710 ASIG5V.n6892 ASIG5V.n6891 0.0200092
R51711 ASIG5V.n6899 ASIG5V.n6898 0.0200092
R51712 ASIG5V.n6906 ASIG5V.n6905 0.0200092
R51713 ASIG5V.n6913 ASIG5V.n6912 0.0200092
R51714 ASIG5V.n6920 ASIG5V.n6919 0.0200092
R51715 ASIG5V.n6927 ASIG5V.n6926 0.0200092
R51716 ASIG5V.n6681 ASIG5V.n6680 0.0200092
R51717 ASIG5V.n6677 ASIG5V.n6676 0.0200092
R51718 ASIG5V.n6669 ASIG5V.n6668 0.0200092
R51719 ASIG5V.n6665 ASIG5V.n6664 0.0200092
R51720 ASIG5V.n6618 ASIG5V.n6617 0.0200092
R51721 ASIG5V.n6621 ASIG5V.n6620 0.0200092
R51722 ASIG5V.n6624 ASIG5V.n6623 0.0200092
R51723 ASIG5V.n6627 ASIG5V.n6626 0.0200092
R51724 ASIG5V.n13519 ASIG5V.n13518 0.0200092
R51725 ASIG5V.n13515 ASIG5V.n13514 0.0200092
R51726 ASIG5V.n13507 ASIG5V.n13506 0.0200092
R51727 ASIG5V.n13503 ASIG5V.n13502 0.0200092
R51728 ASIG5V.n13416 ASIG5V.n13415 0.0200092
R51729 ASIG5V.n13431 ASIG5V.n13430 0.0200092
R51730 ASIG5V.n13438 ASIG5V.n13437 0.0200092
R51731 ASIG5V.n13445 ASIG5V.n13444 0.0200092
R51732 ASIG5V.n13452 ASIG5V.n13451 0.0200092
R51733 ASIG5V.n13459 ASIG5V.n13458 0.0200092
R51734 ASIG5V.n13466 ASIG5V.n13465 0.0200092
R51735 ASIG5V.n13473 ASIG5V.n13472 0.0200092
R51736 ASIG5V.n13480 ASIG5V.n13479 0.0200092
R51737 ASIG5V.n13487 ASIG5V.n13486 0.0200092
R51738 ASIG5V.n13494 ASIG5V.n13493 0.0200092
R51739 ASIG5V.n355 ASIG5V.n354 0.0200092
R51740 ASIG5V.n351 ASIG5V.n350 0.0200092
R51741 ASIG5V.n343 ASIG5V.n342 0.0200092
R51742 ASIG5V.n339 ASIG5V.n338 0.0200092
R51743 ASIG5V.n234 ASIG5V.n233 0.0200092
R51744 ASIG5V.n237 ASIG5V.n236 0.0200092
R51745 ASIG5V.n240 ASIG5V.n239 0.0200092
R51746 ASIG5V.n243 ASIG5V.n242 0.0200092
R51747 ASIG5V.n247 ASIG5V.n246 0.0200092
R51748 ASIG5V.n252 ASIG5V.n251 0.0200092
R51749 ASIG5V.n257 ASIG5V.n256 0.0200092
R51750 ASIG5V.n262 ASIG5V.n261 0.0200092
R51751 ASIG5V.n268 ASIG5V.n267 0.0200092
R51752 ASIG5V.n275 ASIG5V.n274 0.0200092
R51753 ASIG5V.n282 ASIG5V.n281 0.0200092
R51754 ASIG5V.n289 ASIG5V.n288 0.0200092
R51755 ASIG5V.n296 ASIG5V.n295 0.0200092
R51756 ASIG5V.n303 ASIG5V.n302 0.0200092
R51757 ASIG5V.n310 ASIG5V.n309 0.0200092
R51758 ASIG5V.n317 ASIG5V.n316 0.0200092
R51759 ASIG5V.n324 ASIG5V.n323 0.0200092
R51760 ASIG5V.n330 ASIG5V.n329 0.0200092
R51761 ASIG5V.n7430 ASIG5V.n7429 0.0200092
R51762 ASIG5V.n7426 ASIG5V.n7425 0.0200092
R51763 ASIG5V.n7418 ASIG5V.n7417 0.0200092
R51764 ASIG5V.n7414 ASIG5V.n7413 0.0200092
R51765 ASIG5V.n7567 ASIG5V.n7566 0.0200092
R51766 ASIG5V.n7582 ASIG5V.n7581 0.0200092
R51767 ASIG5V.n7590 ASIG5V.n7589 0.0200092
R51768 ASIG5V.n7601 ASIG5V.n7600 0.0200092
R51769 ASIG5V.n7847 ASIG5V.n7846 0.0200092
R51770 ASIG5V.n7843 ASIG5V.n7842 0.0200092
R51771 ASIG5V.n7835 ASIG5V.n7834 0.0200092
R51772 ASIG5V.n7831 ASIG5V.n7830 0.0200092
R51773 ASIG5V.n7265 ASIG5V.n7264 0.0200092
R51774 ASIG5V.n7261 ASIG5V.n7260 0.0200092
R51775 ASIG5V.n7253 ASIG5V.n7252 0.0200092
R51776 ASIG5V.n7249 ASIG5V.n7248 0.0200092
R51777 ASIG5V.n12605 ASIG5V.n12604 0.0200092
R51778 ASIG5V.n12601 ASIG5V.n12600 0.0200092
R51779 ASIG5V.n12593 ASIG5V.n12592 0.0200092
R51780 ASIG5V.n12589 ASIG5V.n12588 0.0200092
R51781 ASIG5V.n12490 ASIG5V.n12489 0.0200092
R51782 ASIG5V.n12493 ASIG5V.n12492 0.0200092
R51783 ASIG5V.n12496 ASIG5V.n12495 0.0200092
R51784 ASIG5V.n12499 ASIG5V.n12498 0.0200092
R51785 ASIG5V.n12503 ASIG5V.n12502 0.0200092
R51786 ASIG5V.n12508 ASIG5V.n12507 0.0200092
R51787 ASIG5V.n12513 ASIG5V.n12512 0.0200092
R51788 ASIG5V.n12518 ASIG5V.n12517 0.0200092
R51789 ASIG5V.n12523 ASIG5V.n12522 0.0200092
R51790 ASIG5V.n12530 ASIG5V.n12529 0.0200092
R51791 ASIG5V.n12537 ASIG5V.n12536 0.0200092
R51792 ASIG5V.n12544 ASIG5V.n12543 0.0200092
R51793 ASIG5V.n12551 ASIG5V.n12550 0.0200092
R51794 ASIG5V.n12558 ASIG5V.n12557 0.0200092
R51795 ASIG5V.n12565 ASIG5V.n12564 0.0200092
R51796 ASIG5V.n12570 ASIG5V.n12569 0.0200092
R51797 ASIG5V.n12575 ASIG5V.n12574 0.0200092
R51798 ASIG5V.n12580 ASIG5V.n12579 0.0200092
R51799 ASIG5V.n12379 ASIG5V.n12378 0.0200092
R51800 ASIG5V.n12375 ASIG5V.n12374 0.0200092
R51801 ASIG5V.n12367 ASIG5V.n12366 0.0200092
R51802 ASIG5V.n12363 ASIG5V.n12362 0.0200092
R51803 ASIG5V.n12262 ASIG5V.n12261 0.0200092
R51804 ASIG5V.n12258 ASIG5V.n12257 0.0200092
R51805 ASIG5V.n12250 ASIG5V.n12249 0.0200092
R51806 ASIG5V.n12246 ASIG5V.n12245 0.0200092
R51807 ASIG5V.n12109 ASIG5V.n12108 0.0200092
R51808 ASIG5V.n12105 ASIG5V.n12104 0.0200092
R51809 ASIG5V.n12097 ASIG5V.n12096 0.0200092
R51810 ASIG5V.n12093 ASIG5V.n12092 0.0200092
R51811 ASIG5V.n11950 ASIG5V.n11949 0.0200092
R51812 ASIG5V.n11946 ASIG5V.n11945 0.0200092
R51813 ASIG5V.n11938 ASIG5V.n11937 0.0200092
R51814 ASIG5V.n11934 ASIG5V.n11933 0.0200092
R51815 ASIG5V.n11917 ASIG5V.n11916 0.0200092
R51816 ASIG5V.n11787 ASIG5V.n11786 0.0200092
R51817 ASIG5V.n11783 ASIG5V.n11782 0.0200092
R51818 ASIG5V.n11775 ASIG5V.n11774 0.0200092
R51819 ASIG5V.n11771 ASIG5V.n11770 0.0200092
R51820 ASIG5V.n11759 ASIG5V.n11758 0.0200092
R51821 ASIG5V.n11658 ASIG5V.n11657 0.0200092
R51822 ASIG5V.n11654 ASIG5V.n11653 0.0200092
R51823 ASIG5V.n11646 ASIG5V.n11645 0.0200092
R51824 ASIG5V.n11642 ASIG5V.n11641 0.0200092
R51825 ASIG5V.n11557 ASIG5V.n11556 0.0200092
R51826 ASIG5V.n11560 ASIG5V.n11559 0.0200092
R51827 ASIG5V.n11563 ASIG5V.n11562 0.0200092
R51828 ASIG5V.n11566 ASIG5V.n11565 0.0200092
R51829 ASIG5V.n11569 ASIG5V.n11568 0.0200092
R51830 ASIG5V.n11574 ASIG5V.n11573 0.0200092
R51831 ASIG5V.n11579 ASIG5V.n11578 0.0200092
R51832 ASIG5V.n11584 ASIG5V.n11583 0.0200092
R51833 ASIG5V.n11589 ASIG5V.n11588 0.0200092
R51834 ASIG5V.n11594 ASIG5V.n11593 0.0200092
R51835 ASIG5V.n11599 ASIG5V.n11598 0.0200092
R51836 ASIG5V.n11604 ASIG5V.n11603 0.0200092
R51837 ASIG5V.n11609 ASIG5V.n11608 0.0200092
R51838 ASIG5V.n11614 ASIG5V.n11613 0.0200092
R51839 ASIG5V.n11619 ASIG5V.n11618 0.0200092
R51840 ASIG5V.n11624 ASIG5V.n11623 0.0200092
R51841 ASIG5V.n11627 ASIG5V.n11626 0.0200092
R51842 ASIG5V.n11630 ASIG5V.n11629 0.0200092
R51843 ASIG5V.n3142 ASIG5V.n3141 0.0200092
R51844 ASIG5V.n3334 ASIG5V.n3333 0.0200092
R51845 ASIG5V.n3628 ASIG5V.n3627 0.0200092
R51846 ASIG5V.n3901 ASIG5V.n3900 0.0200092
R51847 ASIG5V.n4166 ASIG5V.n4165 0.0200092
R51848 ASIG5V.n4449 ASIG5V.n4448 0.0200092
R51849 ASIG5V.n4701 ASIG5V.n4700 0.0200092
R51850 ASIG5V.n4976 ASIG5V.n4975 0.0200092
R51851 ASIG5V.n5401 ASIG5V.n5400 0.0200092
R51852 ASIG5V.n5681 ASIG5V.n5680 0.0200092
R51853 ASIG5V.n5977 ASIG5V.n5976 0.0200092
R51854 ASIG5V.n6334 ASIG5V.n6333 0.0200092
R51855 ASIG5V.n6548 ASIG5V.n6547 0.0200092
R51856 ASIG5V.n103 ASIG5V.n102 0.0200092
R51857 ASIG5V.n144 ASIG5V.n143 0.0200092
R51858 ASIG5V.n7522 ASIG5V.n7521 0.0200092
R51859 ASIG5V.n7944 ASIG5V.n7943 0.0200092
R51860 ASIG5V.n8125 ASIG5V.n8124 0.0200092
R51861 ASIG5V.n8190 ASIG5V.n8189 0.0200092
R51862 ASIG5V.n8365 ASIG5V.n8364 0.0200092
R51863 ASIG5V.n8491 ASIG5V.n8490 0.0200092
R51864 ASIG5V.n8611 ASIG5V.n8610 0.0200092
R51865 ASIG5V.n8715 ASIG5V.n8714 0.0200092
R51866 ASIG5V.n8816 ASIG5V.n8815 0.0200092
R51867 ASIG5V.n8853 ASIG5V.n8852 0.0200092
R51868 ASIG5V.n3133 ASIG5V.n3132 0.0200092
R51869 ASIG5V.n3328 ASIG5V.n3327 0.0200092
R51870 ASIG5V.n3587 ASIG5V.n3586 0.0200092
R51871 ASIG5V.n3862 ASIG5V.n3861 0.0200092
R51872 ASIG5V.n4128 ASIG5V.n4127 0.0200092
R51873 ASIG5V.n4404 ASIG5V.n4403 0.0200092
R51874 ASIG5V.n4662 ASIG5V.n4661 0.0200092
R51875 ASIG5V.n4930 ASIG5V.n4929 0.0200092
R51876 ASIG5V.n5357 ASIG5V.n5356 0.0200092
R51877 ASIG5V.n5588 ASIG5V.n5587 0.0200092
R51878 ASIG5V.n5889 ASIG5V.n5888 0.0200092
R51879 ASIG5V.n511 ASIG5V.n510 0.0200092
R51880 ASIG5V.n6964 ASIG5V.n6963 0.0200092
R51881 ASIG5V.n6686 ASIG5V.n6685 0.0200092
R51882 ASIG5V.n13524 ASIG5V.n13523 0.0200092
R51883 ASIG5V.n360 ASIG5V.n359 0.0200092
R51884 ASIG5V.n7435 ASIG5V.n7434 0.0200092
R51885 ASIG5V.n7852 ASIG5V.n7851 0.0200092
R51886 ASIG5V.n7270 ASIG5V.n7269 0.0200092
R51887 ASIG5V.n12610 ASIG5V.n12609 0.0200092
R51888 ASIG5V.n12384 ASIG5V.n12383 0.0200092
R51889 ASIG5V.n12267 ASIG5V.n12266 0.0200092
R51890 ASIG5V.n12114 ASIG5V.n12113 0.0200092
R51891 ASIG5V.n11955 ASIG5V.n11954 0.0200092
R51892 ASIG5V.n11792 ASIG5V.n11791 0.0200092
R51893 ASIG5V.n11663 ASIG5V.n11662 0.0200092
R51894 ASIG5V.n11660 ASIG5V.n11659 0.0200092
R51895 ASIG5V.n11789 ASIG5V.n11788 0.0200092
R51896 ASIG5V.n11952 ASIG5V.n11951 0.0200092
R51897 ASIG5V.n12111 ASIG5V.n12110 0.0200092
R51898 ASIG5V.n12264 ASIG5V.n12263 0.0200092
R51899 ASIG5V.n12381 ASIG5V.n12380 0.0200092
R51900 ASIG5V.n12607 ASIG5V.n12606 0.0200092
R51901 ASIG5V.n7267 ASIG5V.n7266 0.0200092
R51902 ASIG5V.n7849 ASIG5V.n7848 0.0200092
R51903 ASIG5V.n7432 ASIG5V.n7431 0.0200092
R51904 ASIG5V.n357 ASIG5V.n356 0.0200092
R51905 ASIG5V.n13521 ASIG5V.n13520 0.0200092
R51906 ASIG5V.n6683 ASIG5V.n6682 0.0200092
R51907 ASIG5V.n6961 ASIG5V.n6960 0.0200092
R51908 ASIG5V.n508 ASIG5V.n507 0.0200092
R51909 ASIG5V.n5886 ASIG5V.n5885 0.0200092
R51910 ASIG5V.n5585 ASIG5V.n5584 0.0200092
R51911 ASIG5V.n5354 ASIG5V.n5353 0.0200092
R51912 ASIG5V.n4927 ASIG5V.n4926 0.0200092
R51913 ASIG5V.n4659 ASIG5V.n4658 0.0200092
R51914 ASIG5V.n4401 ASIG5V.n4400 0.0200092
R51915 ASIG5V.n4125 ASIG5V.n4124 0.0200092
R51916 ASIG5V.n3859 ASIG5V.n3858 0.0200092
R51917 ASIG5V.n3584 ASIG5V.n3583 0.0200092
R51918 ASIG5V.n3325 ASIG5V.n3324 0.0200092
R51919 ASIG5V.n3130 ASIG5V.n3129 0.0200092
R51920 ASIG5V.n11656 ASIG5V.n11655 0.0200092
R51921 ASIG5V.n11785 ASIG5V.n11784 0.0200092
R51922 ASIG5V.n11948 ASIG5V.n11947 0.0200092
R51923 ASIG5V.n12107 ASIG5V.n12106 0.0200092
R51924 ASIG5V.n12260 ASIG5V.n12259 0.0200092
R51925 ASIG5V.n12377 ASIG5V.n12376 0.0200092
R51926 ASIG5V.n12603 ASIG5V.n12602 0.0200092
R51927 ASIG5V.n7263 ASIG5V.n7262 0.0200092
R51928 ASIG5V.n7845 ASIG5V.n7844 0.0200092
R51929 ASIG5V.n7428 ASIG5V.n7427 0.0200092
R51930 ASIG5V.n353 ASIG5V.n352 0.0200092
R51931 ASIG5V.n13517 ASIG5V.n13516 0.0200092
R51932 ASIG5V.n6679 ASIG5V.n6678 0.0200092
R51933 ASIG5V.n6957 ASIG5V.n6956 0.0200092
R51934 ASIG5V.n504 ASIG5V.n503 0.0200092
R51935 ASIG5V.n5882 ASIG5V.n5881 0.0200092
R51936 ASIG5V.n5581 ASIG5V.n5580 0.0200092
R51937 ASIG5V.n5350 ASIG5V.n5349 0.0200092
R51938 ASIG5V.n4923 ASIG5V.n4922 0.0200092
R51939 ASIG5V.n4655 ASIG5V.n4654 0.0200092
R51940 ASIG5V.n4397 ASIG5V.n4396 0.0200092
R51941 ASIG5V.n4121 ASIG5V.n4120 0.0200092
R51942 ASIG5V.n3855 ASIG5V.n3854 0.0200092
R51943 ASIG5V.n3580 ASIG5V.n3579 0.0200092
R51944 ASIG5V.n3321 ASIG5V.n3320 0.0200092
R51945 ASIG5V.n3126 ASIG5V.n3125 0.0200092
R51946 ASIG5V.n3122 ASIG5V.n3121 0.0200092
R51947 ASIG5V.n3317 ASIG5V.n3316 0.0200092
R51948 ASIG5V.n3576 ASIG5V.n3575 0.0200092
R51949 ASIG5V.n3851 ASIG5V.n3850 0.0200092
R51950 ASIG5V.n4117 ASIG5V.n4116 0.0200092
R51951 ASIG5V.n4393 ASIG5V.n4392 0.0200092
R51952 ASIG5V.n4651 ASIG5V.n4650 0.0200092
R51953 ASIG5V.n4919 ASIG5V.n4918 0.0200092
R51954 ASIG5V.n5346 ASIG5V.n5345 0.0200092
R51955 ASIG5V.n5577 ASIG5V.n5576 0.0200092
R51956 ASIG5V.n5878 ASIG5V.n5877 0.0200092
R51957 ASIG5V.n500 ASIG5V.n499 0.0200092
R51958 ASIG5V.n6953 ASIG5V.n6952 0.0200092
R51959 ASIG5V.n6675 ASIG5V.n6674 0.0200092
R51960 ASIG5V.n13513 ASIG5V.n13512 0.0200092
R51961 ASIG5V.n349 ASIG5V.n348 0.0200092
R51962 ASIG5V.n7424 ASIG5V.n7423 0.0200092
R51963 ASIG5V.n7841 ASIG5V.n7840 0.0200092
R51964 ASIG5V.n7259 ASIG5V.n7258 0.0200092
R51965 ASIG5V.n12599 ASIG5V.n12598 0.0200092
R51966 ASIG5V.n12373 ASIG5V.n12372 0.0200092
R51967 ASIG5V.n12256 ASIG5V.n12255 0.0200092
R51968 ASIG5V.n12103 ASIG5V.n12102 0.0200092
R51969 ASIG5V.n11944 ASIG5V.n11943 0.0200092
R51970 ASIG5V.n11781 ASIG5V.n11780 0.0200092
R51971 ASIG5V.n11652 ASIG5V.n11651 0.0200092
R51972 ASIG5V.n11648 ASIG5V.n11647 0.0200092
R51973 ASIG5V.n11777 ASIG5V.n11776 0.0200092
R51974 ASIG5V.n11940 ASIG5V.n11939 0.0200092
R51975 ASIG5V.n12099 ASIG5V.n12098 0.0200092
R51976 ASIG5V.n12252 ASIG5V.n12251 0.0200092
R51977 ASIG5V.n12369 ASIG5V.n12368 0.0200092
R51978 ASIG5V.n12595 ASIG5V.n12594 0.0200092
R51979 ASIG5V.n7255 ASIG5V.n7254 0.0200092
R51980 ASIG5V.n7837 ASIG5V.n7836 0.0200092
R51981 ASIG5V.n7420 ASIG5V.n7419 0.0200092
R51982 ASIG5V.n345 ASIG5V.n344 0.0200092
R51983 ASIG5V.n13509 ASIG5V.n13508 0.0200092
R51984 ASIG5V.n6671 ASIG5V.n6670 0.0200092
R51985 ASIG5V.n6949 ASIG5V.n6948 0.0200092
R51986 ASIG5V.n496 ASIG5V.n495 0.0200092
R51987 ASIG5V.n5874 ASIG5V.n5873 0.0200092
R51988 ASIG5V.n5573 ASIG5V.n5572 0.0200092
R51989 ASIG5V.n5342 ASIG5V.n5341 0.0200092
R51990 ASIG5V.n4915 ASIG5V.n4914 0.0200092
R51991 ASIG5V.n4647 ASIG5V.n4646 0.0200092
R51992 ASIG5V.n4389 ASIG5V.n4388 0.0200092
R51993 ASIG5V.n4113 ASIG5V.n4112 0.0200092
R51994 ASIG5V.n3847 ASIG5V.n3846 0.0200092
R51995 ASIG5V.n3572 ASIG5V.n3571 0.0200092
R51996 ASIG5V.n3313 ASIG5V.n3312 0.0200092
R51997 ASIG5V.n3118 ASIG5V.n3117 0.0200092
R51998 ASIG5V.n11644 ASIG5V.n11643 0.0200092
R51999 ASIG5V.n11773 ASIG5V.n11772 0.0200092
R52000 ASIG5V.n11936 ASIG5V.n11935 0.0200092
R52001 ASIG5V.n12095 ASIG5V.n12094 0.0200092
R52002 ASIG5V.n12248 ASIG5V.n12247 0.0200092
R52003 ASIG5V.n12365 ASIG5V.n12364 0.0200092
R52004 ASIG5V.n12591 ASIG5V.n12590 0.0200092
R52005 ASIG5V.n7251 ASIG5V.n7250 0.0200092
R52006 ASIG5V.n7833 ASIG5V.n7832 0.0200092
R52007 ASIG5V.n7416 ASIG5V.n7415 0.0200092
R52008 ASIG5V.n341 ASIG5V.n340 0.0200092
R52009 ASIG5V.n13505 ASIG5V.n13504 0.0200092
R52010 ASIG5V.n6667 ASIG5V.n6666 0.0200092
R52011 ASIG5V.n6945 ASIG5V.n6944 0.0200092
R52012 ASIG5V.n492 ASIG5V.n491 0.0200092
R52013 ASIG5V.n5870 ASIG5V.n5869 0.0200092
R52014 ASIG5V.n5569 ASIG5V.n5568 0.0200092
R52015 ASIG5V.n5338 ASIG5V.n5337 0.0200092
R52016 ASIG5V.n4911 ASIG5V.n4910 0.0200092
R52017 ASIG5V.n4643 ASIG5V.n4642 0.0200092
R52018 ASIG5V.n4385 ASIG5V.n4384 0.0200092
R52019 ASIG5V.n4109 ASIG5V.n4108 0.0200092
R52020 ASIG5V.n3843 ASIG5V.n3842 0.0200092
R52021 ASIG5V.n3568 ASIG5V.n3567 0.0200092
R52022 ASIG5V.n3309 ASIG5V.n3308 0.0200092
R52023 ASIG5V.n3114 ASIG5V.n3113 0.0200092
R52024 ASIG5V.n3110 ASIG5V.n3109 0.0200092
R52025 ASIG5V.n3305 ASIG5V.n3304 0.0200092
R52026 ASIG5V.n3564 ASIG5V.n3563 0.0200092
R52027 ASIG5V.n3839 ASIG5V.n3838 0.0200092
R52028 ASIG5V.n4105 ASIG5V.n4104 0.0200092
R52029 ASIG5V.n4381 ASIG5V.n4380 0.0200092
R52030 ASIG5V.n4639 ASIG5V.n4638 0.0200092
R52031 ASIG5V.n4907 ASIG5V.n4906 0.0200092
R52032 ASIG5V.n5334 ASIG5V.n5333 0.0200092
R52033 ASIG5V.n5565 ASIG5V.n5564 0.0200092
R52034 ASIG5V.n5866 ASIG5V.n5865 0.0200092
R52035 ASIG5V.n488 ASIG5V.n487 0.0200092
R52036 ASIG5V.n6941 ASIG5V.n6940 0.0200092
R52037 ASIG5V.n6663 ASIG5V.n6662 0.0200092
R52038 ASIG5V.n13501 ASIG5V.n13500 0.0200092
R52039 ASIG5V.n337 ASIG5V.n336 0.0200092
R52040 ASIG5V.n7412 ASIG5V.n7411 0.0200092
R52041 ASIG5V.n7829 ASIG5V.n7828 0.0200092
R52042 ASIG5V.n7247 ASIG5V.n7246 0.0200092
R52043 ASIG5V.n12587 ASIG5V.n12586 0.0200092
R52044 ASIG5V.n12361 ASIG5V.n12360 0.0200092
R52045 ASIG5V.n12244 ASIG5V.n12243 0.0200092
R52046 ASIG5V.n12091 ASIG5V.n12090 0.0200092
R52047 ASIG5V.n11932 ASIG5V.n11931 0.0200092
R52048 ASIG5V.n11769 ASIG5V.n11768 0.0200092
R52049 ASIG5V.n11640 ASIG5V.n11639 0.0200092
R52050 ASIG5V.n3106 ASIG5V.n3105 0.0200092
R52051 ASIG5V.n3301 ASIG5V.n3300 0.0200092
R52052 ASIG5V.n3560 ASIG5V.n3559 0.0200092
R52053 ASIG5V.n3835 ASIG5V.n3834 0.0200092
R52054 ASIG5V.n4101 ASIG5V.n4100 0.0200092
R52055 ASIG5V.n4377 ASIG5V.n4376 0.0200092
R52056 ASIG5V.n4635 ASIG5V.n4634 0.0200092
R52057 ASIG5V.n4903 ASIG5V.n4902 0.0200092
R52058 ASIG5V.n5330 ASIG5V.n5329 0.0200092
R52059 ASIG5V.n5561 ASIG5V.n5560 0.0200092
R52060 ASIG5V.n5862 ASIG5V.n5861 0.0200092
R52061 ASIG5V.n484 ASIG5V.n483 0.0200092
R52062 ASIG5V.n6937 ASIG5V.n6936 0.0200092
R52063 ASIG5V.n6659 ASIG5V.n6658 0.0200092
R52064 ASIG5V.n13497 ASIG5V.n13496 0.0200092
R52065 ASIG5V.n333 ASIG5V.n332 0.0200092
R52066 ASIG5V.n7408 ASIG5V.n7407 0.0200092
R52067 ASIG5V.n7825 ASIG5V.n7824 0.0200092
R52068 ASIG5V.n7243 ASIG5V.n7242 0.0200092
R52069 ASIG5V.n12583 ASIG5V.n12582 0.0200092
R52070 ASIG5V.n12357 ASIG5V.n12356 0.0200092
R52071 ASIG5V.n12240 ASIG5V.n12239 0.0200092
R52072 ASIG5V.n12087 ASIG5V.n12086 0.0200092
R52073 ASIG5V.n11928 ASIG5V.n11927 0.0200092
R52074 ASIG5V.n11765 ASIG5V.n11764 0.0200092
R52075 ASIG5V.n11636 ASIG5V.n11635 0.0200092
R52076 ASIG5V.n8712 ASIG5V.n8711 0.0200092
R52077 ASIG5V.n8609 ASIG5V.n8608 0.0200092
R52078 ASIG5V.n8363 ASIG5V.n8362 0.0200092
R52079 ASIG5V.n8116 ASIG5V.n8115 0.0200092
R52080 ASIG5V.n7817 ASIG5V.n7816 0.0200092
R52081 ASIG5V.n98 ASIG5V.n97 0.0200092
R52082 ASIG5V.n6320 ASIG5V.n6319 0.0200092
R52083 ASIG5V.n5322 ASIG5V.n5321 0.0200092
R52084 ASIG5V.n8709 ASIG5V.n8708 0.0200092
R52085 ASIG5V.n8360 ASIG5V.n8359 0.0200092
R52086 ASIG5V.n8113 ASIG5V.n8112 0.0200092
R52087 ASIG5V.n7814 ASIG5V.n7813 0.0200092
R52088 ASIG5V.n95 ASIG5V.n94 0.0200092
R52089 ASIG5V.n6317 ASIG5V.n6316 0.0200092
R52090 ASIG5V.n5319 ASIG5V.n5318 0.0200092
R52091 ASIG5V.n3552 ASIG5V.n3551 0.0200092
R52092 ASIG5V.n5316 ASIG5V.n5315 0.0200092
R52093 ASIG5V.n6314 ASIG5V.n6313 0.0200092
R52094 ASIG5V.n6412 ASIG5V.n6411 0.0200092
R52095 ASIG5V.n6542 ASIG5V.n6541 0.0200092
R52096 ASIG5V.n92 ASIG5V.n91 0.0200092
R52097 ASIG5V.n7392 ASIG5V.n7391 0.0200092
R52098 ASIG5V.n7811 ASIG5V.n7810 0.0200092
R52099 ASIG5V.n8357 ASIG5V.n8356 0.0200092
R52100 ASIG5V.n8485 ASIG5V.n8484 0.0200092
R52101 ASIG5V.n8354 ASIG5V.n8353 0.0200092
R52102 ASIG5V.n7808 ASIG5V.n7807 0.0200092
R52103 ASIG5V.n7389 ASIG5V.n7388 0.0200092
R52104 ASIG5V.n89 ASIG5V.n88 0.0200092
R52105 ASIG5V.n6311 ASIG5V.n6310 0.0200092
R52106 ASIG5V.n5313 ASIG5V.n5312 0.0200092
R52107 ASIG5V.n3549 ASIG5V.n3548 0.0200092
R52108 ASIG5V.n8480 ASIG5V.n8479 0.0200092
R52109 ASIG5V.n8351 ASIG5V.n8350 0.0200092
R52110 ASIG5V.n7805 ASIG5V.n7804 0.0200092
R52111 ASIG5V.n86 ASIG5V.n85 0.0200092
R52112 ASIG5V.n6308 ASIG5V.n6307 0.0200092
R52113 ASIG5V.n5310 ASIG5V.n5309 0.0200092
R52114 ASIG5V.n3546 ASIG5V.n3545 0.0200092
R52115 ASIG5V.n5307 ASIG5V.n5306 0.0200092
R52116 ASIG5V.n5548 ASIG5V.n5547 0.0200092
R52117 ASIG5V.n6305 ASIG5V.n6304 0.0200092
R52118 ASIG5V.n83 ASIG5V.n82 0.0200092
R52119 ASIG5V.n7385 ASIG5V.n7384 0.0200092
R52120 ASIG5V.n7802 ASIG5V.n7801 0.0200092
R52121 ASIG5V.n8348 ASIG5V.n8347 0.0200092
R52122 ASIG5V.n8477 ASIG5V.n8476 0.0200092
R52123 ASIG5V.n8598 ASIG5V.n8597 0.0200092
R52124 ASIG5V.n5304 ASIG5V.n5303 0.0200092
R52125 ASIG5V.n5545 ASIG5V.n5544 0.0200092
R52126 ASIG5V.n6302 ASIG5V.n6301 0.0200092
R52127 ASIG5V.n6536 ASIG5V.n6535 0.0200092
R52128 ASIG5V.n7382 ASIG5V.n7381 0.0200092
R52129 ASIG5V.n7799 ASIG5V.n7798 0.0200092
R52130 ASIG5V.n8345 ASIG5V.n8344 0.0200092
R52131 ASIG5V.n8801 ASIG5V.n8800 0.0200092
R52132 ASIG5V.n8696 ASIG5V.n8695 0.0200092
R52133 ASIG5V.n8342 ASIG5V.n8341 0.0200092
R52134 ASIG5V.n7796 ASIG5V.n7795 0.0200092
R52135 ASIG5V.n6299 ASIG5V.n6298 0.0200092
R52136 ASIG5V.n5301 ASIG5V.n5300 0.0200092
R52137 ASIG5V.n3541 ASIG5V.n3540 0.0200092
R52138 ASIG5V.n5298 ASIG5V.n5297 0.0200092
R52139 ASIG5V.n6296 ASIG5V.n6295 0.0200092
R52140 ASIG5V.n6402 ASIG5V.n6401 0.0200092
R52141 ASIG5V.n7793 ASIG5V.n7792 0.0200092
R52142 ASIG5V.n8339 ASIG5V.n8338 0.0200092
R52143 ASIG5V.n8470 ASIG5V.n8469 0.0200092
R52144 ASIG5V.n5293 ASIG5V.n5292 0.0200092
R52145 ASIG5V.n6291 ASIG5V.n6290 0.0200092
R52146 ASIG5V.n6528 ASIG5V.n6527 0.0200092
R52147 ASIG5V.n7788 ASIG5V.n7787 0.0200092
R52148 ASIG5V.n8334 ASIG5V.n8333 0.0200092
R52149 ASIG5V.n8793 ASIG5V.n8792 0.0200092
R52150 ASIG5V.n8329 ASIG5V.n8328 0.0200092
R52151 ASIG5V.n7783 ASIG5V.n7782 0.0200092
R52152 ASIG5V.n6286 ASIG5V.n6285 0.0200092
R52153 ASIG5V.n8582 ASIG5V.n8581 0.0200092
R52154 ASIG5V.n8459 ASIG5V.n8458 0.0200092
R52155 ASIG5V.n8324 ASIG5V.n8323 0.0200092
R52156 ASIG5V.n7778 ASIG5V.n7777 0.0200092
R52157 ASIG5V.n6281 ASIG5V.n6280 0.0200092
R52158 ASIG5V.n5285 ASIG5V.n5284 0.0200092
R52159 ASIG5V.n3536 ASIG5V.n3535 0.0200092
R52160 ASIG5V.n3531 ASIG5V.n3530 0.0200092
R52161 ASIG5V.n3809 ASIG5V.n3808 0.0200092
R52162 ASIG5V.n5280 ASIG5V.n5279 0.0200092
R52163 ASIG5V.n6276 ASIG5V.n6275 0.0200092
R52164 ASIG5V.n6392 ASIG5V.n6391 0.0200092
R52165 ASIG5V.n7773 ASIG5V.n7772 0.0200092
R52166 ASIG5V.n8319 ASIG5V.n8318 0.0200092
R52167 ASIG5V.n8577 ASIG5V.n8576 0.0200092
R52168 ASIG5V.n8451 ASIG5V.n8450 0.0200092
R52169 ASIG5V.n8314 ASIG5V.n8313 0.0200092
R52170 ASIG5V.n7768 ASIG5V.n7767 0.0200092
R52171 ASIG5V.n6271 ASIG5V.n6270 0.0200092
R52172 ASIG5V.n5275 ASIG5V.n5274 0.0200092
R52173 ASIG5V.n8569 ASIG5V.n8568 0.0200092
R52174 ASIG5V.n8309 ASIG5V.n8308 0.0200092
R52175 ASIG5V.n7763 ASIG5V.n7762 0.0200092
R52176 ASIG5V.n6511 ASIG5V.n6510 0.0200092
R52177 ASIG5V.n6266 ASIG5V.n6265 0.0200092
R52178 ASIG5V.n5270 ASIG5V.n5269 0.0200092
R52179 ASIG5V.n3527 ASIG5V.n3526 0.0200092
R52180 ASIG5V.n5265 ASIG5V.n5264 0.0200092
R52181 ASIG5V.n6261 ASIG5V.n6260 0.0200092
R52182 ASIG5V.n57 ASIG5V.n56 0.0200092
R52183 ASIG5V.n7758 ASIG5V.n7757 0.0200092
R52184 ASIG5V.n8304 ASIG5V.n8303 0.0200092
R52185 ASIG5V.n5259 ASIG5V.n5258 0.0200092
R52186 ASIG5V.n6254 ASIG5V.n6253 0.0200092
R52187 ASIG5V.n7752 ASIG5V.n7751 0.0200092
R52188 ASIG5V.n8299 ASIG5V.n8298 0.0200092
R52189 ASIG5V.n8669 ASIG5V.n8668 0.0200092
R52190 ASIG5V.n8664 ASIG5V.n8663 0.0200092
R52191 ASIG5V.n8293 ASIG5V.n8292 0.0200092
R52192 ASIG5V.n8072 ASIG5V.n8071 0.0200092
R52193 ASIG5V.n7745 ASIG5V.n7744 0.0200092
R52194 ASIG5V.n6498 ASIG5V.n6497 0.0200092
R52195 ASIG5V.n6247 ASIG5V.n6246 0.0200092
R52196 ASIG5V.n5252 ASIG5V.n5251 0.0200092
R52197 ASIG5V.n3522 ASIG5V.n3521 0.0200092
R52198 ASIG5V.n8764 ASIG5V.n8763 0.0200092
R52199 ASIG5V.n8434 ASIG5V.n8433 0.0200092
R52200 ASIG5V.n8286 ASIG5V.n8285 0.0200092
R52201 ASIG5V.n8065 ASIG5V.n8064 0.0200092
R52202 ASIG5V.n7738 ASIG5V.n7737 0.0200092
R52203 ASIG5V.n6491 ASIG5V.n6490 0.0200092
R52204 ASIG5V.n6240 ASIG5V.n6239 0.0200092
R52205 ASIG5V.n5245 ASIG5V.n5244 0.0200092
R52206 ASIG5V.n3518 ASIG5V.n3517 0.0200092
R52207 ASIG5V.n4604 ASIG5V.n4603 0.0200092
R52208 ASIG5V.n5238 ASIG5V.n5237 0.0200092
R52209 ASIG5V.n6233 ASIG5V.n6232 0.0200092
R52210 ASIG5V.n44 ASIG5V.n43 0.0200092
R52211 ASIG5V.n7345 ASIG5V.n7344 0.0200092
R52212 ASIG5V.n7731 ASIG5V.n7730 0.0200092
R52213 ASIG5V.n8279 ASIG5V.n8278 0.0200092
R52214 ASIG5V.n8427 ASIG5V.n8426 0.0200092
R52215 ASIG5V.n8551 ASIG5V.n8550 0.0200092
R52216 ASIG5V.n8272 ASIG5V.n8271 0.0200092
R52217 ASIG5V.n7724 ASIG5V.n7723 0.0200092
R52218 ASIG5V.n6226 ASIG5V.n6225 0.0200092
R52219 ASIG5V.n5231 ASIG5V.n5230 0.0200092
R52220 ASIG5V.n3514 ASIG5V.n3513 0.0200092
R52221 ASIG5V.n8265 ASIG5V.n8264 0.0200092
R52222 ASIG5V.n7717 ASIG5V.n7716 0.0200092
R52223 ASIG5V.n6479 ASIG5V.n6478 0.0200092
R52224 ASIG5V.n6219 ASIG5V.n6218 0.0200092
R52225 ASIG5V.n5224 ASIG5V.n5223 0.0200092
R52226 ASIG5V.n5217 ASIG5V.n5216 0.0200092
R52227 ASIG5V.n6212 ASIG5V.n6211 0.0200092
R52228 ASIG5V.n7333 ASIG5V.n7332 0.0200092
R52229 ASIG5V.n7710 ASIG5V.n7709 0.0200092
R52230 ASIG5V.n8046 ASIG5V.n8045 0.0200092
R52231 ASIG5V.n8148 ASIG5V.n8147 0.0200092
R52232 ASIG5V.n8258 ASIG5V.n8257 0.0200092
R52233 ASIG5V.n8536 ASIG5V.n8535 0.0200092
R52234 ASIG5V.n3508 ASIG5V.n3507 0.0200092
R52235 ASIG5V.n5210 ASIG5V.n5209 0.0200092
R52236 ASIG5V.n6205 ASIG5V.n6204 0.0200092
R52237 ASIG5V.n6368 ASIG5V.n6367 0.0200092
R52238 ASIG5V.n7703 ASIG5V.n7702 0.0200092
R52239 ASIG5V.n8039 ASIG5V.n8038 0.0200092
R52240 ASIG5V.n8251 ASIG5V.n8250 0.0200092
R52241 ASIG5V.n8408 ASIG5V.n8407 0.0200092
R52242 ASIG5V.n8244 ASIG5V.n8243 0.0200092
R52243 ASIG5V.n7696 ASIG5V.n7695 0.0200092
R52244 ASIG5V.n6467 ASIG5V.n6466 0.0200092
R52245 ASIG5V.n5489 ASIG5V.n5488 0.0200092
R52246 ASIG5V.n5203 ASIG5V.n5202 0.0200092
R52247 ASIG5V.n3768 ASIG5V.n3767 0.0200092
R52248 ASIG5V.n8522 ASIG5V.n8521 0.0200092
R52249 ASIG5V.n8237 ASIG5V.n8236 0.0200092
R52250 ASIG5V.n7689 ASIG5V.n7688 0.0200092
R52251 ASIG5V.n6463 ASIG5V.n6462 0.0200092
R52252 ASIG5V.n5828 ASIG5V.n5827 0.0200092
R52253 ASIG5V.n5196 ASIG5V.n5195 0.0200092
R52254 ASIG5V.n3502 ASIG5V.n3501 0.0200092
R52255 ASIG5V.n3499 ASIG5V.n3498 0.0200092
R52256 ASIG5V.n5189 ASIG5V.n5188 0.0200092
R52257 ASIG5V.n6356 ASIG5V.n6355 0.0200092
R52258 ASIG5V.n28 ASIG5V.n27 0.0200092
R52259 ASIG5V.n7682 ASIG5V.n7681 0.0200092
R52260 ASIG5V.n8024 ASIG5V.n8023 0.0200092
R52261 ASIG5V.n8230 ASIG5V.n8229 0.0200092
R52262 ASIG5V.n8391 ASIG5V.n8390 0.0200092
R52263 ASIG5V.n8225 ASIG5V.n8224 0.0200092
R52264 ASIG5V.n7675 ASIG5V.n7674 0.0200092
R52265 ASIG5V.n6452 ASIG5V.n6451 0.0200092
R52266 ASIG5V.n6189 ASIG5V.n6188 0.0200092
R52267 ASIG5V.n5182 ASIG5V.n5181 0.0200092
R52268 ASIG5V.n3761 ASIG5V.n3760 0.0200092
R52269 ASIG5V.n3496 ASIG5V.n3495 0.0200092
R52270 ASIG5V.n8511 ASIG5V.n8510 0.0200092
R52271 ASIG5V.n8220 ASIG5V.n8219 0.0200092
R52272 ASIG5V.n7668 ASIG5V.n7667 0.0200092
R52273 ASIG5V.n7306 ASIG5V.n7305 0.0200092
R52274 ASIG5V.n6448 ASIG5V.n6447 0.0200092
R52275 ASIG5V.n6185 ASIG5V.n6184 0.0200092
R52276 ASIG5V.n5819 ASIG5V.n5818 0.0200092
R52277 ASIG5V.n5470 ASIG5V.n5469 0.0200092
R52278 ASIG5V.n5175 ASIG5V.n5174 0.0200092
R52279 ASIG5V.n3493 ASIG5V.n3492 0.0200092
R52280 ASIG5V.n5170 ASIG5V.n5169 0.0200092
R52281 ASIG5V.n19 ASIG5V.n18 0.0200092
R52282 ASIG5V.n7661 ASIG5V.n7660 0.0200092
R52283 ASIG5V.n8009 ASIG5V.n8008 0.0200092
R52284 ASIG5V.n8215 ASIG5V.n8214 0.0200092
R52285 ASIG5V.n8383 ASIG5V.n8382 0.0200092
R52286 ASIG5V.n3489 ASIG5V.n3488 0.0200092
R52287 ASIG5V.n5165 ASIG5V.n5164 0.0200092
R52288 ASIG5V.n6437 ASIG5V.n6436 0.0200092
R52289 ASIG5V.n7655 ASIG5V.n7654 0.0200092
R52290 ASIG5V.n8004 ASIG5V.n8003 0.0200092
R52291 ASIG5V.n8210 ASIG5V.n8209 0.0200092
R52292 ASIG5V.n8378 ASIG5V.n8377 0.0200092
R52293 ASIG5V.n8503 ASIG5V.n8502 0.0200092
R52294 ASIG5V.n8621 ASIG5V.n8620 0.0200092
R52295 ASIG5V.n8723 ASIG5V.n8722 0.0200092
R52296 ASIG5V.n8498 ASIG5V.n8497 0.0200092
R52297 ASIG5V.n8205 ASIG5V.n8204 0.0200092
R52298 ASIG5V.n7650 ASIG5V.n7649 0.0200092
R52299 ASIG5V.n6433 ASIG5V.n6432 0.0200092
R52300 ASIG5V.n5160 ASIG5V.n5159 0.0200092
R52301 ASIG5V.n3487 ASIG5V.n3486 0.0200092
R52302 ASIG5V.n11485 ASIG5V.n11484 0.0200092
R52303 ASIG5V.n8720 ASIG5V.n8719 0.0200092
R52304 ASIG5V.n8370 ASIG5V.n8369 0.0200092
R52305 ASIG5V.n8200 ASIG5V.n8199 0.0200092
R52306 ASIG5V.n7645 ASIG5V.n7644 0.0200092
R52307 ASIG5V.n7 ASIG5V.n6 0.0200092
R52308 ASIG5V.n6429 ASIG5V.n6428 0.0200092
R52309 ASIG5V.n3750 ASIG5V.n3749 0.0200092
R52310 ASIG5V.n3485 ASIG5V.n3484 0.0200092
R52311 ASIG5V.n3120 ASIG5V.n3119 0.0200092
R52312 ASIG5V.n3108 ASIG5V.n3107 0.0200092
R52313 ASIG5V.n3147 ASIG5V.n3146 0.0200092
R52314 ASIG5V.n3150 ASIG5V.n3149 0.0200092
R52315 ASIG5V.n3153 ASIG5V.n3152 0.0200092
R52316 ASIG5V.n3162 ASIG5V.n3161 0.0200092
R52317 ASIG5V.n3167 ASIG5V.n3166 0.0200092
R52318 ASIG5V.n3175 ASIG5V.n3174 0.0200092
R52319 ASIG5V.n3186 ASIG5V.n3185 0.0200092
R52320 ASIG5V.n3192 ASIG5V.n3191 0.0200092
R52321 ASIG5V.n3315 ASIG5V.n3314 0.0200092
R52322 ASIG5V.n3303 ASIG5V.n3302 0.0200092
R52323 ASIG5V.n3339 ASIG5V.n3338 0.0200092
R52324 ASIG5V.n3342 ASIG5V.n3341 0.0200092
R52325 ASIG5V.n3345 ASIG5V.n3344 0.0200092
R52326 ASIG5V.n3348 ASIG5V.n3347 0.0200092
R52327 ASIG5V.n3353 ASIG5V.n3352 0.0200092
R52328 ASIG5V.n3358 ASIG5V.n3357 0.0200092
R52329 ASIG5V.n3363 ASIG5V.n3362 0.0200092
R52330 ASIG5V.n3368 ASIG5V.n3367 0.0200092
R52331 ASIG5V.n3373 ASIG5V.n3372 0.0200092
R52332 ASIG5V.n3378 ASIG5V.n3377 0.0200092
R52333 ASIG5V.n3383 ASIG5V.n3382 0.0200092
R52334 ASIG5V.n3388 ASIG5V.n3387 0.0200092
R52335 ASIG5V.n3393 ASIG5V.n3392 0.0200092
R52336 ASIG5V.n3396 ASIG5V.n3395 0.0200092
R52337 ASIG5V.n3399 ASIG5V.n3398 0.0200092
R52338 ASIG5V.n3574 ASIG5V.n3573 0.0200092
R52339 ASIG5V.n3562 ASIG5V.n3561 0.0200092
R52340 ASIG5V.n3631 ASIG5V.n3630 0.0200092
R52341 ASIG5V.n3635 ASIG5V.n3634 0.0200092
R52342 ASIG5V.n3638 ASIG5V.n3637 0.0200092
R52343 ASIG5V.n3643 ASIG5V.n3642 0.0200092
R52344 ASIG5V.n3648 ASIG5V.n3647 0.0200092
R52345 ASIG5V.n3651 ASIG5V.n3650 0.0200092
R52346 ASIG5V.n3656 ASIG5V.n3655 0.0200092
R52347 ASIG5V.n3661 ASIG5V.n3660 0.0200092
R52348 ASIG5V.n3665 ASIG5V.n3664 0.0200092
R52349 ASIG5V.n3670 ASIG5V.n3669 0.0200092
R52350 ASIG5V.n3674 ASIG5V.n3673 0.0200092
R52351 ASIG5V.n3677 ASIG5V.n3676 0.0200092
R52352 ASIG5V.n3679 ASIG5V.n3678 0.0200092
R52353 ASIG5V.n3849 ASIG5V.n3848 0.0200092
R52354 ASIG5V.n3837 ASIG5V.n3836 0.0200092
R52355 ASIG5V.n3915 ASIG5V.n3914 0.0200092
R52356 ASIG5V.n3937 ASIG5V.n3936 0.0200092
R52357 ASIG5V.n3942 ASIG5V.n3941 0.0200092
R52358 ASIG5V.n3948 ASIG5V.n3947 0.0200092
R52359 ASIG5V.n4115 ASIG5V.n4114 0.0200092
R52360 ASIG5V.n4103 ASIG5V.n4102 0.0200092
R52361 ASIG5V.n4171 ASIG5V.n4170 0.0200092
R52362 ASIG5V.n4174 ASIG5V.n4173 0.0200092
R52363 ASIG5V.n4177 ASIG5V.n4176 0.0200092
R52364 ASIG5V.n4180 ASIG5V.n4179 0.0200092
R52365 ASIG5V.n4188 ASIG5V.n4187 0.0200092
R52366 ASIG5V.n4391 ASIG5V.n4390 0.0200092
R52367 ASIG5V.n4379 ASIG5V.n4378 0.0200092
R52368 ASIG5V.n4454 ASIG5V.n4453 0.0200092
R52369 ASIG5V.n4468 ASIG5V.n4467 0.0200092
R52370 ASIG5V.n4497 ASIG5V.n4496 0.0200092
R52371 ASIG5V.n4649 ASIG5V.n4648 0.0200092
R52372 ASIG5V.n4637 ASIG5V.n4636 0.0200092
R52373 ASIG5V.n4708 ASIG5V.n4707 0.0200092
R52374 ASIG5V.n4711 ASIG5V.n4710 0.0200092
R52375 ASIG5V.n4714 ASIG5V.n4713 0.0200092
R52376 ASIG5V.n4717 ASIG5V.n4716 0.0200092
R52377 ASIG5V.n4722 ASIG5V.n4721 0.0200092
R52378 ASIG5V.n4727 ASIG5V.n4726 0.0200092
R52379 ASIG5V.n4732 ASIG5V.n4731 0.0200092
R52380 ASIG5V.n4737 ASIG5V.n4736 0.0200092
R52381 ASIG5V.n4748 ASIG5V.n4747 0.0200092
R52382 ASIG5V.n4757 ASIG5V.n4756 0.0200092
R52383 ASIG5V.n4762 ASIG5V.n4761 0.0200092
R52384 ASIG5V.n4767 ASIG5V.n4766 0.0200092
R52385 ASIG5V.n4917 ASIG5V.n4916 0.0200092
R52386 ASIG5V.n4905 ASIG5V.n4904 0.0200092
R52387 ASIG5V.n4983 ASIG5V.n4982 0.0200092
R52388 ASIG5V.n4986 ASIG5V.n4985 0.0200092
R52389 ASIG5V.n4989 ASIG5V.n4988 0.0200092
R52390 ASIG5V.n4992 ASIG5V.n4991 0.0200092
R52391 ASIG5V.n4997 ASIG5V.n4996 0.0200092
R52392 ASIG5V.n5002 ASIG5V.n5001 0.0200092
R52393 ASIG5V.n5007 ASIG5V.n5006 0.0200092
R52394 ASIG5V.n5013 ASIG5V.n5012 0.0200092
R52395 ASIG5V.n5020 ASIG5V.n5019 0.0200092
R52396 ASIG5V.n5027 ASIG5V.n5026 0.0200092
R52397 ASIG5V.n5034 ASIG5V.n5033 0.0200092
R52398 ASIG5V.n5041 ASIG5V.n5040 0.0200092
R52399 ASIG5V.n5047 ASIG5V.n5046 0.0200092
R52400 ASIG5V.n5052 ASIG5V.n5051 0.0200092
R52401 ASIG5V.n5057 ASIG5V.n5056 0.0200092
R52402 ASIG5V.n5344 ASIG5V.n5343 0.0200092
R52403 ASIG5V.n5332 ASIG5V.n5331 0.0200092
R52404 ASIG5V.n5575 ASIG5V.n5574 0.0200092
R52405 ASIG5V.n5563 ASIG5V.n5562 0.0200092
R52406 ASIG5V.n5690 ASIG5V.n5689 0.0200092
R52407 ASIG5V.n5730 ASIG5V.n5729 0.0200092
R52408 ASIG5V.n5735 ASIG5V.n5734 0.0200092
R52409 ASIG5V.n5876 ASIG5V.n5875 0.0200092
R52410 ASIG5V.n5864 ASIG5V.n5863 0.0200092
R52411 ASIG5V.n5984 ASIG5V.n5983 0.0200092
R52412 ASIG5V.n5987 ASIG5V.n5986 0.0200092
R52413 ASIG5V.n5990 ASIG5V.n5989 0.0200092
R52414 ASIG5V.n5993 ASIG5V.n5992 0.0200092
R52415 ASIG5V.n5998 ASIG5V.n5997 0.0200092
R52416 ASIG5V.n6003 ASIG5V.n6002 0.0200092
R52417 ASIG5V.n6008 ASIG5V.n6007 0.0200092
R52418 ASIG5V.n6015 ASIG5V.n6014 0.0200092
R52419 ASIG5V.n6022 ASIG5V.n6021 0.0200092
R52420 ASIG5V.n6029 ASIG5V.n6028 0.0200092
R52421 ASIG5V.n6036 ASIG5V.n6035 0.0200092
R52422 ASIG5V.n6043 ASIG5V.n6042 0.0200092
R52423 ASIG5V.n6050 ASIG5V.n6049 0.0200092
R52424 ASIG5V.n6057 ASIG5V.n6056 0.0200092
R52425 ASIG5V.n6062 ASIG5V.n6061 0.0200092
R52426 ASIG5V.n498 ASIG5V.n497 0.0200092
R52427 ASIG5V.n486 ASIG5V.n485 0.0200092
R52428 ASIG5V.n7081 ASIG5V.n7080 0.0200092
R52429 ASIG5V.n7088 ASIG5V.n7087 0.0200092
R52430 ASIG5V.n6951 ASIG5V.n6950 0.0200092
R52431 ASIG5V.n6939 ASIG5V.n6938 0.0200092
R52432 ASIG5V.n6673 ASIG5V.n6672 0.0200092
R52433 ASIG5V.n6661 ASIG5V.n6660 0.0200092
R52434 ASIG5V.n6583 ASIG5V.n6582 0.0200092
R52435 ASIG5V.n6590 ASIG5V.n6589 0.0200092
R52436 ASIG5V.n6597 ASIG5V.n6596 0.0200092
R52437 ASIG5V.n6604 ASIG5V.n6603 0.0200092
R52438 ASIG5V.n6611 ASIG5V.n6610 0.0200092
R52439 ASIG5V.n6615 ASIG5V.n6614 0.0200092
R52440 ASIG5V.n13511 ASIG5V.n13510 0.0200092
R52441 ASIG5V.n13499 ASIG5V.n13498 0.0200092
R52442 ASIG5V.n13398 ASIG5V.n13397 0.0200092
R52443 ASIG5V.n347 ASIG5V.n346 0.0200092
R52444 ASIG5V.n335 ASIG5V.n334 0.0200092
R52445 ASIG5V.n151 ASIG5V.n150 0.0200092
R52446 ASIG5V.n154 ASIG5V.n153 0.0200092
R52447 ASIG5V.n157 ASIG5V.n156 0.0200092
R52448 ASIG5V.n160 ASIG5V.n159 0.0200092
R52449 ASIG5V.n165 ASIG5V.n164 0.0200092
R52450 ASIG5V.n170 ASIG5V.n169 0.0200092
R52451 ASIG5V.n175 ASIG5V.n174 0.0200092
R52452 ASIG5V.n182 ASIG5V.n181 0.0200092
R52453 ASIG5V.n189 ASIG5V.n188 0.0200092
R52454 ASIG5V.n196 ASIG5V.n195 0.0200092
R52455 ASIG5V.n203 ASIG5V.n202 0.0200092
R52456 ASIG5V.n210 ASIG5V.n209 0.0200092
R52457 ASIG5V.n217 ASIG5V.n216 0.0200092
R52458 ASIG5V.n224 ASIG5V.n223 0.0200092
R52459 ASIG5V.n231 ASIG5V.n230 0.0200092
R52460 ASIG5V.n7422 ASIG5V.n7421 0.0200092
R52461 ASIG5V.n7410 ASIG5V.n7409 0.0200092
R52462 ASIG5V.n7528 ASIG5V.n7527 0.0200092
R52463 ASIG5V.n7839 ASIG5V.n7838 0.0200092
R52464 ASIG5V.n7827 ASIG5V.n7826 0.0200092
R52465 ASIG5V.n7257 ASIG5V.n7256 0.0200092
R52466 ASIG5V.n7245 ASIG5V.n7244 0.0200092
R52467 ASIG5V.n12683 ASIG5V.n12682 0.0200092
R52468 ASIG5V.n12597 ASIG5V.n12596 0.0200092
R52469 ASIG5V.n12585 ASIG5V.n12584 0.0200092
R52470 ASIG5V.n12443 ASIG5V.n12442 0.0200092
R52471 ASIG5V.n12458 ASIG5V.n12457 0.0200092
R52472 ASIG5V.n12477 ASIG5V.n12476 0.0200092
R52473 ASIG5V.n12482 ASIG5V.n12481 0.0200092
R52474 ASIG5V.n12487 ASIG5V.n12486 0.0200092
R52475 ASIG5V.n12371 ASIG5V.n12370 0.0200092
R52476 ASIG5V.n12359 ASIG5V.n12358 0.0200092
R52477 ASIG5V.n12254 ASIG5V.n12253 0.0200092
R52478 ASIG5V.n12242 ASIG5V.n12241 0.0200092
R52479 ASIG5V.n12101 ASIG5V.n12100 0.0200092
R52480 ASIG5V.n12089 ASIG5V.n12088 0.0200092
R52481 ASIG5V.n11942 ASIG5V.n11941 0.0200092
R52482 ASIG5V.n11930 ASIG5V.n11929 0.0200092
R52483 ASIG5V.n11779 ASIG5V.n11778 0.0200092
R52484 ASIG5V.n11767 ASIG5V.n11766 0.0200092
R52485 ASIG5V.n11650 ASIG5V.n11649 0.0200092
R52486 ASIG5V.n11638 ASIG5V.n11637 0.0200092
R52487 ASIG5V.n11494 ASIG5V.n11493 0.0200092
R52488 ASIG5V.n11497 ASIG5V.n11496 0.0200092
R52489 ASIG5V.n11500 ASIG5V.n11499 0.0200092
R52490 ASIG5V.n11503 ASIG5V.n11502 0.0200092
R52491 ASIG5V.n11508 ASIG5V.n11507 0.0200092
R52492 ASIG5V.n11513 ASIG5V.n11512 0.0200092
R52493 ASIG5V.n11518 ASIG5V.n11517 0.0200092
R52494 ASIG5V.n11523 ASIG5V.n11522 0.0200092
R52495 ASIG5V.n11528 ASIG5V.n11527 0.0200092
R52496 ASIG5V.n11533 ASIG5V.n11532 0.0200092
R52497 ASIG5V.n11538 ASIG5V.n11537 0.0200092
R52498 ASIG5V.n11543 ASIG5V.n11542 0.0200092
R52499 ASIG5V.n11548 ASIG5V.n11547 0.0200092
R52500 ASIG5V.n11551 ASIG5V.n11550 0.0200092
R52501 ASIG5V.n11554 ASIG5V.n11553 0.0200092
R52502 ASIG5V.n8856 ASIG5V.n8855 0.0200092
R52503 ASIG5V.n11830 ASIG5V.n11829 0.0200092
R52504 ASIG5V.n8718 ASIG5V.n8717 0.0200092
R52505 ASIG5V.n12153 ASIG5V.n12152 0.0200092
R52506 ASIG5V.n12309 ASIG5V.n12308 0.0200092
R52507 ASIG5V.n12424 ASIG5V.n12423 0.0200092
R52508 ASIG5V.n8195 ASIG5V.n8194 0.0200092
R52509 ASIG5V.n8119 ASIG5V.n8118 0.0200092
R52510 ASIG5V.n7822 ASIG5V.n7821 0.0200092
R52511 ASIG5V.n7400 ASIG5V.n7399 0.0200092
R52512 ASIG5V.n149 ASIG5V.n148 0.0200092
R52513 ASIG5V.n106 ASIG5V.n105 0.0200092
R52514 ASIG5V.n6776 ASIG5V.n6775 0.0200092
R52515 ASIG5V.n7051 ASIG5V.n7050 0.0200092
R52516 ASIG5V.n6325 ASIG5V.n6324 0.0200092
R52517 ASIG5V.n5982 ASIG5V.n5981 0.0200092
R52518 ASIG5V.n5686 ASIG5V.n5685 0.0200092
R52519 ASIG5V.n5327 ASIG5V.n5326 0.0200092
R52520 ASIG5V.n4981 ASIG5V.n4980 0.0200092
R52521 ASIG5V.n4706 ASIG5V.n4705 0.0200092
R52522 ASIG5V.n4452 ASIG5V.n4451 0.0200092
R52523 ASIG5V.n4169 ASIG5V.n4168 0.0200092
R52524 ASIG5V.n3903 ASIG5V.n3902 0.0200092
R52525 ASIG5V.n3557 ASIG5V.n3556 0.0200092
R52526 ASIG5V.n3337 ASIG5V.n3336 0.0200092
R52527 ASIG5V.n3145 ASIG5V.n3144 0.0200092
R52528 ASIG5V.n8861 ASIG5V.n8860 0.0200092
R52529 ASIG5V.n11422 ASIG5V.n11421 0.0200092
R52530 ASIG5V.n11410 ASIG5V.n11409 0.019716
R52531 ASIG5V.n11408 ASIG5V.n11407 0.019716
R52532 ASIG5V.n11406 ASIG5V.n11405 0.019716
R52533 ASIG5V.n11404 ASIG5V.n11403 0.019716
R52534 ASIG5V.n11402 ASIG5V.n11401 0.019716
R52535 ASIG5V.n11400 ASIG5V.n11399 0.019716
R52536 ASIG5V.n11398 ASIG5V.n11397 0.019716
R52537 ASIG5V.n11396 ASIG5V.n11395 0.019716
R52538 ASIG5V.n11394 ASIG5V.n11393 0.019716
R52539 ASIG5V.n11392 ASIG5V.n11391 0.019716
R52540 ASIG5V.n11390 ASIG5V.n11389 0.019716
R52541 ASIG5V.n11388 ASIG5V.n11387 0.019716
R52542 ASIG5V.n11386 ASIG5V.n11385 0.019716
R52543 ASIG5V.n11384 ASIG5V.n11383 0.019716
R52544 ASIG5V.n11382 ASIG5V.n11381 0.019716
R52545 ASIG5V.n11380 ASIG5V.n11379 0.019716
R52546 ASIG5V.n11378 ASIG5V.n11377 0.019716
R52547 ASIG5V.n11376 ASIG5V.n11375 0.019716
R52548 ASIG5V.n11374 ASIG5V.n11373 0.019716
R52549 ASIG5V.n11372 ASIG5V.n11371 0.019716
R52550 ASIG5V.n11370 ASIG5V.n11369 0.019716
R52551 ASIG5V.n11368 ASIG5V.n11367 0.019716
R52552 ASIG5V.n11366 ASIG5V.n11365 0.019716
R52553 ASIG5V.n11364 ASIG5V.n11363 0.019716
R52554 ASIG5V.n11362 ASIG5V.n11361 0.019716
R52555 ASIG5V.n11360 ASIG5V.n11359 0.019716
R52556 ASIG5V.n11358 ASIG5V.n11357 0.019716
R52557 ASIG5V.n11356 ASIG5V.n11355 0.019716
R52558 ASIG5V.n11354 ASIG5V.n11353 0.019716
R52559 ASIG5V.n11352 ASIG5V.n11351 0.019716
R52560 ASIG5V.n11350 ASIG5V.n11349 0.019716
R52561 ASIG5V.n11348 ASIG5V.n11347 0.019716
R52562 ASIG5V.n11346 ASIG5V.n11345 0.019716
R52563 ASIG5V.n11344 ASIG5V.n11343 0.019716
R52564 ASIG5V.n11342 ASIG5V.n11341 0.019716
R52565 ASIG5V.n11340 ASIG5V.n11339 0.019716
R52566 ASIG5V.n11338 ASIG5V.n11337 0.019716
R52567 ASIG5V.n11336 ASIG5V.n11335 0.019716
R52568 ASIG5V.n11334 ASIG5V.n11333 0.019716
R52569 ASIG5V.n11332 ASIG5V.n11331 0.019716
R52570 ASIG5V.n11330 ASIG5V.n11329 0.019716
R52571 ASIG5V.n11328 ASIG5V.n11327 0.019716
R52572 ASIG5V.n11326 ASIG5V.n11325 0.019716
R52573 ASIG5V.n11427 ASIG5V.n11426 0.019716
R52574 ASIG5V.n11429 ASIG5V.n11428 0.019716
R52575 ASIG5V.n11431 ASIG5V.n11430 0.019716
R52576 ASIG5V.n11433 ASIG5V.n11432 0.019716
R52577 ASIG5V.n11435 ASIG5V.n11434 0.019716
R52578 ASIG5V.n11437 ASIG5V.n11436 0.019716
R52579 ASIG5V.n11439 ASIG5V.n11438 0.019716
R52580 ASIG5V.n11441 ASIG5V.n11440 0.019716
R52581 ASIG5V.n11443 ASIG5V.n11442 0.019716
R52582 ASIG5V.n11445 ASIG5V.n11444 0.019716
R52583 ASIG5V.n11447 ASIG5V.n11446 0.019716
R52584 ASIG5V.n11449 ASIG5V.n11448 0.019716
R52585 ASIG5V.n11451 ASIG5V.n11450 0.019716
R52586 ASIG5V.n11453 ASIG5V.n11452 0.019716
R52587 ASIG5V.n11455 ASIG5V.n11454 0.019716
R52588 ASIG5V.n11457 ASIG5V.n11456 0.019716
R52589 ASIG5V.n11459 ASIG5V.n11458 0.019716
R52590 ASIG5V.n11461 ASIG5V.n11460 0.019716
R52591 ASIG5V.n11463 ASIG5V.n11462 0.019716
R52592 ASIG5V.n11465 ASIG5V.n11464 0.019716
R52593 ASIG5V.n11467 ASIG5V.n11466 0.019716
R52594 ASIG5V.n11469 ASIG5V.n11468 0.019716
R52595 ASIG5V.n11471 ASIG5V.n11470 0.019716
R52596 ASIG5V.n11473 ASIG5V.n11472 0.019716
R52597 ASIG5V.n11475 ASIG5V.n11474 0.019716
R52598 ASIG5V.n11477 ASIG5V.n11476 0.019716
R52599 ASIG5V.n11479 ASIG5V.n11478 0.019716
R52600 ASIG5V.n11481 ASIG5V.n11480 0.019716
R52601 ASIG5V.n11411 ASIG5V.n11410 0.019716
R52602 ASIG5V.n11409 ASIG5V.n11408 0.019716
R52603 ASIG5V.n11407 ASIG5V.n11406 0.019716
R52604 ASIG5V.n11405 ASIG5V.n11404 0.019716
R52605 ASIG5V.n11403 ASIG5V.n11402 0.019716
R52606 ASIG5V.n11401 ASIG5V.n11400 0.019716
R52607 ASIG5V.n11399 ASIG5V.n11398 0.019716
R52608 ASIG5V.n11397 ASIG5V.n11396 0.019716
R52609 ASIG5V.n11395 ASIG5V.n11394 0.019716
R52610 ASIG5V.n11393 ASIG5V.n11392 0.019716
R52611 ASIG5V.n11391 ASIG5V.n11390 0.019716
R52612 ASIG5V.n11389 ASIG5V.n11388 0.019716
R52613 ASIG5V.n11387 ASIG5V.n11386 0.019716
R52614 ASIG5V.n11385 ASIG5V.n11384 0.019716
R52615 ASIG5V.n11383 ASIG5V.n11382 0.019716
R52616 ASIG5V.n11381 ASIG5V.n11380 0.019716
R52617 ASIG5V.n11379 ASIG5V.n11378 0.019716
R52618 ASIG5V.n11377 ASIG5V.n11376 0.019716
R52619 ASIG5V.n11375 ASIG5V.n11374 0.019716
R52620 ASIG5V.n11373 ASIG5V.n11372 0.019716
R52621 ASIG5V.n11371 ASIG5V.n11370 0.019716
R52622 ASIG5V.n11369 ASIG5V.n11368 0.019716
R52623 ASIG5V.n11367 ASIG5V.n11366 0.019716
R52624 ASIG5V.n11365 ASIG5V.n11364 0.019716
R52625 ASIG5V.n11363 ASIG5V.n11362 0.019716
R52626 ASIG5V.n11361 ASIG5V.n11360 0.019716
R52627 ASIG5V.n11359 ASIG5V.n11358 0.019716
R52628 ASIG5V.n11357 ASIG5V.n11356 0.019716
R52629 ASIG5V.n11355 ASIG5V.n11354 0.019716
R52630 ASIG5V.n11353 ASIG5V.n11352 0.019716
R52631 ASIG5V.n11351 ASIG5V.n11350 0.019716
R52632 ASIG5V.n11349 ASIG5V.n11348 0.019716
R52633 ASIG5V.n11347 ASIG5V.n11346 0.019716
R52634 ASIG5V.n11345 ASIG5V.n11344 0.019716
R52635 ASIG5V.n11343 ASIG5V.n11342 0.019716
R52636 ASIG5V.n11341 ASIG5V.n11340 0.019716
R52637 ASIG5V.n11339 ASIG5V.n11338 0.019716
R52638 ASIG5V.n11337 ASIG5V.n11336 0.019716
R52639 ASIG5V.n11335 ASIG5V.n11334 0.019716
R52640 ASIG5V.n11333 ASIG5V.n11332 0.019716
R52641 ASIG5V.n11331 ASIG5V.n11330 0.019716
R52642 ASIG5V.n11329 ASIG5V.n11328 0.019716
R52643 ASIG5V.n11327 ASIG5V.n11326 0.019716
R52644 ASIG5V.n11426 ASIG5V.n11425 0.019716
R52645 ASIG5V.n11428 ASIG5V.n11427 0.019716
R52646 ASIG5V.n11430 ASIG5V.n11429 0.019716
R52647 ASIG5V.n11432 ASIG5V.n11431 0.019716
R52648 ASIG5V.n11434 ASIG5V.n11433 0.019716
R52649 ASIG5V.n11436 ASIG5V.n11435 0.019716
R52650 ASIG5V.n11438 ASIG5V.n11437 0.019716
R52651 ASIG5V.n11440 ASIG5V.n11439 0.019716
R52652 ASIG5V.n11442 ASIG5V.n11441 0.019716
R52653 ASIG5V.n11444 ASIG5V.n11443 0.019716
R52654 ASIG5V.n11446 ASIG5V.n11445 0.019716
R52655 ASIG5V.n11448 ASIG5V.n11447 0.019716
R52656 ASIG5V.n11450 ASIG5V.n11449 0.019716
R52657 ASIG5V.n11452 ASIG5V.n11451 0.019716
R52658 ASIG5V.n11454 ASIG5V.n11453 0.019716
R52659 ASIG5V.n11456 ASIG5V.n11455 0.019716
R52660 ASIG5V.n11458 ASIG5V.n11457 0.019716
R52661 ASIG5V.n11460 ASIG5V.n11459 0.019716
R52662 ASIG5V.n11462 ASIG5V.n11461 0.019716
R52663 ASIG5V.n11464 ASIG5V.n11463 0.019716
R52664 ASIG5V.n11466 ASIG5V.n11465 0.019716
R52665 ASIG5V.n11468 ASIG5V.n11467 0.019716
R52666 ASIG5V.n11470 ASIG5V.n11469 0.019716
R52667 ASIG5V.n11472 ASIG5V.n11471 0.019716
R52668 ASIG5V.n11474 ASIG5V.n11473 0.019716
R52669 ASIG5V.n11476 ASIG5V.n11475 0.019716
R52670 ASIG5V.n11478 ASIG5V.n11477 0.019716
R52671 ASIG5V.n11480 ASIG5V.n11479 0.019716
R52672 ASIG5V.n11185 ASIG5V.n11184 0.0196384
R52673 ASIG5V.n11184 ASIG5V.n11183 0.0196384
R52674 ASIG5V.n11181 ASIG5V.n11180 0.0196384
R52675 ASIG5V.n11180 ASIG5V.n11179 0.0196384
R52676 ASIG5V.n11177 ASIG5V.n11176 0.0196384
R52677 ASIG5V.n11176 ASIG5V.n11175 0.0196384
R52678 ASIG5V.n11173 ASIG5V.n11172 0.0196384
R52679 ASIG5V.n11172 ASIG5V.n11171 0.0196384
R52680 ASIG5V.n11169 ASIG5V.n11168 0.0196384
R52681 ASIG5V.n11168 ASIG5V.n11167 0.0196384
R52682 ASIG5V.n11165 ASIG5V.n11164 0.0196384
R52683 ASIG5V.n11164 ASIG5V.n11163 0.0196384
R52684 ASIG5V.n11161 ASIG5V.n11160 0.0196384
R52685 ASIG5V.n11160 ASIG5V.n11159 0.0196384
R52686 ASIG5V.n11192 ASIG5V.n11190 0.0196384
R52687 ASIG5V.n11195 ASIG5V.n11193 0.0196384
R52688 ASIG5V.n11198 ASIG5V.n11196 0.0196384
R52689 ASIG5V.n11201 ASIG5V.n11199 0.0196384
R52690 ASIG5V.n11204 ASIG5V.n11202 0.0196384
R52691 ASIG5V.n11206 ASIG5V.n11205 0.0196384
R52692 ASIG5V.n11208 ASIG5V.n11207 0.0196384
R52693 ASIG5V.n11210 ASIG5V.n11209 0.0196384
R52694 ASIG5V.n11119 ASIG5V.n11117 0.0196384
R52695 ASIG5V.n11216 ASIG5V.n11213 0.0196384
R52696 ASIG5V.n11221 ASIG5V.n11218 0.0196384
R52697 ASIG5V.n11226 ASIG5V.n11223 0.0196384
R52698 ASIG5V.n11231 ASIG5V.n11228 0.0196384
R52699 ASIG5V.n11236 ASIG5V.n11233 0.0196384
R52700 ASIG5V.n11241 ASIG5V.n11238 0.0196384
R52701 ASIG5V.n11246 ASIG5V.n11243 0.0196384
R52702 ASIG5V.n11129 ASIG5V.n11128 0.0196384
R52703 ASIG5V.n11252 ASIG5V.n11249 0.0196384
R52704 ASIG5V.n11257 ASIG5V.n11254 0.0196384
R52705 ASIG5V.n11262 ASIG5V.n11259 0.0196384
R52706 ASIG5V.n11137 ASIG5V.n11136 0.0196384
R52707 ASIG5V.n11270 ASIG5V.n11267 0.0196384
R52708 ASIG5V.n11275 ASIG5V.n11272 0.0196384
R52709 ASIG5V.n11280 ASIG5V.n11277 0.0196384
R52710 ASIG5V.n11285 ASIG5V.n11282 0.0196384
R52711 ASIG5V.n11290 ASIG5V.n11287 0.0196384
R52712 ASIG5V.n11293 ASIG5V.n11292 0.0196384
R52713 ASIG5V.n11296 ASIG5V.n11294 0.0196384
R52714 ASIG5V.n11299 ASIG5V.n11297 0.0196384
R52715 ASIG5V.n11302 ASIG5V.n11300 0.0196384
R52716 ASIG5V.n11305 ASIG5V.n11303 0.0196384
R52717 ASIG5V.n11307 ASIG5V.n11306 0.0196384
R52718 ASIG5V.n11310 ASIG5V.n11308 0.0196384
R52719 ASIG5V.n11153 ASIG5V.n11152 0.0196384
R52720 ASIG5V.n8867 ASIG5V.n8865 0.0196384
R52721 ASIG5V.n2912 ASIG5V.n2911 0.0196384
R52722 ASIG5V.n2910 ASIG5V.n2909 0.0196384
R52723 ASIG5V.n2907 ASIG5V.n2906 0.0196384
R52724 ASIG5V.n2906 ASIG5V.n2905 0.0196384
R52725 ASIG5V.n2903 ASIG5V.n2902 0.0196384
R52726 ASIG5V.n2902 ASIG5V.n2901 0.0196384
R52727 ASIG5V.n2899 ASIG5V.n2898 0.0196384
R52728 ASIG5V.n2898 ASIG5V.n2897 0.0196384
R52729 ASIG5V.n2895 ASIG5V.n2894 0.0196384
R52730 ASIG5V.n2894 ASIG5V.n2893 0.0196384
R52731 ASIG5V.n2891 ASIG5V.n2890 0.0196384
R52732 ASIG5V.n2890 ASIG5V.n2889 0.0196384
R52733 ASIG5V.n2887 ASIG5V.n2886 0.0196384
R52734 ASIG5V.n2886 ASIG5V.n2885 0.0196384
R52735 ASIG5V.n2829 ASIG5V.n2828 0.0196384
R52736 ASIG5V.n3030 ASIG5V.n3028 0.0196384
R52737 ASIG5V.n3027 ASIG5V.n3025 0.0196384
R52738 ASIG5V.n3024 ASIG5V.n3022 0.0196384
R52739 ASIG5V.n3021 ASIG5V.n3019 0.0196384
R52740 ASIG5V.n3018 ASIG5V.n3016 0.0196384
R52741 ASIG5V.n3015 ASIG5V.n3013 0.0196384
R52742 ASIG5V.n3012 ASIG5V.n3011 0.0196384
R52743 ASIG5V.n3010 ASIG5V.n3008 0.0196384
R52744 ASIG5V.n3007 ASIG5V.n3005 0.0196384
R52745 ASIG5V.n3004 ASIG5V.n3003 0.0196384
R52746 ASIG5V.n3001 ASIG5V.n2998 0.0196384
R52747 ASIG5V.n2996 ASIG5V.n2993 0.0196384
R52748 ASIG5V.n2991 ASIG5V.n2990 0.0196384
R52749 ASIG5V.n2988 ASIG5V.n2985 0.0196384
R52750 ASIG5V.n2983 ASIG5V.n2980 0.0196384
R52751 ASIG5V.n2978 ASIG5V.n2977 0.0196384
R52752 ASIG5V.n2855 ASIG5V.n2854 0.0196384
R52753 ASIG5V.n2972 ASIG5V.n2969 0.0196384
R52754 ASIG5V.n2967 ASIG5V.n2964 0.0196384
R52755 ASIG5V.n2962 ASIG5V.n2959 0.0196384
R52756 ASIG5V.n2957 ASIG5V.n2954 0.0196384
R52757 ASIG5V.n2952 ASIG5V.n2951 0.0196384
R52758 ASIG5V.n2949 ASIG5V.n2948 0.0196384
R52759 ASIG5V.n2946 ASIG5V.n2943 0.0196384
R52760 ASIG5V.n2941 ASIG5V.n2940 0.0196384
R52761 ASIG5V.n2938 ASIG5V.n2935 0.0196384
R52762 ASIG5V.n2934 ASIG5V.n2933 0.0196384
R52763 ASIG5V.n2932 ASIG5V.n2930 0.0196384
R52764 ASIG5V.n2929 ASIG5V.n2927 0.0196384
R52765 ASIG5V.n2926 ASIG5V.n2924 0.0196384
R52766 ASIG5V.n2877 ASIG5V.n2876 0.0196384
R52767 ASIG5V.n2921 ASIG5V.n2919 0.0196384
R52768 ASIG5V.n2918 ASIG5V.n2916 0.0196384
R52769 ASIG5V.n2827 ASIG5V.n2826 0.0196384
R52770 ASIG5V.n2918 ASIG5V.n2917 0.0196384
R52771 ASIG5V.n2908 ASIG5V.n2907 0.0196384
R52772 ASIG5V.n2904 ASIG5V.n2903 0.0196384
R52773 ASIG5V.n2900 ASIG5V.n2899 0.0196384
R52774 ASIG5V.n2896 ASIG5V.n2895 0.0196384
R52775 ASIG5V.n2892 ASIG5V.n2891 0.0196384
R52776 ASIG5V.n2888 ASIG5V.n2887 0.0196384
R52777 ASIG5V.n3030 ASIG5V.n3029 0.0196384
R52778 ASIG5V.n3027 ASIG5V.n3026 0.0196384
R52779 ASIG5V.n3024 ASIG5V.n3023 0.0196384
R52780 ASIG5V.n3021 ASIG5V.n3020 0.0196384
R52781 ASIG5V.n3018 ASIG5V.n3017 0.0196384
R52782 ASIG5V.n3015 ASIG5V.n3014 0.0196384
R52783 ASIG5V.n3010 ASIG5V.n3009 0.0196384
R52784 ASIG5V.n3007 ASIG5V.n3006 0.0196384
R52785 ASIG5V.n3001 ASIG5V.n3000 0.0196384
R52786 ASIG5V.n2996 ASIG5V.n2995 0.0196384
R52787 ASIG5V.n2988 ASIG5V.n2987 0.0196384
R52788 ASIG5V.n2983 ASIG5V.n2982 0.0196384
R52789 ASIG5V.n2975 ASIG5V.n2974 0.0196384
R52790 ASIG5V.n2972 ASIG5V.n2971 0.0196384
R52791 ASIG5V.n2967 ASIG5V.n2966 0.0196384
R52792 ASIG5V.n2962 ASIG5V.n2961 0.0196384
R52793 ASIG5V.n2957 ASIG5V.n2956 0.0196384
R52794 ASIG5V.n2946 ASIG5V.n2945 0.0196384
R52795 ASIG5V.n2938 ASIG5V.n2937 0.0196384
R52796 ASIG5V.n2932 ASIG5V.n2931 0.0196384
R52797 ASIG5V.n2929 ASIG5V.n2928 0.0196384
R52798 ASIG5V.n2926 ASIG5V.n2925 0.0196384
R52799 ASIG5V.n2923 ASIG5V.n2922 0.0196384
R52800 ASIG5V.n2921 ASIG5V.n2920 0.0196384
R52801 ASIG5V.n2911 ASIG5V.n2910 0.0196384
R52802 ASIG5V.n2909 ASIG5V.n2908 0.0196384
R52803 ASIG5V.n2905 ASIG5V.n2904 0.0196384
R52804 ASIG5V.n2901 ASIG5V.n2900 0.0196384
R52805 ASIG5V.n2897 ASIG5V.n2896 0.0196384
R52806 ASIG5V.n2893 ASIG5V.n2892 0.0196384
R52807 ASIG5V.n2889 ASIG5V.n2888 0.0196384
R52808 ASIG5V.n2885 ASIG5V.n2884 0.0196384
R52809 ASIG5V.n2836 ASIG5V.n2835 0.0196384
R52810 ASIG5V.n2841 ASIG5V.n2840 0.0196384
R52811 ASIG5V.n2846 ASIG5V.n2845 0.0196384
R52812 ASIG5V.n2851 ASIG5V.n2850 0.0196384
R52813 ASIG5V.n2861 ASIG5V.n2860 0.0196384
R52814 ASIG5V.n2864 ASIG5V.n2863 0.0196384
R52815 ASIG5V.n2868 ASIG5V.n2867 0.0196384
R52816 ASIG5V.n2871 ASIG5V.n2870 0.0196384
R52817 ASIG5V.n2879 ASIG5V.n2878 0.0196384
R52818 ASIG5V.n8867 ASIG5V.n8866 0.0196384
R52819 ASIG5V.n11310 ASIG5V.n11309 0.0196384
R52820 ASIG5V.n11151 ASIG5V.n11150 0.0196384
R52821 ASIG5V.n11305 ASIG5V.n11304 0.0196384
R52822 ASIG5V.n11302 ASIG5V.n11301 0.0196384
R52823 ASIG5V.n11299 ASIG5V.n11298 0.0196384
R52824 ASIG5V.n11296 ASIG5V.n11295 0.0196384
R52825 ASIG5V.n11145 ASIG5V.n11144 0.0196384
R52826 ASIG5V.n11290 ASIG5V.n11289 0.0196384
R52827 ASIG5V.n11285 ASIG5V.n11284 0.0196384
R52828 ASIG5V.n11280 ASIG5V.n11279 0.0196384
R52829 ASIG5V.n11275 ASIG5V.n11274 0.0196384
R52830 ASIG5V.n11270 ASIG5V.n11269 0.0196384
R52831 ASIG5V.n11265 ASIG5V.n11264 0.0196384
R52832 ASIG5V.n11262 ASIG5V.n11261 0.0196384
R52833 ASIG5V.n11257 ASIG5V.n11256 0.0196384
R52834 ASIG5V.n11252 ASIG5V.n11251 0.0196384
R52835 ASIG5V.n11132 ASIG5V.n11131 0.0196384
R52836 ASIG5V.n11246 ASIG5V.n11245 0.0196384
R52837 ASIG5V.n11241 ASIG5V.n11240 0.0196384
R52838 ASIG5V.n11236 ASIG5V.n11235 0.0196384
R52839 ASIG5V.n11231 ASIG5V.n11230 0.0196384
R52840 ASIG5V.n11226 ASIG5V.n11225 0.0196384
R52841 ASIG5V.n11221 ASIG5V.n11220 0.0196384
R52842 ASIG5V.n11216 ASIG5V.n11215 0.0196384
R52843 ASIG5V.n11212 ASIG5V.n11211 0.0196384
R52844 ASIG5V.n11119 ASIG5V.n11118 0.0196384
R52845 ASIG5V.n11116 ASIG5V.n11115 0.0196384
R52846 ASIG5V.n11114 ASIG5V.n11113 0.0196384
R52847 ASIG5V.n11204 ASIG5V.n11203 0.0196384
R52848 ASIG5V.n11201 ASIG5V.n11200 0.0196384
R52849 ASIG5V.n11198 ASIG5V.n11197 0.0196384
R52850 ASIG5V.n11195 ASIG5V.n11194 0.0196384
R52851 ASIG5V.n11192 ASIG5V.n11191 0.0196384
R52852 ASIG5V.n11159 ASIG5V.n11158 0.0196384
R52853 ASIG5V.n11163 ASIG5V.n11162 0.0196384
R52854 ASIG5V.n11162 ASIG5V.n11161 0.0196384
R52855 ASIG5V.n11167 ASIG5V.n11166 0.0196384
R52856 ASIG5V.n11166 ASIG5V.n11165 0.0196384
R52857 ASIG5V.n11171 ASIG5V.n11170 0.0196384
R52858 ASIG5V.n11170 ASIG5V.n11169 0.0196384
R52859 ASIG5V.n11175 ASIG5V.n11174 0.0196384
R52860 ASIG5V.n11174 ASIG5V.n11173 0.0196384
R52861 ASIG5V.n11179 ASIG5V.n11178 0.0196384
R52862 ASIG5V.n11178 ASIG5V.n11177 0.0196384
R52863 ASIG5V.n11183 ASIG5V.n11182 0.0196384
R52864 ASIG5V.n11182 ASIG5V.n11181 0.0196384
R52865 ASIG5V.n11186 ASIG5V.n11185 0.0196384
R52866 ASIG5V.n9969 ASIG5V 0.0196322
R52867 ASIG5V.n13254 ASIG5V 0.0196322
R52868 ASIG5V ASIG5V.n401 0.0196322
R52869 ASIG5V.n9374 ASIG5V.n9373 0.019625
R52870 ASIG5V.n9421 ASIG5V.n9420 0.019625
R52871 ASIG5V.n9069 ASIG5V.n9068 0.0195611
R52872 ASIG5V.n9379 ASIG5V.n9378 0.019175
R52873 ASIG5V.n9416 ASIG5V.n9415 0.019175
R52874 ASIG5V.n733 ASIG5V.n732 0.0187751
R52875 ASIG5V.n1010 ASIG5V.n1009 0.018725
R52876 ASIG5V.n9769 ASIG5V.n9768 0.0176434
R52877 ASIG5V.n9777 ASIG5V.n9776 0.0176434
R52878 ASIG5V.n719 ASIG5V.n718 0.0175961
R52879 ASIG5V.n2496 ASIG5V.n2495 0.017282
R52880 ASIG5V.n2495 ASIG5V.n2494 0.017282
R52881 ASIG5V.n2492 ASIG5V.n2491 0.017282
R52882 ASIG5V.n2491 ASIG5V.n2490 0.017282
R52883 ASIG5V.n2488 ASIG5V.n2487 0.017282
R52884 ASIG5V.n2487 ASIG5V.n2486 0.017282
R52885 ASIG5V.n2484 ASIG5V.n2483 0.017282
R52886 ASIG5V.n2483 ASIG5V.n2482 0.017282
R52887 ASIG5V.n2480 ASIG5V.n2479 0.017282
R52888 ASIG5V.n2477 ASIG5V.n2476 0.017282
R52889 ASIG5V.n2476 ASIG5V.n2475 0.017282
R52890 ASIG5V.n2475 ASIG5V.n2474 0.017282
R52891 ASIG5V.n2474 ASIG5V.n2473 0.017282
R52892 ASIG5V.n2471 ASIG5V.n2470 0.017282
R52893 ASIG5V.n2470 ASIG5V.n2469 0.017282
R52894 ASIG5V.n2467 ASIG5V.n2466 0.017282
R52895 ASIG5V.n2185 ASIG5V.n2184 0.017282
R52896 ASIG5V.n2184 ASIG5V.n2183 0.017282
R52897 ASIG5V.n2181 ASIG5V.n2180 0.017282
R52898 ASIG5V.n2180 ASIG5V.n2179 0.017282
R52899 ASIG5V.n2179 ASIG5V.n2178 0.017282
R52900 ASIG5V.n10716 ASIG5V.n10715 0.017282
R52901 ASIG5V.n10717 ASIG5V.n10716 0.017282
R52902 ASIG5V.n10720 ASIG5V.n10719 0.017282
R52903 ASIG5V.n10721 ASIG5V.n10720 0.017282
R52904 ASIG5V.n10724 ASIG5V.n10723 0.017282
R52905 ASIG5V.n10725 ASIG5V.n10724 0.017282
R52906 ASIG5V.n10730 ASIG5V.n10729 0.017282
R52907 ASIG5V.n10731 ASIG5V.n10730 0.017282
R52908 ASIG5V.n10734 ASIG5V.n10733 0.017282
R52909 ASIG5V.n10735 ASIG5V.n10734 0.017282
R52910 ASIG5V.n10738 ASIG5V.n10737 0.017282
R52911 ASIG5V.n10743 ASIG5V.n10742 0.017282
R52912 ASIG5V.n10744 ASIG5V.n10743 0.017282
R52913 ASIG5V.n10747 ASIG5V.n10746 0.017282
R52914 ASIG5V.n10748 ASIG5V.n10747 0.017282
R52915 ASIG5V.n10749 ASIG5V.n10748 0.017282
R52916 ASIG5V.n10752 ASIG5V.n10751 0.017282
R52917 ASIG5V.n10753 ASIG5V.n10752 0.017282
R52918 ASIG5V.n10756 ASIG5V.n10755 0.017282
R52919 ASIG5V.n10757 ASIG5V.n10756 0.017282
R52920 ASIG5V.n9088 ASIG5V.n9087 0.0172031
R52921 ASIG5V.n10478 ASIG5V.n10477 0.0171683
R52922 ASIG5V.n992 ASIG5V.n991 0.016925
R52923 ASIG5V.n9866 ASIG5V.n9865 0.0168133
R52924 ASIG5V.n9838 ASIG5V.n9837 0.0168133
R52925 ASIG5V.n9811 ASIG5V.n9810 0.0168133
R52926 ASIG5V.n9083 ASIG5V.n9082 0.01681
R52927 ASIG5V.n2465 ASIG5V.n2187 0.0167406
R52928 ASIG5V.n10745 ASIG5V.n10744 0.0167406
R52929 ASIG5V.n10097 ASIG5V.n10096 0.0165881
R52930 ASIG5V.n9397 ASIG5V.n9396 0.016475
R52931 ASIG5V.n9398 ASIG5V.n9397 0.016475
R52932 ASIG5V.n10758 ASIG5V.n10757 0.0164699
R52933 ASIG5V.n1448 ASIG5V.n1447 0.0164246
R52934 ASIG5V.n714 ASIG5V.n713 0.016417
R52935 ASIG5V.n10729 ASIG5V.n10728 0.0161992
R52936 ASIG5V.n991 ASIG5V.n990 0.016025
R52937 ASIG5V.n13258 ASIG5V.n13257 0.0159671
R52938 ASIG5V.n13256 ASIG5V.n13255 0.0159671
R52939 ASIG5V.n13248 ASIG5V.n13247 0.0159671
R52940 ASIG5V.n2191 ASIG5V.n2190 0.0159671
R52941 ASIG5V.n2193 ASIG5V.n2192 0.0159671
R52942 ASIG5V.n1540 ASIG5V.n1539 0.0157064
R52943 ASIG5V.n1409 ASIG5V.n1408 0.0157064
R52944 ASIG5V.n1407 ASIG5V.n1406 0.0157064
R52945 ASIG5V.n2231 ASIG5V.n2230 0.0157064
R52946 ASIG5V.n2229 ASIG5V.n2228 0.0157064
R52947 ASIG5V.n2227 ASIG5V.n2226 0.0157064
R52948 ASIG5V.n13155 ASIG5V.n13154 0.0157064
R52949 ASIG5V.n13157 ASIG5V.n13156 0.0157064
R52950 ASIG5V.n9976 ASIG5V.n9975 0.0157064
R52951 ASIG5V.n9978 ASIG5V.n9977 0.0157064
R52952 ASIG5V.n10002 ASIG5V.n10001 0.0157064
R52953 ASIG5V.n12889 ASIG5V.n12888 0.0157064
R52954 ASIG5V.n10311 ASIG5V.n10310 0.0157064
R52955 ASIG5V.n1510 ASIG5V.n1509 0.0157064
R52956 ASIG5V.n1418 ASIG5V.n1417 0.0157064
R52957 ASIG5V.n1416 ASIG5V.n1415 0.0157064
R52958 ASIG5V.n2240 ASIG5V.n2239 0.0157064
R52959 ASIG5V.n2238 ASIG5V.n2237 0.0157064
R52960 ASIG5V.n2236 ASIG5V.n2235 0.0157064
R52961 ASIG5V.n7178 ASIG5V.n7177 0.0157064
R52962 ASIG5V.n7181 ASIG5V.n7180 0.0157064
R52963 ASIG5V.n13125 ASIG5V.n13124 0.0157064
R52964 ASIG5V.n13123 ASIG5V.n13122 0.0157064
R52965 ASIG5V.n13118 ASIG5V.n13117 0.0157064
R52966 ASIG5V.n10316 ASIG5V.n10315 0.0157064
R52967 ASIG5V.n10318 ASIG5V.n10317 0.0157064
R52968 ASIG5V.n10320 ASIG5V.n10319 0.0157064
R52969 ASIG5V.n10324 ASIG5V.n10323 0.0157064
R52970 ASIG5V.n1426 ASIG5V.n1425 0.0157064
R52971 ASIG5V.n1478 ASIG5V.n1477 0.0157064
R52972 ASIG5V.n2252 ASIG5V.n2243 0.0157064
R52973 ASIG5V.n2250 ASIG5V.n2249 0.0157064
R52974 ASIG5V.n2248 ASIG5V.n2247 0.0157064
R52975 ASIG5V.n2246 ASIG5V.n2245 0.0157064
R52976 ASIG5V.n13039 ASIG5V.n13038 0.0157064
R52977 ASIG5V.n13041 ASIG5V.n13040 0.0157064
R52978 ASIG5V.n13049 ASIG5V.n13048 0.0157064
R52979 ASIG5V.n13051 ASIG5V.n13050 0.0157064
R52980 ASIG5V.n13090 ASIG5V.n13089 0.0157064
R52981 ASIG5V.n10329 ASIG5V.n10328 0.0157064
R52982 ASIG5V.n10331 ASIG5V.n10330 0.0157064
R52983 ASIG5V.n10333 ASIG5V.n10332 0.0157064
R52984 ASIG5V.n10337 ASIG5V.n10336 0.0157064
R52985 ASIG5V.n2262 ASIG5V.n2261 0.0157064
R52986 ASIG5V.n2257 ASIG5V.n2256 0.0157064
R52987 ASIG5V.n2255 ASIG5V.n2254 0.0157064
R52988 ASIG5V.n12998 ASIG5V.n12997 0.0157064
R52989 ASIG5V.n12996 ASIG5V.n12995 0.0157064
R52990 ASIG5V.n12992 ASIG5V.n12991 0.0157064
R52991 ASIG5V.n12990 ASIG5V.n12989 0.0157064
R52992 ASIG5V.n12988 ASIG5V.n12987 0.0157064
R52993 ASIG5V.n12984 ASIG5V.n12983 0.0157064
R52994 ASIG5V.n12982 ASIG5V.n7208 0.0157064
R52995 ASIG5V.n12978 ASIG5V.n12977 0.0157064
R52996 ASIG5V.n9797 ASIG5V.n9796 0.0157064
R52997 ASIG5V.n9799 ASIG5V.n9798 0.0157064
R52998 ASIG5V.n9801 ASIG5V.n9800 0.0157064
R52999 ASIG5V.n2493 ASIG5V.n2492 0.0156579
R53000 ASIG5V.n2183 ASIG5V.n2182 0.0156579
R53001 ASIG5V.n10727 ASIG5V.n10726 0.0156579
R53002 ASIG5V.n2745 ASIG5V.n2744 0.0154799
R53003 ASIG5V.n2744 ASIG5V.n2743 0.0154799
R53004 ASIG5V.n2741 ASIG5V.n2740 0.0154799
R53005 ASIG5V.n2740 ASIG5V.n2739 0.0154799
R53006 ASIG5V.n2737 ASIG5V.n2736 0.0154799
R53007 ASIG5V.n2736 ASIG5V.n2735 0.0154799
R53008 ASIG5V.n2733 ASIG5V.n2732 0.0154799
R53009 ASIG5V.n2732 ASIG5V.n2731 0.0154799
R53010 ASIG5V.n10924 ASIG5V.n10923 0.0154799
R53011 ASIG5V.n10927 ASIG5V.n10926 0.0154799
R53012 ASIG5V.n10928 ASIG5V.n10927 0.0154799
R53013 ASIG5V.n10929 ASIG5V.n10928 0.0154799
R53014 ASIG5V.n10983 ASIG5V.n10982 0.0154799
R53015 ASIG5V.n10984 ASIG5V.n10983 0.0154799
R53016 ASIG5V.n11021 ASIG5V.n11020 0.0154799
R53017 ASIG5V.n11022 ASIG5V.n11021 0.0154799
R53018 ASIG5V.n12862 ASIG5V.n12857 0.015443
R53019 ASIG5V.n12891 ASIG5V.n12886 0.015443
R53020 ASIG5V.n12836 ASIG5V.n12835 0.015443
R53021 ASIG5V.n10061 ASIG5V.n10055 0.015443
R53022 ASIG5V.n10034 ASIG5V.n10033 0.015443
R53023 ASIG5V.n10006 ASIG5V.n10005 0.015443
R53024 ASIG5V.n12916 ASIG5V.n12915 0.015443
R53025 ASIG5V.n13121 ASIG5V.n7184 0.015443
R53026 ASIG5V.n13220 ASIG5V.n13214 0.015443
R53027 ASIG5V.n13193 ASIG5V.n13192 0.015443
R53028 ASIG5V.n13162 ASIG5V.n13161 0.015443
R53029 ASIG5V.n13131 ASIG5V.n13130 0.015443
R53030 ASIG5V.n12808 ASIG5V.n12803 0.015443
R53031 ASIG5V.n13263 ASIG5V.n13262 0.015443
R53032 ASIG5V.n13252 ASIG5V.n7169 0.015443
R53033 ASIG5V.n2111 ASIG5V.n2110 0.015443
R53034 ASIG5V.n2089 ASIG5V.n2088 0.015443
R53035 ASIG5V.n2064 ASIG5V.n2063 0.015443
R53036 ASIG5V.n2039 ASIG5V.n2038 0.015443
R53037 ASIG5V.n12941 ASIG5V.n12940 0.015443
R53038 ASIG5V.n13094 ASIG5V.n13093 0.015443
R53039 ASIG5V.n13045 ASIG5V.n7206 0.015443
R53040 ASIG5V.n2014 ASIG5V.n2013 0.015443
R53041 ASIG5V.n1602 ASIG5V.n1596 0.015443
R53042 ASIG5V.n1575 ASIG5V.n1574 0.015443
R53043 ASIG5V.n1545 ASIG5V.n1544 0.015443
R53044 ASIG5V.n1515 ASIG5V.n1514 0.015443
R53045 ASIG5V.n1485 ASIG5V.n1484 0.015443
R53046 ASIG5V.n1635 ASIG5V.n1634 0.015443
R53047 ASIG5V.n7145 ASIG5V.n7139 0.015443
R53048 ASIG5V.n2164 ASIG5V.n2163 0.015443
R53049 ASIG5V.n1665 ASIG5V.n1664 0.015443
R53050 ASIG5V.n12779 ASIG5V.n12773 0.015443
R53051 ASIG5V.n10454 ASIG5V.n10453 0.015443
R53052 ASIG5V.n10429 ASIG5V.n10428 0.015443
R53053 ASIG5V.n10404 ASIG5V.n10403 0.015443
R53054 ASIG5V.n10379 ASIG5V.n10378 0.015443
R53055 ASIG5V.n10485 ASIG5V.n10475 0.015443
R53056 ASIG5V.n10488 ASIG5V.n10487 0.015443
R53057 ASIG5V.n10516 ASIG5V.n10509 0.015443
R53058 ASIG5V.n1453 ASIG5V.n1452 0.015443
R53059 ASIG5V.n12981 ASIG5V.n12965 0.015443
R53060 ASIG5V.n13015 ASIG5V.n13014 0.015443
R53061 ASIG5V.n10100 ASIG5V.n10094 0.015443
R53062 ASIG5V.n9926 ASIG5V.n9925 0.015443
R53063 ASIG5V.n9898 ASIG5V.n9897 0.015443
R53064 ASIG5V.n9870 ASIG5V.n9869 0.015443
R53065 ASIG5V.n9842 ASIG5V.n9841 0.015443
R53066 ASIG5V.n10070 ASIG5V.n9947 0.015443
R53067 ASIG5V.n2401 ASIG5V.n2400 0.015443
R53068 ASIG5V.n2278 ASIG5V.n2277 0.015443
R53069 ASIG5V.n2379 ASIG5V.n2378 0.015443
R53070 ASIG5V.n2354 ASIG5V.n2353 0.015443
R53071 ASIG5V.n2329 ASIG5V.n2328 0.015443
R53072 ASIG5V.n2304 ASIG5V.n2303 0.015443
R53073 ASIG5V.n2429 ASIG5V.n2428 0.015443
R53074 ASIG5V.n2454 ASIG5V.n2453 0.015443
R53075 ASIG5V.n1400 ASIG5V.n1399 0.0152665
R53076 ASIG5V.n1398 ASIG5V.n1397 0.0152665
R53077 ASIG5V.n1389 ASIG5V.n1388 0.0152665
R53078 ASIG5V.n1380 ASIG5V.n1379 0.0152665
R53079 ASIG5V.n1570 ASIG5V.n1569 0.0152665
R53080 ASIG5V.n2222 ASIG5V.n2221 0.0152665
R53081 ASIG5V.n2220 ASIG5V.n2219 0.0152665
R53082 ASIG5V.n2218 ASIG5V.n2217 0.0152665
R53083 ASIG5V.n13186 ASIG5V.n13185 0.0152665
R53084 ASIG5V.n13188 ASIG5V.n13187 0.0152665
R53085 ASIG5V.n9971 ASIG5V.n9970 0.0152665
R53086 ASIG5V.n9973 ASIG5V.n9972 0.0152665
R53087 ASIG5V.n10030 ASIG5V.n10029 0.0152665
R53088 ASIG5V.n12860 ASIG5V.n12859 0.0152665
R53089 ASIG5V.n10302 ASIG5V.n10301 0.0152665
R53090 ASIG5V.n1600 ASIG5V.n1599 0.0152665
R53091 ASIG5V.n2211 ASIG5V.n2210 0.0152665
R53092 ASIG5V.n2209 ASIG5V.n2208 0.0152665
R53093 ASIG5V.n13218 ASIG5V.n13217 0.0152665
R53094 ASIG5V.n10060 ASIG5V.n10059 0.0152665
R53095 ASIG5V.n10481 ASIG5V.n10480 0.0152665
R53096 ASIG5V.n9744 ASIG5V.n9743 0.0152665
R53097 ASIG5V.n1630 ASIG5V.n1629 0.0152665
R53098 ASIG5V.n2201 ASIG5V.n2200 0.0152665
R53099 ASIG5V.n2199 ASIG5V.n2198 0.0152665
R53100 ASIG5V.n12806 ASIG5V.n12805 0.0152665
R53101 ASIG5V.n10512 ASIG5V.n10511 0.0152665
R53102 ASIG5V.n9736 ASIG5V.n9735 0.0152665
R53103 ASIG5V.n1660 ASIG5V.n1659 0.0152665
R53104 ASIG5V.n1372 ASIG5V.n1371 0.0152665
R53105 ASIG5V.n7142 ASIG5V.n7141 0.0152665
R53106 ASIG5V.n7144 ASIG5V.n7143 0.0152665
R53107 ASIG5V.n404 ASIG5V.n403 0.0152665
R53108 ASIG5V.n396 ASIG5V.n395 0.0152665
R53109 ASIG5V.n13288 ASIG5V.n13287 0.0152665
R53110 ASIG5V.n12776 ASIG5V.n12775 0.0152665
R53111 ASIG5V.n12778 ASIG5V.n12777 0.0152665
R53112 ASIG5V.n10545 ASIG5V.n10544 0.0152665
R53113 ASIG5V.n10560 ASIG5V.n10551 0.0152665
R53114 ASIG5V.n2479 ASIG5V.n2478 0.0151165
R53115 ASIG5V.n2177 ASIG5V.n2176 0.0151165
R53116 ASIG5V.n10925 ASIG5V.n10924 0.0149966
R53117 ASIG5V.n12894 ASIG5V.n12893 0.0147766
R53118 ASIG5V.n12865 ASIG5V.n12864 0.0147766
R53119 ASIG5V.n12833 ASIG5V.n12832 0.0147766
R53120 ASIG5V.n10063 ASIG5V.n9968 0.0147766
R53121 ASIG5V.n10031 ASIG5V.n10027 0.0147766
R53122 ASIG5V.n10003 ASIG5V.n9999 0.0147766
R53123 ASIG5V.n13119 ASIG5V.n13115 0.0147766
R53124 ASIG5V.n12919 ASIG5V.n12918 0.0147766
R53125 ASIG5V.n13128 ASIG5V.n7182 0.0147766
R53126 ASIG5V.n13223 ASIG5V.n13222 0.0147766
R53127 ASIG5V.n13190 ASIG5V.n13183 0.0147766
R53128 ASIG5V.n13159 ASIG5V.n13152 0.0147766
R53129 ASIG5V.n13250 ASIG5V.n13244 0.0147766
R53130 ASIG5V.n13260 ASIG5V.n399 0.0147766
R53131 ASIG5V.n12811 ASIG5V.n12810 0.0147766
R53132 ASIG5V.n2139 ASIG5V.n2138 0.0147766
R53133 ASIG5V.n2086 ASIG5V.n2085 0.0147766
R53134 ASIG5V.n2061 ASIG5V.n2060 0.0147766
R53135 ASIG5V.n2036 ASIG5V.n2035 0.0147766
R53136 ASIG5V.n2114 ASIG5V.n2113 0.0147766
R53137 ASIG5V.n2136 ASIG5V.n2135 0.0147766
R53138 ASIG5V.n2011 ASIG5V.n2010 0.0147766
R53139 ASIG5V.n13043 ASIG5V.n13036 0.0147766
R53140 ASIG5V.n13091 ASIG5V.n13087 0.0147766
R53141 ASIG5V.n12944 ASIG5V.n12943 0.0147766
R53142 ASIG5V.n1482 ASIG5V.n1474 0.0147766
R53143 ASIG5V.n1605 ASIG5V.n1604 0.0147766
R53144 ASIG5V.n1572 ASIG5V.n1566 0.0147766
R53145 ASIG5V.n1542 ASIG5V.n1536 0.0147766
R53146 ASIG5V.n1512 ASIG5V.n1506 0.0147766
R53147 ASIG5V.n1632 ASIG5V.n1626 0.0147766
R53148 ASIG5V.n13292 ASIG5V.n13291 0.0147766
R53149 ASIG5V.n13289 ASIG5V.n13284 0.0147766
R53150 ASIG5V.n12782 ASIG5V.n12781 0.0147766
R53151 ASIG5V.n1662 ASIG5V.n1656 0.0147766
R53152 ASIG5V.n2161 ASIG5V.n2160 0.0147766
R53153 ASIG5V.n7148 ASIG5V.n7147 0.0147766
R53154 ASIG5V.n10451 ASIG5V.n10450 0.0147766
R53155 ASIG5V.n10426 ASIG5V.n10425 0.0147766
R53156 ASIG5V.n10401 ASIG5V.n10400 0.0147766
R53157 ASIG5V.n10376 ASIG5V.n10375 0.0147766
R53158 ASIG5V.n10519 ASIG5V.n10518 0.0147766
R53159 ASIG5V.n10562 ASIG5V.n10561 0.0147766
R53160 ASIG5V.n10549 ASIG5V.n10540 0.0147766
R53161 ASIG5V.n1450 ASIG5V.n1444 0.0147766
R53162 ASIG5V.n13012 ASIG5V.n13009 0.0147766
R53163 ASIG5V.n12979 ASIG5V.n12976 0.0147766
R53164 ASIG5V.n9814 ASIG5V.n9813 0.0147766
R53165 ASIG5V.n10103 ASIG5V.n10102 0.0147766
R53166 ASIG5V.n9923 ASIG5V.n9919 0.0147766
R53167 ASIG5V.n9895 ASIG5V.n9891 0.0147766
R53168 ASIG5V.n9867 ASIG5V.n9863 0.0147766
R53169 ASIG5V.n9839 ASIG5V.n9835 0.0147766
R53170 ASIG5V.n10073 ASIG5V.n10072 0.0147766
R53171 ASIG5V.n9808 ASIG5V.n9793 0.0147766
R53172 ASIG5V.n2404 ASIG5V.n2403 0.0147766
R53173 ASIG5V.n2376 ASIG5V.n2375 0.0147766
R53174 ASIG5V.n2351 ASIG5V.n2350 0.0147766
R53175 ASIG5V.n2326 ASIG5V.n2325 0.0147766
R53176 ASIG5V.n2301 ASIG5V.n2299 0.0147766
R53177 ASIG5V.n2426 ASIG5V.n2425 0.0147766
R53178 ASIG5V.n2451 ASIG5V.n2450 0.0147766
R53179 ASIG5V.n2275 ASIG5V.n2274 0.0147766
R53180 ASIG5V.n11097 ASIG5V.n11096 0.014755
R53181 ASIG5V.n11023 ASIG5V.n11022 0.014755
R53182 ASIG5V.n10722 ASIG5V.n10721 0.0145752
R53183 ASIG5V.n12354 ASIG5V.n12353 0.014452
R53184 ASIG5V.n9064 ASIG5V.n9063 0.014452
R53185 ASIG5V.n9065 ASIG5V.n9064 0.014452
R53186 ASIG5V.n1150 ASIG5V.n1149 0.01445
R53187 ASIG5V.n1148 ASIG5V.n1147 0.01445
R53188 ASIG5V.n1147 ASIG5V.n1146 0.01445
R53189 ASIG5V.n1146 ASIG5V.n1145 0.01445
R53190 ASIG5V.n1145 ASIG5V.n1144 0.01445
R53191 ASIG5V.n1144 ASIG5V.n1143 0.01445
R53192 ASIG5V.n1143 ASIG5V.n1142 0.01445
R53193 ASIG5V.n1142 ASIG5V.n1141 0.01445
R53194 ASIG5V.n1141 ASIG5V.n1140 0.01445
R53195 ASIG5V.n1140 ASIG5V.n1139 0.01445
R53196 ASIG5V.n1139 ASIG5V.n1138 0.01445
R53197 ASIG5V.n1138 ASIG5V.n1137 0.01445
R53198 ASIG5V.n1137 ASIG5V.n1136 0.01445
R53199 ASIG5V.n1136 ASIG5V.n1135 0.01445
R53200 ASIG5V.n1135 ASIG5V.n1134 0.01445
R53201 ASIG5V.n1134 ASIG5V.n1133 0.01445
R53202 ASIG5V.n1133 ASIG5V.n1132 0.01445
R53203 ASIG5V.n1132 ASIG5V.n1131 0.01445
R53204 ASIG5V.n1131 ASIG5V.n1130 0.01445
R53205 ASIG5V.n1130 ASIG5V.n1129 0.01445
R53206 ASIG5V.n1129 ASIG5V.n1128 0.01445
R53207 ASIG5V.n1128 ASIG5V.n1127 0.01445
R53208 ASIG5V.n1127 ASIG5V.n1126 0.01445
R53209 ASIG5V.n1126 ASIG5V.n1125 0.01445
R53210 ASIG5V.n1125 ASIG5V.n1124 0.01445
R53211 ASIG5V.n1124 ASIG5V.n1123 0.01445
R53212 ASIG5V.n1123 ASIG5V.n1122 0.01445
R53213 ASIG5V.n1122 ASIG5V.n1121 0.01445
R53214 ASIG5V.n1121 ASIG5V.n1120 0.01445
R53215 ASIG5V.n1120 ASIG5V.n1119 0.01445
R53216 ASIG5V.n1119 ASIG5V.n1118 0.01445
R53217 ASIG5V.n1118 ASIG5V.n1117 0.01445
R53218 ASIG5V.n1117 ASIG5V.n1116 0.01445
R53219 ASIG5V.n1116 ASIG5V.n1115 0.01445
R53220 ASIG5V.n1115 ASIG5V.n1114 0.01445
R53221 ASIG5V.n1114 ASIG5V.n1113 0.01445
R53222 ASIG5V.n1113 ASIG5V.n1112 0.01445
R53223 ASIG5V.n1112 ASIG5V.n1111 0.01445
R53224 ASIG5V.n1111 ASIG5V.n1110 0.01445
R53225 ASIG5V.n1110 ASIG5V.n1109 0.01445
R53226 ASIG5V.n1109 ASIG5V.n1108 0.01445
R53227 ASIG5V.n1108 ASIG5V.n1107 0.01445
R53228 ASIG5V.n1107 ASIG5V.n1106 0.01445
R53229 ASIG5V.n1106 ASIG5V.n1105 0.01445
R53230 ASIG5V.n1105 ASIG5V.n1104 0.01445
R53231 ASIG5V.n1104 ASIG5V.n1103 0.01445
R53232 ASIG5V.n1103 ASIG5V.n1102 0.01445
R53233 ASIG5V.n1102 ASIG5V.n1101 0.01445
R53234 ASIG5V.n1101 ASIG5V.n1100 0.01445
R53235 ASIG5V.n1100 ASIG5V.n1099 0.01445
R53236 ASIG5V.n1099 ASIG5V.n1098 0.01445
R53237 ASIG5V.n1098 ASIG5V.n1097 0.01445
R53238 ASIG5V.n1097 ASIG5V.n1096 0.01445
R53239 ASIG5V.n1096 ASIG5V.n1095 0.01445
R53240 ASIG5V.n1095 ASIG5V.n1094 0.01445
R53241 ASIG5V.n1094 ASIG5V.n1093 0.01445
R53242 ASIG5V.n1093 ASIG5V.n1092 0.01445
R53243 ASIG5V.n1092 ASIG5V.n1091 0.01445
R53244 ASIG5V.n1091 ASIG5V.n1090 0.01445
R53245 ASIG5V.n1090 ASIG5V.n1089 0.01445
R53246 ASIG5V.n1089 ASIG5V.n1088 0.01445
R53247 ASIG5V.n1088 ASIG5V.n1087 0.01445
R53248 ASIG5V.n1087 ASIG5V.n1086 0.01445
R53249 ASIG5V.n1086 ASIG5V.n1085 0.01445
R53250 ASIG5V.n1085 ASIG5V.n1084 0.01445
R53251 ASIG5V.n1084 ASIG5V.n1083 0.01445
R53252 ASIG5V.n1083 ASIG5V.n1082 0.01445
R53253 ASIG5V.n1082 ASIG5V.n1081 0.01445
R53254 ASIG5V.n1081 ASIG5V.n1080 0.01445
R53255 ASIG5V.n1080 ASIG5V.n1079 0.01445
R53256 ASIG5V.n1079 ASIG5V.n1078 0.01445
R53257 ASIG5V.n1078 ASIG5V.n1077 0.01445
R53258 ASIG5V.n1077 ASIG5V.n1076 0.01445
R53259 ASIG5V.n1076 ASIG5V.n1075 0.01445
R53260 ASIG5V.n1075 ASIG5V.n1074 0.01445
R53261 ASIG5V.n1074 ASIG5V.n1073 0.01445
R53262 ASIG5V.n1073 ASIG5V.n1072 0.01445
R53263 ASIG5V.n1072 ASIG5V.n1071 0.01445
R53264 ASIG5V.n592 ASIG5V.n591 0.01445
R53265 ASIG5V.n597 ASIG5V.n596 0.01445
R53266 ASIG5V.n598 ASIG5V.n597 0.01445
R53267 ASIG5V.n607 ASIG5V.n606 0.01445
R53268 ASIG5V.n608 ASIG5V.n607 0.01445
R53269 ASIG5V.n609 ASIG5V.n608 0.01445
R53270 ASIG5V.n610 ASIG5V.n609 0.01445
R53271 ASIG5V.n614 ASIG5V.n613 0.01445
R53272 ASIG5V.n2817 ASIG5V.n2816 0.01445
R53273 ASIG5V.n2815 ASIG5V.n2814 0.01445
R53274 ASIG5V.n2814 ASIG5V.n2813 0.01445
R53275 ASIG5V.n2813 ASIG5V.n2812 0.01445
R53276 ASIG5V.n2812 ASIG5V.n2811 0.01445
R53277 ASIG5V.n2811 ASIG5V.n2810 0.01445
R53278 ASIG5V.n2810 ASIG5V.n2809 0.01445
R53279 ASIG5V.n2809 ASIG5V.n2808 0.01445
R53280 ASIG5V.n2808 ASIG5V.n2807 0.01445
R53281 ASIG5V.n2807 ASIG5V.n2806 0.01445
R53282 ASIG5V.n2806 ASIG5V.n2805 0.01445
R53283 ASIG5V.n2805 ASIG5V.n2804 0.01445
R53284 ASIG5V.n2804 ASIG5V.n2803 0.01445
R53285 ASIG5V.n2803 ASIG5V.n2802 0.01445
R53286 ASIG5V.n2802 ASIG5V.n2801 0.01445
R53287 ASIG5V.n2801 ASIG5V.n2800 0.01445
R53288 ASIG5V.n2800 ASIG5V.n2799 0.01445
R53289 ASIG5V.n2799 ASIG5V.n2798 0.01445
R53290 ASIG5V.n2798 ASIG5V.n2797 0.01445
R53291 ASIG5V.n2797 ASIG5V.n2796 0.01445
R53292 ASIG5V.n2796 ASIG5V.n2795 0.01445
R53293 ASIG5V.n2795 ASIG5V.n2794 0.01445
R53294 ASIG5V.n2794 ASIG5V.n2793 0.01445
R53295 ASIG5V.n2793 ASIG5V.n2792 0.01445
R53296 ASIG5V.n2792 ASIG5V.n2791 0.01445
R53297 ASIG5V.n2791 ASIG5V.n2790 0.01445
R53298 ASIG5V.n2790 ASIG5V.n2789 0.01445
R53299 ASIG5V.n2789 ASIG5V.n2788 0.01445
R53300 ASIG5V.n2788 ASIG5V.n2787 0.01445
R53301 ASIG5V.n2787 ASIG5V.n2786 0.01445
R53302 ASIG5V.n2786 ASIG5V.n2785 0.01445
R53303 ASIG5V.n2785 ASIG5V.n2784 0.01445
R53304 ASIG5V.n2784 ASIG5V.n2783 0.01445
R53305 ASIG5V.n2783 ASIG5V.n2782 0.01445
R53306 ASIG5V.n2782 ASIG5V.n2781 0.01445
R53307 ASIG5V.n2781 ASIG5V.n2780 0.01445
R53308 ASIG5V.n2780 ASIG5V.n2779 0.01445
R53309 ASIG5V.n2779 ASIG5V.n2778 0.01445
R53310 ASIG5V.n2778 ASIG5V.n2777 0.01445
R53311 ASIG5V.n2777 ASIG5V.n2776 0.01445
R53312 ASIG5V.n2776 ASIG5V.n2775 0.01445
R53313 ASIG5V.n2775 ASIG5V.n2774 0.01445
R53314 ASIG5V.n2774 ASIG5V.n2773 0.01445
R53315 ASIG5V.n2773 ASIG5V.n2772 0.01445
R53316 ASIG5V.n2772 ASIG5V.n2771 0.01445
R53317 ASIG5V.n2771 ASIG5V.n2770 0.01445
R53318 ASIG5V.n2770 ASIG5V.n2769 0.01445
R53319 ASIG5V.n2769 ASIG5V.n2768 0.01445
R53320 ASIG5V.n2768 ASIG5V.n2767 0.01445
R53321 ASIG5V.n2767 ASIG5V.n2766 0.01445
R53322 ASIG5V.n2766 ASIG5V.n2765 0.01445
R53323 ASIG5V.n2765 ASIG5V.n2764 0.01445
R53324 ASIG5V.n2764 ASIG5V.n2763 0.01445
R53325 ASIG5V.n2763 ASIG5V.n2762 0.01445
R53326 ASIG5V.n2762 ASIG5V.n2761 0.01445
R53327 ASIG5V.n2761 ASIG5V.n2760 0.01445
R53328 ASIG5V.n2760 ASIG5V.n2759 0.01445
R53329 ASIG5V.n2759 ASIG5V.n2758 0.01445
R53330 ASIG5V.n2758 ASIG5V.n2757 0.01445
R53331 ASIG5V.n2757 ASIG5V.n2756 0.01445
R53332 ASIG5V.n2756 ASIG5V.n2755 0.01445
R53333 ASIG5V.n2755 ASIG5V.n2754 0.01445
R53334 ASIG5V.n2754 ASIG5V.n2753 0.01445
R53335 ASIG5V.n2753 ASIG5V.n2752 0.01445
R53336 ASIG5V.n2752 ASIG5V.n2751 0.01445
R53337 ASIG5V.n2751 ASIG5V.n2750 0.01445
R53338 ASIG5V.n2750 ASIG5V.n2749 0.01445
R53339 ASIG5V.n2749 ASIG5V.n2748 0.01445
R53340 ASIG5V.n2748 ASIG5V.n2747 0.01445
R53341 ASIG5V.n578 ASIG5V.n577 0.01445
R53342 ASIG5V.n579 ASIG5V.n578 0.01445
R53343 ASIG5V.n580 ASIG5V.n579 0.01445
R53344 ASIG5V.n581 ASIG5V.n580 0.01445
R53345 ASIG5V.n582 ASIG5V.n581 0.01445
R53346 ASIG5V.n583 ASIG5V.n582 0.01445
R53347 ASIG5V.n584 ASIG5V.n583 0.01445
R53348 ASIG5V.n585 ASIG5V.n584 0.01445
R53349 ASIG5V.n587 ASIG5V.n585 0.01445
R53350 ASIG5V.n589 ASIG5V.n587 0.01445
R53351 ASIG5V.n590 ASIG5V.n589 0.01445
R53352 ASIG5V.n593 ASIG5V.n590 0.01445
R53353 ASIG5V.n594 ASIG5V.n593 0.01445
R53354 ASIG5V.n595 ASIG5V.n594 0.01445
R53355 ASIG5V.n599 ASIG5V.n595 0.01445
R53356 ASIG5V.n601 ASIG5V.n599 0.01445
R53357 ASIG5V.n602 ASIG5V.n601 0.01445
R53358 ASIG5V.n603 ASIG5V.n602 0.01445
R53359 ASIG5V.n604 ASIG5V.n603 0.01445
R53360 ASIG5V.n605 ASIG5V.n604 0.01445
R53361 ASIG5V.n611 ASIG5V.n605 0.01445
R53362 ASIG5V.n612 ASIG5V.n611 0.01445
R53363 ASIG5V.n615 ASIG5V.n612 0.01445
R53364 ASIG5V.n9515 ASIG5V.n9514 0.01445
R53365 ASIG5V.n9513 ASIG5V.n9512 0.01445
R53366 ASIG5V.n9512 ASIG5V.n9511 0.01445
R53367 ASIG5V.n9511 ASIG5V.n9510 0.01445
R53368 ASIG5V.n9510 ASIG5V.n9509 0.01445
R53369 ASIG5V.n9509 ASIG5V.n9508 0.01445
R53370 ASIG5V.n9508 ASIG5V.n9507 0.01445
R53371 ASIG5V.n9507 ASIG5V.n9506 0.01445
R53372 ASIG5V.n9506 ASIG5V.n9505 0.01445
R53373 ASIG5V.n9505 ASIG5V.n9504 0.01445
R53374 ASIG5V.n9504 ASIG5V.n9503 0.01445
R53375 ASIG5V.n9503 ASIG5V.n9502 0.01445
R53376 ASIG5V.n9502 ASIG5V.n9501 0.01445
R53377 ASIG5V.n9501 ASIG5V.n9500 0.01445
R53378 ASIG5V.n9500 ASIG5V.n9499 0.01445
R53379 ASIG5V.n9499 ASIG5V.n9498 0.01445
R53380 ASIG5V.n9498 ASIG5V.n9497 0.01445
R53381 ASIG5V.n9497 ASIG5V.n9496 0.01445
R53382 ASIG5V.n9496 ASIG5V.n9495 0.01445
R53383 ASIG5V.n9495 ASIG5V.n9494 0.01445
R53384 ASIG5V.n9494 ASIG5V.n9493 0.01445
R53385 ASIG5V.n9493 ASIG5V.n9492 0.01445
R53386 ASIG5V.n9492 ASIG5V.n9491 0.01445
R53387 ASIG5V.n9491 ASIG5V.n9490 0.01445
R53388 ASIG5V.n9490 ASIG5V.n9489 0.01445
R53389 ASIG5V.n9489 ASIG5V.n9488 0.01445
R53390 ASIG5V.n9488 ASIG5V.n9487 0.01445
R53391 ASIG5V.n9487 ASIG5V.n9486 0.01445
R53392 ASIG5V.n9486 ASIG5V.n9485 0.01445
R53393 ASIG5V.n9485 ASIG5V.n9484 0.01445
R53394 ASIG5V.n9484 ASIG5V.n9483 0.01445
R53395 ASIG5V.n9483 ASIG5V.n9482 0.01445
R53396 ASIG5V.n9482 ASIG5V.n9481 0.01445
R53397 ASIG5V.n9481 ASIG5V.n9480 0.01445
R53398 ASIG5V.n9480 ASIG5V.n9479 0.01445
R53399 ASIG5V.n9479 ASIG5V.n9478 0.01445
R53400 ASIG5V.n9478 ASIG5V.n9477 0.01445
R53401 ASIG5V.n9477 ASIG5V.n9476 0.01445
R53402 ASIG5V.n9476 ASIG5V.n9475 0.01445
R53403 ASIG5V.n9475 ASIG5V.n9474 0.01445
R53404 ASIG5V.n9474 ASIG5V.n9473 0.01445
R53405 ASIG5V.n9473 ASIG5V.n9472 0.01445
R53406 ASIG5V.n9472 ASIG5V.n9471 0.01445
R53407 ASIG5V.n9471 ASIG5V.n9470 0.01445
R53408 ASIG5V.n9470 ASIG5V.n9469 0.01445
R53409 ASIG5V.n9469 ASIG5V.n9468 0.01445
R53410 ASIG5V.n9468 ASIG5V.n9467 0.01445
R53411 ASIG5V.n9467 ASIG5V.n9466 0.01445
R53412 ASIG5V.n9466 ASIG5V.n9465 0.01445
R53413 ASIG5V.n9465 ASIG5V.n9464 0.01445
R53414 ASIG5V.n9464 ASIG5V.n9463 0.01445
R53415 ASIG5V.n9463 ASIG5V.n9462 0.01445
R53416 ASIG5V.n9462 ASIG5V.n9461 0.01445
R53417 ASIG5V.n9461 ASIG5V.n9460 0.01445
R53418 ASIG5V.n9460 ASIG5V.n9459 0.01445
R53419 ASIG5V.n9459 ASIG5V.n9458 0.01445
R53420 ASIG5V.n9458 ASIG5V.n9457 0.01445
R53421 ASIG5V.n9457 ASIG5V.n9456 0.01445
R53422 ASIG5V.n9456 ASIG5V.n9455 0.01445
R53423 ASIG5V.n9455 ASIG5V.n9454 0.01445
R53424 ASIG5V.n9454 ASIG5V.n9453 0.01445
R53425 ASIG5V.n9453 ASIG5V.n9452 0.01445
R53426 ASIG5V.n9452 ASIG5V.n9451 0.01445
R53427 ASIG5V.n9451 ASIG5V.n9450 0.01445
R53428 ASIG5V.n9450 ASIG5V.n9449 0.01445
R53429 ASIG5V.n9449 ASIG5V.n9448 0.01445
R53430 ASIG5V.n9448 ASIG5V.n9447 0.01445
R53431 ASIG5V.n9447 ASIG5V.n9446 0.01445
R53432 ASIG5V.n9446 ASIG5V.n9445 0.01445
R53433 ASIG5V.n9445 ASIG5V.n9444 0.01445
R53434 ASIG5V.n9444 ASIG5V.n9443 0.01445
R53435 ASIG5V.n9443 ASIG5V.n9442 0.01445
R53436 ASIG5V.n9442 ASIG5V.n9441 0.01445
R53437 ASIG5V.n9441 ASIG5V.n9440 0.01445
R53438 ASIG5V.n9440 ASIG5V.n9439 0.01445
R53439 ASIG5V.n9439 ASIG5V.n9438 0.01445
R53440 ASIG5V.n9438 ASIG5V.n9437 0.01445
R53441 ASIG5V.n9437 ASIG5V.n9436 0.01445
R53442 ASIG5V.n8950 ASIG5V.n8949 0.01445
R53443 ASIG5V.n8951 ASIG5V.n8950 0.01445
R53444 ASIG5V.n8955 ASIG5V.n8954 0.01445
R53445 ASIG5V.n8967 ASIG5V.n8966 0.01445
R53446 ASIG5V.n8968 ASIG5V.n8967 0.01445
R53447 ASIG5V.n8969 ASIG5V.n8968 0.01445
R53448 ASIG5V.n11094 ASIG5V.n11093 0.01445
R53449 ASIG5V.n11092 ASIG5V.n11091 0.01445
R53450 ASIG5V.n11091 ASIG5V.n11090 0.01445
R53451 ASIG5V.n11090 ASIG5V.n11089 0.01445
R53452 ASIG5V.n11089 ASIG5V.n11088 0.01445
R53453 ASIG5V.n11088 ASIG5V.n11087 0.01445
R53454 ASIG5V.n11087 ASIG5V.n11086 0.01445
R53455 ASIG5V.n11086 ASIG5V.n11085 0.01445
R53456 ASIG5V.n11085 ASIG5V.n11084 0.01445
R53457 ASIG5V.n11084 ASIG5V.n11083 0.01445
R53458 ASIG5V.n11083 ASIG5V.n11082 0.01445
R53459 ASIG5V.n11082 ASIG5V.n11081 0.01445
R53460 ASIG5V.n11081 ASIG5V.n11080 0.01445
R53461 ASIG5V.n11080 ASIG5V.n11079 0.01445
R53462 ASIG5V.n11079 ASIG5V.n11078 0.01445
R53463 ASIG5V.n11078 ASIG5V.n11077 0.01445
R53464 ASIG5V.n11077 ASIG5V.n11076 0.01445
R53465 ASIG5V.n11076 ASIG5V.n11075 0.01445
R53466 ASIG5V.n11075 ASIG5V.n11074 0.01445
R53467 ASIG5V.n11074 ASIG5V.n11073 0.01445
R53468 ASIG5V.n11073 ASIG5V.n11072 0.01445
R53469 ASIG5V.n11072 ASIG5V.n11071 0.01445
R53470 ASIG5V.n11071 ASIG5V.n11070 0.01445
R53471 ASIG5V.n11070 ASIG5V.n11069 0.01445
R53472 ASIG5V.n11069 ASIG5V.n11068 0.01445
R53473 ASIG5V.n11068 ASIG5V.n11067 0.01445
R53474 ASIG5V.n11067 ASIG5V.n11066 0.01445
R53475 ASIG5V.n11066 ASIG5V.n11065 0.01445
R53476 ASIG5V.n11065 ASIG5V.n11064 0.01445
R53477 ASIG5V.n11064 ASIG5V.n11063 0.01445
R53478 ASIG5V.n11063 ASIG5V.n11062 0.01445
R53479 ASIG5V.n11062 ASIG5V.n11061 0.01445
R53480 ASIG5V.n11061 ASIG5V.n11060 0.01445
R53481 ASIG5V.n11060 ASIG5V.n11059 0.01445
R53482 ASIG5V.n11059 ASIG5V.n11058 0.01445
R53483 ASIG5V.n11058 ASIG5V.n11057 0.01445
R53484 ASIG5V.n11057 ASIG5V.n11056 0.01445
R53485 ASIG5V.n11056 ASIG5V.n11055 0.01445
R53486 ASIG5V.n11055 ASIG5V.n11054 0.01445
R53487 ASIG5V.n11054 ASIG5V.n11053 0.01445
R53488 ASIG5V.n11053 ASIG5V.n11052 0.01445
R53489 ASIG5V.n11052 ASIG5V.n11051 0.01445
R53490 ASIG5V.n11051 ASIG5V.n11050 0.01445
R53491 ASIG5V.n11050 ASIG5V.n11049 0.01445
R53492 ASIG5V.n11049 ASIG5V.n11048 0.01445
R53493 ASIG5V.n11048 ASIG5V.n11047 0.01445
R53494 ASIG5V.n11047 ASIG5V.n11046 0.01445
R53495 ASIG5V.n11046 ASIG5V.n11045 0.01445
R53496 ASIG5V.n11045 ASIG5V.n11044 0.01445
R53497 ASIG5V.n11044 ASIG5V.n11043 0.01445
R53498 ASIG5V.n11043 ASIG5V.n11042 0.01445
R53499 ASIG5V.n11042 ASIG5V.n11041 0.01445
R53500 ASIG5V.n11041 ASIG5V.n11040 0.01445
R53501 ASIG5V.n11040 ASIG5V.n11039 0.01445
R53502 ASIG5V.n11039 ASIG5V.n11038 0.01445
R53503 ASIG5V.n11038 ASIG5V.n11037 0.01445
R53504 ASIG5V.n11037 ASIG5V.n11036 0.01445
R53505 ASIG5V.n11036 ASIG5V.n11035 0.01445
R53506 ASIG5V.n11035 ASIG5V.n11034 0.01445
R53507 ASIG5V.n11034 ASIG5V.n11033 0.01445
R53508 ASIG5V.n11033 ASIG5V.n11032 0.01445
R53509 ASIG5V.n11032 ASIG5V.n11031 0.01445
R53510 ASIG5V.n11031 ASIG5V.n11030 0.01445
R53511 ASIG5V.n11030 ASIG5V.n11029 0.01445
R53512 ASIG5V.n11029 ASIG5V.n11028 0.01445
R53513 ASIG5V.n11028 ASIG5V.n11027 0.01445
R53514 ASIG5V.n11027 ASIG5V.n11026 0.01445
R53515 ASIG5V.n11026 ASIG5V.n11025 0.01445
R53516 ASIG5V.n11025 ASIG5V.n11024 0.01445
R53517 ASIG5V.n8937 ASIG5V.n8936 0.01445
R53518 ASIG5V.n8938 ASIG5V.n8937 0.01445
R53519 ASIG5V.n8939 ASIG5V.n8938 0.01445
R53520 ASIG5V.n8940 ASIG5V.n8939 0.01445
R53521 ASIG5V.n8941 ASIG5V.n8940 0.01445
R53522 ASIG5V.n8942 ASIG5V.n8941 0.01445
R53523 ASIG5V.n8943 ASIG5V.n8942 0.01445
R53524 ASIG5V.n8944 ASIG5V.n8943 0.01445
R53525 ASIG5V.n8946 ASIG5V.n8944 0.01445
R53526 ASIG5V.n8947 ASIG5V.n8946 0.01445
R53527 ASIG5V.n8948 ASIG5V.n8947 0.01445
R53528 ASIG5V.n8952 ASIG5V.n8948 0.01445
R53529 ASIG5V.n8953 ASIG5V.n8952 0.01445
R53530 ASIG5V.n8956 ASIG5V.n8953 0.01445
R53531 ASIG5V.n8958 ASIG5V.n8956 0.01445
R53532 ASIG5V.n8960 ASIG5V.n8958 0.01445
R53533 ASIG5V.n8962 ASIG5V.n8960 0.01445
R53534 ASIG5V.n8963 ASIG5V.n8962 0.01445
R53535 ASIG5V.n8964 ASIG5V.n8963 0.01445
R53536 ASIG5V.n8965 ASIG5V.n8964 0.01445
R53537 ASIG5V.n8970 ASIG5V.n8965 0.01445
R53538 ASIG5V.n8972 ASIG5V.n8970 0.01445
R53539 ASIG5V.n2497 ASIG5V.n2496 0.0143045
R53540 ASIG5V.n1011 ASIG5V.n1010 0.014225
R53541 ASIG5V.n5675 ASIG5V.n5672 0.014059
R53542 ASIG5V.n5674 ASIG5V.n5673 0.014059
R53543 ASIG5V.n10751 ASIG5V.n10750 0.0140338
R53544 ASIG5V.n2742 ASIG5V.n2741 0.0140302
R53545 ASIG5V.n11413 ASIG5V.n11412 0.013791
R53546 ASIG5V.n9378 ASIG5V.n9377 0.013775
R53547 ASIG5V.n9417 ASIG5V.n9416 0.013775
R53548 ASIG5V.n2482 ASIG5V.n2481 0.0134925
R53549 ASIG5V.n2472 ASIG5V.n2471 0.0134925
R53550 ASIG5V.n11483 ASIG5V.n11482 0.01346
R53551 ASIG5V.n9375 ASIG5V.n9374 0.013325
R53552 ASIG5V.n9420 ASIG5V.n9419 0.013325
R53553 ASIG5V.n13246 ASIG5V.n13245 0.0132748
R53554 ASIG5V.n1447 ASIG5V.n1446 0.0130845
R53555 ASIG5V.n9922 ASIG5V.n9921 0.0130199
R53556 ASIG5V.n10069 ASIG5V.n10068 0.0130199
R53557 ASIG5V.n10554 ASIG5V.n10553 0.0130199
R53558 ASIG5V.n10740 ASIG5V.n10739 0.0129511
R53559 ASIG5V.n10741 ASIG5V.n10740 0.0129511
R53560 ASIG5V.n1014 ASIG5V.n1013 0.012875
R53561 ASIG5V.n2820 ASIG5V.n2819 0.0128221
R53562 ASIG5V.n2746 ASIG5V.n2745 0.0128221
R53563 ASIG5V.n9894 ASIG5V.n9893 0.0128209
R53564 ASIG5V.n9760 ASIG5V.n9759 0.0126672
R53565 ASIG5V.n9752 ASIG5V.n9751 0.0126436
R53566 ASIG5V.n1374 ASIG5V.n1373 0.0126436
R53567 ASIG5V.n1569 ASIG5V.n1568 0.0126296
R53568 ASIG5V.n1599 ASIG5V.n1598 0.0126296
R53569 ASIG5V.n1629 ASIG5V.n1628 0.0126296
R53570 ASIG5V.n1659 ASIG5V.n1658 0.0126296
R53571 ASIG5V.n10982 ASIG5V.n10981 0.0125805
R53572 ASIG5V.n4098 ASIG5V.n4097 0.0124869
R53573 ASIG5V.n715 ASIG5V.n714 0.0124869
R53574 ASIG5V.n1539 ASIG5V.n1538 0.0124187
R53575 ASIG5V.n1509 ASIG5V.n1508 0.0124187
R53576 ASIG5V.n1426 ASIG5V.n1423 0.0124187
R53577 ASIG5V.n10733 ASIG5V.n10732 0.0124098
R53578 ASIG5V.n11096 ASIG5V.n10761 0.0123125
R53579 ASIG5V.n2819 ASIG5V.n2500 0.0123125
R53580 ASIG5V.n13247 ASIG5V.n13246 0.0121168
R53581 ASIG5V.n13357 ASIG5V.n13354 0.0120939
R53582 ASIG5V.n11633 ASIG5V.n11632 0.0120939
R53583 ASIG5V.n13356 ASIG5V.n13355 0.0120939
R53584 ASIG5V.n9084 ASIG5V.n9083 0.0120939
R53585 ASIG5V.n2489 ASIG5V.n2488 0.0118684
R53586 ASIG5V.n2187 ASIG5V.n2186 0.0118684
R53587 ASIG5V.n9753 ASIG5V.n9752 0.0117553
R53588 ASIG5V.n1373 ASIG5V.n1372 0.0117553
R53589 ASIG5V.n9761 ASIG5V.n9760 0.0117317
R53590 ASIG5V.n13611 ASIG5V.n13608 0.0117009
R53591 ASIG5V.n11418 ASIG5V.n11417 0.0117009
R53592 ASIG5V.n13610 ASIG5V.n13609 0.0117009
R53593 ASIG5V.n9087 ASIG5V.n9086 0.0117009
R53594 ASIG5V.n1060 ASIG5V.n1059 0.011525
R53595 ASIG5V.n13064 ASIG5V.n13063 0.0113404
R53596 ASIG5V.n13066 ASIG5V.n13065 0.0113404
R53597 ASIG5V.n1987 ASIG5V.n1986 0.0113404
R53598 ASIG5V.n1989 ASIG5V.n1988 0.0113404
R53599 ASIG5V.n10352 ASIG5V.n10351 0.0113404
R53600 ASIG5V.n10354 ASIG5V.n10353 0.0113404
R53601 ASIG5V.n10353 ASIG5V.n10352 0.0113404
R53602 ASIG5V.n13065 ASIG5V.n13064 0.0113404
R53603 ASIG5V.n1988 ASIG5V.n1987 0.0113404
R53604 ASIG5V.n1986 ASIG5V.n1985 0.0113404
R53605 ASIG5V.n13063 ASIG5V.n13062 0.0113404
R53606 ASIG5V.n10351 ASIG5V.n10350 0.0113404
R53607 ASIG5V.n10126 ASIG5V.n10125 0.0113404
R53608 ASIG5V.n10128 ASIG5V.n10127 0.0113404
R53609 ASIG5V.n10127 ASIG5V.n10126 0.0113404
R53610 ASIG5V.n10125 ASIG5V.n10124 0.0113404
R53611 ASIG5V.n3898 ASIG5V.n3897 0.0113079
R53612 ASIG5V.n718 ASIG5V.n717 0.0113079
R53613 ASIG5V.n988 ASIG5V.n987 0.011075
R53614 ASIG5V.n10887 ASIG5V.n10886 0.0109473
R53615 ASIG5V.n2628 ASIG5V.n2627 0.0109473
R53616 ASIG5V.n10883 ASIG5V.n10882 0.0109473
R53617 ASIG5V.n10877 ASIG5V.n10876 0.0109473
R53618 ASIG5V.n10869 ASIG5V.n10868 0.0109473
R53619 ASIG5V.n10861 ASIG5V.n10860 0.0109473
R53620 ASIG5V.n10853 ASIG5V.n10852 0.0109473
R53621 ASIG5V.n10847 ASIG5V.n10846 0.0109473
R53622 ASIG5V.n10837 ASIG5V.n10836 0.0109473
R53623 ASIG5V.n10831 ASIG5V.n10830 0.0109473
R53624 ASIG5V.n10821 ASIG5V.n10820 0.0109473
R53625 ASIG5V.n10815 ASIG5V.n10814 0.0109473
R53626 ASIG5V.n10805 ASIG5V.n10804 0.0109473
R53627 ASIG5V.n10799 ASIG5V.n10798 0.0109473
R53628 ASIG5V.n10789 ASIG5V.n10788 0.0109473
R53629 ASIG5V.n10783 ASIG5V.n10782 0.0109473
R53630 ASIG5V.n10773 ASIG5V.n10772 0.0109473
R53631 ASIG5V.n10767 ASIG5V.n10766 0.0109473
R53632 ASIG5V.n8886 ASIG5V.n8885 0.0109473
R53633 ASIG5V.n8892 ASIG5V.n8891 0.0109473
R53634 ASIG5V.n8902 ASIG5V.n8901 0.0109473
R53635 ASIG5V.n8908 ASIG5V.n8907 0.0109473
R53636 ASIG5V.n8916 ASIG5V.n8915 0.0109473
R53637 ASIG5V.n8924 ASIG5V.n8923 0.0109473
R53638 ASIG5V.n8932 ASIG5V.n8931 0.0109473
R53639 ASIG5V.n2259 ASIG5V.n2258 0.0109072
R53640 ASIG5V.n9764 ASIG5V.n9763 0.0109072
R53641 ASIG5V.n9774 ASIG5V.n9773 0.0109072
R53642 ASIG5V.n9782 ASIG5V.n9781 0.0109072
R53643 ASIG5V.n9807 ASIG5V.n9806 0.0109072
R53644 ASIG5V.n10479 ASIG5V.n10478 0.0108977
R53645 ASIG5V.n10066 ASIG5V.n10065 0.0108977
R53646 ASIG5V.n13216 ASIG5V.n13215 0.0108977
R53647 ASIG5V.n2203 ASIG5V.n2202 0.0108977
R53648 ASIG5V.n2213 ASIG5V.n2212 0.0108977
R53649 ASIG5V.n10295 ASIG5V.n10294 0.0108977
R53650 ASIG5V.n9756 ASIG5V.n9755 0.0108977
R53651 ASIG5V.n9748 ASIG5V.n9747 0.0108977
R53652 ASIG5V.n10099 ASIG5V.n10098 0.0108977
R53653 ASIG5V.n10558 ASIG5V.n10557 0.0108977
R53654 ASIG5V.n10715 ASIG5V.n10714 0.0107857
R53655 ASIG5V.n10718 ASIG5V.n10717 0.0107857
R53656 ASIG5V.n2738 ASIG5V.n2737 0.0106477
R53657 ASIG5V.n9394 ASIG5V.n9393 0.010625
R53658 ASIG5V.n9401 ASIG5V.n9400 0.010625
R53659 ASIG5V.n2738 ASIG5V.n2698 0.0105588
R53660 ASIG5V.n729 ASIG5V.n661 0.0105588
R53661 ASIG5V.n3134 ASIG5V.n3133 0.0105588
R53662 ASIG5V.n2734 ASIG5V.n2730 0.0105588
R53663 ASIG5V.n726 ASIG5V.n673 0.0105588
R53664 ASIG5V.n3329 ASIG5V.n3328 0.0105588
R53665 ASIG5V.n3620 ASIG5V.n3619 0.0105588
R53666 ASIG5V.n722 ASIG5V.n683 0.0105588
R53667 ASIG5V.n3588 ASIG5V.n3587 0.0105588
R53668 ASIG5V.n3894 ASIG5V.n3893 0.0105588
R53669 ASIG5V.n718 ASIG5V.n691 0.0105588
R53670 ASIG5V.n3895 ASIG5V.n3862 0.0105588
R53671 ASIG5V.n4161 ASIG5V.n4160 0.0105588
R53672 ASIG5V.n714 ASIG5V.n697 0.0105588
R53673 ASIG5V.n4129 ASIG5V.n4128 0.0105588
R53674 ASIG5V.n4437 ASIG5V.n4436 0.0105588
R53675 ASIG5V.n710 ASIG5V.n701 0.0105588
R53676 ASIG5V.n4405 ASIG5V.n4404 0.0105588
R53677 ASIG5V.n4695 ASIG5V.n4694 0.0105588
R53678 ASIG5V.n706 ASIG5V.n703 0.0105588
R53679 ASIG5V.n4663 ASIG5V.n4662 0.0105588
R53680 ASIG5V.n4963 ASIG5V.n4962 0.0105588
R53681 ASIG5V.n4931 ASIG5V.n4930 0.0105588
R53682 ASIG5V.n5390 ASIG5V.n5389 0.0105588
R53683 ASIG5V.n5358 ASIG5V.n5357 0.0105588
R53684 ASIG5V.n5621 ASIG5V.n5620 0.0105588
R53685 ASIG5V.n5589 ASIG5V.n5588 0.0105588
R53686 ASIG5V.n5922 ASIG5V.n5921 0.0105588
R53687 ASIG5V.n5890 ASIG5V.n5889 0.0105588
R53688 ASIG5V.n482 ASIG5V.n481 0.0105588
R53689 ASIG5V.n512 ASIG5V.n511 0.0105588
R53690 ASIG5V.n6997 ASIG5V.n6996 0.0105588
R53691 ASIG5V.n6932 ASIG5V.n6931 0.0105588
R53692 ASIG5V.n6965 ASIG5V.n6964 0.0105588
R53693 ASIG5V.n6930 ASIG5V.n6929 0.0105588
R53694 ASIG5V.n6719 ASIG5V.n6718 0.0105588
R53695 ASIG5V.n6687 ASIG5V.n6686 0.0105588
R53696 ASIG5V.n13557 ASIG5V.n13556 0.0105588
R53697 ASIG5V.n13525 ASIG5V.n13524 0.0105588
R53698 ASIG5V.n393 ASIG5V.n392 0.0105588
R53699 ASIG5V.n361 ASIG5V.n360 0.0105588
R53700 ASIG5V.n7468 ASIG5V.n7467 0.0105588
R53701 ASIG5V.n7436 ASIG5V.n7435 0.0105588
R53702 ASIG5V.n7885 ASIG5V.n7884 0.0105588
R53703 ASIG5V.n7853 ASIG5V.n7852 0.0105588
R53704 ASIG5V.n7241 ASIG5V.n7240 0.0105588
R53705 ASIG5V.n7271 ASIG5V.n7270 0.0105588
R53706 ASIG5V.n12643 ASIG5V.n12642 0.0105588
R53707 ASIG5V.n12611 ASIG5V.n12610 0.0105588
R53708 ASIG5V.n12417 ASIG5V.n12416 0.0105588
R53709 ASIG5V.n9064 ASIG5V.n9061 0.0105588
R53710 ASIG5V.n12385 ASIG5V.n12384 0.0105588
R53711 ASIG5V.n12300 ASIG5V.n12299 0.0105588
R53712 ASIG5V.n9068 ASIG5V.n9059 0.0105588
R53713 ASIG5V.n12268 ASIG5V.n12267 0.0105588
R53714 ASIG5V.n12147 ASIG5V.n12146 0.0105588
R53715 ASIG5V.n9072 ASIG5V.n9055 0.0105588
R53716 ASIG5V.n12115 ASIG5V.n12114 0.0105588
R53717 ASIG5V.n11994 ASIG5V.n11993 0.0105588
R53718 ASIG5V.n9075 ASIG5V.n9049 0.0105588
R53719 ASIG5V.n11956 ASIG5V.n11955 0.0105588
R53720 ASIG5V.n11825 ASIG5V.n11824 0.0105588
R53721 ASIG5V.n9079 ASIG5V.n9041 0.0105588
R53722 ASIG5V.n11793 ASIG5V.n11792 0.0105588
R53723 ASIG5V.n10925 ASIG5V.n10922 0.0105588
R53724 ASIG5V.n9083 ASIG5V.n9031 0.0105588
R53725 ASIG5V.n11664 ASIG5V.n11663 0.0105588
R53726 ASIG5V.n11414 ASIG5V.n11413 0.0105588
R53727 ASIG5V.n11187 ASIG5V.n11186 0.0105588
R53728 ASIG5V.n2913 ASIG5V.n2912 0.0105588
R53729 ASIG5V.n2742 ASIG5V.n2665 0.0105588
R53730 ASIG5V.n733 ASIG5V.n646 0.0105588
R53731 ASIG5V.n10981 ASIG5V.n10980 0.0105588
R53732 ASIG5V.n9087 ASIG5V.n9019 0.0105588
R53733 ASIG5V.n11019 ASIG5V.n11018 0.0105588
R53734 ASIG5V.n9107 ASIG5V.n9106 0.0105588
R53735 ASIG5V.n9758 ASIG5V.n9756 0.0105415
R53736 ASIG5V.n2212 ASIG5V.n2211 0.0105415
R53737 ASIG5V.n13217 ASIG5V.n13216 0.0105415
R53738 ASIG5V.n10065 ASIG5V.n10064 0.0105415
R53739 ASIG5V.n10480 ASIG5V.n10479 0.0105415
R53740 ASIG5V.n9750 ASIG5V.n9748 0.0105415
R53741 ASIG5V.n2202 ASIG5V.n2201 0.0105415
R53742 ASIG5V.n10098 ASIG5V.n10097 0.0105415
R53743 ASIG5V.n10557 ASIG5V.n10556 0.0105415
R53744 ASIG5V.n9766 ASIG5V.n9764 0.010532
R53745 ASIG5V.n2258 ASIG5V.n2257 0.010532
R53746 ASIG5V.n8935 ASIG5V.n8934 0.0102808
R53747 ASIG5V.n8929 ASIG5V.n8928 0.0102808
R53748 ASIG5V.n8921 ASIG5V.n8920 0.0102808
R53749 ASIG5V.n8913 ASIG5V.n8912 0.0102808
R53750 ASIG5V.n8905 ASIG5V.n8904 0.0102808
R53751 ASIG5V.n8899 ASIG5V.n8898 0.0102808
R53752 ASIG5V.n8889 ASIG5V.n8888 0.0102808
R53753 ASIG5V.n8883 ASIG5V.n8882 0.0102808
R53754 ASIG5V.n10770 ASIG5V.n10769 0.0102808
R53755 ASIG5V.n10776 ASIG5V.n10775 0.0102808
R53756 ASIG5V.n10786 ASIG5V.n10785 0.0102808
R53757 ASIG5V.n10792 ASIG5V.n10791 0.0102808
R53758 ASIG5V.n10802 ASIG5V.n10801 0.0102808
R53759 ASIG5V.n10808 ASIG5V.n10807 0.0102808
R53760 ASIG5V.n10818 ASIG5V.n10817 0.0102808
R53761 ASIG5V.n10824 ASIG5V.n10823 0.0102808
R53762 ASIG5V.n10834 ASIG5V.n10833 0.0102808
R53763 ASIG5V.n10840 ASIG5V.n10839 0.0102808
R53764 ASIG5V.n10850 ASIG5V.n10849 0.0102808
R53765 ASIG5V.n10856 ASIG5V.n10855 0.0102808
R53766 ASIG5V.n10864 ASIG5V.n10863 0.0102808
R53767 ASIG5V.n10872 ASIG5V.n10871 0.0102808
R53768 ASIG5V.n10880 ASIG5V.n10879 0.0102808
R53769 ASIG5V.n10886 ASIG5V.n10885 0.0102808
R53770 ASIG5V.n576 ASIG5V.n575 0.0102808
R53771 ASIG5V.n10755 ASIG5V.n10754 0.0102444
R53772 ASIG5V.n995 ASIG5V.n994 0.010175
R53773 ASIG5V.n9428 ASIG5V.n9427 0.010175
R53774 ASIG5V.n2882 ASIG5V.n2881 0.0101288
R53775 ASIG5V.n734 ASIG5V.n733 0.0101288
R53776 ASIG5V.n10298 ASIG5V.n10297 0.0098
R53777 ASIG5V.n10299 ASIG5V.n10298 0.0098
R53778 ASIG5V.n10304 ASIG5V.n10303 0.0098
R53779 ASIG5V.n9758 ASIG5V.n9757 0.0098
R53780 ASIG5V.n10307 ASIG5V.n10306 0.0098
R53781 ASIG5V.n10308 ASIG5V.n10307 0.0098
R53782 ASIG5V.n10313 ASIG5V.n10312 0.0098
R53783 ASIG5V.n9766 ASIG5V.n9765 0.0098
R53784 ASIG5V.n1392 ASIG5V.n1391 0.0098
R53785 ASIG5V.n1391 ASIG5V.n1390 0.0098
R53786 ASIG5V.n10295 ASIG5V.n10293 0.0098
R53787 ASIG5V.n9750 ASIG5V.n9749 0.0098
R53788 ASIG5V.n10326 ASIG5V.n10325 0.0098
R53789 ASIG5V.n9772 ASIG5V.n9771 0.0098
R53790 ASIG5V.n9774 ASIG5V.n9772 0.0098
R53791 ASIG5V.n1383 ASIG5V.n1382 0.0098
R53792 ASIG5V.n1382 ASIG5V.n1381 0.0098
R53793 ASIG5V.n9738 ASIG5V.n9737 0.0098
R53794 ASIG5V.n9739 ASIG5V.n9738 0.0098
R53795 ASIG5V.n9742 ASIG5V.n9741 0.0098
R53796 ASIG5V.n1481 ASIG5V.n1475 0.0098
R53797 ASIG5V.n10339 ASIG5V.n10338 0.0098
R53798 ASIG5V.n9780 ASIG5V.n9779 0.0098
R53799 ASIG5V.n9782 ASIG5V.n9780 0.0098
R53800 ASIG5V.n10547 ASIG5V.n10546 0.0098
R53801 ASIG5V.n10548 ASIG5V.n10547 0.0098
R53802 ASIG5V.n10556 ASIG5V.n10555 0.0098
R53803 ASIG5V.n10555 ASIG5V.n10554 0.0098
R53804 ASIG5V.n1431 ASIG5V.n1430 0.0098
R53805 ASIG5V.n1430 ASIG5V.n1429 0.0098
R53806 ASIG5V.n9805 ASIG5V.n9804 0.0098
R53807 ASIG5V.n9807 ASIG5V.n9805 0.0098
R53808 ASIG5V.n5859 ASIG5V.n5856 0.00973581
R53809 ASIG5V.n5858 ASIG5V.n5857 0.00973581
R53810 ASIG5V.n2486 ASIG5V.n2485 0.00970301
R53811 ASIG5V.n2468 ASIG5V.n2467 0.00970301
R53812 ASIG5V.n12650 ASIG5V.n12647 0.00934279
R53813 ASIG5V.n12305 ASIG5V.n12304 0.00934279
R53814 ASIG5V.n12649 ASIG5V.n12648 0.00934279
R53815 ASIG5V.n9068 ASIG5V.n9067 0.00934279
R53816 ASIG5V.n1446 ASIG5V.n1445 0.00929472
R53817 ASIG5V.n11020 ASIG5V.n11019 0.00919799
R53818 ASIG5V.n13604 ASIG5V.n13603 0.00916165
R53819 ASIG5V.n10736 ASIG5V.n10735 0.00916165
R53820 ASIG5V.n1538 ASIG5V.n1537 0.00897723
R53821 ASIG5V.n1508 ASIG5V.n1507 0.00897723
R53822 ASIG5V.n1423 ASIG5V.n1422 0.00897723
R53823 ASIG5V.n5397 ASIG5V.n5394 0.00894978
R53824 ASIG5V.n9432 ASIG5V.n9431 0.00894978
R53825 ASIG5V.n5396 ASIG5V.n5395 0.00894978
R53826 ASIG5V.n9111 ASIG5V.n9110 0.00894978
R53827 ASIG5V.n12960 ASIG5V.n12959 0.00887007
R53828 ASIG5V.n12935 ASIG5V.n12934 0.00887007
R53829 ASIG5V.n12910 ASIG5V.n12909 0.00887007
R53830 ASIG5V.n12881 ASIG5V.n12880 0.00887007
R53831 ASIG5V.n12852 ASIG5V.n12851 0.00887007
R53832 ASIG5V.n12827 ASIG5V.n12826 0.00887007
R53833 ASIG5V.n12798 ASIG5V.n12797 0.00887007
R53834 ASIG5V.n12768 ASIG5V.n12767 0.00887007
R53835 ASIG5V.n12853 ASIG5V.n12852 0.00887007
R53836 ASIG5V.n12882 ASIG5V.n12881 0.00887007
R53837 ASIG5V.n12828 ASIG5V.n12827 0.00887007
R53838 ASIG5V.n13072 ASIG5V.n13071 0.00887007
R53839 ASIG5V.n13099 ASIG5V.n13098 0.00887007
R53840 ASIG5V.n9984 ASIG5V.n9983 0.00887007
R53841 ASIG5V.n10011 ASIG5V.n10010 0.00887007
R53842 ASIG5V.n10039 ASIG5V.n10038 0.00887007
R53843 ASIG5V.n9964 ASIG5V.n9963 0.00887007
R53844 ASIG5V.n13269 ASIG5V.n13268 0.00887007
R53845 ASIG5V.n13298 ASIG5V.n13297 0.00887007
R53846 ASIG5V.n10040 ASIG5V.n10039 0.00887007
R53847 ASIG5V.n10012 ASIG5V.n10011 0.00887007
R53848 ASIG5V.n9963 ASIG5V.n9962 0.00887007
R53849 ASIG5V.n9983 ASIG5V.n9982 0.00887007
R53850 ASIG5V.n12911 ASIG5V.n12910 0.00887007
R53851 ASIG5V.n13021 ASIG5V.n13020 0.00887007
R53852 ASIG5V.n7201 ASIG5V.n7200 0.00887007
R53853 ASIG5V.n13137 ASIG5V.n13136 0.00887007
R53854 ASIG5V.n13168 ASIG5V.n13167 0.00887007
R53855 ASIG5V.n13199 ASIG5V.n13198 0.00887007
R53856 ASIG5V.n13229 ASIG5V.n13228 0.00887007
R53857 ASIG5V.n7164 ASIG5V.n7163 0.00887007
R53858 ASIG5V.n7134 ASIG5V.n7133 0.00887007
R53859 ASIG5V.n13198 ASIG5V.n13197 0.00887007
R53860 ASIG5V.n13167 ASIG5V.n13166 0.00887007
R53861 ASIG5V.n13136 ASIG5V.n13135 0.00887007
R53862 ASIG5V.n13228 ASIG5V.n13227 0.00887007
R53863 ASIG5V.n7165 ASIG5V.n7164 0.00887007
R53864 ASIG5V.n13268 ASIG5V.n13267 0.00887007
R53865 ASIG5V.n12799 ASIG5V.n12798 0.00887007
R53866 ASIG5V.n1995 ASIG5V.n1994 0.00887007
R53867 ASIG5V.n2020 ASIG5V.n2019 0.00887007
R53868 ASIG5V.n2044 ASIG5V.n2043 0.00887007
R53869 ASIG5V.n2069 ASIG5V.n2068 0.00887007
R53870 ASIG5V.n2094 ASIG5V.n2093 0.00887007
R53871 ASIG5V.n2120 ASIG5V.n2119 0.00887007
R53872 ASIG5V.n2144 ASIG5V.n2143 0.00887007
R53873 ASIG5V.n2170 ASIG5V.n2169 0.00887007
R53874 ASIG5V.n2095 ASIG5V.n2094 0.00887007
R53875 ASIG5V.n2070 ASIG5V.n2069 0.00887007
R53876 ASIG5V.n2045 ASIG5V.n2044 0.00887007
R53877 ASIG5V.n2119 ASIG5V.n2118 0.00887007
R53878 ASIG5V.n2145 ASIG5V.n2144 0.00887007
R53879 ASIG5V.n2019 ASIG5V.n2018 0.00887007
R53880 ASIG5V.n7202 ASIG5V.n7201 0.00887007
R53881 ASIG5V.n12936 ASIG5V.n12935 0.00887007
R53882 ASIG5V.n13100 ASIG5V.n13099 0.00887007
R53883 ASIG5V.n1459 ASIG5V.n1458 0.00887007
R53884 ASIG5V.n1491 ASIG5V.n1490 0.00887007
R53885 ASIG5V.n1521 ASIG5V.n1520 0.00887007
R53886 ASIG5V.n1551 ASIG5V.n1550 0.00887007
R53887 ASIG5V.n1581 ASIG5V.n1580 0.00887007
R53888 ASIG5V.n1611 ASIG5V.n1610 0.00887007
R53889 ASIG5V.n1641 ASIG5V.n1640 0.00887007
R53890 ASIG5V.n1671 ASIG5V.n1670 0.00887007
R53891 ASIG5V.n1580 ASIG5V.n1579 0.00887007
R53892 ASIG5V.n1550 ASIG5V.n1549 0.00887007
R53893 ASIG5V.n1520 ASIG5V.n1519 0.00887007
R53894 ASIG5V.n1490 ASIG5V.n1489 0.00887007
R53895 ASIG5V.n1610 ASIG5V.n1609 0.00887007
R53896 ASIG5V.n1640 ASIG5V.n1639 0.00887007
R53897 ASIG5V.n12769 ASIG5V.n12768 0.00887007
R53898 ASIG5V.n13297 ASIG5V.n13296 0.00887007
R53899 ASIG5V.n1670 ASIG5V.n1669 0.00887007
R53900 ASIG5V.n2169 ASIG5V.n2168 0.00887007
R53901 ASIG5V.n7135 ASIG5V.n7134 0.00887007
R53902 ASIG5V.n10360 ASIG5V.n10359 0.00887007
R53903 ASIG5V.n10384 ASIG5V.n10383 0.00887007
R53904 ASIG5V.n10409 ASIG5V.n10408 0.00887007
R53905 ASIG5V.n10434 ASIG5V.n10433 0.00887007
R53906 ASIG5V.n10459 ASIG5V.n10458 0.00887007
R53907 ASIG5V.n10494 ASIG5V.n10493 0.00887007
R53908 ASIG5V.n10525 ASIG5V.n10524 0.00887007
R53909 ASIG5V.n10568 ASIG5V.n10567 0.00887007
R53910 ASIG5V.n10460 ASIG5V.n10459 0.00887007
R53911 ASIG5V.n10435 ASIG5V.n10434 0.00887007
R53912 ASIG5V.n10410 ASIG5V.n10409 0.00887007
R53913 ASIG5V.n10385 ASIG5V.n10384 0.00887007
R53914 ASIG5V.n10493 ASIG5V.n10492 0.00887007
R53915 ASIG5V.n10524 ASIG5V.n10523 0.00887007
R53916 ASIG5V.n10567 ASIG5V.n10566 0.00887007
R53917 ASIG5V.n13020 ASIG5V.n13019 0.00887007
R53918 ASIG5V.n13071 ASIG5V.n13070 0.00887007
R53919 ASIG5V.n12961 ASIG5V.n12960 0.00887007
R53920 ASIG5V.n10359 ASIG5V.n10358 0.00887007
R53921 ASIG5V.n1994 ASIG5V.n1993 0.00887007
R53922 ASIG5V.n1458 ASIG5V.n1457 0.00887007
R53923 ASIG5V.n9819 ASIG5V.n9818 0.00887007
R53924 ASIG5V.n9847 ASIG5V.n9846 0.00887007
R53925 ASIG5V.n9875 ASIG5V.n9874 0.00887007
R53926 ASIG5V.n9903 ASIG5V.n9902 0.00887007
R53927 ASIG5V.n9931 ASIG5V.n9930 0.00887007
R53928 ASIG5V.n10079 ASIG5V.n10078 0.00887007
R53929 ASIG5V.n10109 ASIG5V.n10108 0.00887007
R53930 ASIG5V.n10134 ASIG5V.n10133 0.00887007
R53931 ASIG5V.n9820 ASIG5V.n9819 0.00887007
R53932 ASIG5V.n9932 ASIG5V.n9931 0.00887007
R53933 ASIG5V.n9904 ASIG5V.n9903 0.00887007
R53934 ASIG5V.n9876 ASIG5V.n9875 0.00887007
R53935 ASIG5V.n9848 ASIG5V.n9847 0.00887007
R53936 ASIG5V.n10078 ASIG5V.n10077 0.00887007
R53937 ASIG5V.n10108 ASIG5V.n10107 0.00887007
R53938 ASIG5V.n10133 ASIG5V.n10132 0.00887007
R53939 ASIG5V.n2284 ASIG5V.n2283 0.00887007
R53940 ASIG5V.n2310 ASIG5V.n2309 0.00887007
R53941 ASIG5V.n2335 ASIG5V.n2334 0.00887007
R53942 ASIG5V.n2360 ASIG5V.n2359 0.00887007
R53943 ASIG5V.n2385 ASIG5V.n2384 0.00887007
R53944 ASIG5V.n2410 ASIG5V.n2409 0.00887007
R53945 ASIG5V.n2435 ASIG5V.n2434 0.00887007
R53946 ASIG5V.n2460 ASIG5V.n2459 0.00887007
R53947 ASIG5V.n2384 ASIG5V.n2383 0.00887007
R53948 ASIG5V.n2359 ASIG5V.n2358 0.00887007
R53949 ASIG5V.n2334 ASIG5V.n2333 0.00887007
R53950 ASIG5V.n2309 ASIG5V.n2308 0.00887007
R53951 ASIG5V.n2409 ASIG5V.n2408 0.00887007
R53952 ASIG5V.n2434 ASIG5V.n2433 0.00887007
R53953 ASIG5V.n2283 ASIG5V.n2282 0.00887007
R53954 ASIG5V.n2459 ASIG5V.n2458 0.00887007
R53955 ASIG5V.n12972 ASIG5V.n12971 0.0087818
R53956 ASIG5V.n12949 ASIG5V.n12948 0.0087818
R53957 ASIG5V.n12924 ASIG5V.n12923 0.0087818
R53958 ASIG5V.n12841 ASIG5V.n12840 0.0087818
R53959 ASIG5V.n12816 ASIG5V.n12815 0.0087818
R53960 ASIG5V.n12787 ASIG5V.n12786 0.0087818
R53961 ASIG5V.n12842 ASIG5V.n12841 0.0087818
R53962 ASIG5V.n13058 ASIG5V.n13057 0.0087818
R53963 ASIG5V.n13083 ASIG5V.n13082 0.0087818
R53964 ASIG5V.n13111 ASIG5V.n13110 0.0087818
R53965 ASIG5V.n9995 ASIG5V.n9994 0.0087818
R53966 ASIG5V.n10023 ASIG5V.n10022 0.0087818
R53967 ASIG5V.n9952 ASIG5V.n9951 0.0087818
R53968 ASIG5V.n13280 ASIG5V.n13279 0.0087818
R53969 ASIG5V.n10022 ASIG5V.n10021 0.0087818
R53970 ASIG5V.n9994 ASIG5V.n9993 0.0087818
R53971 ASIG5V.n13110 ASIG5V.n13109 0.0087818
R53972 ASIG5V.n12925 ASIG5V.n12924 0.0087818
R53973 ASIG5V.n13005 ASIG5V.n13004 0.0087818
R53974 ASIG5V.n13032 ASIG5V.n13031 0.0087818
R53975 ASIG5V.n13148 ASIG5V.n13147 0.0087818
R53976 ASIG5V.n13179 ASIG5V.n13178 0.0087818
R53977 ASIG5V.n13210 ASIG5V.n13209 0.0087818
R53978 ASIG5V.n13240 ASIG5V.n13239 0.0087818
R53979 ASIG5V.n7153 ASIG5V.n7152 0.0087818
R53980 ASIG5V.n13178 ASIG5V.n13177 0.0087818
R53981 ASIG5V.n13147 ASIG5V.n13146 0.0087818
R53982 ASIG5V.n13209 ASIG5V.n13208 0.0087818
R53983 ASIG5V.n13239 ASIG5V.n13238 0.0087818
R53984 ASIG5V.n9953 ASIG5V.n9952 0.0087818
R53985 ASIG5V.n12817 ASIG5V.n12816 0.0087818
R53986 ASIG5V.n1981 ASIG5V.n1980 0.0087818
R53987 ASIG5V.n2006 ASIG5V.n2005 0.0087818
R53988 ASIG5V.n2031 ASIG5V.n2030 0.0087818
R53989 ASIG5V.n2056 ASIG5V.n2055 0.0087818
R53990 ASIG5V.n2081 ASIG5V.n2080 0.0087818
R53991 ASIG5V.n2106 ASIG5V.n2105 0.0087818
R53992 ASIG5V.n2156 ASIG5V.n2155 0.0087818
R53993 ASIG5V.n2080 ASIG5V.n2079 0.0087818
R53994 ASIG5V.n2055 ASIG5V.n2054 0.0087818
R53995 ASIG5V.n2030 ASIG5V.n2029 0.0087818
R53996 ASIG5V.n2105 ASIG5V.n2104 0.0087818
R53997 ASIG5V.n2005 ASIG5V.n2004 0.0087818
R53998 ASIG5V.n13031 ASIG5V.n13030 0.0087818
R53999 ASIG5V.n13082 ASIG5V.n13081 0.0087818
R54000 ASIG5V.n12950 ASIG5V.n12949 0.0087818
R54001 ASIG5V.n1440 ASIG5V.n1439 0.0087818
R54002 ASIG5V.n1502 ASIG5V.n1501 0.0087818
R54003 ASIG5V.n1532 ASIG5V.n1531 0.0087818
R54004 ASIG5V.n1562 ASIG5V.n1561 0.0087818
R54005 ASIG5V.n1592 ASIG5V.n1591 0.0087818
R54006 ASIG5V.n1622 ASIG5V.n1621 0.0087818
R54007 ASIG5V.n1652 ASIG5V.n1651 0.0087818
R54008 ASIG5V.n1561 ASIG5V.n1560 0.0087818
R54009 ASIG5V.n1531 ASIG5V.n1530 0.0087818
R54010 ASIG5V.n1501 ASIG5V.n1500 0.0087818
R54011 ASIG5V.n1591 ASIG5V.n1590 0.0087818
R54012 ASIG5V.n1621 ASIG5V.n1620 0.0087818
R54013 ASIG5V.n1651 ASIG5V.n1650 0.0087818
R54014 ASIG5V.n2155 ASIG5V.n2154 0.0087818
R54015 ASIG5V.n7154 ASIG5V.n7153 0.0087818
R54016 ASIG5V.n13279 ASIG5V.n13278 0.0087818
R54017 ASIG5V.n12788 ASIG5V.n12787 0.0087818
R54018 ASIG5V.n10346 ASIG5V.n10345 0.0087818
R54019 ASIG5V.n10371 ASIG5V.n10370 0.0087818
R54020 ASIG5V.n10396 ASIG5V.n10395 0.0087818
R54021 ASIG5V.n10421 ASIG5V.n10420 0.0087818
R54022 ASIG5V.n10446 ASIG5V.n10445 0.0087818
R54023 ASIG5V.n10471 ASIG5V.n10470 0.0087818
R54024 ASIG5V.n10505 ASIG5V.n10504 0.0087818
R54025 ASIG5V.n10445 ASIG5V.n10444 0.0087818
R54026 ASIG5V.n10420 ASIG5V.n10419 0.0087818
R54027 ASIG5V.n10395 ASIG5V.n10394 0.0087818
R54028 ASIG5V.n10370 ASIG5V.n10369 0.0087818
R54029 ASIG5V.n10470 ASIG5V.n10469 0.0087818
R54030 ASIG5V.n10504 ASIG5V.n10503 0.0087818
R54031 ASIG5V.n1439 ASIG5V.n1438 0.0087818
R54032 ASIG5V.n1980 ASIG5V.n1979 0.0087818
R54033 ASIG5V.n13004 ASIG5V.n13003 0.0087818
R54034 ASIG5V.n13057 ASIG5V.n13056 0.0087818
R54035 ASIG5V.n12971 ASIG5V.n12970 0.0087818
R54036 ASIG5V.n10345 ASIG5V.n10344 0.0087818
R54037 ASIG5V.n9831 ASIG5V.n9830 0.0087818
R54038 ASIG5V.n9859 ASIG5V.n9858 0.0087818
R54039 ASIG5V.n9887 ASIG5V.n9886 0.0087818
R54040 ASIG5V.n9915 ASIG5V.n9914 0.0087818
R54041 ASIG5V.n9943 ASIG5V.n9942 0.0087818
R54042 ASIG5V.n10090 ASIG5V.n10089 0.0087818
R54043 ASIG5V.n10120 ASIG5V.n10119 0.0087818
R54044 ASIG5V.n10119 ASIG5V.n10118 0.0087818
R54045 ASIG5V.n10089 ASIG5V.n10088 0.0087818
R54046 ASIG5V.n9942 ASIG5V.n9941 0.0087818
R54047 ASIG5V.n9914 ASIG5V.n9913 0.0087818
R54048 ASIG5V.n9886 ASIG5V.n9885 0.0087818
R54049 ASIG5V.n9858 ASIG5V.n9857 0.0087818
R54050 ASIG5V.n9830 ASIG5V.n9829 0.0087818
R54051 ASIG5V.n2270 ASIG5V.n2269 0.0087818
R54052 ASIG5V.n2295 ASIG5V.n2294 0.0087818
R54053 ASIG5V.n2321 ASIG5V.n2320 0.0087818
R54054 ASIG5V.n2346 ASIG5V.n2345 0.0087818
R54055 ASIG5V.n2371 ASIG5V.n2370 0.0087818
R54056 ASIG5V.n2396 ASIG5V.n2395 0.0087818
R54057 ASIG5V.n2421 ASIG5V.n2420 0.0087818
R54058 ASIG5V.n2446 ASIG5V.n2445 0.0087818
R54059 ASIG5V.n2370 ASIG5V.n2369 0.0087818
R54060 ASIG5V.n2345 ASIG5V.n2344 0.0087818
R54061 ASIG5V.n2320 ASIG5V.n2319 0.0087818
R54062 ASIG5V.n2294 ASIG5V.n2293 0.0087818
R54063 ASIG5V.n2395 ASIG5V.n2394 0.0087818
R54064 ASIG5V.n2420 ASIG5V.n2419 0.0087818
R54065 ASIG5V.n2445 ASIG5V.n2444 0.0087818
R54066 ASIG5V.n2269 ASIG5V.n2268 0.0087818
R54067 ASIG5V.n12900 ASIG5V.n12899 0.0087818
R54068 ASIG5V.n12871 ASIG5V.n12870 0.0087818
R54069 ASIG5V.n12870 ASIG5V.n12869 0.0087818
R54070 ASIG5V.n12899 ASIG5V.n12898 0.0087818
R54071 ASIG5V.n10050 ASIG5V.n10049 0.0087818
R54072 ASIG5V.n10051 ASIG5V.n10050 0.0087818
R54073 ASIG5V.n7191 ASIG5V.n7190 0.0087818
R54074 ASIG5V.n7190 ASIG5V.n7189 0.0087818
R54075 ASIG5V.n2130 ASIG5V.n2129 0.0087818
R54076 ASIG5V.n2131 ASIG5V.n2130 0.0087818
R54077 ASIG5V.n1469 ASIG5V.n1468 0.0087818
R54078 ASIG5V.n1470 ASIG5V.n1469 0.0087818
R54079 ASIG5V.n10536 ASIG5V.n10535 0.0087818
R54080 ASIG5V.n10535 ASIG5V.n10534 0.0087818
R54081 ASIG5V.n9789 ASIG5V.n9788 0.0087818
R54082 ASIG5V.n9788 ASIG5V.n9787 0.0087818
R54083 ASIG5V.n1568 ASIG5V.n1567 0.00875907
R54084 ASIG5V.n1598 ASIG5V.n1597 0.00875907
R54085 ASIG5V.n1628 ASIG5V.n1627 0.00875907
R54086 ASIG5V.n1658 ASIG5V.n1657 0.00875907
R54087 ASIG5V.n2735 ASIG5V.n2734 0.00871477
R54088 ASIG5V.n738 ASIG5V.n737 0.0087125
R54089 ASIG5V.n9113 ASIG5V.n9111 0.0087125
R54090 ASIG5V.n10737 ASIG5V.n10736 0.0086203
R54091 ASIG5V.n521 ASIG5V.n517 0.00857847
R54092 ASIG5V.n8986 ASIG5V.n8985 0.00857847
R54093 ASIG5V.n2631 ASIG5V.n2630 0.00857847
R54094 ASIG5V.n10761 ASIG5V.n9435 0.00857847
R54095 ASIG5V.n11095 ASIG5V.n10890 0.00857847
R54096 ASIG5V.n2500 ASIG5V.n1070 0.00857847
R54097 ASIG5V.n8874 ASIG5V.n8870 0.00857847
R54098 ASIG5V.n620 ASIG5V.n616 0.00857847
R54099 ASIG5V.n9893 ASIG5V.n9892 0.0085739
R54100 ASIG5V.n1007 ASIG5V.n1006 0.008375
R54101 ASIG5V.n9921 ASIG5V.n9920 0.00836718
R54102 ASIG5V.n10068 ASIG5V.n10067 0.00836718
R54103 ASIG5V.n10553 ASIG5V.n10552 0.00836718
R54104 ASIG5V.n10890 ASIG5V.n10889 0.00832684
R54105 ASIG5V.n8980 ASIG5V.n8979 0.00832684
R54106 ASIG5V.n626 ASIG5V.n625 0.00832684
R54107 ASIG5V.n521 ASIG5V.n520 0.00832684
R54108 ASIG5V.n1070 ASIG5V.n1069 0.00832684
R54109 ASIG5V.n2818 ASIG5V.n2631 0.00832684
R54110 ASIG5V.n9435 ASIG5V.n9434 0.00832684
R54111 ASIG5V.n8874 ASIG5V.n8873 0.00832684
R54112 ASIG5V.n8974 ASIG5V.n8973 0.00832684
R54113 ASIG5V.n620 ASIG5V.n619 0.00832684
R54114 ASIG5V.n8878 ASIG5V.n8877 0.00832684
R54115 ASIG5V.n9115 ASIG5V.n9114 0.00832684
R54116 ASIG5V.n740 ASIG5V.n739 0.00832684
R54117 ASIG5V.n13606 ASIG5V.n13525 0.00823154
R54118 ASIG5V.n13605 ASIG5V.n13557 0.00823154
R54119 ASIG5V.n11995 ASIG5V.n11994 0.00823154
R54120 ASIG5V.n12835 ASIG5V.n12834 0.00822031
R54121 ASIG5V.n12892 ASIG5V.n12891 0.00822031
R54122 ASIG5V.n12863 ASIG5V.n12862 0.00822031
R54123 ASIG5V.n10062 ASIG5V.n10061 0.00822031
R54124 ASIG5V.n10033 ASIG5V.n10032 0.00822031
R54125 ASIG5V.n10005 ASIG5V.n10004 0.00822031
R54126 ASIG5V.n13121 ASIG5V.n13120 0.00822031
R54127 ASIG5V.n12917 ASIG5V.n12916 0.00822031
R54128 ASIG5V.n13221 ASIG5V.n13220 0.00822031
R54129 ASIG5V.n13130 ASIG5V.n13129 0.00822031
R54130 ASIG5V.n13161 ASIG5V.n13160 0.00822031
R54131 ASIG5V.n13192 ASIG5V.n13191 0.00822031
R54132 ASIG5V.n13252 ASIG5V.n13251 0.00822031
R54133 ASIG5V.n13262 ASIG5V.n13261 0.00822031
R54134 ASIG5V.n12809 ASIG5V.n12808 0.00822031
R54135 ASIG5V.n2112 ASIG5V.n2111 0.00822031
R54136 ASIG5V.n2088 ASIG5V.n2087 0.00822031
R54137 ASIG5V.n2063 ASIG5V.n2062 0.00822031
R54138 ASIG5V.n2038 ASIG5V.n2037 0.00822031
R54139 ASIG5V.n2013 ASIG5V.n2012 0.00822031
R54140 ASIG5V.n13045 ASIG5V.n13044 0.00822031
R54141 ASIG5V.n13093 ASIG5V.n13092 0.00822031
R54142 ASIG5V.n12942 ASIG5V.n12941 0.00822031
R54143 ASIG5V.n1603 ASIG5V.n1602 0.00822031
R54144 ASIG5V.n1484 ASIG5V.n1483 0.00822031
R54145 ASIG5V.n1514 ASIG5V.n1513 0.00822031
R54146 ASIG5V.n1544 ASIG5V.n1543 0.00822031
R54147 ASIG5V.n1574 ASIG5V.n1573 0.00822031
R54148 ASIG5V.n1634 ASIG5V.n1633 0.00822031
R54149 ASIG5V.n1664 ASIG5V.n1663 0.00822031
R54150 ASIG5V.n2163 ASIG5V.n2162 0.00822031
R54151 ASIG5V.n7146 ASIG5V.n7145 0.00822031
R54152 ASIG5V.n12780 ASIG5V.n12779 0.00822031
R54153 ASIG5V.n10486 ASIG5V.n10485 0.00822031
R54154 ASIG5V.n10517 ASIG5V.n10516 0.00822031
R54155 ASIG5V.n10453 ASIG5V.n10452 0.00822031
R54156 ASIG5V.n10428 ASIG5V.n10427 0.00822031
R54157 ASIG5V.n10403 ASIG5V.n10402 0.00822031
R54158 ASIG5V.n10378 ASIG5V.n10377 0.00822031
R54159 ASIG5V.n10487 ASIG5V.n10486 0.00822031
R54160 ASIG5V.n1452 ASIG5V.n1451 0.00822031
R54161 ASIG5V.n12981 ASIG5V.n12980 0.00822031
R54162 ASIG5V.n13014 ASIG5V.n13013 0.00822031
R54163 ASIG5V.n10071 ASIG5V.n10070 0.00822031
R54164 ASIG5V.n10101 ASIG5V.n10100 0.00822031
R54165 ASIG5V.n9925 ASIG5V.n9924 0.00822031
R54166 ASIG5V.n9897 ASIG5V.n9896 0.00822031
R54167 ASIG5V.n9869 ASIG5V.n9868 0.00822031
R54168 ASIG5V.n9841 ASIG5V.n9840 0.00822031
R54169 ASIG5V.n2402 ASIG5V.n2401 0.00822031
R54170 ASIG5V.n2303 ASIG5V.n2302 0.00822031
R54171 ASIG5V.n2328 ASIG5V.n2327 0.00822031
R54172 ASIG5V.n2353 ASIG5V.n2352 0.00822031
R54173 ASIG5V.n2378 ASIG5V.n2377 0.00822031
R54174 ASIG5V.n2428 ASIG5V.n2427 0.00822031
R54175 ASIG5V.n2453 ASIG5V.n2452 0.00822031
R54176 ASIG5V.n2277 ASIG5V.n2276 0.00822031
R54177 ASIG5V.n2485 ASIG5V.n2484 0.00807895
R54178 ASIG5V.n2469 ASIG5V.n2468 0.00807895
R54179 ASIG5V.n10881 ASIG5V.n10880 0.00796421
R54180 ASIG5V.n10875 ASIG5V.n10874 0.00796421
R54181 ASIG5V.n10873 ASIG5V.n10872 0.00796421
R54182 ASIG5V.n10867 ASIG5V.n10866 0.00796421
R54183 ASIG5V.n10865 ASIG5V.n10864 0.00796421
R54184 ASIG5V.n10859 ASIG5V.n10858 0.00796421
R54185 ASIG5V.n10857 ASIG5V.n10856 0.00796421
R54186 ASIG5V.n10851 ASIG5V.n10850 0.00796421
R54187 ASIG5V.n10845 ASIG5V.n10844 0.00796421
R54188 ASIG5V.n10843 ASIG5V.n10842 0.00796421
R54189 ASIG5V.n10841 ASIG5V.n10840 0.00796421
R54190 ASIG5V.n10835 ASIG5V.n10834 0.00796421
R54191 ASIG5V.n10829 ASIG5V.n10828 0.00796421
R54192 ASIG5V.n10827 ASIG5V.n10826 0.00796421
R54193 ASIG5V.n10825 ASIG5V.n10824 0.00796421
R54194 ASIG5V.n10819 ASIG5V.n10818 0.00796421
R54195 ASIG5V.n10813 ASIG5V.n10812 0.00796421
R54196 ASIG5V.n10811 ASIG5V.n10810 0.00796421
R54197 ASIG5V.n10809 ASIG5V.n10808 0.00796421
R54198 ASIG5V.n10803 ASIG5V.n10802 0.00796421
R54199 ASIG5V.n10797 ASIG5V.n10796 0.00796421
R54200 ASIG5V.n10795 ASIG5V.n10794 0.00796421
R54201 ASIG5V.n10793 ASIG5V.n10792 0.00796421
R54202 ASIG5V.n10787 ASIG5V.n10786 0.00796421
R54203 ASIG5V.n10781 ASIG5V.n10780 0.00796421
R54204 ASIG5V.n10779 ASIG5V.n10778 0.00796421
R54205 ASIG5V.n10777 ASIG5V.n10776 0.00796421
R54206 ASIG5V.n10771 ASIG5V.n10770 0.00796421
R54207 ASIG5V.n10765 ASIG5V.n10764 0.00796421
R54208 ASIG5V.n10763 ASIG5V.n10762 0.00796421
R54209 ASIG5V.n8882 ASIG5V.n8881 0.00796421
R54210 ASIG5V.n8888 ASIG5V.n8887 0.00796421
R54211 ASIG5V.n8894 ASIG5V.n8893 0.00796421
R54212 ASIG5V.n8896 ASIG5V.n8895 0.00796421
R54213 ASIG5V.n8898 ASIG5V.n8897 0.00796421
R54214 ASIG5V.n8904 ASIG5V.n8903 0.00796421
R54215 ASIG5V.n8910 ASIG5V.n8909 0.00796421
R54216 ASIG5V.n8912 ASIG5V.n8911 0.00796421
R54217 ASIG5V.n8918 ASIG5V.n8917 0.00796421
R54218 ASIG5V.n8920 ASIG5V.n8919 0.00796421
R54219 ASIG5V.n8926 ASIG5V.n8925 0.00796421
R54220 ASIG5V.n8928 ASIG5V.n8927 0.00796421
R54221 ASIG5V.n8934 ASIG5V.n8933 0.00796421
R54222 ASIG5V.n2626 ASIG5V.n2625 0.00796421
R54223 ASIG5V.n2624 ASIG5V.n2623 0.00796421
R54224 ASIG5V.n2622 ASIG5V.n2621 0.00796421
R54225 ASIG5V.n2620 ASIG5V.n2619 0.00796421
R54226 ASIG5V.n2618 ASIG5V.n2617 0.00796421
R54227 ASIG5V.n2616 ASIG5V.n2615 0.00796421
R54228 ASIG5V.n2614 ASIG5V.n2613 0.00796421
R54229 ASIG5V.n2612 ASIG5V.n2611 0.00796421
R54230 ASIG5V.n2610 ASIG5V.n2609 0.00796421
R54231 ASIG5V.n2608 ASIG5V.n2607 0.00796421
R54232 ASIG5V.n2606 ASIG5V.n2605 0.00796421
R54233 ASIG5V.n2604 ASIG5V.n2603 0.00796421
R54234 ASIG5V.n2602 ASIG5V.n2601 0.00796421
R54235 ASIG5V.n2600 ASIG5V.n2599 0.00796421
R54236 ASIG5V.n2598 ASIG5V.n2597 0.00796421
R54237 ASIG5V.n2596 ASIG5V.n2595 0.00796421
R54238 ASIG5V.n2594 ASIG5V.n2593 0.00796421
R54239 ASIG5V.n2592 ASIG5V.n2591 0.00796421
R54240 ASIG5V.n2590 ASIG5V.n2589 0.00796421
R54241 ASIG5V.n2588 ASIG5V.n2587 0.00796421
R54242 ASIG5V.n2586 ASIG5V.n2585 0.00796421
R54243 ASIG5V.n2584 ASIG5V.n2583 0.00796421
R54244 ASIG5V.n2582 ASIG5V.n2581 0.00796421
R54245 ASIG5V.n2580 ASIG5V.n2579 0.00796421
R54246 ASIG5V.n2578 ASIG5V.n2577 0.00796421
R54247 ASIG5V.n2576 ASIG5V.n2575 0.00796421
R54248 ASIG5V.n2574 ASIG5V.n2573 0.00796421
R54249 ASIG5V.n2572 ASIG5V.n2571 0.00796421
R54250 ASIG5V.n2570 ASIG5V.n2569 0.00796421
R54251 ASIG5V.n2568 ASIG5V.n2567 0.00796421
R54252 ASIG5V.n2566 ASIG5V.n2565 0.00796421
R54253 ASIG5V.n2564 ASIG5V.n2563 0.00796421
R54254 ASIG5V.n2562 ASIG5V.n2561 0.00796421
R54255 ASIG5V.n2560 ASIG5V.n2559 0.00796421
R54256 ASIG5V.n2558 ASIG5V.n2557 0.00796421
R54257 ASIG5V.n2556 ASIG5V.n2555 0.00796421
R54258 ASIG5V.n2554 ASIG5V.n2553 0.00796421
R54259 ASIG5V.n2552 ASIG5V.n2551 0.00796421
R54260 ASIG5V.n2550 ASIG5V.n2549 0.00796421
R54261 ASIG5V.n2548 ASIG5V.n2547 0.00796421
R54262 ASIG5V.n2546 ASIG5V.n2545 0.00796421
R54263 ASIG5V.n2544 ASIG5V.n2543 0.00796421
R54264 ASIG5V.n2542 ASIG5V.n2541 0.00796421
R54265 ASIG5V.n2540 ASIG5V.n2539 0.00796421
R54266 ASIG5V.n2538 ASIG5V.n2537 0.00796421
R54267 ASIG5V.n2536 ASIG5V.n2535 0.00796421
R54268 ASIG5V.n2534 ASIG5V.n2533 0.00796421
R54269 ASIG5V.n2532 ASIG5V.n2531 0.00796421
R54270 ASIG5V.n2530 ASIG5V.n2529 0.00796421
R54271 ASIG5V.n2528 ASIG5V.n2527 0.00796421
R54272 ASIG5V.n2526 ASIG5V.n2525 0.00796421
R54273 ASIG5V.n2524 ASIG5V.n2523 0.00796421
R54274 ASIG5V.n2522 ASIG5V.n2521 0.00796421
R54275 ASIG5V.n2520 ASIG5V.n2519 0.00796421
R54276 ASIG5V.n2518 ASIG5V.n2517 0.00796421
R54277 ASIG5V.n2516 ASIG5V.n2515 0.00796421
R54278 ASIG5V.n2514 ASIG5V.n2513 0.00796421
R54279 ASIG5V.n2512 ASIG5V.n2511 0.00796421
R54280 ASIG5V.n2510 ASIG5V.n2509 0.00796421
R54281 ASIG5V.n2508 ASIG5V.n2507 0.00796421
R54282 ASIG5V.n2506 ASIG5V.n2505 0.00796421
R54283 ASIG5V.n2504 ASIG5V.n2503 0.00796421
R54284 ASIG5V.n2502 ASIG5V.n2501 0.00796421
R54285 ASIG5V.n523 ASIG5V.n522 0.00796421
R54286 ASIG5V.n525 ASIG5V.n524 0.00796421
R54287 ASIG5V.n527 ASIG5V.n526 0.00796421
R54288 ASIG5V.n529 ASIG5V.n528 0.00796421
R54289 ASIG5V.n531 ASIG5V.n530 0.00796421
R54290 ASIG5V.n533 ASIG5V.n532 0.00796421
R54291 ASIG5V.n535 ASIG5V.n534 0.00796421
R54292 ASIG5V.n537 ASIG5V.n536 0.00796421
R54293 ASIG5V.n539 ASIG5V.n538 0.00796421
R54294 ASIG5V.n541 ASIG5V.n540 0.00796421
R54295 ASIG5V.n543 ASIG5V.n542 0.00796421
R54296 ASIG5V.n545 ASIG5V.n544 0.00796421
R54297 ASIG5V.n547 ASIG5V.n546 0.00796421
R54298 ASIG5V.n549 ASIG5V.n548 0.00796421
R54299 ASIG5V.n551 ASIG5V.n550 0.00796421
R54300 ASIG5V.n553 ASIG5V.n552 0.00796421
R54301 ASIG5V.n555 ASIG5V.n554 0.00796421
R54302 ASIG5V.n557 ASIG5V.n556 0.00796421
R54303 ASIG5V.n559 ASIG5V.n558 0.00796421
R54304 ASIG5V.n561 ASIG5V.n560 0.00796421
R54305 ASIG5V.n563 ASIG5V.n562 0.00796421
R54306 ASIG5V.n565 ASIG5V.n564 0.00796421
R54307 ASIG5V.n567 ASIG5V.n566 0.00796421
R54308 ASIG5V.n569 ASIG5V.n568 0.00796421
R54309 ASIG5V.n571 ASIG5V.n570 0.00796421
R54310 ASIG5V.n573 ASIG5V.n572 0.00796421
R54311 ASIG5V.n575 ASIG5V.n574 0.00796421
R54312 ASIG5V.n8933 ASIG5V.n8932 0.00796421
R54313 ASIG5V.n8927 ASIG5V.n8926 0.00796421
R54314 ASIG5V.n8925 ASIG5V.n8924 0.00796421
R54315 ASIG5V.n8919 ASIG5V.n8918 0.00796421
R54316 ASIG5V.n8917 ASIG5V.n8916 0.00796421
R54317 ASIG5V.n8911 ASIG5V.n8910 0.00796421
R54318 ASIG5V.n8909 ASIG5V.n8908 0.00796421
R54319 ASIG5V.n8903 ASIG5V.n8902 0.00796421
R54320 ASIG5V.n8897 ASIG5V.n8896 0.00796421
R54321 ASIG5V.n8895 ASIG5V.n8894 0.00796421
R54322 ASIG5V.n8893 ASIG5V.n8892 0.00796421
R54323 ASIG5V.n8887 ASIG5V.n8886 0.00796421
R54324 ASIG5V.n10764 ASIG5V.n10763 0.00796421
R54325 ASIG5V.n10766 ASIG5V.n10765 0.00796421
R54326 ASIG5V.n10772 ASIG5V.n10771 0.00796421
R54327 ASIG5V.n10778 ASIG5V.n10777 0.00796421
R54328 ASIG5V.n10780 ASIG5V.n10779 0.00796421
R54329 ASIG5V.n10782 ASIG5V.n10781 0.00796421
R54330 ASIG5V.n10788 ASIG5V.n10787 0.00796421
R54331 ASIG5V.n10794 ASIG5V.n10793 0.00796421
R54332 ASIG5V.n10796 ASIG5V.n10795 0.00796421
R54333 ASIG5V.n10798 ASIG5V.n10797 0.00796421
R54334 ASIG5V.n10804 ASIG5V.n10803 0.00796421
R54335 ASIG5V.n10810 ASIG5V.n10809 0.00796421
R54336 ASIG5V.n10812 ASIG5V.n10811 0.00796421
R54337 ASIG5V.n10814 ASIG5V.n10813 0.00796421
R54338 ASIG5V.n10820 ASIG5V.n10819 0.00796421
R54339 ASIG5V.n10826 ASIG5V.n10825 0.00796421
R54340 ASIG5V.n10828 ASIG5V.n10827 0.00796421
R54341 ASIG5V.n10830 ASIG5V.n10829 0.00796421
R54342 ASIG5V.n10836 ASIG5V.n10835 0.00796421
R54343 ASIG5V.n10842 ASIG5V.n10841 0.00796421
R54344 ASIG5V.n10844 ASIG5V.n10843 0.00796421
R54345 ASIG5V.n10846 ASIG5V.n10845 0.00796421
R54346 ASIG5V.n10852 ASIG5V.n10851 0.00796421
R54347 ASIG5V.n10858 ASIG5V.n10857 0.00796421
R54348 ASIG5V.n10860 ASIG5V.n10859 0.00796421
R54349 ASIG5V.n10866 ASIG5V.n10865 0.00796421
R54350 ASIG5V.n10868 ASIG5V.n10867 0.00796421
R54351 ASIG5V.n10874 ASIG5V.n10873 0.00796421
R54352 ASIG5V.n10876 ASIG5V.n10875 0.00796421
R54353 ASIG5V.n10882 ASIG5V.n10881 0.00796421
R54354 ASIG5V.n574 ASIG5V.n573 0.00796421
R54355 ASIG5V.n572 ASIG5V.n571 0.00796421
R54356 ASIG5V.n570 ASIG5V.n569 0.00796421
R54357 ASIG5V.n568 ASIG5V.n567 0.00796421
R54358 ASIG5V.n566 ASIG5V.n565 0.00796421
R54359 ASIG5V.n564 ASIG5V.n563 0.00796421
R54360 ASIG5V.n562 ASIG5V.n561 0.00796421
R54361 ASIG5V.n560 ASIG5V.n559 0.00796421
R54362 ASIG5V.n558 ASIG5V.n557 0.00796421
R54363 ASIG5V.n556 ASIG5V.n555 0.00796421
R54364 ASIG5V.n554 ASIG5V.n553 0.00796421
R54365 ASIG5V.n552 ASIG5V.n551 0.00796421
R54366 ASIG5V.n550 ASIG5V.n549 0.00796421
R54367 ASIG5V.n548 ASIG5V.n547 0.00796421
R54368 ASIG5V.n546 ASIG5V.n545 0.00796421
R54369 ASIG5V.n544 ASIG5V.n543 0.00796421
R54370 ASIG5V.n542 ASIG5V.n541 0.00796421
R54371 ASIG5V.n540 ASIG5V.n539 0.00796421
R54372 ASIG5V.n538 ASIG5V.n537 0.00796421
R54373 ASIG5V.n536 ASIG5V.n535 0.00796421
R54374 ASIG5V.n534 ASIG5V.n533 0.00796421
R54375 ASIG5V.n532 ASIG5V.n531 0.00796421
R54376 ASIG5V.n530 ASIG5V.n529 0.00796421
R54377 ASIG5V.n528 ASIG5V.n527 0.00796421
R54378 ASIG5V.n526 ASIG5V.n525 0.00796421
R54379 ASIG5V.n524 ASIG5V.n523 0.00796421
R54380 ASIG5V.n2503 ASIG5V.n2502 0.00796421
R54381 ASIG5V.n2505 ASIG5V.n2504 0.00796421
R54382 ASIG5V.n2507 ASIG5V.n2506 0.00796421
R54383 ASIG5V.n2509 ASIG5V.n2508 0.00796421
R54384 ASIG5V.n2511 ASIG5V.n2510 0.00796421
R54385 ASIG5V.n2513 ASIG5V.n2512 0.00796421
R54386 ASIG5V.n2515 ASIG5V.n2514 0.00796421
R54387 ASIG5V.n2517 ASIG5V.n2516 0.00796421
R54388 ASIG5V.n2519 ASIG5V.n2518 0.00796421
R54389 ASIG5V.n2521 ASIG5V.n2520 0.00796421
R54390 ASIG5V.n2523 ASIG5V.n2522 0.00796421
R54391 ASIG5V.n2525 ASIG5V.n2524 0.00796421
R54392 ASIG5V.n2527 ASIG5V.n2526 0.00796421
R54393 ASIG5V.n2529 ASIG5V.n2528 0.00796421
R54394 ASIG5V.n2531 ASIG5V.n2530 0.00796421
R54395 ASIG5V.n2533 ASIG5V.n2532 0.00796421
R54396 ASIG5V.n2535 ASIG5V.n2534 0.00796421
R54397 ASIG5V.n2537 ASIG5V.n2536 0.00796421
R54398 ASIG5V.n2539 ASIG5V.n2538 0.00796421
R54399 ASIG5V.n2541 ASIG5V.n2540 0.00796421
R54400 ASIG5V.n2543 ASIG5V.n2542 0.00796421
R54401 ASIG5V.n2545 ASIG5V.n2544 0.00796421
R54402 ASIG5V.n2547 ASIG5V.n2546 0.00796421
R54403 ASIG5V.n2549 ASIG5V.n2548 0.00796421
R54404 ASIG5V.n2551 ASIG5V.n2550 0.00796421
R54405 ASIG5V.n2553 ASIG5V.n2552 0.00796421
R54406 ASIG5V.n2555 ASIG5V.n2554 0.00796421
R54407 ASIG5V.n2557 ASIG5V.n2556 0.00796421
R54408 ASIG5V.n2559 ASIG5V.n2558 0.00796421
R54409 ASIG5V.n2561 ASIG5V.n2560 0.00796421
R54410 ASIG5V.n2563 ASIG5V.n2562 0.00796421
R54411 ASIG5V.n2565 ASIG5V.n2564 0.00796421
R54412 ASIG5V.n2567 ASIG5V.n2566 0.00796421
R54413 ASIG5V.n2569 ASIG5V.n2568 0.00796421
R54414 ASIG5V.n2571 ASIG5V.n2570 0.00796421
R54415 ASIG5V.n2573 ASIG5V.n2572 0.00796421
R54416 ASIG5V.n2575 ASIG5V.n2574 0.00796421
R54417 ASIG5V.n2577 ASIG5V.n2576 0.00796421
R54418 ASIG5V.n2579 ASIG5V.n2578 0.00796421
R54419 ASIG5V.n2581 ASIG5V.n2580 0.00796421
R54420 ASIG5V.n2583 ASIG5V.n2582 0.00796421
R54421 ASIG5V.n2585 ASIG5V.n2584 0.00796421
R54422 ASIG5V.n2587 ASIG5V.n2586 0.00796421
R54423 ASIG5V.n2589 ASIG5V.n2588 0.00796421
R54424 ASIG5V.n2591 ASIG5V.n2590 0.00796421
R54425 ASIG5V.n2593 ASIG5V.n2592 0.00796421
R54426 ASIG5V.n2595 ASIG5V.n2594 0.00796421
R54427 ASIG5V.n2597 ASIG5V.n2596 0.00796421
R54428 ASIG5V.n2599 ASIG5V.n2598 0.00796421
R54429 ASIG5V.n2601 ASIG5V.n2600 0.00796421
R54430 ASIG5V.n2603 ASIG5V.n2602 0.00796421
R54431 ASIG5V.n2605 ASIG5V.n2604 0.00796421
R54432 ASIG5V.n2607 ASIG5V.n2606 0.00796421
R54433 ASIG5V.n2609 ASIG5V.n2608 0.00796421
R54434 ASIG5V.n2611 ASIG5V.n2610 0.00796421
R54435 ASIG5V.n2613 ASIG5V.n2612 0.00796421
R54436 ASIG5V.n2615 ASIG5V.n2614 0.00796421
R54437 ASIG5V.n2617 ASIG5V.n2616 0.00796421
R54438 ASIG5V.n2619 ASIG5V.n2618 0.00796421
R54439 ASIG5V.n2621 ASIG5V.n2620 0.00796421
R54440 ASIG5V.n2623 ASIG5V.n2622 0.00796421
R54441 ASIG5V.n2625 ASIG5V.n2624 0.00796421
R54442 ASIG5V.n2627 ASIG5V.n2626 0.00796421
R54443 ASIG5V.n9382 ASIG5V.n9381 0.007925
R54444 ASIG5V.n9413 ASIG5V.n9412 0.007925
R54445 ASIG5V.n12980 ASIG5V.n12979 0.0078883
R54446 ASIG5V.n12943 ASIG5V.n12942 0.0078883
R54447 ASIG5V.n12918 ASIG5V.n12917 0.0078883
R54448 ASIG5V.n12810 ASIG5V.n12809 0.0078883
R54449 ASIG5V.n12781 ASIG5V.n12780 0.0078883
R54450 ASIG5V.n12893 ASIG5V.n12892 0.0078883
R54451 ASIG5V.n12864 ASIG5V.n12863 0.0078883
R54452 ASIG5V.n12834 ASIG5V.n12833 0.0078883
R54453 ASIG5V.n13092 ASIG5V.n13091 0.0078883
R54454 ASIG5V.n13120 ASIG5V.n13119 0.0078883
R54455 ASIG5V.n10004 ASIG5V.n10003 0.0078883
R54456 ASIG5V.n10032 ASIG5V.n10031 0.0078883
R54457 ASIG5V.n13261 ASIG5V.n13260 0.0078883
R54458 ASIG5V.n13290 ASIG5V.n13289 0.0078883
R54459 ASIG5V.n13291 ASIG5V.n13290 0.0078883
R54460 ASIG5V.n10063 ASIG5V.n10062 0.0078883
R54461 ASIG5V.n13013 ASIG5V.n13012 0.0078883
R54462 ASIG5V.n13044 ASIG5V.n13043 0.0078883
R54463 ASIG5V.n13160 ASIG5V.n13159 0.0078883
R54464 ASIG5V.n13191 ASIG5V.n13190 0.0078883
R54465 ASIG5V.n13251 ASIG5V.n13250 0.0078883
R54466 ASIG5V.n7147 ASIG5V.n7146 0.0078883
R54467 ASIG5V.n13129 ASIG5V.n13128 0.0078883
R54468 ASIG5V.n13222 ASIG5V.n13221 0.0078883
R54469 ASIG5V.n2012 ASIG5V.n2011 0.0078883
R54470 ASIG5V.n2037 ASIG5V.n2036 0.0078883
R54471 ASIG5V.n2062 ASIG5V.n2061 0.0078883
R54472 ASIG5V.n2087 ASIG5V.n2086 0.0078883
R54473 ASIG5V.n2113 ASIG5V.n2112 0.0078883
R54474 ASIG5V.n2137 ASIG5V.n2136 0.0078883
R54475 ASIG5V.n2162 ASIG5V.n2161 0.0078883
R54476 ASIG5V.n2138 ASIG5V.n2137 0.0078883
R54477 ASIG5V.n1451 ASIG5V.n1450 0.0078883
R54478 ASIG5V.n1513 ASIG5V.n1512 0.0078883
R54479 ASIG5V.n1543 ASIG5V.n1542 0.0078883
R54480 ASIG5V.n1573 ASIG5V.n1572 0.0078883
R54481 ASIG5V.n1633 ASIG5V.n1632 0.0078883
R54482 ASIG5V.n1663 ASIG5V.n1662 0.0078883
R54483 ASIG5V.n1483 ASIG5V.n1482 0.0078883
R54484 ASIG5V.n1604 ASIG5V.n1603 0.0078883
R54485 ASIG5V.n10377 ASIG5V.n10376 0.0078883
R54486 ASIG5V.n10402 ASIG5V.n10401 0.0078883
R54487 ASIG5V.n10427 ASIG5V.n10426 0.0078883
R54488 ASIG5V.n10452 ASIG5V.n10451 0.0078883
R54489 ASIG5V.n10518 ASIG5V.n10517 0.0078883
R54490 ASIG5V.n10550 ASIG5V.n10549 0.0078883
R54491 ASIG5V.n10561 ASIG5V.n10550 0.0078883
R54492 ASIG5V.n9809 ASIG5V.n9808 0.0078883
R54493 ASIG5V.n9840 ASIG5V.n9839 0.0078883
R54494 ASIG5V.n9868 ASIG5V.n9867 0.0078883
R54495 ASIG5V.n9896 ASIG5V.n9895 0.0078883
R54496 ASIG5V.n9924 ASIG5V.n9923 0.0078883
R54497 ASIG5V.n10072 ASIG5V.n10071 0.0078883
R54498 ASIG5V.n10102 ASIG5V.n10101 0.0078883
R54499 ASIG5V.n9813 ASIG5V.n9809 0.0078883
R54500 ASIG5V.n2276 ASIG5V.n2275 0.0078883
R54501 ASIG5V.n2302 ASIG5V.n2301 0.0078883
R54502 ASIG5V.n2327 ASIG5V.n2326 0.0078883
R54503 ASIG5V.n2352 ASIG5V.n2351 0.0078883
R54504 ASIG5V.n2377 ASIG5V.n2376 0.0078883
R54505 ASIG5V.n2427 ASIG5V.n2426 0.0078883
R54506 ASIG5V.n2452 ASIG5V.n2451 0.0078883
R54507 ASIG5V.n2403 ASIG5V.n2402 0.0078883
R54508 ASIG5V.n11958 ASIG5V.n11956 0.00774832
R54509 ASIG5V.n10760 ASIG5V.n10759 0.00772484
R54510 ASIG5V.n2499 ASIG5V.n2498 0.00772484
R54511 ASIG5V.n5969 ASIG5V.n5968 0.00753759
R54512 ASIG5V.n10754 ASIG5V.n10753 0.00753759
R54513 ASIG5V.n976 ASIG5V.n975 0.007475
R54514 ASIG5V.n9424 ASIG5V.n9423 0.007475
R54515 ASIG5V.n4442 ASIG5V.n4441 0.00737773
R54516 ASIG5V.n711 ASIG5V.n710 0.00737773
R54517 ASIG5V.n3330 ASIG5V.n3329 0.0072651
R54518 ASIG5V.n4439 ASIG5V.n4405 0.0072651
R54519 ASIG5V.n2734 ASIG5V.n2733 0.0072651
R54520 ASIG5V.n4438 ASIG5V.n4437 0.0072651
R54521 ASIG5V.n2497 ASIG5V.n1150 0.0071375
R54522 ASIG5V.n10758 ASIG5V.n9515 0.0071375
R54523 ASIG5V.n1063 ASIG5V.n1062 0.007025
R54524 ASIG5V.n1018 ASIG5V.n1017 0.007025
R54525 ASIG5V.n10719 ASIG5V.n10718 0.00699624
R54526 ASIG5V.n7405 ASIG5V.n7402 0.00698472
R54527 ASIG5V.n11762 ASIG5V.n11761 0.00698472
R54528 ASIG5V.n7404 ASIG5V.n7403 0.00698472
R54529 ASIG5V.n9080 ASIG5V.n9079 0.00698472
R54530 ASIG5V.n5971 ASIG5V.n5890 0.00678188
R54531 ASIG5V.n11188 ASIG5V.n11187 0.00678188
R54532 ASIG5V.n5970 ASIG5V.n5922 0.00678188
R54533 ASIG5V.n11019 ASIG5V.n10984 0.00678188
R54534 ASIG5V.n6656 ASIG5V.n6653 0.0065917
R54535 ASIG5V.n11156 ASIG5V.n11155 0.0065917
R54536 ASIG5V.n6655 ASIG5V.n6654 0.0065917
R54537 ASIG5V.n9107 ASIG5V.n9090 0.0065917
R54538 ASIG5V.n5668 ASIG5V.n5667 0.00645489
R54539 ASIG5V.n7128 ASIG5V.n7127 0.00645489
R54540 ASIG5V.n10477 ASIG5V.n10476 0.00638991
R54541 ASIG5V.n12759 ASIG5V.n7271 0.00629866
R54542 ASIG5V.n12645 ASIG5V.n12611 0.00629866
R54543 ASIG5V.n12760 ASIG5V.n7241 0.00629866
R54544 ASIG5V.n12644 ASIG5V.n12643 0.00629866
R54545 ASIG5V.n9431 ASIG5V.n9430 0.0062375
R54546 ASIG5V.n1066 ASIG5V.n1065 0.0062375
R54547 ASIG5V.n1067 ASIG5V.n1066 0.00619869
R54548 ASIG5V.n3625 ASIG5V.n3624 0.00619869
R54549 ASIG5V.n737 ASIG5V.n736 0.00619869
R54550 ASIG5V.n722 ASIG5V.n721 0.00619869
R54551 ASIG5V.n8931 ASIG5V.n8930 0.00597283
R54552 ASIG5V.n8923 ASIG5V.n8922 0.00597283
R54553 ASIG5V.n8915 ASIG5V.n8914 0.00597283
R54554 ASIG5V.n8907 ASIG5V.n8906 0.00597283
R54555 ASIG5V.n8901 ASIG5V.n8900 0.00597283
R54556 ASIG5V.n8891 ASIG5V.n8890 0.00597283
R54557 ASIG5V.n8885 ASIG5V.n8884 0.00597283
R54558 ASIG5V.n10768 ASIG5V.n10767 0.00597283
R54559 ASIG5V.n10774 ASIG5V.n10773 0.00597283
R54560 ASIG5V.n10784 ASIG5V.n10783 0.00597283
R54561 ASIG5V.n10790 ASIG5V.n10789 0.00597283
R54562 ASIG5V.n10800 ASIG5V.n10799 0.00597283
R54563 ASIG5V.n10806 ASIG5V.n10805 0.00597283
R54564 ASIG5V.n10816 ASIG5V.n10815 0.00597283
R54565 ASIG5V.n10822 ASIG5V.n10821 0.00597283
R54566 ASIG5V.n10832 ASIG5V.n10831 0.00597283
R54567 ASIG5V.n10838 ASIG5V.n10837 0.00597283
R54568 ASIG5V.n10848 ASIG5V.n10847 0.00597283
R54569 ASIG5V.n10854 ASIG5V.n10853 0.00597283
R54570 ASIG5V.n10862 ASIG5V.n10861 0.00597283
R54571 ASIG5V.n10870 ASIG5V.n10869 0.00597283
R54572 ASIG5V.n10878 ASIG5V.n10877 0.00597283
R54573 ASIG5V.n10884 ASIG5V.n10883 0.00597283
R54574 ASIG5V.n10888 ASIG5V.n10887 0.00597283
R54575 ASIG5V.n2629 ASIG5V.n2628 0.00597283
R54576 ASIG5V.n9768 ASIG5V.n9767 0.00591907
R54577 ASIG5V.n9776 ASIG5V.n9775 0.00591907
R54578 ASIG5V.n2490 ASIG5V.n2489 0.00591353
R54579 ASIG5V.n2186 ASIG5V.n2185 0.00591353
R54580 ASIG5V.n5670 ASIG5V.n5589 0.00581544
R54581 ASIG5V.n5669 ASIG5V.n5621 0.00581544
R54582 ASIG5V.n1026 ASIG5V.n1025 0.005675
R54583 ASIG5V.n10885 ASIG5V.n10884 0.00564041
R54584 ASIG5V.n10879 ASIG5V.n10878 0.00564041
R54585 ASIG5V.n10871 ASIG5V.n10870 0.00564041
R54586 ASIG5V.n10863 ASIG5V.n10862 0.00564041
R54587 ASIG5V.n10855 ASIG5V.n10854 0.00564041
R54588 ASIG5V.n10849 ASIG5V.n10848 0.00564041
R54589 ASIG5V.n10839 ASIG5V.n10838 0.00564041
R54590 ASIG5V.n10833 ASIG5V.n10832 0.00564041
R54591 ASIG5V.n10823 ASIG5V.n10822 0.00564041
R54592 ASIG5V.n10817 ASIG5V.n10816 0.00564041
R54593 ASIG5V.n10807 ASIG5V.n10806 0.00564041
R54594 ASIG5V.n10801 ASIG5V.n10800 0.00564041
R54595 ASIG5V.n10791 ASIG5V.n10790 0.00564041
R54596 ASIG5V.n10785 ASIG5V.n10784 0.00564041
R54597 ASIG5V.n10775 ASIG5V.n10774 0.00564041
R54598 ASIG5V.n10769 ASIG5V.n10768 0.00564041
R54599 ASIG5V.n8890 ASIG5V.n8889 0.00564041
R54600 ASIG5V.n8900 ASIG5V.n8899 0.00564041
R54601 ASIG5V.n8906 ASIG5V.n8905 0.00564041
R54602 ASIG5V.n8914 ASIG5V.n8913 0.00564041
R54603 ASIG5V.n8922 ASIG5V.n8921 0.00564041
R54604 ASIG5V.n8930 ASIG5V.n8929 0.00564041
R54605 ASIG5V.n8973 ASIG5V.n8935 0.00564041
R54606 ASIG5V.n616 ASIG5V.n576 0.00564041
R54607 ASIG5V.n398 ASIG5V.n397 0.00559443
R54608 ASIG5V.n13257 ASIG5V.n13256 0.00559443
R54609 ASIG5V.n13259 ASIG5V.n13258 0.00559443
R54610 ASIG5V.n13253 ASIG5V.n400 0.00559443
R54611 ASIG5V.n13249 ASIG5V.n13248 0.00559443
R54612 ASIG5V.n1974 ASIG5V.n1973 0.00559443
R54613 ASIG5V.n2192 ASIG5V.n2191 0.00559443
R54614 ASIG5V.n2190 ASIG5V.n2189 0.00559443
R54615 ASIG5V.n10732 ASIG5V.n10731 0.00537218
R54616 ASIG5V.n3135 ASIG5V.n3134 0.00533221
R54617 ASIG5V.n4697 ASIG5V.n4663 0.00533221
R54618 ASIG5V.n2739 ASIG5V.n2738 0.00533221
R54619 ASIG5V.n4696 ASIG5V.n4695 0.00533221
R54620 ASIG5V.n1401 ASIG5V.n1400 0.00529795
R54621 ASIG5V.n1397 ASIG5V.n1396 0.00529795
R54622 ASIG5V.n1390 ASIG5V.n1389 0.00529795
R54623 ASIG5V.n1381 ASIG5V.n1380 0.00529795
R54624 ASIG5V.n1399 ASIG5V.n1398 0.00529795
R54625 ASIG5V.n1388 ASIG5V.n1387 0.00529795
R54626 ASIG5V.n1379 ASIG5V.n1378 0.00529795
R54627 ASIG5V.n1571 ASIG5V.n1570 0.00529795
R54628 ASIG5V.n1403 ASIG5V.n1395 0.00529795
R54629 ASIG5V.n2221 ASIG5V.n2220 0.00529795
R54630 ASIG5V.n2219 ASIG5V.n2218 0.00529795
R54631 ASIG5V.n2217 ASIG5V.n2216 0.00529795
R54632 ASIG5V.n13187 ASIG5V.n13186 0.00529795
R54633 ASIG5V.n13189 ASIG5V.n13188 0.00529795
R54634 ASIG5V.n7173 ASIG5V.n7172 0.00529795
R54635 ASIG5V.n9973 ASIG5V.n9971 0.00529795
R54636 ASIG5V.n10029 ASIG5V.n10028 0.00529795
R54637 ASIG5V.n12861 ASIG5V.n12860 0.00529795
R54638 ASIG5V.n10297 ASIG5V.n10296 0.00529795
R54639 ASIG5V.n10304 ASIG5V.n10302 0.00529795
R54640 ASIG5V.n1601 ASIG5V.n1600 0.00529795
R54641 ASIG5V.n1394 ASIG5V.n1386 0.00529795
R54642 ASIG5V.n2210 ASIG5V.n2209 0.00529795
R54643 ASIG5V.n2208 ASIG5V.n2207 0.00529795
R54644 ASIG5V.n13219 ASIG5V.n13218 0.00529795
R54645 ASIG5V.n7171 ASIG5V.n7170 0.00529795
R54646 ASIG5V.n10060 ASIG5V.n10056 0.00529795
R54647 ASIG5V.n10059 ASIG5V.n10058 0.00529795
R54648 ASIG5V.n10482 ASIG5V.n10481 0.00529795
R54649 ASIG5V.n9745 ASIG5V.n9744 0.00529795
R54650 ASIG5V.n1631 ASIG5V.n1630 0.00529795
R54651 ASIG5V.n1385 ASIG5V.n1377 0.00529795
R54652 ASIG5V.n2200 ASIG5V.n2199 0.00529795
R54653 ASIG5V.n2198 ASIG5V.n2197 0.00529795
R54654 ASIG5V.n12807 ASIG5V.n12806 0.00529795
R54655 ASIG5V.n10511 ASIG5V.n10510 0.00529795
R54656 ASIG5V.n10513 ASIG5V.n10512 0.00529795
R54657 ASIG5V.n9735 ASIG5V.n9734 0.00529795
R54658 ASIG5V.n9737 ASIG5V.n9736 0.00529795
R54659 ASIG5V.n1661 ASIG5V.n1660 0.00529795
R54660 ASIG5V.n1376 ASIG5V.n1369 0.00529795
R54661 ASIG5V.n1371 ASIG5V.n1370 0.00529795
R54662 ASIG5V.n2195 ASIG5V.n2188 0.00529795
R54663 ASIG5V.n7144 ASIG5V.n7142 0.00529795
R54664 ASIG5V.n403 ASIG5V.n402 0.00529795
R54665 ASIG5V.n395 ASIG5V.n394 0.00529795
R54666 ASIG5V.n13288 ASIG5V.n13285 0.00529795
R54667 ASIG5V.n13287 ASIG5V.n13286 0.00529795
R54668 ASIG5V.n12778 ASIG5V.n12776 0.00529795
R54669 ASIG5V.n10542 ASIG5V.n10541 0.00529795
R54670 ASIG5V.n10546 ASIG5V.n10545 0.00529795
R54671 ASIG5V.n984 ASIG5V.n983 0.005225
R54672 ASIG5V.n1449 ASIG5V.n1448 0.00514086
R54673 ASIG5V.n1433 ASIG5V.n1427 0.00514086
R54674 ASIG5V.n3138 ASIG5V.n3137 0.00501965
R54675 ASIG5V.n730 ASIG5V.n729 0.00501965
R54676 ASIG5V.n1541 ASIG5V.n1540 0.0048617
R54677 ASIG5V.n1412 ASIG5V.n1404 0.0048617
R54678 ASIG5V.n1410 ASIG5V.n1409 0.0048617
R54679 ASIG5V.n1406 ASIG5V.n1405 0.0048617
R54680 ASIG5V.n2230 ASIG5V.n2229 0.0048617
R54681 ASIG5V.n2228 ASIG5V.n2227 0.0048617
R54682 ASIG5V.n2226 ASIG5V.n2225 0.0048617
R54683 ASIG5V.n13156 ASIG5V.n13155 0.0048617
R54684 ASIG5V.n13158 ASIG5V.n13157 0.0048617
R54685 ASIG5V.n7175 ASIG5V.n7174 0.0048617
R54686 ASIG5V.n9978 ASIG5V.n9976 0.0048617
R54687 ASIG5V.n10001 ASIG5V.n10000 0.0048617
R54688 ASIG5V.n12890 ASIG5V.n12889 0.0048617
R54689 ASIG5V.n10306 ASIG5V.n10305 0.0048617
R54690 ASIG5V.n10313 ASIG5V.n10311 0.0048617
R54691 ASIG5V.n1511 ASIG5V.n1510 0.0048617
R54692 ASIG5V.n1421 ASIG5V.n1413 0.0048617
R54693 ASIG5V.n1419 ASIG5V.n1418 0.0048617
R54694 ASIG5V.n1415 ASIG5V.n1414 0.0048617
R54695 ASIG5V.n2239 ASIG5V.n2238 0.0048617
R54696 ASIG5V.n2237 ASIG5V.n2236 0.0048617
R54697 ASIG5V.n2235 ASIG5V.n2234 0.0048617
R54698 ASIG5V.n7181 ASIG5V.n7178 0.0048617
R54699 ASIG5V.n7180 ASIG5V.n7179 0.0048617
R54700 ASIG5V.n13124 ASIG5V.n13123 0.0048617
R54701 ASIG5V.n13117 ASIG5V.n13116 0.0048617
R54702 ASIG5V.n10317 ASIG5V.n10316 0.0048617
R54703 ASIG5V.n10319 ASIG5V.n10318 0.0048617
R54704 ASIG5V.n10321 ASIG5V.n10320 0.0048617
R54705 ASIG5V.n10326 ASIG5V.n10324 0.0048617
R54706 ASIG5V.n13127 ASIG5V.n7183 0.0048617
R54707 ASIG5V.n1425 ASIG5V.n1424 0.0048617
R54708 ASIG5V.n1479 ASIG5V.n1478 0.0048617
R54709 ASIG5V.n2249 ASIG5V.n2248 0.0048617
R54710 ASIG5V.n2247 ASIG5V.n2246 0.0048617
R54711 ASIG5V.n2245 ASIG5V.n2244 0.0048617
R54712 ASIG5V.n13040 ASIG5V.n13039 0.0048617
R54713 ASIG5V.n13042 ASIG5V.n13041 0.0048617
R54714 ASIG5V.n13046 ASIG5V.n7185 0.0048617
R54715 ASIG5V.n13051 ASIG5V.n13049 0.0048617
R54716 ASIG5V.n13089 ASIG5V.n13088 0.0048617
R54717 ASIG5V.n10330 ASIG5V.n10329 0.0048617
R54718 ASIG5V.n10332 ASIG5V.n10331 0.0048617
R54719 ASIG5V.n10334 ASIG5V.n10333 0.0048617
R54720 ASIG5V.n10339 ASIG5V.n10337 0.0048617
R54721 ASIG5V.n1429 ASIG5V.n1428 0.0048617
R54722 ASIG5V.n2256 ASIG5V.n2255 0.0048617
R54723 ASIG5V.n2254 ASIG5V.n2253 0.0048617
R54724 ASIG5V.n12998 ASIG5V.n7207 0.0048617
R54725 ASIG5V.n12997 ASIG5V.n12996 0.0048617
R54726 ASIG5V.n12995 ASIG5V.n12994 0.0048617
R54727 ASIG5V.n12991 ASIG5V.n12990 0.0048617
R54728 ASIG5V.n12989 ASIG5V.n12988 0.0048617
R54729 ASIG5V.n12987 ASIG5V.n12986 0.0048617
R54730 ASIG5V.n12983 ASIG5V.n12982 0.0048617
R54731 ASIG5V.n9798 ASIG5V.n9797 0.0048617
R54732 ASIG5V.n9800 ASIG5V.n9799 0.0048617
R54733 ASIG5V.n9802 ASIG5V.n9801 0.0048617
R54734 ASIG5V.n1408 ASIG5V.n1407 0.0048617
R54735 ASIG5V.n1417 ASIG5V.n1416 0.0048617
R54736 ASIG5V.n1477 ASIG5V.n1476 0.0048617
R54737 ASIG5V.n2263 ASIG5V.n2262 0.0048617
R54738 ASIG5V.n13352 ASIG5V.n361 0.00484899
R54739 ASIG5V.n12149 ASIG5V.n12115 0.00484899
R54740 ASIG5V.n13351 ASIG5V.n393 0.00484899
R54741 ASIG5V.n12148 ASIG5V.n12147 0.00484899
R54742 ASIG5V.n6766 ASIG5V.n6765 0.00483083
R54743 ASIG5V.n10739 ASIG5V.n10738 0.00483083
R54744 ASIG5V.n10742 ASIG5V.n10741 0.00483083
R54745 ASIG5V.n9390 ASIG5V.n9389 0.004775
R54746 ASIG5V.n9405 ASIG5V.n9404 0.004775
R54747 ASIG5V.n6330 ASIG5V.n6327 0.00462664
R54748 ASIG5V.n6329 ASIG5V.n6328 0.00462664
R54749 ASIG5V.n6768 ASIG5V.n6687 0.00436577
R54750 ASIG5V.n11827 ASIG5V.n11793 0.00436577
R54751 ASIG5V.n6767 ASIG5V.n6719 0.00436577
R54752 ASIG5V.n11826 ASIG5V.n11825 0.00436577
R54753 ASIG5V.n999 ASIG5V.n998 0.004325
R54754 ASIG5V.n2481 ASIG5V.n2480 0.00428947
R54755 ASIG5V.n2473 ASIG5V.n2472 0.00428947
R54756 ASIG5V.n13350 ASIG5V.n13349 0.00428947
R54757 ASIG5V.n12756 ASIG5V.n12753 0.00423362
R54758 ASIG5V.n12084 ASIG5V.n12083 0.00423362
R54759 ASIG5V.n12755 ASIG5V.n12754 0.00423362
R54760 ASIG5V.n9072 ASIG5V.n9071 0.00423362
R54761 ASIG5V.n10096 ASIG5V.n10095 0.00396691
R54762 ASIG5V.n3622 ASIG5V.n3588 0.00388255
R54763 ASIG5V.n4163 ASIG5V.n4129 0.00388255
R54764 ASIG5V.n3621 ASIG5V.n3620 0.00388255
R54765 ASIG5V.n4162 ASIG5V.n4161 0.00388255
R54766 ASIG5V.n4970 ASIG5V.n4967 0.00384061
R54767 ASIG5V.n4969 ASIG5V.n4968 0.00384061
R54768 ASIG5V.n9865 ASIG5V.n9864 0.00374825
R54769 ASIG5V.n9837 ASIG5V.n9836 0.00374825
R54770 ASIG5V.n9812 ASIG5V.n9811 0.00374825
R54771 ASIG5V.n2176 ASIG5V.n2175 0.00374812
R54772 ASIG5V.n7127 ASIG5V.n450 0.00374812
R54773 ASIG5V.n10750 ASIG5V.n10749 0.00374812
R54774 ASIG5V.n7125 ASIG5V.n512 0.00339933
R54775 ASIG5V.n11415 ASIG5V.n11414 0.00339933
R54776 ASIG5V.n7126 ASIG5V.n482 0.00339933
R54777 ASIG5V.n10981 ASIG5V.n10929 0.00339933
R54778 ASIG5V.n7933 ASIG5V.n7932 0.00320677
R54779 ASIG5V.n10723 ASIG5V.n10722 0.00320677
R54780 ASIG5V.n7935 ASIG5V.n7853 0.00291611
R54781 ASIG5V.n12419 ASIG5V.n12385 0.00291611
R54782 ASIG5V.n7934 ASIG5V.n7885 0.00291611
R54783 ASIG5V.n12418 ASIG5V.n12417 0.00291611
R54784 ASIG5V.n12974 ASIG5V.n12973 0.00268244
R54785 ASIG5V.n12963 ASIG5V.n12962 0.00268244
R54786 ASIG5V.n12947 ASIG5V.n12946 0.00268244
R54787 ASIG5V.n12937 ASIG5V.n12936 0.00268244
R54788 ASIG5V.n12922 ASIG5V.n12921 0.00268244
R54789 ASIG5V.n12912 ASIG5V.n12911 0.00268244
R54790 ASIG5V.n12897 ASIG5V.n12896 0.00268244
R54791 ASIG5V.n12883 ASIG5V.n12882 0.00268244
R54792 ASIG5V.n12868 ASIG5V.n12867 0.00268244
R54793 ASIG5V.n12854 ASIG5V.n12853 0.00268244
R54794 ASIG5V.n12839 ASIG5V.n12838 0.00268244
R54795 ASIG5V.n12829 ASIG5V.n12828 0.00268244
R54796 ASIG5V.n12814 ASIG5V.n12813 0.00268244
R54797 ASIG5V.n12800 ASIG5V.n12799 0.00268244
R54798 ASIG5V.n12785 ASIG5V.n12784 0.00268244
R54799 ASIG5V.n12771 ASIG5V.n12770 0.00268244
R54800 ASIG5V.n12884 ASIG5V.n12883 0.00268244
R54801 ASIG5V.n12855 ASIG5V.n12854 0.00268244
R54802 ASIG5V.n12869 ASIG5V.n12868 0.00268244
R54803 ASIG5V.n12898 ASIG5V.n12897 0.00268244
R54804 ASIG5V.n12830 ASIG5V.n12829 0.00268244
R54805 ASIG5V.n12840 ASIG5V.n12839 0.00268244
R54806 ASIG5V.n13060 ASIG5V.n13059 0.00268244
R54807 ASIG5V.n13070 ASIG5V.n13069 0.00268244
R54808 ASIG5V.n13085 ASIG5V.n13084 0.00268244
R54809 ASIG5V.n13098 ASIG5V.n13097 0.00268244
R54810 ASIG5V.n13113 ASIG5V.n13112 0.00268244
R54811 ASIG5V.n9982 ASIG5V.n9981 0.00268244
R54812 ASIG5V.n9997 ASIG5V.n9996 0.00268244
R54813 ASIG5V.n10010 ASIG5V.n10009 0.00268244
R54814 ASIG5V.n10025 ASIG5V.n10024 0.00268244
R54815 ASIG5V.n10038 ASIG5V.n10037 0.00268244
R54816 ASIG5V.n10053 ASIG5V.n10052 0.00268244
R54817 ASIG5V.n9966 ASIG5V.n9965 0.00268244
R54818 ASIG5V.n9950 ASIG5V.n9949 0.00268244
R54819 ASIG5V.n13267 ASIG5V.n13266 0.00268244
R54820 ASIG5V.n13282 ASIG5V.n13281 0.00268244
R54821 ASIG5V.n13296 ASIG5V.n13295 0.00268244
R54822 ASIG5V.n10037 ASIG5V.n10036 0.00268244
R54823 ASIG5V.n10009 ASIG5V.n10008 0.00268244
R54824 ASIG5V.n10024 ASIG5V.n10023 0.00268244
R54825 ASIG5V.n9996 ASIG5V.n9995 0.00268244
R54826 ASIG5V.n10052 ASIG5V.n10051 0.00268244
R54827 ASIG5V.n9965 ASIG5V.n9964 0.00268244
R54828 ASIG5V.n9981 ASIG5V.n9980 0.00268244
R54829 ASIG5V.n12913 ASIG5V.n12912 0.00268244
R54830 ASIG5V.n12923 ASIG5V.n12922 0.00268244
R54831 ASIG5V.n13112 ASIG5V.n13111 0.00268244
R54832 ASIG5V.n13007 ASIG5V.n13006 0.00268244
R54833 ASIG5V.n13018 ASIG5V.n13017 0.00268244
R54834 ASIG5V.n13034 ASIG5V.n13033 0.00268244
R54835 ASIG5V.n7203 ASIG5V.n7202 0.00268244
R54836 ASIG5V.n7188 ASIG5V.n7187 0.00268244
R54837 ASIG5V.n13135 ASIG5V.n13134 0.00268244
R54838 ASIG5V.n13150 ASIG5V.n13149 0.00268244
R54839 ASIG5V.n13166 ASIG5V.n13165 0.00268244
R54840 ASIG5V.n13181 ASIG5V.n13180 0.00268244
R54841 ASIG5V.n13197 ASIG5V.n13196 0.00268244
R54842 ASIG5V.n13212 ASIG5V.n13211 0.00268244
R54843 ASIG5V.n13227 ASIG5V.n13226 0.00268244
R54844 ASIG5V.n13242 ASIG5V.n13241 0.00268244
R54845 ASIG5V.n7166 ASIG5V.n7165 0.00268244
R54846 ASIG5V.n7151 ASIG5V.n7150 0.00268244
R54847 ASIG5V.n7136 ASIG5V.n7135 0.00268244
R54848 ASIG5V.n13134 ASIG5V.n13133 0.00268244
R54849 ASIG5V.n13165 ASIG5V.n13164 0.00268244
R54850 ASIG5V.n13196 ASIG5V.n13195 0.00268244
R54851 ASIG5V.n13226 ASIG5V.n13225 0.00268244
R54852 ASIG5V.n13180 ASIG5V.n13179 0.00268244
R54853 ASIG5V.n13149 ASIG5V.n13148 0.00268244
R54854 ASIG5V.n7189 ASIG5V.n7188 0.00268244
R54855 ASIG5V.n13211 ASIG5V.n13210 0.00268244
R54856 ASIG5V.n7167 ASIG5V.n7166 0.00268244
R54857 ASIG5V.n13266 ASIG5V.n13265 0.00268244
R54858 ASIG5V.n12801 ASIG5V.n12800 0.00268244
R54859 ASIG5V.n12815 ASIG5V.n12814 0.00268244
R54860 ASIG5V.n9951 ASIG5V.n9950 0.00268244
R54861 ASIG5V.n13241 ASIG5V.n13240 0.00268244
R54862 ASIG5V.n1983 ASIG5V.n1982 0.00268244
R54863 ASIG5V.n1993 ASIG5V.n1992 0.00268244
R54864 ASIG5V.n2008 ASIG5V.n2007 0.00268244
R54865 ASIG5V.n2018 ASIG5V.n2017 0.00268244
R54866 ASIG5V.n2033 ASIG5V.n2032 0.00268244
R54867 ASIG5V.n2043 ASIG5V.n2042 0.00268244
R54868 ASIG5V.n2058 ASIG5V.n2057 0.00268244
R54869 ASIG5V.n2068 ASIG5V.n2067 0.00268244
R54870 ASIG5V.n2083 ASIG5V.n2082 0.00268244
R54871 ASIG5V.n2093 ASIG5V.n2092 0.00268244
R54872 ASIG5V.n2108 ASIG5V.n2107 0.00268244
R54873 ASIG5V.n2118 ASIG5V.n2117 0.00268244
R54874 ASIG5V.n2133 ASIG5V.n2132 0.00268244
R54875 ASIG5V.n2142 ASIG5V.n2141 0.00268244
R54876 ASIG5V.n2158 ASIG5V.n2157 0.00268244
R54877 ASIG5V.n2168 ASIG5V.n2167 0.00268244
R54878 ASIG5V.n2117 ASIG5V.n2116 0.00268244
R54879 ASIG5V.n2092 ASIG5V.n2091 0.00268244
R54880 ASIG5V.n2067 ASIG5V.n2066 0.00268244
R54881 ASIG5V.n2042 ASIG5V.n2041 0.00268244
R54882 ASIG5V.n2082 ASIG5V.n2081 0.00268244
R54883 ASIG5V.n2057 ASIG5V.n2056 0.00268244
R54884 ASIG5V.n2032 ASIG5V.n2031 0.00268244
R54885 ASIG5V.n2107 ASIG5V.n2106 0.00268244
R54886 ASIG5V.n2132 ASIG5V.n2131 0.00268244
R54887 ASIG5V.n2143 ASIG5V.n2142 0.00268244
R54888 ASIG5V.n2017 ASIG5V.n2016 0.00268244
R54889 ASIG5V.n7204 ASIG5V.n7203 0.00268244
R54890 ASIG5V.n13097 ASIG5V.n13096 0.00268244
R54891 ASIG5V.n12938 ASIG5V.n12937 0.00268244
R54892 ASIG5V.n12948 ASIG5V.n12947 0.00268244
R54893 ASIG5V.n13084 ASIG5V.n13083 0.00268244
R54894 ASIG5V.n13033 ASIG5V.n13032 0.00268244
R54895 ASIG5V.n2007 ASIG5V.n2006 0.00268244
R54896 ASIG5V.n1442 ASIG5V.n1441 0.00268244
R54897 ASIG5V.n1457 ASIG5V.n1456 0.00268244
R54898 ASIG5V.n1472 ASIG5V.n1471 0.00268244
R54899 ASIG5V.n1489 ASIG5V.n1488 0.00268244
R54900 ASIG5V.n1504 ASIG5V.n1503 0.00268244
R54901 ASIG5V.n1519 ASIG5V.n1518 0.00268244
R54902 ASIG5V.n1534 ASIG5V.n1533 0.00268244
R54903 ASIG5V.n1549 ASIG5V.n1548 0.00268244
R54904 ASIG5V.n1564 ASIG5V.n1563 0.00268244
R54905 ASIG5V.n1579 ASIG5V.n1578 0.00268244
R54906 ASIG5V.n1594 ASIG5V.n1593 0.00268244
R54907 ASIG5V.n1609 ASIG5V.n1608 0.00268244
R54908 ASIG5V.n1624 ASIG5V.n1623 0.00268244
R54909 ASIG5V.n1639 ASIG5V.n1638 0.00268244
R54910 ASIG5V.n1654 ASIG5V.n1653 0.00268244
R54911 ASIG5V.n1669 ASIG5V.n1668 0.00268244
R54912 ASIG5V.n1488 ASIG5V.n1487 0.00268244
R54913 ASIG5V.n1518 ASIG5V.n1517 0.00268244
R54914 ASIG5V.n1548 ASIG5V.n1547 0.00268244
R54915 ASIG5V.n1578 ASIG5V.n1577 0.00268244
R54916 ASIG5V.n1608 ASIG5V.n1607 0.00268244
R54917 ASIG5V.n1638 ASIG5V.n1637 0.00268244
R54918 ASIG5V.n1563 ASIG5V.n1562 0.00268244
R54919 ASIG5V.n1533 ASIG5V.n1532 0.00268244
R54920 ASIG5V.n1503 ASIG5V.n1502 0.00268244
R54921 ASIG5V.n1471 ASIG5V.n1470 0.00268244
R54922 ASIG5V.n1593 ASIG5V.n1592 0.00268244
R54923 ASIG5V.n1623 ASIG5V.n1622 0.00268244
R54924 ASIG5V.n1668 ASIG5V.n1667 0.00268244
R54925 ASIG5V.n2167 ASIG5V.n2166 0.00268244
R54926 ASIG5V.n7137 ASIG5V.n7136 0.00268244
R54927 ASIG5V.n7152 ASIG5V.n7151 0.00268244
R54928 ASIG5V.n2157 ASIG5V.n2156 0.00268244
R54929 ASIG5V.n1653 ASIG5V.n1652 0.00268244
R54930 ASIG5V.n12786 ASIG5V.n12785 0.00268244
R54931 ASIG5V.n13281 ASIG5V.n13280 0.00268244
R54932 ASIG5V.n13295 ASIG5V.n13294 0.00268244
R54933 ASIG5V.n12770 ASIG5V.n12769 0.00268244
R54934 ASIG5V.n10348 ASIG5V.n10347 0.00268244
R54935 ASIG5V.n10358 ASIG5V.n10357 0.00268244
R54936 ASIG5V.n10373 ASIG5V.n10372 0.00268244
R54937 ASIG5V.n10383 ASIG5V.n10382 0.00268244
R54938 ASIG5V.n10398 ASIG5V.n10397 0.00268244
R54939 ASIG5V.n10408 ASIG5V.n10407 0.00268244
R54940 ASIG5V.n10423 ASIG5V.n10422 0.00268244
R54941 ASIG5V.n10433 ASIG5V.n10432 0.00268244
R54942 ASIG5V.n10448 ASIG5V.n10447 0.00268244
R54943 ASIG5V.n10458 ASIG5V.n10457 0.00268244
R54944 ASIG5V.n10473 ASIG5V.n10472 0.00268244
R54945 ASIG5V.n10492 ASIG5V.n10491 0.00268244
R54946 ASIG5V.n10507 ASIG5V.n10506 0.00268244
R54947 ASIG5V.n10523 ASIG5V.n10522 0.00268244
R54948 ASIG5V.n10538 ASIG5V.n10537 0.00268244
R54949 ASIG5V.n10565 ASIG5V.n10564 0.00268244
R54950 ASIG5V.n10457 ASIG5V.n10456 0.00268244
R54951 ASIG5V.n10447 ASIG5V.n10446 0.00268244
R54952 ASIG5V.n10432 ASIG5V.n10431 0.00268244
R54953 ASIG5V.n10422 ASIG5V.n10421 0.00268244
R54954 ASIG5V.n10407 ASIG5V.n10406 0.00268244
R54955 ASIG5V.n10397 ASIG5V.n10396 0.00268244
R54956 ASIG5V.n10382 ASIG5V.n10381 0.00268244
R54957 ASIG5V.n10372 ASIG5V.n10371 0.00268244
R54958 ASIG5V.n10472 ASIG5V.n10471 0.00268244
R54959 ASIG5V.n10491 ASIG5V.n10490 0.00268244
R54960 ASIG5V.n10506 ASIG5V.n10505 0.00268244
R54961 ASIG5V.n10522 ASIG5V.n10521 0.00268244
R54962 ASIG5V.n10537 ASIG5V.n10536 0.00268244
R54963 ASIG5V.n10566 ASIG5V.n10565 0.00268244
R54964 ASIG5V.n1456 ASIG5V.n1455 0.00268244
R54965 ASIG5V.n10347 ASIG5V.n10346 0.00268244
R54966 ASIG5V.n12973 ASIG5V.n12972 0.00268244
R54967 ASIG5V.n13059 ASIG5V.n13058 0.00268244
R54968 ASIG5V.n13006 ASIG5V.n13005 0.00268244
R54969 ASIG5V.n1982 ASIG5V.n1981 0.00268244
R54970 ASIG5V.n1441 ASIG5V.n1440 0.00268244
R54971 ASIG5V.n1992 ASIG5V.n1991 0.00268244
R54972 ASIG5V.n13069 ASIG5V.n13068 0.00268244
R54973 ASIG5V.n10357 ASIG5V.n10356 0.00268244
R54974 ASIG5V.n13019 ASIG5V.n13018 0.00268244
R54975 ASIG5V.n12962 ASIG5V.n12961 0.00268244
R54976 ASIG5V.n9791 ASIG5V.n9790 0.00268244
R54977 ASIG5V.n9818 ASIG5V.n9817 0.00268244
R54978 ASIG5V.n9833 ASIG5V.n9832 0.00268244
R54979 ASIG5V.n9846 ASIG5V.n9845 0.00268244
R54980 ASIG5V.n9861 ASIG5V.n9860 0.00268244
R54981 ASIG5V.n9874 ASIG5V.n9873 0.00268244
R54982 ASIG5V.n9889 ASIG5V.n9888 0.00268244
R54983 ASIG5V.n9902 ASIG5V.n9901 0.00268244
R54984 ASIG5V.n9917 ASIG5V.n9916 0.00268244
R54985 ASIG5V.n9930 ASIG5V.n9929 0.00268244
R54986 ASIG5V.n9945 ASIG5V.n9944 0.00268244
R54987 ASIG5V.n10077 ASIG5V.n10076 0.00268244
R54988 ASIG5V.n10092 ASIG5V.n10091 0.00268244
R54989 ASIG5V.n10107 ASIG5V.n10106 0.00268244
R54990 ASIG5V.n10122 ASIG5V.n10121 0.00268244
R54991 ASIG5V.n10132 ASIG5V.n10131 0.00268244
R54992 ASIG5V.n10131 ASIG5V.n10130 0.00268244
R54993 ASIG5V.n10106 ASIG5V.n10105 0.00268244
R54994 ASIG5V.n10076 ASIG5V.n10075 0.00268244
R54995 ASIG5V.n9929 ASIG5V.n9928 0.00268244
R54996 ASIG5V.n9901 ASIG5V.n9900 0.00268244
R54997 ASIG5V.n9873 ASIG5V.n9872 0.00268244
R54998 ASIG5V.n9845 ASIG5V.n9844 0.00268244
R54999 ASIG5V.n9817 ASIG5V.n9816 0.00268244
R55000 ASIG5V.n9790 ASIG5V.n9789 0.00268244
R55001 ASIG5V.n9916 ASIG5V.n9915 0.00268244
R55002 ASIG5V.n9888 ASIG5V.n9887 0.00268244
R55003 ASIG5V.n9860 ASIG5V.n9859 0.00268244
R55004 ASIG5V.n9832 ASIG5V.n9831 0.00268244
R55005 ASIG5V.n9944 ASIG5V.n9943 0.00268244
R55006 ASIG5V.n10091 ASIG5V.n10090 0.00268244
R55007 ASIG5V.n10121 ASIG5V.n10120 0.00268244
R55008 ASIG5V.n2272 ASIG5V.n2271 0.00268244
R55009 ASIG5V.n2282 ASIG5V.n2281 0.00268244
R55010 ASIG5V.n2297 ASIG5V.n2296 0.00268244
R55011 ASIG5V.n2308 ASIG5V.n2307 0.00268244
R55012 ASIG5V.n2323 ASIG5V.n2322 0.00268244
R55013 ASIG5V.n2333 ASIG5V.n2332 0.00268244
R55014 ASIG5V.n2348 ASIG5V.n2347 0.00268244
R55015 ASIG5V.n2358 ASIG5V.n2357 0.00268244
R55016 ASIG5V.n2373 ASIG5V.n2372 0.00268244
R55017 ASIG5V.n2383 ASIG5V.n2382 0.00268244
R55018 ASIG5V.n2398 ASIG5V.n2397 0.00268244
R55019 ASIG5V.n2408 ASIG5V.n2407 0.00268244
R55020 ASIG5V.n2423 ASIG5V.n2422 0.00268244
R55021 ASIG5V.n2433 ASIG5V.n2432 0.00268244
R55022 ASIG5V.n2448 ASIG5V.n2447 0.00268244
R55023 ASIG5V.n2458 ASIG5V.n2457 0.00268244
R55024 ASIG5V.n2271 ASIG5V.n2270 0.00268244
R55025 ASIG5V.n2307 ASIG5V.n2306 0.00268244
R55026 ASIG5V.n2332 ASIG5V.n2331 0.00268244
R55027 ASIG5V.n2357 ASIG5V.n2356 0.00268244
R55028 ASIG5V.n2382 ASIG5V.n2381 0.00268244
R55029 ASIG5V.n2407 ASIG5V.n2406 0.00268244
R55030 ASIG5V.n2432 ASIG5V.n2431 0.00268244
R55031 ASIG5V.n2457 ASIG5V.n2456 0.00268244
R55032 ASIG5V.n2281 ASIG5V.n2280 0.00268244
R55033 ASIG5V.n2372 ASIG5V.n2371 0.00268244
R55034 ASIG5V.n2347 ASIG5V.n2346 0.00268244
R55035 ASIG5V.n2322 ASIG5V.n2321 0.00268244
R55036 ASIG5V.n2296 ASIG5V.n2295 0.00268244
R55037 ASIG5V.n2397 ASIG5V.n2396 0.00268244
R55038 ASIG5V.n2422 ASIG5V.n2421 0.00268244
R55039 ASIG5V.n2447 ASIG5V.n2446 0.00268244
R55040 ASIG5V.n2478 ASIG5V.n2477 0.00266541
R55041 ASIG5V.n2178 ASIG5V.n2177 0.00266541
R55042 ASIG5V.n2817 ASIG5V.n2746 0.0026375
R55043 ASIG5V.n11094 ASIG5V.n11023 0.0026375
R55044 ASIG5V.n11096 ASIG5V.n11095 0.0026375
R55045 ASIG5V.n2819 ASIG5V.n2818 0.0026375
R55046 ASIG5V.n1003 ASIG5V.n1002 0.002525
R55047 ASIG5V.n12970 ASIG5V.n12969 0.0025054
R55048 ASIG5V.n12951 ASIG5V.n12950 0.0025054
R55049 ASIG5V.n12926 ASIG5V.n12925 0.0025054
R55050 ASIG5V.n12901 ASIG5V.n12900 0.0025054
R55051 ASIG5V.n12872 ASIG5V.n12871 0.0025054
R55052 ASIG5V.n12843 ASIG5V.n12842 0.0025054
R55053 ASIG5V.n12818 ASIG5V.n12817 0.0025054
R55054 ASIG5V.n12789 ASIG5V.n12788 0.0025054
R55055 ASIG5V.n12902 ASIG5V.n12901 0.0025054
R55056 ASIG5V.n12873 ASIG5V.n12872 0.0025054
R55057 ASIG5V.n12844 ASIG5V.n12843 0.0025054
R55058 ASIG5V.n13056 ASIG5V.n13055 0.0025054
R55059 ASIG5V.n13081 ASIG5V.n13080 0.0025054
R55060 ASIG5V.n13109 ASIG5V.n13108 0.0025054
R55061 ASIG5V.n9993 ASIG5V.n9992 0.0025054
R55062 ASIG5V.n10021 ASIG5V.n10020 0.0025054
R55063 ASIG5V.n10049 ASIG5V.n10048 0.0025054
R55064 ASIG5V.n9954 ASIG5V.n9953 0.0025054
R55065 ASIG5V.n13278 ASIG5V.n13277 0.0025054
R55066 ASIG5V.n10048 ASIG5V.n10047 0.0025054
R55067 ASIG5V.n10020 ASIG5V.n10019 0.0025054
R55068 ASIG5V.n9992 ASIG5V.n9991 0.0025054
R55069 ASIG5V.n13108 ASIG5V.n13107 0.0025054
R55070 ASIG5V.n12927 ASIG5V.n12926 0.0025054
R55071 ASIG5V.n13003 ASIG5V.n13002 0.0025054
R55072 ASIG5V.n13030 ASIG5V.n13029 0.0025054
R55073 ASIG5V.n7192 ASIG5V.n7191 0.0025054
R55074 ASIG5V.n13146 ASIG5V.n13145 0.0025054
R55075 ASIG5V.n13177 ASIG5V.n13176 0.0025054
R55076 ASIG5V.n13208 ASIG5V.n13207 0.0025054
R55077 ASIG5V.n13238 ASIG5V.n13237 0.0025054
R55078 ASIG5V.n7155 ASIG5V.n7154 0.0025054
R55079 ASIG5V.n7193 ASIG5V.n7192 0.0025054
R55080 ASIG5V.n13145 ASIG5V.n13144 0.0025054
R55081 ASIG5V.n13176 ASIG5V.n13175 0.0025054
R55082 ASIG5V.n13207 ASIG5V.n13206 0.0025054
R55083 ASIG5V.n13237 ASIG5V.n13236 0.0025054
R55084 ASIG5V.n9955 ASIG5V.n9954 0.0025054
R55085 ASIG5V.n12819 ASIG5V.n12818 0.0025054
R55086 ASIG5V.n1979 ASIG5V.n1978 0.0025054
R55087 ASIG5V.n2004 ASIG5V.n2003 0.0025054
R55088 ASIG5V.n2029 ASIG5V.n2028 0.0025054
R55089 ASIG5V.n2054 ASIG5V.n2053 0.0025054
R55090 ASIG5V.n2079 ASIG5V.n2078 0.0025054
R55091 ASIG5V.n2104 ASIG5V.n2103 0.0025054
R55092 ASIG5V.n2129 ASIG5V.n2128 0.0025054
R55093 ASIG5V.n2154 ASIG5V.n2153 0.0025054
R55094 ASIG5V.n2128 ASIG5V.n2127 0.0025054
R55095 ASIG5V.n2103 ASIG5V.n2102 0.0025054
R55096 ASIG5V.n2078 ASIG5V.n2077 0.0025054
R55097 ASIG5V.n2053 ASIG5V.n2052 0.0025054
R55098 ASIG5V.n2028 ASIG5V.n2027 0.0025054
R55099 ASIG5V.n2003 ASIG5V.n2002 0.0025054
R55100 ASIG5V.n13029 ASIG5V.n13028 0.0025054
R55101 ASIG5V.n13080 ASIG5V.n13079 0.0025054
R55102 ASIG5V.n12952 ASIG5V.n12951 0.0025054
R55103 ASIG5V.n1438 ASIG5V.n1437 0.0025054
R55104 ASIG5V.n1468 ASIG5V.n1467 0.0025054
R55105 ASIG5V.n1500 ASIG5V.n1499 0.0025054
R55106 ASIG5V.n1530 ASIG5V.n1529 0.0025054
R55107 ASIG5V.n1560 ASIG5V.n1559 0.0025054
R55108 ASIG5V.n1590 ASIG5V.n1589 0.0025054
R55109 ASIG5V.n1620 ASIG5V.n1619 0.0025054
R55110 ASIG5V.n1650 ASIG5V.n1649 0.0025054
R55111 ASIG5V.n1467 ASIG5V.n1466 0.0025054
R55112 ASIG5V.n1499 ASIG5V.n1498 0.0025054
R55113 ASIG5V.n1529 ASIG5V.n1528 0.0025054
R55114 ASIG5V.n1559 ASIG5V.n1558 0.0025054
R55115 ASIG5V.n1589 ASIG5V.n1588 0.0025054
R55116 ASIG5V.n1619 ASIG5V.n1618 0.0025054
R55117 ASIG5V.n1649 ASIG5V.n1648 0.0025054
R55118 ASIG5V.n2153 ASIG5V.n2152 0.0025054
R55119 ASIG5V.n7156 ASIG5V.n7155 0.0025054
R55120 ASIG5V.n13277 ASIG5V.n13276 0.0025054
R55121 ASIG5V.n12790 ASIG5V.n12789 0.0025054
R55122 ASIG5V.n10344 ASIG5V.n10343 0.0025054
R55123 ASIG5V.n10368 ASIG5V.n10367 0.0025054
R55124 ASIG5V.n10393 ASIG5V.n10392 0.0025054
R55125 ASIG5V.n10418 ASIG5V.n10417 0.0025054
R55126 ASIG5V.n10443 ASIG5V.n10442 0.0025054
R55127 ASIG5V.n10469 ASIG5V.n10468 0.0025054
R55128 ASIG5V.n10503 ASIG5V.n10502 0.0025054
R55129 ASIG5V.n10534 ASIG5V.n10533 0.0025054
R55130 ASIG5V.n10444 ASIG5V.n10443 0.0025054
R55131 ASIG5V.n10419 ASIG5V.n10418 0.0025054
R55132 ASIG5V.n10394 ASIG5V.n10393 0.0025054
R55133 ASIG5V.n10369 ASIG5V.n10368 0.0025054
R55134 ASIG5V.n10468 ASIG5V.n10467 0.0025054
R55135 ASIG5V.n10502 ASIG5V.n10501 0.0025054
R55136 ASIG5V.n10533 ASIG5V.n10532 0.0025054
R55137 ASIG5V.n1437 ASIG5V.n1436 0.0025054
R55138 ASIG5V.n1978 ASIG5V.n1977 0.0025054
R55139 ASIG5V.n13002 ASIG5V.n13001 0.0025054
R55140 ASIG5V.n13055 ASIG5V.n13054 0.0025054
R55141 ASIG5V.n12969 ASIG5V.n12968 0.0025054
R55142 ASIG5V.n10343 ASIG5V.n10342 0.0025054
R55143 ASIG5V.n9787 ASIG5V.n9786 0.0025054
R55144 ASIG5V.n9829 ASIG5V.n9828 0.0025054
R55145 ASIG5V.n9857 ASIG5V.n9856 0.0025054
R55146 ASIG5V.n9885 ASIG5V.n9884 0.0025054
R55147 ASIG5V.n9913 ASIG5V.n9912 0.0025054
R55148 ASIG5V.n9941 ASIG5V.n9940 0.0025054
R55149 ASIG5V.n10088 ASIG5V.n10087 0.0025054
R55150 ASIG5V.n10118 ASIG5V.n10117 0.0025054
R55151 ASIG5V.n10117 ASIG5V.n10116 0.0025054
R55152 ASIG5V.n10087 ASIG5V.n10086 0.0025054
R55153 ASIG5V.n9940 ASIG5V.n9939 0.0025054
R55154 ASIG5V.n9912 ASIG5V.n9911 0.0025054
R55155 ASIG5V.n9884 ASIG5V.n9883 0.0025054
R55156 ASIG5V.n9856 ASIG5V.n9855 0.0025054
R55157 ASIG5V.n9828 ASIG5V.n9827 0.0025054
R55158 ASIG5V.n9786 ASIG5V.n9785 0.0025054
R55159 ASIG5V.n2268 ASIG5V.n2267 0.0025054
R55160 ASIG5V.n2293 ASIG5V.n2292 0.0025054
R55161 ASIG5V.n2319 ASIG5V.n2318 0.0025054
R55162 ASIG5V.n2344 ASIG5V.n2343 0.0025054
R55163 ASIG5V.n2369 ASIG5V.n2368 0.0025054
R55164 ASIG5V.n2394 ASIG5V.n2393 0.0025054
R55165 ASIG5V.n2419 ASIG5V.n2418 0.0025054
R55166 ASIG5V.n2444 ASIG5V.n2443 0.0025054
R55167 ASIG5V.n2292 ASIG5V.n2291 0.0025054
R55168 ASIG5V.n2318 ASIG5V.n2317 0.0025054
R55169 ASIG5V.n2343 ASIG5V.n2342 0.0025054
R55170 ASIG5V.n2368 ASIG5V.n2367 0.0025054
R55171 ASIG5V.n2393 ASIG5V.n2392 0.0025054
R55172 ASIG5V.n2418 ASIG5V.n2417 0.0025054
R55173 ASIG5V.n2443 ASIG5V.n2442 0.0025054
R55174 ASIG5V.n2267 ASIG5V.n2266 0.0025054
R55175 ASIG5V.n5392 ASIG5V.n5358 0.00243289
R55176 ASIG5V.n5391 ASIG5V.n5390 0.00243289
R55177 ASIG5V.n12958 ASIG5V.n12957 0.00241688
R55178 ASIG5V.n12933 ASIG5V.n12932 0.00241688
R55179 ASIG5V.n12908 ASIG5V.n12907 0.00241688
R55180 ASIG5V.n12879 ASIG5V.n12878 0.00241688
R55181 ASIG5V.n12850 ASIG5V.n12849 0.00241688
R55182 ASIG5V.n12825 ASIG5V.n12824 0.00241688
R55183 ASIG5V.n12796 ASIG5V.n12795 0.00241688
R55184 ASIG5V.n12766 ASIG5V.n12765 0.00241688
R55185 ASIG5V.n12851 ASIG5V.n12850 0.00241688
R55186 ASIG5V.n12880 ASIG5V.n12879 0.00241688
R55187 ASIG5V.n12826 ASIG5V.n12825 0.00241688
R55188 ASIG5V.n13074 ASIG5V.n13073 0.00241688
R55189 ASIG5V.n13102 ASIG5V.n13101 0.00241688
R55190 ASIG5V.n9986 ASIG5V.n9985 0.00241688
R55191 ASIG5V.n10014 ASIG5V.n10013 0.00241688
R55192 ASIG5V.n10042 ASIG5V.n10041 0.00241688
R55193 ASIG5V.n9961 ASIG5V.n9960 0.00241688
R55194 ASIG5V.n13271 ASIG5V.n13270 0.00241688
R55195 ASIG5V.n13300 ASIG5V.n13299 0.00241688
R55196 ASIG5V.n10041 ASIG5V.n10040 0.00241688
R55197 ASIG5V.n10013 ASIG5V.n10012 0.00241688
R55198 ASIG5V.n9962 ASIG5V.n9961 0.00241688
R55199 ASIG5V.n12909 ASIG5V.n12908 0.00241688
R55200 ASIG5V.n9985 ASIG5V.n9984 0.00241688
R55201 ASIG5V.n13023 ASIG5V.n13022 0.00241688
R55202 ASIG5V.n7199 ASIG5V.n7198 0.00241688
R55203 ASIG5V.n13139 ASIG5V.n13138 0.00241688
R55204 ASIG5V.n13170 ASIG5V.n13169 0.00241688
R55205 ASIG5V.n13201 ASIG5V.n13200 0.00241688
R55206 ASIG5V.n13231 ASIG5V.n13230 0.00241688
R55207 ASIG5V.n7162 ASIG5V.n7161 0.00241688
R55208 ASIG5V.n7132 ASIG5V.n7131 0.00241688
R55209 ASIG5V.n13200 ASIG5V.n13199 0.00241688
R55210 ASIG5V.n13169 ASIG5V.n13168 0.00241688
R55211 ASIG5V.n13138 ASIG5V.n13137 0.00241688
R55212 ASIG5V.n13230 ASIG5V.n13229 0.00241688
R55213 ASIG5V.n7163 ASIG5V.n7162 0.00241688
R55214 ASIG5V.n13270 ASIG5V.n13269 0.00241688
R55215 ASIG5V.n12797 ASIG5V.n12796 0.00241688
R55216 ASIG5V.n1997 ASIG5V.n1996 0.00241688
R55217 ASIG5V.n2022 ASIG5V.n2021 0.00241688
R55218 ASIG5V.n2047 ASIG5V.n2046 0.00241688
R55219 ASIG5V.n2072 ASIG5V.n2071 0.00241688
R55220 ASIG5V.n2097 ASIG5V.n2096 0.00241688
R55221 ASIG5V.n2122 ASIG5V.n2121 0.00241688
R55222 ASIG5V.n2147 ASIG5V.n2146 0.00241688
R55223 ASIG5V.n2172 ASIG5V.n2171 0.00241688
R55224 ASIG5V.n2096 ASIG5V.n2095 0.00241688
R55225 ASIG5V.n2071 ASIG5V.n2070 0.00241688
R55226 ASIG5V.n2046 ASIG5V.n2045 0.00241688
R55227 ASIG5V.n2121 ASIG5V.n2120 0.00241688
R55228 ASIG5V.n2146 ASIG5V.n2145 0.00241688
R55229 ASIG5V.n12934 ASIG5V.n12933 0.00241688
R55230 ASIG5V.n13101 ASIG5V.n13100 0.00241688
R55231 ASIG5V.n7200 ASIG5V.n7199 0.00241688
R55232 ASIG5V.n2021 ASIG5V.n2020 0.00241688
R55233 ASIG5V.n1461 ASIG5V.n1460 0.00241688
R55234 ASIG5V.n1493 ASIG5V.n1492 0.00241688
R55235 ASIG5V.n1523 ASIG5V.n1522 0.00241688
R55236 ASIG5V.n1553 ASIG5V.n1552 0.00241688
R55237 ASIG5V.n1583 ASIG5V.n1582 0.00241688
R55238 ASIG5V.n1613 ASIG5V.n1612 0.00241688
R55239 ASIG5V.n1643 ASIG5V.n1642 0.00241688
R55240 ASIG5V.n1673 ASIG5V.n1672 0.00241688
R55241 ASIG5V.n1582 ASIG5V.n1581 0.00241688
R55242 ASIG5V.n1552 ASIG5V.n1551 0.00241688
R55243 ASIG5V.n1522 ASIG5V.n1521 0.00241688
R55244 ASIG5V.n1492 ASIG5V.n1491 0.00241688
R55245 ASIG5V.n1612 ASIG5V.n1611 0.00241688
R55246 ASIG5V.n1642 ASIG5V.n1641 0.00241688
R55247 ASIG5V.n2171 ASIG5V.n2170 0.00241688
R55248 ASIG5V.n12767 ASIG5V.n12766 0.00241688
R55249 ASIG5V.n13299 ASIG5V.n13298 0.00241688
R55250 ASIG5V.n7133 ASIG5V.n7132 0.00241688
R55251 ASIG5V.n1672 ASIG5V.n1671 0.00241688
R55252 ASIG5V.n10362 ASIG5V.n10361 0.00241688
R55253 ASIG5V.n10387 ASIG5V.n10386 0.00241688
R55254 ASIG5V.n10412 ASIG5V.n10411 0.00241688
R55255 ASIG5V.n10437 ASIG5V.n10436 0.00241688
R55256 ASIG5V.n10462 ASIG5V.n10461 0.00241688
R55257 ASIG5V.n10496 ASIG5V.n10495 0.00241688
R55258 ASIG5V.n10527 ASIG5V.n10526 0.00241688
R55259 ASIG5V.n10569 ASIG5V.n10568 0.00241688
R55260 ASIG5V.n10461 ASIG5V.n10460 0.00241688
R55261 ASIG5V.n10436 ASIG5V.n10435 0.00241688
R55262 ASIG5V.n10411 ASIG5V.n10410 0.00241688
R55263 ASIG5V.n10386 ASIG5V.n10385 0.00241688
R55264 ASIG5V.n10495 ASIG5V.n10494 0.00241688
R55265 ASIG5V.n10526 ASIG5V.n10525 0.00241688
R55266 ASIG5V.n10570 ASIG5V.n10569 0.00241688
R55267 ASIG5V.n10361 ASIG5V.n10360 0.00241688
R55268 ASIG5V.n12959 ASIG5V.n12958 0.00241688
R55269 ASIG5V.n13073 ASIG5V.n13072 0.00241688
R55270 ASIG5V.n13022 ASIG5V.n13021 0.00241688
R55271 ASIG5V.n1996 ASIG5V.n1995 0.00241688
R55272 ASIG5V.n1460 ASIG5V.n1459 0.00241688
R55273 ASIG5V.n9822 ASIG5V.n9821 0.00241688
R55274 ASIG5V.n9850 ASIG5V.n9849 0.00241688
R55275 ASIG5V.n9878 ASIG5V.n9877 0.00241688
R55276 ASIG5V.n9906 ASIG5V.n9905 0.00241688
R55277 ASIG5V.n9934 ASIG5V.n9933 0.00241688
R55278 ASIG5V.n10081 ASIG5V.n10080 0.00241688
R55279 ASIG5V.n10111 ASIG5V.n10110 0.00241688
R55280 ASIG5V.n10136 ASIG5V.n10135 0.00241688
R55281 ASIG5V.n9821 ASIG5V.n9820 0.00241688
R55282 ASIG5V.n9933 ASIG5V.n9932 0.00241688
R55283 ASIG5V.n9905 ASIG5V.n9904 0.00241688
R55284 ASIG5V.n9877 ASIG5V.n9876 0.00241688
R55285 ASIG5V.n9849 ASIG5V.n9848 0.00241688
R55286 ASIG5V.n10080 ASIG5V.n10079 0.00241688
R55287 ASIG5V.n10110 ASIG5V.n10109 0.00241688
R55288 ASIG5V.n10135 ASIG5V.n10134 0.00241688
R55289 ASIG5V.n2286 ASIG5V.n2285 0.00241688
R55290 ASIG5V.n2312 ASIG5V.n2311 0.00241688
R55291 ASIG5V.n2337 ASIG5V.n2336 0.00241688
R55292 ASIG5V.n2362 ASIG5V.n2361 0.00241688
R55293 ASIG5V.n2387 ASIG5V.n2386 0.00241688
R55294 ASIG5V.n2412 ASIG5V.n2411 0.00241688
R55295 ASIG5V.n2437 ASIG5V.n2436 0.00241688
R55296 ASIG5V.n2462 ASIG5V.n2461 0.00241688
R55297 ASIG5V.n2285 ASIG5V.n2284 0.00241688
R55298 ASIG5V.n2461 ASIG5V.n2460 0.00241688
R55299 ASIG5V.n2386 ASIG5V.n2385 0.00241688
R55300 ASIG5V.n2361 ASIG5V.n2360 0.00241688
R55301 ASIG5V.n2336 ASIG5V.n2335 0.00241688
R55302 ASIG5V.n2311 ASIG5V.n2310 0.00241688
R55303 ASIG5V.n2411 ASIG5V.n2410 0.00241688
R55304 ASIG5V.n2436 ASIG5V.n2435 0.00241688
R55305 ASIG5V.n4632 ASIG5V.n4631 0.00226856
R55306 ASIG5V.n707 ASIG5V.n706 0.00226856
R55307 ASIG5V.n2494 ASIG5V.n2493 0.00212406
R55308 ASIG5V.n2182 ASIG5V.n2181 0.00212406
R55309 ASIG5V.n10726 ASIG5V.n10725 0.00212406
R55310 ASIG5V.n9386 ASIG5V.n9385 0.002075
R55311 ASIG5V.n9409 ASIG5V.n9408 0.002075
R55312 ASIG5V.n2914 ASIG5V.n2913 0.00194966
R55313 ASIG5V.n4965 ASIG5V.n4931 0.00194966
R55314 ASIG5V.n2743 ASIG5V.n2742 0.00194966
R55315 ASIG5V.n4964 ASIG5V.n4963 0.00194966
R55316 ASIG5V.n12956 ASIG5V.n12955 0.00188565
R55317 ASIG5V.n12931 ASIG5V.n12930 0.00188565
R55318 ASIG5V.n12906 ASIG5V.n12905 0.00188565
R55319 ASIG5V.n12877 ASIG5V.n12876 0.00188565
R55320 ASIG5V.n12848 ASIG5V.n12847 0.00188565
R55321 ASIG5V.n12824 ASIG5V.n12823 0.00188565
R55322 ASIG5V.n12794 ASIG5V.n12793 0.00188565
R55323 ASIG5V.n12764 ASIG5V.n12763 0.00188565
R55324 ASIG5V.n12878 ASIG5V.n12877 0.00188565
R55325 ASIG5V.n12849 ASIG5V.n12848 0.00188565
R55326 ASIG5V.n12823 ASIG5V.n12822 0.00188565
R55327 ASIG5V.n13076 ASIG5V.n13075 0.00188565
R55328 ASIG5V.n13104 ASIG5V.n13103 0.00188565
R55329 ASIG5V.n9988 ASIG5V.n9987 0.00188565
R55330 ASIG5V.n10016 ASIG5V.n10015 0.00188565
R55331 ASIG5V.n10044 ASIG5V.n10043 0.00188565
R55332 ASIG5V.n9959 ASIG5V.n9958 0.00188565
R55333 ASIG5V.n13273 ASIG5V.n13272 0.00188565
R55334 ASIG5V.n13302 ASIG5V.n13301 0.00188565
R55335 ASIG5V.n9960 ASIG5V.n9959 0.00188565
R55336 ASIG5V.n10043 ASIG5V.n10042 0.00188565
R55337 ASIG5V.n10015 ASIG5V.n10014 0.00188565
R55338 ASIG5V.n9987 ASIG5V.n9986 0.00188565
R55339 ASIG5V.n12907 ASIG5V.n12906 0.00188565
R55340 ASIG5V.n13025 ASIG5V.n13024 0.00188565
R55341 ASIG5V.n7197 ASIG5V.n7196 0.00188565
R55342 ASIG5V.n13141 ASIG5V.n13140 0.00188565
R55343 ASIG5V.n13172 ASIG5V.n13171 0.00188565
R55344 ASIG5V.n13203 ASIG5V.n13202 0.00188565
R55345 ASIG5V.n13233 ASIG5V.n13232 0.00188565
R55346 ASIG5V.n7161 ASIG5V.n7160 0.00188565
R55347 ASIG5V.n7130 ASIG5V.n7129 0.00188565
R55348 ASIG5V.n13140 ASIG5V.n13139 0.00188565
R55349 ASIG5V.n13171 ASIG5V.n13170 0.00188565
R55350 ASIG5V.n13202 ASIG5V.n13201 0.00188565
R55351 ASIG5V.n13232 ASIG5V.n13231 0.00188565
R55352 ASIG5V.n13272 ASIG5V.n13271 0.00188565
R55353 ASIG5V.n12795 ASIG5V.n12794 0.00188565
R55354 ASIG5V.n7160 ASIG5V.n7159 0.00188565
R55355 ASIG5V.n1999 ASIG5V.n1998 0.00188565
R55356 ASIG5V.n2024 ASIG5V.n2023 0.00188565
R55357 ASIG5V.n2049 ASIG5V.n2048 0.00188565
R55358 ASIG5V.n2074 ASIG5V.n2073 0.00188565
R55359 ASIG5V.n2099 ASIG5V.n2098 0.00188565
R55360 ASIG5V.n2124 ASIG5V.n2123 0.00188565
R55361 ASIG5V.n2149 ASIG5V.n2148 0.00188565
R55362 ASIG5V.n2174 ASIG5V.n2173 0.00188565
R55363 ASIG5V.n2148 ASIG5V.n2147 0.00188565
R55364 ASIG5V.n2123 ASIG5V.n2122 0.00188565
R55365 ASIG5V.n2098 ASIG5V.n2097 0.00188565
R55366 ASIG5V.n2073 ASIG5V.n2072 0.00188565
R55367 ASIG5V.n2048 ASIG5V.n2047 0.00188565
R55368 ASIG5V.n2023 ASIG5V.n2022 0.00188565
R55369 ASIG5V.n7198 ASIG5V.n7197 0.00188565
R55370 ASIG5V.n13103 ASIG5V.n13102 0.00188565
R55371 ASIG5V.n12932 ASIG5V.n12931 0.00188565
R55372 ASIG5V.n1463 ASIG5V.n1462 0.00188565
R55373 ASIG5V.n1495 ASIG5V.n1494 0.00188565
R55374 ASIG5V.n1525 ASIG5V.n1524 0.00188565
R55375 ASIG5V.n1555 ASIG5V.n1554 0.00188565
R55376 ASIG5V.n1585 ASIG5V.n1584 0.00188565
R55377 ASIG5V.n1615 ASIG5V.n1614 0.00188565
R55378 ASIG5V.n1645 ASIG5V.n1644 0.00188565
R55379 ASIG5V.n1675 ASIG5V.n1674 0.00188565
R55380 ASIG5V.n1494 ASIG5V.n1493 0.00188565
R55381 ASIG5V.n1524 ASIG5V.n1523 0.00188565
R55382 ASIG5V.n1554 ASIG5V.n1553 0.00188565
R55383 ASIG5V.n1584 ASIG5V.n1583 0.00188565
R55384 ASIG5V.n1614 ASIG5V.n1613 0.00188565
R55385 ASIG5V.n1644 ASIG5V.n1643 0.00188565
R55386 ASIG5V.n1674 ASIG5V.n1673 0.00188565
R55387 ASIG5V.n2173 ASIG5V.n2172 0.00188565
R55388 ASIG5V.n7131 ASIG5V.n7130 0.00188565
R55389 ASIG5V.n13301 ASIG5V.n13300 0.00188565
R55390 ASIG5V.n12765 ASIG5V.n12764 0.00188565
R55391 ASIG5V.n10364 ASIG5V.n10363 0.00188565
R55392 ASIG5V.n10389 ASIG5V.n10388 0.00188565
R55393 ASIG5V.n10414 ASIG5V.n10413 0.00188565
R55394 ASIG5V.n10439 ASIG5V.n10438 0.00188565
R55395 ASIG5V.n10464 ASIG5V.n10463 0.00188565
R55396 ASIG5V.n10498 ASIG5V.n10497 0.00188565
R55397 ASIG5V.n10529 ASIG5V.n10528 0.00188565
R55398 ASIG5V.n10572 ASIG5V.n10571 0.00188565
R55399 ASIG5V.n10463 ASIG5V.n10462 0.00188565
R55400 ASIG5V.n10438 ASIG5V.n10437 0.00188565
R55401 ASIG5V.n10413 ASIG5V.n10412 0.00188565
R55402 ASIG5V.n10388 ASIG5V.n10387 0.00188565
R55403 ASIG5V.n10497 ASIG5V.n10496 0.00188565
R55404 ASIG5V.n10528 ASIG5V.n10527 0.00188565
R55405 ASIG5V.n10571 ASIG5V.n10570 0.00188565
R55406 ASIG5V.n1462 ASIG5V.n1461 0.00188565
R55407 ASIG5V.n1998 ASIG5V.n1997 0.00188565
R55408 ASIG5V.n13024 ASIG5V.n13023 0.00188565
R55409 ASIG5V.n13075 ASIG5V.n13074 0.00188565
R55410 ASIG5V.n12957 ASIG5V.n12956 0.00188565
R55411 ASIG5V.n10363 ASIG5V.n10362 0.00188565
R55412 ASIG5V.n9824 ASIG5V.n9823 0.00188565
R55413 ASIG5V.n9852 ASIG5V.n9851 0.00188565
R55414 ASIG5V.n9880 ASIG5V.n9879 0.00188565
R55415 ASIG5V.n9908 ASIG5V.n9907 0.00188565
R55416 ASIG5V.n9936 ASIG5V.n9935 0.00188565
R55417 ASIG5V.n10083 ASIG5V.n10082 0.00188565
R55418 ASIG5V.n10113 ASIG5V.n10112 0.00188565
R55419 ASIG5V.n10138 ASIG5V.n10137 0.00188565
R55420 ASIG5V.n10137 ASIG5V.n10136 0.00188565
R55421 ASIG5V.n10112 ASIG5V.n10111 0.00188565
R55422 ASIG5V.n10082 ASIG5V.n10081 0.00188565
R55423 ASIG5V.n9935 ASIG5V.n9934 0.00188565
R55424 ASIG5V.n9907 ASIG5V.n9906 0.00188565
R55425 ASIG5V.n9879 ASIG5V.n9878 0.00188565
R55426 ASIG5V.n9851 ASIG5V.n9850 0.00188565
R55427 ASIG5V.n9823 ASIG5V.n9822 0.00188565
R55428 ASIG5V.n2288 ASIG5V.n2287 0.00188565
R55429 ASIG5V.n2314 ASIG5V.n2313 0.00188565
R55430 ASIG5V.n2339 ASIG5V.n2338 0.00188565
R55431 ASIG5V.n2364 ASIG5V.n2363 0.00188565
R55432 ASIG5V.n2389 ASIG5V.n2388 0.00188565
R55433 ASIG5V.n2414 ASIG5V.n2413 0.00188565
R55434 ASIG5V.n2439 ASIG5V.n2438 0.00188565
R55435 ASIG5V.n2463 ASIG5V.n2462 0.00188565
R55436 ASIG5V.n2287 ASIG5V.n2286 0.00188565
R55437 ASIG5V.n2313 ASIG5V.n2312 0.00188565
R55438 ASIG5V.n2338 ASIG5V.n2337 0.00188565
R55439 ASIG5V.n2363 ASIG5V.n2362 0.00188565
R55440 ASIG5V.n2388 ASIG5V.n2387 0.00188565
R55441 ASIG5V.n2413 ASIG5V.n2412 0.00188565
R55442 ASIG5V.n2438 ASIG5V.n2437 0.00188565
R55443 ASIG5V.n2464 ASIG5V.n2463 0.00188565
R55444 ASIG5V.n7940 ASIG5V.n7937 0.00187555
R55445 ASIG5V.n11961 ASIG5V.n11960 0.00187555
R55446 ASIG5V.n7939 ASIG5V.n7938 0.00187555
R55447 ASIG5V.n9076 ASIG5V.n9075 0.00187555
R55448 ASIG5V.n12968 ASIG5V.n12967 0.0017971
R55449 ASIG5V.n12953 ASIG5V.n12952 0.0017971
R55450 ASIG5V.n12928 ASIG5V.n12927 0.0017971
R55451 ASIG5V.n12904 ASIG5V.n12903 0.0017971
R55452 ASIG5V.n12875 ASIG5V.n12874 0.0017971
R55453 ASIG5V.n12845 ASIG5V.n12844 0.0017971
R55454 ASIG5V.n12820 ASIG5V.n12819 0.0017971
R55455 ASIG5V.n12791 ASIG5V.n12790 0.0017971
R55456 ASIG5V.n12903 ASIG5V.n12902 0.0017971
R55457 ASIG5V.n12874 ASIG5V.n12873 0.0017971
R55458 ASIG5V.n12846 ASIG5V.n12845 0.0017971
R55459 ASIG5V.n13054 ASIG5V.n13053 0.0017971
R55460 ASIG5V.n13079 ASIG5V.n13078 0.0017971
R55461 ASIG5V.n13107 ASIG5V.n13106 0.0017971
R55462 ASIG5V.n9991 ASIG5V.n9990 0.0017971
R55463 ASIG5V.n10019 ASIG5V.n10018 0.0017971
R55464 ASIG5V.n10046 ASIG5V.n10045 0.0017971
R55465 ASIG5V.n9956 ASIG5V.n9955 0.0017971
R55466 ASIG5V.n13276 ASIG5V.n13275 0.0017971
R55467 ASIG5V.n10047 ASIG5V.n10046 0.0017971
R55468 ASIG5V.n10018 ASIG5V.n10017 0.0017971
R55469 ASIG5V.n9990 ASIG5V.n9989 0.0017971
R55470 ASIG5V.n12929 ASIG5V.n12928 0.0017971
R55471 ASIG5V.n13106 ASIG5V.n13105 0.0017971
R55472 ASIG5V.n13001 ASIG5V.n13000 0.0017971
R55473 ASIG5V.n13028 ASIG5V.n13027 0.0017971
R55474 ASIG5V.n7195 ASIG5V.n7194 0.0017971
R55475 ASIG5V.n13144 ASIG5V.n13143 0.0017971
R55476 ASIG5V.n13175 ASIG5V.n13174 0.0017971
R55477 ASIG5V.n13206 ASIG5V.n13205 0.0017971
R55478 ASIG5V.n13236 ASIG5V.n13235 0.0017971
R55479 ASIG5V.n7157 ASIG5V.n7156 0.0017971
R55480 ASIG5V.n7194 ASIG5V.n7193 0.0017971
R55481 ASIG5V.n13174 ASIG5V.n13173 0.0017971
R55482 ASIG5V.n13143 ASIG5V.n13142 0.0017971
R55483 ASIG5V.n13205 ASIG5V.n13204 0.0017971
R55484 ASIG5V.n12821 ASIG5V.n12820 0.0017971
R55485 ASIG5V.n9957 ASIG5V.n9956 0.0017971
R55486 ASIG5V.n13235 ASIG5V.n13234 0.0017971
R55487 ASIG5V.n1977 ASIG5V.n1976 0.0017971
R55488 ASIG5V.n2002 ASIG5V.n2001 0.0017971
R55489 ASIG5V.n2027 ASIG5V.n2026 0.0017971
R55490 ASIG5V.n2052 ASIG5V.n2051 0.0017971
R55491 ASIG5V.n2077 ASIG5V.n2076 0.0017971
R55492 ASIG5V.n2102 ASIG5V.n2101 0.0017971
R55493 ASIG5V.n2126 ASIG5V.n2125 0.0017971
R55494 ASIG5V.n2152 ASIG5V.n2151 0.0017971
R55495 ASIG5V.n2127 ASIG5V.n2126 0.0017971
R55496 ASIG5V.n2076 ASIG5V.n2075 0.0017971
R55497 ASIG5V.n2051 ASIG5V.n2050 0.0017971
R55498 ASIG5V.n2026 ASIG5V.n2025 0.0017971
R55499 ASIG5V.n2101 ASIG5V.n2100 0.0017971
R55500 ASIG5V.n12954 ASIG5V.n12953 0.0017971
R55501 ASIG5V.n13078 ASIG5V.n13077 0.0017971
R55502 ASIG5V.n13027 ASIG5V.n13026 0.0017971
R55503 ASIG5V.n2001 ASIG5V.n2000 0.0017971
R55504 ASIG5V.n1436 ASIG5V.n1435 0.0017971
R55505 ASIG5V.n1465 ASIG5V.n1464 0.0017971
R55506 ASIG5V.n1498 ASIG5V.n1497 0.0017971
R55507 ASIG5V.n1528 ASIG5V.n1527 0.0017971
R55508 ASIG5V.n1558 ASIG5V.n1557 0.0017971
R55509 ASIG5V.n1588 ASIG5V.n1587 0.0017971
R55510 ASIG5V.n1618 ASIG5V.n1617 0.0017971
R55511 ASIG5V.n1648 ASIG5V.n1647 0.0017971
R55512 ASIG5V.n1466 ASIG5V.n1465 0.0017971
R55513 ASIG5V.n1557 ASIG5V.n1556 0.0017971
R55514 ASIG5V.n1527 ASIG5V.n1526 0.0017971
R55515 ASIG5V.n1497 ASIG5V.n1496 0.0017971
R55516 ASIG5V.n1587 ASIG5V.n1586 0.0017971
R55517 ASIG5V.n1617 ASIG5V.n1616 0.0017971
R55518 ASIG5V.n12792 ASIG5V.n12791 0.0017971
R55519 ASIG5V.n13275 ASIG5V.n13274 0.0017971
R55520 ASIG5V.n7158 ASIG5V.n7157 0.0017971
R55521 ASIG5V.n2151 ASIG5V.n2150 0.0017971
R55522 ASIG5V.n1647 ASIG5V.n1646 0.0017971
R55523 ASIG5V.n10342 ASIG5V.n10341 0.0017971
R55524 ASIG5V.n10367 ASIG5V.n10366 0.0017971
R55525 ASIG5V.n10392 ASIG5V.n10391 0.0017971
R55526 ASIG5V.n10417 ASIG5V.n10416 0.0017971
R55527 ASIG5V.n10442 ASIG5V.n10441 0.0017971
R55528 ASIG5V.n10467 ASIG5V.n10466 0.0017971
R55529 ASIG5V.n10501 ASIG5V.n10500 0.0017971
R55530 ASIG5V.n10531 ASIG5V.n10530 0.0017971
R55531 ASIG5V.n10500 ASIG5V.n10499 0.0017971
R55532 ASIG5V.n10441 ASIG5V.n10440 0.0017971
R55533 ASIG5V.n10416 ASIG5V.n10415 0.0017971
R55534 ASIG5V.n10391 ASIG5V.n10390 0.0017971
R55535 ASIG5V.n10366 ASIG5V.n10365 0.0017971
R55536 ASIG5V.n10466 ASIG5V.n10465 0.0017971
R55537 ASIG5V.n10532 ASIG5V.n10531 0.0017971
R55538 ASIG5V.n10341 ASIG5V.n10340 0.0017971
R55539 ASIG5V.n12967 ASIG5V.n12966 0.0017971
R55540 ASIG5V.n13053 ASIG5V.n13052 0.0017971
R55541 ASIG5V.n13000 ASIG5V.n12999 0.0017971
R55542 ASIG5V.n1976 ASIG5V.n1975 0.0017971
R55543 ASIG5V.n1435 ASIG5V.n1434 0.0017971
R55544 ASIG5V.n9784 ASIG5V.n9783 0.0017971
R55545 ASIG5V.n9827 ASIG5V.n9826 0.0017971
R55546 ASIG5V.n9855 ASIG5V.n9854 0.0017971
R55547 ASIG5V.n9883 ASIG5V.n9882 0.0017971
R55548 ASIG5V.n9911 ASIG5V.n9910 0.0017971
R55549 ASIG5V.n9939 ASIG5V.n9938 0.0017971
R55550 ASIG5V.n10086 ASIG5V.n10085 0.0017971
R55551 ASIG5V.n10116 ASIG5V.n10115 0.0017971
R55552 ASIG5V.n9910 ASIG5V.n9909 0.0017971
R55553 ASIG5V.n9882 ASIG5V.n9881 0.0017971
R55554 ASIG5V.n9854 ASIG5V.n9853 0.0017971
R55555 ASIG5V.n9826 ASIG5V.n9825 0.0017971
R55556 ASIG5V.n9938 ASIG5V.n9937 0.0017971
R55557 ASIG5V.n10085 ASIG5V.n10084 0.0017971
R55558 ASIG5V.n10115 ASIG5V.n10114 0.0017971
R55559 ASIG5V.n9785 ASIG5V.n9784 0.0017971
R55560 ASIG5V.n2266 ASIG5V.n2265 0.0017971
R55561 ASIG5V.n2291 ASIG5V.n2290 0.0017971
R55562 ASIG5V.n2317 ASIG5V.n2316 0.0017971
R55563 ASIG5V.n2342 ASIG5V.n2341 0.0017971
R55564 ASIG5V.n2367 ASIG5V.n2366 0.0017971
R55565 ASIG5V.n2392 ASIG5V.n2391 0.0017971
R55566 ASIG5V.n2417 ASIG5V.n2416 0.0017971
R55567 ASIG5V.n2442 ASIG5V.n2441 0.0017971
R55568 ASIG5V.n2265 ASIG5V.n2264 0.0017971
R55569 ASIG5V.n2366 ASIG5V.n2365 0.0017971
R55570 ASIG5V.n2341 ASIG5V.n2340 0.0017971
R55571 ASIG5V.n2316 ASIG5V.n2315 0.0017971
R55572 ASIG5V.n2290 ASIG5V.n2289 0.0017971
R55573 ASIG5V.n2391 ASIG5V.n2390 0.0017971
R55574 ASIG5V.n2416 ASIG5V.n2415 0.0017971
R55575 ASIG5V.n2441 ASIG5V.n2440 0.0017971
R55576 ASIG5V.n980 ASIG5V.n979 0.001625
R55577 ASIG5V.n12976 ASIG5V.n12975 0.00161999
R55578 ASIG5V.n12964 ASIG5V.n12963 0.00161999
R55579 ASIG5V.n12945 ASIG5V.n12944 0.00161999
R55580 ASIG5V.n12939 ASIG5V.n12938 0.00161999
R55581 ASIG5V.n12920 ASIG5V.n12919 0.00161999
R55582 ASIG5V.n12914 ASIG5V.n12913 0.00161999
R55583 ASIG5V.n12896 ASIG5V.n12895 0.00161999
R55584 ASIG5V.n12886 ASIG5V.n12885 0.00161999
R55585 ASIG5V.n12867 ASIG5V.n12866 0.00161999
R55586 ASIG5V.n12857 ASIG5V.n12856 0.00161999
R55587 ASIG5V.n12837 ASIG5V.n12836 0.00161999
R55588 ASIG5V.n12831 ASIG5V.n12830 0.00161999
R55589 ASIG5V.n12812 ASIG5V.n12811 0.00161999
R55590 ASIG5V.n12802 ASIG5V.n12801 0.00161999
R55591 ASIG5V.n12783 ASIG5V.n12782 0.00161999
R55592 ASIG5V.n12772 ASIG5V.n12771 0.00161999
R55593 ASIG5V.n12885 ASIG5V.n12884 0.00161999
R55594 ASIG5V.n12856 ASIG5V.n12855 0.00161999
R55595 ASIG5V.n12866 ASIG5V.n12865 0.00161999
R55596 ASIG5V.n12895 ASIG5V.n12894 0.00161999
R55597 ASIG5V.n12838 ASIG5V.n12837 0.00161999
R55598 ASIG5V.n12832 ASIG5V.n12831 0.00161999
R55599 ASIG5V.n13062 ASIG5V.n13061 0.00161999
R55600 ASIG5V.n13068 ASIG5V.n13067 0.00161999
R55601 ASIG5V.n13087 ASIG5V.n13086 0.00161999
R55602 ASIG5V.n13096 ASIG5V.n13095 0.00161999
R55603 ASIG5V.n13115 ASIG5V.n13114 0.00161999
R55604 ASIG5V.n9980 ASIG5V.n9979 0.00161999
R55605 ASIG5V.n9999 ASIG5V.n9998 0.00161999
R55606 ASIG5V.n10008 ASIG5V.n10007 0.00161999
R55607 ASIG5V.n10027 ASIG5V.n10026 0.00161999
R55608 ASIG5V.n10036 ASIG5V.n10035 0.00161999
R55609 ASIG5V.n10055 ASIG5V.n10054 0.00161999
R55610 ASIG5V.n9967 ASIG5V.n9966 0.00161999
R55611 ASIG5V.n9948 ASIG5V.n399 0.00161999
R55612 ASIG5V.n13265 ASIG5V.n13264 0.00161999
R55613 ASIG5V.n13284 ASIG5V.n13283 0.00161999
R55614 ASIG5V.n13294 ASIG5V.n13293 0.00161999
R55615 ASIG5V.n10054 ASIG5V.n10053 0.00161999
R55616 ASIG5V.n10026 ASIG5V.n10025 0.00161999
R55617 ASIG5V.n9998 ASIG5V.n9997 0.00161999
R55618 ASIG5V.n10035 ASIG5V.n10034 0.00161999
R55619 ASIG5V.n10007 ASIG5V.n10006 0.00161999
R55620 ASIG5V.n9968 ASIG5V.n9967 0.00161999
R55621 ASIG5V.n13114 ASIG5V.n13113 0.00161999
R55622 ASIG5V.n12921 ASIG5V.n12920 0.00161999
R55623 ASIG5V.n12915 ASIG5V.n12914 0.00161999
R55624 ASIG5V.n9979 ASIG5V.n7184 0.00161999
R55625 ASIG5V.n13009 ASIG5V.n13008 0.00161999
R55626 ASIG5V.n13017 ASIG5V.n13016 0.00161999
R55627 ASIG5V.n13036 ASIG5V.n13035 0.00161999
R55628 ASIG5V.n7205 ASIG5V.n7204 0.00161999
R55629 ASIG5V.n7187 ASIG5V.n7186 0.00161999
R55630 ASIG5V.n13132 ASIG5V.n13131 0.00161999
R55631 ASIG5V.n13152 ASIG5V.n13151 0.00161999
R55632 ASIG5V.n13164 ASIG5V.n13163 0.00161999
R55633 ASIG5V.n13183 ASIG5V.n13182 0.00161999
R55634 ASIG5V.n13195 ASIG5V.n13194 0.00161999
R55635 ASIG5V.n13214 ASIG5V.n13213 0.00161999
R55636 ASIG5V.n13225 ASIG5V.n13224 0.00161999
R55637 ASIG5V.n13244 ASIG5V.n13243 0.00161999
R55638 ASIG5V.n7168 ASIG5V.n7167 0.00161999
R55639 ASIG5V.n7149 ASIG5V.n7148 0.00161999
R55640 ASIG5V.n7138 ASIG5V.n7137 0.00161999
R55641 ASIG5V.n13133 ASIG5V.n13132 0.00161999
R55642 ASIG5V.n13151 ASIG5V.n13150 0.00161999
R55643 ASIG5V.n13182 ASIG5V.n13181 0.00161999
R55644 ASIG5V.n13213 ASIG5V.n13212 0.00161999
R55645 ASIG5V.n13194 ASIG5V.n13193 0.00161999
R55646 ASIG5V.n13163 ASIG5V.n13162 0.00161999
R55647 ASIG5V.n7186 ASIG5V.n7182 0.00161999
R55648 ASIG5V.n13224 ASIG5V.n13223 0.00161999
R55649 ASIG5V.n13243 ASIG5V.n13242 0.00161999
R55650 ASIG5V.n9949 ASIG5V.n9948 0.00161999
R55651 ASIG5V.n12813 ASIG5V.n12812 0.00161999
R55652 ASIG5V.n12803 ASIG5V.n12802 0.00161999
R55653 ASIG5V.n13264 ASIG5V.n13263 0.00161999
R55654 ASIG5V.n7169 ASIG5V.n7168 0.00161999
R55655 ASIG5V.n1985 ASIG5V.n1984 0.00161999
R55656 ASIG5V.n1991 ASIG5V.n1990 0.00161999
R55657 ASIG5V.n2010 ASIG5V.n2009 0.00161999
R55658 ASIG5V.n2016 ASIG5V.n2015 0.00161999
R55659 ASIG5V.n2035 ASIG5V.n2034 0.00161999
R55660 ASIG5V.n2041 ASIG5V.n2040 0.00161999
R55661 ASIG5V.n2060 ASIG5V.n2059 0.00161999
R55662 ASIG5V.n2066 ASIG5V.n2065 0.00161999
R55663 ASIG5V.n2085 ASIG5V.n2084 0.00161999
R55664 ASIG5V.n2091 ASIG5V.n2090 0.00161999
R55665 ASIG5V.n2110 ASIG5V.n2109 0.00161999
R55666 ASIG5V.n2116 ASIG5V.n2115 0.00161999
R55667 ASIG5V.n2135 ASIG5V.n2134 0.00161999
R55668 ASIG5V.n2141 ASIG5V.n2140 0.00161999
R55669 ASIG5V.n2160 ASIG5V.n2159 0.00161999
R55670 ASIG5V.n2166 ASIG5V.n2165 0.00161999
R55671 ASIG5V.n2134 ASIG5V.n2133 0.00161999
R55672 ASIG5V.n2109 ASIG5V.n2108 0.00161999
R55673 ASIG5V.n2084 ASIG5V.n2083 0.00161999
R55674 ASIG5V.n2059 ASIG5V.n2058 0.00161999
R55675 ASIG5V.n2034 ASIG5V.n2033 0.00161999
R55676 ASIG5V.n2090 ASIG5V.n2089 0.00161999
R55677 ASIG5V.n2065 ASIG5V.n2064 0.00161999
R55678 ASIG5V.n2040 ASIG5V.n2039 0.00161999
R55679 ASIG5V.n2115 ASIG5V.n2114 0.00161999
R55680 ASIG5V.n2140 ASIG5V.n2139 0.00161999
R55681 ASIG5V.n2009 ASIG5V.n2008 0.00161999
R55682 ASIG5V.n13035 ASIG5V.n13034 0.00161999
R55683 ASIG5V.n13086 ASIG5V.n13085 0.00161999
R55684 ASIG5V.n12946 ASIG5V.n12945 0.00161999
R55685 ASIG5V.n12940 ASIG5V.n12939 0.00161999
R55686 ASIG5V.n13095 ASIG5V.n13094 0.00161999
R55687 ASIG5V.n7206 ASIG5V.n7205 0.00161999
R55688 ASIG5V.n2015 ASIG5V.n2014 0.00161999
R55689 ASIG5V.n1444 ASIG5V.n1443 0.00161999
R55690 ASIG5V.n1455 ASIG5V.n1454 0.00161999
R55691 ASIG5V.n1473 ASIG5V.n1472 0.00161999
R55692 ASIG5V.n1486 ASIG5V.n1485 0.00161999
R55693 ASIG5V.n1506 ASIG5V.n1505 0.00161999
R55694 ASIG5V.n1517 ASIG5V.n1516 0.00161999
R55695 ASIG5V.n1536 ASIG5V.n1535 0.00161999
R55696 ASIG5V.n1547 ASIG5V.n1546 0.00161999
R55697 ASIG5V.n1566 ASIG5V.n1565 0.00161999
R55698 ASIG5V.n1577 ASIG5V.n1576 0.00161999
R55699 ASIG5V.n1596 ASIG5V.n1595 0.00161999
R55700 ASIG5V.n1607 ASIG5V.n1606 0.00161999
R55701 ASIG5V.n1626 ASIG5V.n1625 0.00161999
R55702 ASIG5V.n1637 ASIG5V.n1636 0.00161999
R55703 ASIG5V.n1656 ASIG5V.n1655 0.00161999
R55704 ASIG5V.n1667 ASIG5V.n1666 0.00161999
R55705 ASIG5V.n1487 ASIG5V.n1486 0.00161999
R55706 ASIG5V.n1505 ASIG5V.n1504 0.00161999
R55707 ASIG5V.n1535 ASIG5V.n1534 0.00161999
R55708 ASIG5V.n1565 ASIG5V.n1564 0.00161999
R55709 ASIG5V.n1595 ASIG5V.n1594 0.00161999
R55710 ASIG5V.n1625 ASIG5V.n1624 0.00161999
R55711 ASIG5V.n1576 ASIG5V.n1575 0.00161999
R55712 ASIG5V.n1546 ASIG5V.n1545 0.00161999
R55713 ASIG5V.n1516 ASIG5V.n1515 0.00161999
R55714 ASIG5V.n1474 ASIG5V.n1473 0.00161999
R55715 ASIG5V.n1606 ASIG5V.n1605 0.00161999
R55716 ASIG5V.n1636 ASIG5V.n1635 0.00161999
R55717 ASIG5V.n1655 ASIG5V.n1654 0.00161999
R55718 ASIG5V.n2159 ASIG5V.n2158 0.00161999
R55719 ASIG5V.n7150 ASIG5V.n7149 0.00161999
R55720 ASIG5V.n7139 ASIG5V.n7138 0.00161999
R55721 ASIG5V.n2165 ASIG5V.n2164 0.00161999
R55722 ASIG5V.n1666 ASIG5V.n1665 0.00161999
R55723 ASIG5V.n12773 ASIG5V.n12772 0.00161999
R55724 ASIG5V.n13293 ASIG5V.n13292 0.00161999
R55725 ASIG5V.n12784 ASIG5V.n12783 0.00161999
R55726 ASIG5V.n13283 ASIG5V.n13282 0.00161999
R55727 ASIG5V.n10350 ASIG5V.n10349 0.00161999
R55728 ASIG5V.n10356 ASIG5V.n10355 0.00161999
R55729 ASIG5V.n10375 ASIG5V.n10374 0.00161999
R55730 ASIG5V.n10381 ASIG5V.n10380 0.00161999
R55731 ASIG5V.n10400 ASIG5V.n10399 0.00161999
R55732 ASIG5V.n10406 ASIG5V.n10405 0.00161999
R55733 ASIG5V.n10425 ASIG5V.n10424 0.00161999
R55734 ASIG5V.n10431 ASIG5V.n10430 0.00161999
R55735 ASIG5V.n10450 ASIG5V.n10449 0.00161999
R55736 ASIG5V.n10456 ASIG5V.n10455 0.00161999
R55737 ASIG5V.n10475 ASIG5V.n10474 0.00161999
R55738 ASIG5V.n10490 ASIG5V.n10489 0.00161999
R55739 ASIG5V.n10509 ASIG5V.n10508 0.00161999
R55740 ASIG5V.n10521 ASIG5V.n10520 0.00161999
R55741 ASIG5V.n10539 ASIG5V.n10538 0.00161999
R55742 ASIG5V.n10564 ASIG5V.n10563 0.00161999
R55743 ASIG5V.n10449 ASIG5V.n10448 0.00161999
R55744 ASIG5V.n10455 ASIG5V.n10454 0.00161999
R55745 ASIG5V.n10424 ASIG5V.n10423 0.00161999
R55746 ASIG5V.n10430 ASIG5V.n10429 0.00161999
R55747 ASIG5V.n10399 ASIG5V.n10398 0.00161999
R55748 ASIG5V.n10405 ASIG5V.n10404 0.00161999
R55749 ASIG5V.n10374 ASIG5V.n10373 0.00161999
R55750 ASIG5V.n10380 ASIG5V.n10379 0.00161999
R55751 ASIG5V.n10489 ASIG5V.n10488 0.00161999
R55752 ASIG5V.n10474 ASIG5V.n10473 0.00161999
R55753 ASIG5V.n10508 ASIG5V.n10507 0.00161999
R55754 ASIG5V.n10520 ASIG5V.n10519 0.00161999
R55755 ASIG5V.n10563 ASIG5V.n10562 0.00161999
R55756 ASIG5V.n10540 ASIG5V.n10539 0.00161999
R55757 ASIG5V.n1443 ASIG5V.n1442 0.00161999
R55758 ASIG5V.n1454 ASIG5V.n1453 0.00161999
R55759 ASIG5V.n10355 ASIG5V.n10354 0.00161999
R55760 ASIG5V.n12965 ASIG5V.n12964 0.00161999
R55761 ASIG5V.n13067 ASIG5V.n13066 0.00161999
R55762 ASIG5V.n13016 ASIG5V.n13015 0.00161999
R55763 ASIG5V.n1990 ASIG5V.n1989 0.00161999
R55764 ASIG5V.n1984 ASIG5V.n1983 0.00161999
R55765 ASIG5V.n13008 ASIG5V.n13007 0.00161999
R55766 ASIG5V.n13061 ASIG5V.n13060 0.00161999
R55767 ASIG5V.n12975 ASIG5V.n12974 0.00161999
R55768 ASIG5V.n10349 ASIG5V.n10348 0.00161999
R55769 ASIG5V.n9792 ASIG5V.n9791 0.00161999
R55770 ASIG5V.n9816 ASIG5V.n9815 0.00161999
R55771 ASIG5V.n9835 ASIG5V.n9834 0.00161999
R55772 ASIG5V.n9844 ASIG5V.n9843 0.00161999
R55773 ASIG5V.n9863 ASIG5V.n9862 0.00161999
R55774 ASIG5V.n9872 ASIG5V.n9871 0.00161999
R55775 ASIG5V.n9891 ASIG5V.n9890 0.00161999
R55776 ASIG5V.n9900 ASIG5V.n9899 0.00161999
R55777 ASIG5V.n9919 ASIG5V.n9918 0.00161999
R55778 ASIG5V.n9928 ASIG5V.n9927 0.00161999
R55779 ASIG5V.n9947 ASIG5V.n9946 0.00161999
R55780 ASIG5V.n10075 ASIG5V.n10074 0.00161999
R55781 ASIG5V.n10094 ASIG5V.n10093 0.00161999
R55782 ASIG5V.n10105 ASIG5V.n10104 0.00161999
R55783 ASIG5V.n10124 ASIG5V.n10123 0.00161999
R55784 ASIG5V.n10130 ASIG5V.n10129 0.00161999
R55785 ASIG5V.n10123 ASIG5V.n10122 0.00161999
R55786 ASIG5V.n10093 ASIG5V.n10092 0.00161999
R55787 ASIG5V.n9946 ASIG5V.n9945 0.00161999
R55788 ASIG5V.n9918 ASIG5V.n9917 0.00161999
R55789 ASIG5V.n9890 ASIG5V.n9889 0.00161999
R55790 ASIG5V.n9862 ASIG5V.n9861 0.00161999
R55791 ASIG5V.n9834 ASIG5V.n9833 0.00161999
R55792 ASIG5V.n9815 ASIG5V.n9814 0.00161999
R55793 ASIG5V.n9927 ASIG5V.n9926 0.00161999
R55794 ASIG5V.n9899 ASIG5V.n9898 0.00161999
R55795 ASIG5V.n9871 ASIG5V.n9870 0.00161999
R55796 ASIG5V.n9843 ASIG5V.n9842 0.00161999
R55797 ASIG5V.n10074 ASIG5V.n10073 0.00161999
R55798 ASIG5V.n10104 ASIG5V.n10103 0.00161999
R55799 ASIG5V.n10129 ASIG5V.n10128 0.00161999
R55800 ASIG5V.n9793 ASIG5V.n9792 0.00161999
R55801 ASIG5V.n2274 ASIG5V.n2273 0.00161999
R55802 ASIG5V.n2280 ASIG5V.n2279 0.00161999
R55803 ASIG5V.n2299 ASIG5V.n2298 0.00161999
R55804 ASIG5V.n2306 ASIG5V.n2305 0.00161999
R55805 ASIG5V.n2325 ASIG5V.n2324 0.00161999
R55806 ASIG5V.n2331 ASIG5V.n2330 0.00161999
R55807 ASIG5V.n2350 ASIG5V.n2349 0.00161999
R55808 ASIG5V.n2356 ASIG5V.n2355 0.00161999
R55809 ASIG5V.n2375 ASIG5V.n2374 0.00161999
R55810 ASIG5V.n2381 ASIG5V.n2380 0.00161999
R55811 ASIG5V.n2400 ASIG5V.n2399 0.00161999
R55812 ASIG5V.n2406 ASIG5V.n2405 0.00161999
R55813 ASIG5V.n2425 ASIG5V.n2424 0.00161999
R55814 ASIG5V.n2431 ASIG5V.n2430 0.00161999
R55815 ASIG5V.n2450 ASIG5V.n2449 0.00161999
R55816 ASIG5V.n2456 ASIG5V.n2455 0.00161999
R55817 ASIG5V.n2298 ASIG5V.n2297 0.00161999
R55818 ASIG5V.n2324 ASIG5V.n2323 0.00161999
R55819 ASIG5V.n2349 ASIG5V.n2348 0.00161999
R55820 ASIG5V.n2374 ASIG5V.n2373 0.00161999
R55821 ASIG5V.n2399 ASIG5V.n2398 0.00161999
R55822 ASIG5V.n2424 ASIG5V.n2423 0.00161999
R55823 ASIG5V.n2449 ASIG5V.n2448 0.00161999
R55824 ASIG5V.n2279 ASIG5V.n2278 0.00161999
R55825 ASIG5V.n2380 ASIG5V.n2379 0.00161999
R55826 ASIG5V.n2355 ASIG5V.n2354 0.00161999
R55827 ASIG5V.n2330 ASIG5V.n2329 0.00161999
R55828 ASIG5V.n2305 ASIG5V.n2304 0.00161999
R55829 ASIG5V.n2405 ASIG5V.n2404 0.00161999
R55830 ASIG5V.n2430 ASIG5V.n2429 0.00161999
R55831 ASIG5V.n2455 ASIG5V.n2454 0.00161999
R55832 ASIG5V.n2273 ASIG5V.n2272 0.00161999
R55833 ASIG5V.n13349 ASIG5V.n13348 0.00158271
R55834 ASIG5V.n7516 ASIG5V.n7515 0.00158271
R55835 ASIG5V.n12762 ASIG5V.n12761 0.00158271
R55836 ASIG5V.n10728 ASIG5V.n10727 0.00158271
R55837 ASIG5V.n6934 ASIG5V.n6930 0.00148253
R55838 ASIG5V.n6933 ASIG5V.n6932 0.00148253
R55839 ASIG5V.n7518 ASIG5V.n7436 0.00146644
R55840 ASIG5V.n12302 ASIG5V.n12268 0.00146644
R55841 ASIG5V.n7517 ASIG5V.n7468 0.00146644
R55842 ASIG5V.n12301 ASIG5V.n12300 0.00146644
R55843 ASIG5V.n747 ASIG5V.n746 0.0011898
R55844 ASIG5V.n9121 ASIG5V.n9120 0.0011898
R55845 ASIG5V.n9120 ASIG5V.n9119 0.0011898
R55846 ASIG5V.n746 ASIG5V.n745 0.0011898
R55847 ASIG5V.n1022 ASIG5V.n1021 0.001175
R55848 ASIG5V.n3298 ASIG5V.n3297 0.00108952
R55849 ASIG5V.n726 ASIG5V.n725 0.00108952
R55850 ASIG5V.n2466 ASIG5V.n2465 0.00104135
R55851 ASIG5V.n7045 ASIG5V.n7044 0.00104135
R55852 ASIG5V.n10746 ASIG5V.n10745 0.00104135
R55853 ASIG5V.n7047 ASIG5V.n6965 0.000983221
R55854 ASIG5V.n11665 ASIG5V.n11664 0.000983221
R55855 ASIG5V.n7046 ASIG5V.n6997 0.000983221
R55856 ASIG5V.n10926 ASIG5V.n10925 0.000983221
R55857 ASIG5V.n4285 ASIG5V.n4282 0.00087964
R55858 ASIG5V.n5801 ASIG5V.n5797 0.00087964
R55859 ASIG5V.n11317 ASIG5V.n11315 0.00087964
R55860 ASIG5V.n3038 ASIG5V.n3036 0.000876579
R55861 ASIG5V.n12162 ASIG5V.n12159 0.000876579
R55862 ASIG5V.n7636 ASIG5V.n7633 0.000864332
R55863 ASIG5V.n5808 ASIG5V.n5804 0.000858209
R55864 ASIG5V.n13616 ASIG5V.n13612 0.000858209
R55865 ASIG5V.n621 ASIG5V.n514 0.000855147
R55866 ASIG5V.n627 ASIG5V.n622 0.000855147
R55867 ASIG5V.n741 ASIG5V.n628 0.000855147
R55868 ASIG5V.n744 ASIG5V.n742 0.000855147
R55869 ASIG5V.n7063 ASIG5V.n7059 0.000852086
R55870 ASIG5V.n13495 ASIG5V.n13371 0.000852086
R55871 ASIG5V.n5676 ASIG5V.n5671 0.000845963
R55872 ASIG5V.n13367 ASIG5V.n13364 0.000845963
R55873 ASIG5V.n4854 ASIG5V.n4852 0.000839839
R55874 ASIG5V.n12653 ASIG5V.n12651 0.000836778
R55875 ASIG5V.n12432 ASIG5V.n12430 0.000833716
R55876 ASIG5V.n3481 ASIG5V.n3479 0.000827593
R55877 ASIG5V.n4375 ASIG5V.n4287 0.000827593
R55878 ASIG5V.n11839 ASIG5V.n11836 0.000827593
R55879 ASIG5V.n3745 ASIG5V.n3742 0.00082147
R55880 ASIG5V.n11674 ASIG5V.n11672 0.00082147
R55881 ASIG5V.n4277 ASIG5V.n4164 0.000818408
R55882 ASIG5V.n4446 ASIG5V.n4443 0.000815346
R55883 ASIG5V.n12662 ASIG5V.n12659 0.000815346
R55884 ASIG5V.n11831 ASIG5V.n11828 0.000815346
R55885 ASIG5V.n5151 ASIG5V.n5148 0.000809223
R55886 ASIG5V.n11313 ASIG5V.n11311 0.000806161
R55887 ASIG5V.n11157 ASIG5V.n11154 0.000806161
R55888 ASIG5V.n5972 ASIG5V.n5860 0.0008031
R55889 ASIG5V.n3251 ASIG5V.n3139 0.000796977
R55890 ASIG5V.n6787 ASIG5V.n6784 0.000796977
R55891 ASIG5V.n3104 ASIG5V.n3040 0.000793915
R55892 ASIG5V.n5455 ASIG5V.n5452 0.000790853
R55893 ASIG5V.n13358 ASIG5V.n13353 0.000790853
R55894 ASIG5V.n12581 ASIG5V.n12435 0.000790853
R55895 ASIG5V.n7990 ASIG5V.n7986 0.00078473
R55896 ASIG5V.n11416 ASIG5V.n11324 0.000781669
R55897 ASIG5V.n9118 ASIG5V.n9117 0.000781669
R55898 ASIG5V.n9116 ASIG5V.n8982 0.000781669
R55899 ASIG5V.n8981 ASIG5V.n8976 0.000781669
R55900 ASIG5V.n8975 ASIG5V.n8880 0.000781669
R55901 ASIG5V.n3623 ASIG5V.n3558 0.000778607
R55902 ASIG5V.n3257 ASIG5V.n3255 0.000772484
R55903 ASIG5V.n12085 ASIG5V.n12082 0.000772484
R55904 ASIG5V.n12006 ASIG5V.n12004 0.000772484
R55905 ASIG5V.n12425 ASIG5V.n12420 0.000769422
R55906 ASIG5V.n12157 ASIG5V.n12154 0.000769422
R55907 ASIG5V ASIG5V.n13621 0.00076636
R55908 ASIG5V.n4096 ASIG5V.n4012 0.000763299
R55909 ASIG5V.n4566 ASIG5V.n4563 0.000760237
R55910 ASIG5V.n12668 ASIG5V.n12665 0.000760237
R55911 ASIG5V.n11760 ASIG5V.n11676 0.000760237
R55912 ASIG5V.n11104 ASIG5V.n11102 0.000760237
R55913 ASIG5V.n12303 ASIG5V.n12238 0.000751052
R55914 ASIG5V.n3032 ASIG5V.n2915 0.000747991
R55915 ASIG5V.n4966 ASIG5V.n4901 0.000747991
R55916 ASIG5V.n6156 ASIG5V.n6152 0.000747991
R55917 ASIG5V.n6556 ASIG5V.n6552 0.000747991
R55918 ASIG5V.n7979 ASIG5V.n7941 0.000741868
R55919 ASIG5V.n11668 ASIG5V.n11666 0.000738806
R55920 ASIG5V.n5448 ASIG5V.n5445 0.000735744
R55921 ASIG5V.n7278 ASIG5V.n7274 0.000735744
R55922 ASIG5V.n11926 ASIG5V.n11841 0.000729621
R55923 ASIG5V.n11098 ASIG5V.n9433 0.000729621
R55924 ASIG5V.n7823 ASIG5V.n7640 0.00072656
R55925 ASIG5V.n11488 ASIG5V.n11486 0.00072656
R55926 ASIG5V.n2821 ASIG5V.n1068 0.000723498
R55927 ASIG5V.n3740 ASIG5V.n3737 0.000723498
R55928 ASIG5V.n4009 ASIG5V.n4007 0.000723498
R55929 ASIG5V.n11492 ASIG5V.n11490 0.000723498
R55930 ASIG5V.n3296 ASIG5V.n3259 0.000717375
R55931 ASIG5V.n3299 ASIG5V.n3296 0.000717375
R55932 ASIG5V.n3477 ASIG5V.n3475 0.000717375
R55933 ASIG5V.n11997 ASIG5V.n11962 0.000717375
R55934 ASIG5V.n7052 ASIG5V.n7048 0.000714313
R55935 ASIG5V.n12352 ASIG5V.n12318 0.000714313
R55936 ASIG5V.n2823 ASIG5V.n2821 0.000711251
R55937 ASIG5V.n12318 ASIG5V.n12315 0.000711251
R55938 ASIG5V.n4571 ASIG5V.n4568 0.000705128
R55939 ASIG5V.n12758 ASIG5V.n12757 0.000705128
R55940 ASIG5V.n12001 ASIG5V.n11999 0.000705128
R55941 ASIG5V.n11100 ASIG5V.n11098 0.000705128
R55942 ASIG5V.n3896 ASIG5V.n3833 0.000702067
R55943 ASIG5V.n7281 ASIG5V.n7278 0.000699005
R55944 ASIG5V.n12313 ASIG5V.n12310 0.000695943
R55945 ASIG5V.n2880 ASIG5V.n2825 0.000692882
R55946 ASIG5V.n5145 ASIG5V.n5142 0.000692882
R55947 ASIG5V.n6163 ASIG5V.n6159 0.000692882
R55948 ASIG5V.n6935 ASIG5V.n6928 0.000692882
R55949 ASIG5V.n6769 ASIG5V.n6657 0.000692882
R55950 ASIG5V.n6159 ASIG5V.n6156 0.000686759
R55951 ASIG5V.n11631 ASIG5V.n11492 0.000683697
R55952 ASIG5V.n5398 ASIG5V.n5393 0.000680635
R55953 ASIG5V.n7285 ASIG5V.n7281 0.000680635
R55954 ASIG5V.n7626 ASIG5V.n7519 0.000680635
R55955 ASIG5V.n4568 ASIG5V.n4566 0.000674512
R55956 ASIG5V.n4633 ASIG5V.n4630 0.000674512
R55957 ASIG5V.n4849 ASIG5V.n4847 0.000674512
R55958 ASIG5V.n11102 ASIG5V.n11100 0.000674512
R55959 ASIG5V.n5142 ASIG5V.n4971 0.00067145
R55960 ASIG5V.n5393 ASIG5V.n5328 0.00067145
R55961 ASIG5V.n6331 ASIG5V.n6326 0.00067145
R55962 ASIG5V.n7123 ASIG5V.n7066 0.00067145
R55963 ASIG5V.n2825 ASIG5V.n2823 0.000668389
R55964 ASIG5V.n3899 ASIG5V.n3896 0.000668389
R55965 ASIG5V.n12315 ASIG5V.n12313 0.000668389
R55966 ASIG5V.n11666 ASIG5V.n11634 0.000668389
R55967 ASIG5V.n7056 ASIG5V.n7052 0.000665327
R55968 ASIG5V.n3259 ASIG5V.n3257 0.000662266
R55969 ASIG5V.n3331 ASIG5V.n3299 0.000662266
R55970 ASIG5V.n8120 ASIG5V.n7993 0.000662266
R55971 ASIG5V.n12757 ASIG5V.n12752 0.000662266
R55972 ASIG5V.n12004 ASIG5V.n12001 0.000662266
R55973 ASIG5V.n11962 ASIG5V.n11959 0.000662266
R55974 ASIG5V.n6928 ASIG5V.n6791 0.000659204
R55975 ASIG5V.n1068 ASIG5V.n747 0.000656142
R55976 ASIG5V.n4012 ASIG5V.n4009 0.000656142
R55977 ASIG5V.n12420 ASIG5V.n12355 0.000656142
R55978 ASIG5V.n11490 ASIG5V.n11488 0.000656142
R55979 ASIG5V.n3737 ASIG5V.n3626 0.000653081
R55980 ASIG5V.n7936 ASIG5V.n7823 0.000653081
R55981 ASIG5V.n4698 ASIG5V.n4633 0.000650019
R55982 ASIG5V.n7993 ASIG5V.n7990 0.000650019
R55983 ASIG5V.n9433 ASIG5V.n9121 0.000650019
R55984 ASIG5V.n4007 ASIG5V.n4004 0.000646958
R55985 ASIG5V.n5452 ASIG5V.n5448 0.000643896
R55986 ASIG5V.n7124 ASIG5V.n6331 0.000637773
R55987 ASIG5V.n6784 ASIG5V.n6780 0.000637773
R55988 ASIG5V.n4901 ASIG5V.n4857 0.000631649
R55989 ASIG5V.n6552 ASIG5V.n3 0.000631649
R55990 ASIG5V.n7406 ASIG5V.n7401 0.000628588
R55991 ASIG5V.n7629 ASIG5V.n7626 0.000628588
R55992 ASIG5V.n5154 ASIG5V.n5151 0.000625526
R55993 ASIG5V.n7124 ASIG5V.n7123 0.000625526
R55994 ASIG5V.n7401 ASIG5V.n7285 0.000625526
R55995 ASIG5V.n7519 ASIG5V.n7406 0.000625526
R55996 ASIG5V.n6777 ASIG5V.n6769 0.000622465
R55997 ASIG5V.n6780 ASIG5V.n6777 0.000619403
R55998 ASIG5V.n6657 ASIG5V.n6652 0.000619403
R55999 ASIG5V.n12665 ASIG5V.n12662 0.000619403
R56000 ASIG5V.n11106 ASIG5V.n11104 0.000619403
R56001 ASIG5V.n5445 ASIG5V.n5442 0.000616341
R56002 ASIG5V.n11763 ASIG5V.n11760 0.000616341
R56003 ASIG5V.n2915 ASIG5V.n2883 0.00061328
R56004 ASIG5V.n3747 ASIG5V.n3745 0.00061328
R56005 ASIG5V.n12306 ASIG5V.n12303 0.00061328
R56006 ASIG5V.n11672 ASIG5V.n11670 0.00061328
R56007 ASIG5V.n4847 ASIG5V.n4698 0.000610218
R56008 ASIG5V.n12154 ASIG5V.n12150 0.000610218
R56009 ASIG5V.n3255 ASIG5V.n3253 0.000607157
R56010 ASIG5V.n3479 ASIG5V.n3477 0.000607157
R56011 ASIG5V.n4563 ASIG5V.n4561 0.000607157
R56012 ASIG5V.n12009 ASIG5V.n12006 0.000607157
R56013 ASIG5V.n11841 ASIG5V.n11839 0.000607157
R56014 ASIG5V.n13353 ASIG5V.n331 0.000604095
R56015 ASIG5V.n3558 ASIG5V.n3483 0.000601033
R56016 ASIG5V.n4164 ASIG5V.n4099 0.000601033
R56017 ASIG5V.n12430 ASIG5V.n12427 0.000601033
R56018 ASIG5V.n11419 ASIG5V.n11416 0.000601033
R56019 ASIG5V.n7983 ASIG5V.n7979 0.000597972
R56020 ASIG5V.n9119 ASIG5V.n9118 0.000597972
R56021 ASIG5V.n9117 ASIG5V.n9116 0.000597972
R56022 ASIG5V.n8982 ASIG5V.n8981 0.000597972
R56023 ASIG5V.n8976 ASIG5V.n8975 0.000597972
R56024 ASIG5V.n8880 ASIG5V.n8879 0.000597972
R56025 ASIG5V.n4852 ASIG5V.n4849 0.00059491
R56026 ASIG5V.n7986 ASIG5V.n7983 0.00059491
R56027 ASIG5V.n12646 ASIG5V.n12581 0.000588787
R56028 ASIG5V.n3136 ASIG5V.n3104 0.000585725
R56029 ASIG5V.n5671 ASIG5V.n5559 0.000585725
R56030 ASIG5V.n5328 ASIG5V.n5154 0.000582664
R56031 ASIG5V.n5442 ASIG5V.n5398 0.000582664
R56032 ASIG5V.n7066 ASIG5V.n7063 0.000582664
R56033 ASIG5V.n6791 ASIG5V.n6787 0.000582664
R56034 ASIG5V.n2883 ASIG5V.n2880 0.000573479
R56035 ASIG5V.n3034 ASIG5V.n3032 0.000573479
R56036 ASIG5V.n5860 ASIG5V.n5855 0.000573479
R56037 ASIG5V.n6152 ASIG5V.n6149 0.000573479
R56038 ASIG5V.n5148 ASIG5V.n5145 0.000570417
R56039 ASIG5V.n6326 ASIG5V.n6163 0.000570417
R56040 ASIG5V.n7633 ASIG5V.n7629 0.000570417
R56041 ASIG5V.n12310 ASIG5V.n12306 0.000570417
R56042 ASIG5V.n12238 ASIG5V.n12164 0.000570417
R56043 ASIG5V.n6652 ASIG5V.n6556 0.000567356
R56044 ASIG5V.n12758 ASIG5V.n8120 0.000567356
R56045 ASIG5V.n3833 ASIG5V.n3747 0.000564294
R56046 ASIG5V.n4004 ASIG5V.n3899 0.000564294
R56047 ASIG5V.n4443 ASIG5V.n4440 0.000564294
R56048 ASIG5V.n12659 ASIG5V.n12656 0.000564294
R56049 ASIG5V.n11834 ASIG5V.n11831 0.000564294
R56050 ASIG5V.n11311 ASIG5V.n11189 0.000564294
R56051 ASIG5V.n11189 ASIG5V.n11157 0.000564294
R56052 ASIG5V.n3036 ASIG5V.n3034 0.000558171
R56053 ASIG5V.n3742 ASIG5V.n3740 0.000558171
R56054 ASIG5V.n6149 ASIG5V.n5972 0.000558171
R56055 ASIG5V.n12164 ASIG5V.n12162 0.000558171
R56056 ASIG5V.n11676 ASIG5V.n11674 0.000558171
R56057 ASIG5V.n3475 ASIG5V.n3331 0.000555109
R56058 ASIG5V.n4630 ASIG5V.n4571 0.000555109
R56059 ASIG5V.n12082 ASIG5V.n12009 0.000555109
R56060 ASIG5V.n3139 ASIG5V.n3136 0.000552047
R56061 ASIG5V.n3483 ASIG5V.n3481 0.000552047
R56062 ASIG5V.n12150 ASIG5V.n12085 0.000552047
R56063 ASIG5V.n11836 ASIG5V.n11834 0.000552047
R56064 ASIG5V.n11486 ASIG5V.n11419 0.000552047
R56065 ASIG5V.n11324 ASIG5V.n11319 0.000552047
R56066 ASIG5V.n13621 ASIG5V.n13618 0.000548986
R56067 ASIG5V.n13364 ASIG5V.n13360 0.000548986
R56068 ASIG5V.n4282 ASIG5V.n4279 0.000545924
R56069 ASIG5V.n12435 ASIG5V.n12432 0.000545924
R56070 ASIG5V.n11319 ASIG5V.n11317 0.000545924
R56071 ASIG5V.n4440 ASIG5V.n4375 0.000542863
R56072 ASIG5V.n11959 ASIG5V.n11926 0.000542863
R56073 ASIG5V.n4857 ASIG5V.n4854 0.000539801
R56074 ASIG5V.n13360 ASIG5V.n13358 0.000539801
R56075 ASIG5V.n7274 ASIG5V.n331 0.000539801
R56076 ASIG5V.n7941 ASIG5V.n7936 0.000539801
R56077 ASIG5V ASIG5V.n3 0.000536739
R56078 ASIG5V.n13371 ASIG5V.n13367 0.000533678
R56079 ASIG5V.n12656 ASIG5V.n12653 0.000533678
R56080 ASIG5V.n3253 ASIG5V.n3251 0.000530616
R56081 ASIG5V.n5797 ASIG5V.n5793 0.000530616
R56082 ASIG5V.n7059 ASIG5V.n7056 0.000527555
R56083 ASIG5V.n7048 ASIG5V.n6935 0.000527555
R56084 ASIG5V.n13618 ASIG5V.n13616 0.000527555
R56085 ASIG5V.n13607 ASIG5V.n13495 0.000527555
R56086 ASIG5V.n11670 ASIG5V.n11668 0.000527555
R56087 ASIG5V.n11634 ASIG5V.n11631 0.000527555
R56088 ASIG5V.n514 ASIG5V.n513 0.000524493
R56089 ASIG5V.n622 ASIG5V.n621 0.000524493
R56090 ASIG5V.n628 ASIG5V.n627 0.000524493
R56091 ASIG5V.n742 ASIG5V.n741 0.000524493
R56092 ASIG5V.n745 ASIG5V.n744 0.000524493
R56093 ASIG5V.n5804 ASIG5V.n5801 0.000521431
R56094 ASIG5V.n13612 ASIG5V.n13607 0.000521431
R56095 ASIG5V.n4099 ASIG5V.n4096 0.000515308
R56096 ASIG5V.n4279 ASIG5V.n4277 0.000515308
R56097 ASIG5V.n4971 ASIG5V.n4966 0.000515308
R56098 ASIG5V.n7640 ASIG5V.n7636 0.000515308
R56099 ASIG5V.n4561 ASIG5V.n4446 0.000512246
R56100 ASIG5V.n12752 ASIG5V.n12668 0.000512246
R56101 ASIG5V.n11999 ASIG5V.n11997 0.000512246
R56102 ASIG5V.n4287 ASIG5V.n4285 0.000509185
R56103 ASIG5V.n12651 ASIG5V.n12646 0.000509185
R56104 ASIG5V.n12427 ASIG5V.n12425 0.000509185
R56105 ASIG5V.n12355 ASIG5V.n12352 0.000509185
R56106 ASIG5V.n11315 ASIG5V.n11313 0.000509185
R56107 ASIG5V.n11154 ASIG5V.n11106 0.000509185
R56108 ASIG5V.n3040 ASIG5V.n3038 0.000503062
R56109 ASIG5V.n3626 ASIG5V.n3623 0.000503062
R56110 ASIG5V.n5559 ASIG5V.n5455 0.000503062
R56111 ASIG5V.n5793 ASIG5V.n5676 0.000503062
R56112 ASIG5V.n5855 ASIG5V.n5808 0.000503062
R56113 ASIG5V.n12159 ASIG5V.n12157 0.000503062
R56114 ASIG5V.n11828 ASIG5V.n11763 0.000503062
R56115 VDD.n15 VDD.n14 4.74241
R56116 VDD.n10 VDD.n9 0.2255
R56117 VDD.n8 VDD.n7 0.2255
R56118 VDD.n14 VDD.n13 0.207672
R56119 VDD.n16 VDD.n15 0.207641
R56120 VDD.n14 VDD.n4 0.207427
R56121 VDD.n6 VDD 0.087472
R56122 VDD.n19 VDD 0.0780816
R56123 VDD.n6 VDD.n5 0.0714207
R56124 VDD.n16 VDD.n2 0.0677462
R56125 VDD.n19 VDD 0.0567182
R56126 VDD.n13 VDD.n12 0.0557908
R56127 VDD.n2 VDD.n1 0.0504883
R56128 VDD.n12 VDD.n9 0.0403484
R56129 VDD.n2 VDD.n0 0.0213316
R56130 VDD.n12 VDD.n11 0.0190982
R56131 VDD.n20 VDD.n19 0.016049
R56132 VDD.n7 VDD.n6 0.0110106
R56133 VDD.n11 VDD 0.00782857
R56134 VDD VDD.n0 0.00782857
R56135 VDD.n4 VDD.n3 0.00467857
R56136 VDD.n18 VDD.n17 0.00467857
R56137 VDD.n9 VDD.n8 0.00455714
R56138 VDD.n1 VDD 0.00455714
R56139 VDD.n17 VDD.n16 0.00429286
R56140 VDD VDD.n4 0.00365
R56141 VDD VDD.n18 0.00365
R56142 VDD VDD.n10 0.0023
R56143 VDD.n5 VDD 0.0023
R56144 VDD VDD.n20 0.0023
R56145 VDD.n8 VDD 0.0011
R56146 VSS.n13649 VSS.n13648 4017.81
R56147 VSS.n14264 VSS.n14263 4017.81
R56148 VSS.n15679 VSS.n15678 99.2437
R56149 VSS.n9837 VSS.n9836 32.468
R56150 VSS.n12643 VSS.n12642 32.468
R56151 VSS.n16296 VSS.n16295 6.79968
R56152 VSS.n1377 VSS.n1376 6.79968
R56153 VSS.n16332 VSS.n16331 6.79968
R56154 VSS.n1421 VSS.n1419 6.79968
R56155 VSS.n13653 VSS.n13651 6.39837
R56156 VSS.n14269 VSS.n14266 6.39837
R56157 VSS.n19411 VSS.n19359 6.3005
R56158 VSS.n19405 VSS.n19361 6.3005
R56159 VSS.n19390 VSS.n19368 6.3005
R56160 VSS.n19393 VSS.n19365 6.3005
R56161 VSS.n19399 VSS.n19363 6.3005
R56162 VSS.n19414 VSS.n19356 6.3005
R56163 VSS.n19419 VSS.n19355 6.3005
R56164 VSS.n19423 VSS.n19353 6.3005
R56165 VSS.n19427 VSS.n19351 6.3005
R56166 VSS.n19431 VSS.n19349 6.3005
R56167 VSS.n19435 VSS.n19347 6.3005
R56168 VSS.n19345 VSS.n19343 6.3005
R56169 VSS.n19331 VSS.n19329 6.3005
R56170 VSS.n19324 VSS.n19322 6.3005
R56171 VSS.n19317 VSS.n19315 6.3005
R56172 VSS.n19310 VSS.n19308 6.3005
R56173 VSS.n19303 VSS.n19301 6.3005
R56174 VSS.n19296 VSS.n19294 6.3005
R56175 VSS.n19289 VSS.n19287 6.3005
R56176 VSS.n19282 VSS.n19280 6.3005
R56177 VSS.n19275 VSS.n19273 6.3005
R56178 VSS.n19267 VSS.n19265 6.3005
R56179 VSS.n19259 VSS.n19257 6.3005
R56180 VSS.n19251 VSS.n19249 6.3005
R56181 VSS.n19414 VSS.n19413 6.3005
R56182 VSS.n19251 VSS.n19250 6.3005
R56183 VSS.n19259 VSS.n19258 6.3005
R56184 VSS.n19267 VSS.n19266 6.3005
R56185 VSS.n19275 VSS.n19274 6.3005
R56186 VSS.n19282 VSS.n19281 6.3005
R56187 VSS.n19289 VSS.n19288 6.3005
R56188 VSS.n19296 VSS.n19295 6.3005
R56189 VSS.n19303 VSS.n19302 6.3005
R56190 VSS.n19310 VSS.n19309 6.3005
R56191 VSS.n19317 VSS.n19316 6.3005
R56192 VSS.n19324 VSS.n19323 6.3005
R56193 VSS.n19331 VSS.n19330 6.3005
R56194 VSS.n19345 VSS.n19344 6.3005
R56195 VSS.n19435 VSS.n19434 6.3005
R56196 VSS.n19431 VSS.n19430 6.3005
R56197 VSS.n19427 VSS.n19426 6.3005
R56198 VSS.n19423 VSS.n19422 6.3005
R56199 VSS.n19419 VSS.n19418 6.3005
R56200 VSS.n19399 VSS.n19398 6.3005
R56201 VSS.n19390 VSS.n19389 6.3005
R56202 VSS.n19393 VSS.n19392 6.3005
R56203 VSS.n19405 VSS.n19404 6.3005
R56204 VSS.n19411 VSS.n19410 6.3005
R56205 VSS.n18479 VSS.n18477 6.3005
R56206 VSS.n18479 VSS.n18478 6.3005
R56207 VSS.n18652 VSS.n18650 6.3005
R56208 VSS.n18645 VSS.n18643 6.3005
R56209 VSS.n18638 VSS.n18636 6.3005
R56210 VSS.n18631 VSS.n18629 6.3005
R56211 VSS.n18624 VSS.n18622 6.3005
R56212 VSS.n18617 VSS.n18615 6.3005
R56213 VSS.n18610 VSS.n18608 6.3005
R56214 VSS.n18603 VSS.n18601 6.3005
R56215 VSS.n18596 VSS.n18594 6.3005
R56216 VSS.n18589 VSS.n18587 6.3005
R56217 VSS.n18582 VSS.n18580 6.3005
R56218 VSS.n18575 VSS.n18573 6.3005
R56219 VSS.n18555 VSS.n18553 6.3005
R56220 VSS.n18562 VSS.n18557 6.3005
R56221 VSS.n18547 VSS.n18545 6.3005
R56222 VSS.n18540 VSS.n18538 6.3005
R56223 VSS.n18533 VSS.n18531 6.3005
R56224 VSS.n18526 VSS.n18524 6.3005
R56225 VSS.n18519 VSS.n18517 6.3005
R56226 VSS.n18512 VSS.n18510 6.3005
R56227 VSS.n18505 VSS.n18503 6.3005
R56228 VSS.n18498 VSS.n18496 6.3005
R56229 VSS.n18491 VSS.n18489 6.3005
R56230 VSS.n18498 VSS.n18497 6.3005
R56231 VSS.n18652 VSS.n18651 6.3005
R56232 VSS.n18645 VSS.n18644 6.3005
R56233 VSS.n18638 VSS.n18637 6.3005
R56234 VSS.n18631 VSS.n18630 6.3005
R56235 VSS.n18624 VSS.n18623 6.3005
R56236 VSS.n18617 VSS.n18616 6.3005
R56237 VSS.n18610 VSS.n18609 6.3005
R56238 VSS.n18603 VSS.n18602 6.3005
R56239 VSS.n18596 VSS.n18595 6.3005
R56240 VSS.n18589 VSS.n18588 6.3005
R56241 VSS.n18582 VSS.n18581 6.3005
R56242 VSS.n18575 VSS.n18574 6.3005
R56243 VSS.n18555 VSS.n18554 6.3005
R56244 VSS.n18562 VSS.n18561 6.3005
R56245 VSS.n18547 VSS.n18546 6.3005
R56246 VSS.n18540 VSS.n18539 6.3005
R56247 VSS.n18533 VSS.n18532 6.3005
R56248 VSS.n18526 VSS.n18525 6.3005
R56249 VSS.n18519 VSS.n18518 6.3005
R56250 VSS.n18512 VSS.n18511 6.3005
R56251 VSS.n18505 VSS.n18504 6.3005
R56252 VSS.n18491 VSS.n18490 6.3005
R56253 VSS.n18254 VSS.n18239 6.3005
R56254 VSS.n18260 VSS.n18237 6.3005
R56255 VSS.n18266 VSS.n18235 6.3005
R56256 VSS.n18272 VSS.n18233 6.3005
R56257 VSS.n18276 VSS.n18231 6.3005
R56258 VSS.n18280 VSS.n18229 6.3005
R56259 VSS.n18284 VSS.n18227 6.3005
R56260 VSS.n18288 VSS.n18225 6.3005
R56261 VSS.n18292 VSS.n18223 6.3005
R56262 VSS.n18296 VSS.n18221 6.3005
R56263 VSS.n18300 VSS.n18219 6.3005
R56264 VSS.n18217 VSS.n18215 6.3005
R56265 VSS.n18313 VSS.n18311 6.3005
R56266 VSS.n18320 VSS.n18318 6.3005
R56267 VSS.n18327 VSS.n18325 6.3005
R56268 VSS.n18334 VSS.n18332 6.3005
R56269 VSS.n18341 VSS.n18339 6.3005
R56270 VSS.n18348 VSS.n18346 6.3005
R56271 VSS.n18355 VSS.n18353 6.3005
R56272 VSS.n18386 VSS.n18384 6.3005
R56273 VSS.n18378 VSS.n18376 6.3005
R56274 VSS.n18370 VSS.n18368 6.3005
R56275 VSS.n18362 VSS.n18360 6.3005
R56276 VSS.n18416 VSS.n18414 6.3005
R56277 VSS.n18254 VSS.n18253 6.3005
R56278 VSS.n18416 VSS.n18415 6.3005
R56279 VSS.n18362 VSS.n18361 6.3005
R56280 VSS.n18370 VSS.n18369 6.3005
R56281 VSS.n18378 VSS.n18377 6.3005
R56282 VSS.n18386 VSS.n18385 6.3005
R56283 VSS.n18355 VSS.n18354 6.3005
R56284 VSS.n18348 VSS.n18347 6.3005
R56285 VSS.n18341 VSS.n18340 6.3005
R56286 VSS.n18334 VSS.n18333 6.3005
R56287 VSS.n18327 VSS.n18326 6.3005
R56288 VSS.n18320 VSS.n18319 6.3005
R56289 VSS.n18313 VSS.n18312 6.3005
R56290 VSS.n18217 VSS.n18216 6.3005
R56291 VSS.n18300 VSS.n18299 6.3005
R56292 VSS.n18296 VSS.n18295 6.3005
R56293 VSS.n18292 VSS.n18291 6.3005
R56294 VSS.n18288 VSS.n18287 6.3005
R56295 VSS.n18284 VSS.n18283 6.3005
R56296 VSS.n18280 VSS.n18279 6.3005
R56297 VSS.n18276 VSS.n18275 6.3005
R56298 VSS.n18272 VSS.n18271 6.3005
R56299 VSS.n18266 VSS.n18265 6.3005
R56300 VSS.n18260 VSS.n18259 6.3005
R56301 VSS.n14955 VSS.n14953 6.3005
R56302 VSS.n16864 VSS.n16862 6.3005
R56303 VSS.n16864 VSS.n16863 6.3005
R56304 VSS.n16853 VSS.n16851 6.3005
R56305 VSS.n16853 VSS.n16852 6.3005
R56306 VSS.n16844 VSS.n16842 6.3005
R56307 VSS.n16844 VSS.n16843 6.3005
R56308 VSS.n16839 VSS.n16837 6.3005
R56309 VSS.n16839 VSS.n16838 6.3005
R56310 VSS.n16830 VSS.n16828 6.3005
R56311 VSS.n16830 VSS.n16829 6.3005
R56312 VSS.n16825 VSS.n16823 6.3005
R56313 VSS.n16825 VSS.n16824 6.3005
R56314 VSS.n16816 VSS.n16814 6.3005
R56315 VSS.n16816 VSS.n16815 6.3005
R56316 VSS.n16811 VSS.n16809 6.3005
R56317 VSS.n16811 VSS.n16810 6.3005
R56318 VSS.n16802 VSS.n16800 6.3005
R56319 VSS.n16802 VSS.n16801 6.3005
R56320 VSS.n16797 VSS.n16795 6.3005
R56321 VSS.n16797 VSS.n16796 6.3005
R56322 VSS.n16788 VSS.n16786 6.3005
R56323 VSS.n16788 VSS.n16787 6.3005
R56324 VSS.n16783 VSS.n16781 6.3005
R56325 VSS.n16783 VSS.n16782 6.3005
R56326 VSS.n16769 VSS.n16767 6.3005
R56327 VSS.n16769 VSS.n16768 6.3005
R56328 VSS.n16760 VSS.n16752 6.3005
R56329 VSS.n16760 VSS.n16759 6.3005
R56330 VSS.n16757 VSS.n16755 6.3005
R56331 VSS.n16757 VSS.n16756 6.3005
R56332 VSS.n16746 VSS.n16744 6.3005
R56333 VSS.n16746 VSS.n16745 6.3005
R56334 VSS.n16741 VSS.n16739 6.3005
R56335 VSS.n16741 VSS.n16740 6.3005
R56336 VSS.n16732 VSS.n16730 6.3005
R56337 VSS.n16732 VSS.n16731 6.3005
R56338 VSS.n16727 VSS.n16725 6.3005
R56339 VSS.n16727 VSS.n16726 6.3005
R56340 VSS.n16718 VSS.n16716 6.3005
R56341 VSS.n16718 VSS.n16717 6.3005
R56342 VSS.n16713 VSS.n16711 6.3005
R56343 VSS.n16713 VSS.n16712 6.3005
R56344 VSS.n16704 VSS.n16702 6.3005
R56345 VSS.n16704 VSS.n16703 6.3005
R56346 VSS.n14949 VSS.n14947 6.3005
R56347 VSS.n14949 VSS.n14948 6.3005
R56348 VSS.n14955 VSS.n14954 6.3005
R56349 VSS.n14678 VSS.n14676 6.3005
R56350 VSS.n14685 VSS.n14683 6.3005
R56351 VSS.n19786 VSS.n19784 6.3005
R56352 VSS.n14693 VSS.n14691 6.3005
R56353 VSS.n19794 VSS.n19792 6.3005
R56354 VSS.n14701 VSS.n14699 6.3005
R56355 VSS.n14708 VSS.n14706 6.3005
R56356 VSS.n14715 VSS.n14713 6.3005
R56357 VSS.n19804 VSS.n19802 6.3005
R56358 VSS.n14723 VSS.n14721 6.3005
R56359 VSS.n19812 VSS.n19810 6.3005
R56360 VSS.n19819 VSS.n19817 6.3005
R56361 VSS.n14733 VSS.n14731 6.3005
R56362 VSS.n14806 VSS.n14736 6.3005
R56363 VSS.n14802 VSS.n14738 6.3005
R56364 VSS.n14799 VSS.n14741 6.3005
R56365 VSS.n14795 VSS.n14743 6.3005
R56366 VSS.n14792 VSS.n14746 6.3005
R56367 VSS.n14788 VSS.n14748 6.3005
R56368 VSS.n14785 VSS.n14751 6.3005
R56369 VSS.n14781 VSS.n14753 6.3005
R56370 VSS.n14778 VSS.n14756 6.3005
R56371 VSS.n14774 VSS.n14758 6.3005
R56372 VSS.n14678 VSS.n14677 6.3005
R56373 VSS.n14685 VSS.n14684 6.3005
R56374 VSS.n19786 VSS.n19785 6.3005
R56375 VSS.n14693 VSS.n14692 6.3005
R56376 VSS.n19794 VSS.n19793 6.3005
R56377 VSS.n14701 VSS.n14700 6.3005
R56378 VSS.n14708 VSS.n14707 6.3005
R56379 VSS.n14715 VSS.n14714 6.3005
R56380 VSS.n19804 VSS.n19803 6.3005
R56381 VSS.n14723 VSS.n14722 6.3005
R56382 VSS.n19812 VSS.n19811 6.3005
R56383 VSS.n19819 VSS.n19818 6.3005
R56384 VSS.n14733 VSS.n14732 6.3005
R56385 VSS.n14806 VSS.n14805 6.3005
R56386 VSS.n14802 VSS.n14801 6.3005
R56387 VSS.n14799 VSS.n14798 6.3005
R56388 VSS.n14795 VSS.n14794 6.3005
R56389 VSS.n14792 VSS.n14791 6.3005
R56390 VSS.n14788 VSS.n14787 6.3005
R56391 VSS.n14785 VSS.n14784 6.3005
R56392 VSS.n14781 VSS.n14780 6.3005
R56393 VSS.n14778 VSS.n14777 6.3005
R56394 VSS.n14774 VSS.n14773 6.3005
R56395 VSS.n14771 VSS.n14761 6.3005
R56396 VSS.n14771 VSS.n14770 6.3005
R56397 VSS.n14473 VSS.n14471 6.3005
R56398 VSS.n14480 VSS.n14478 6.3005
R56399 VSS.n14487 VSS.n14485 6.3005
R56400 VSS.n14494 VSS.n14492 6.3005
R56401 VSS.n14501 VSS.n14499 6.3005
R56402 VSS.n14508 VSS.n14506 6.3005
R56403 VSS.n14515 VSS.n14513 6.3005
R56404 VSS.n14522 VSS.n14520 6.3005
R56405 VSS.n14529 VSS.n14527 6.3005
R56406 VSS.n14536 VSS.n14534 6.3005
R56407 VSS.n14543 VSS.n14541 6.3005
R56408 VSS.n14550 VSS.n14548 6.3005
R56409 VSS.n14450 VSS.n14448 6.3005
R56410 VSS.n14590 VSS.n14588 6.3005
R56411 VSS.n14596 VSS.n14594 6.3005
R56412 VSS.n14602 VSS.n14600 6.3005
R56413 VSS.n14608 VSS.n14606 6.3005
R56414 VSS.n14614 VSS.n14612 6.3005
R56415 VSS.n14620 VSS.n14618 6.3005
R56416 VSS.n14626 VSS.n14624 6.3005
R56417 VSS.n14632 VSS.n14630 6.3005
R56418 VSS.n14638 VSS.n14636 6.3005
R56419 VSS.n14644 VSS.n14642 6.3005
R56420 VSS.n14473 VSS.n14472 6.3005
R56421 VSS.n14480 VSS.n14479 6.3005
R56422 VSS.n14487 VSS.n14486 6.3005
R56423 VSS.n14494 VSS.n14493 6.3005
R56424 VSS.n14501 VSS.n14500 6.3005
R56425 VSS.n14508 VSS.n14507 6.3005
R56426 VSS.n14515 VSS.n14514 6.3005
R56427 VSS.n14522 VSS.n14521 6.3005
R56428 VSS.n14529 VSS.n14528 6.3005
R56429 VSS.n14536 VSS.n14535 6.3005
R56430 VSS.n14543 VSS.n14542 6.3005
R56431 VSS.n14550 VSS.n14549 6.3005
R56432 VSS.n14450 VSS.n14449 6.3005
R56433 VSS.n14590 VSS.n14589 6.3005
R56434 VSS.n14596 VSS.n14595 6.3005
R56435 VSS.n14602 VSS.n14601 6.3005
R56436 VSS.n14608 VSS.n14607 6.3005
R56437 VSS.n14614 VSS.n14613 6.3005
R56438 VSS.n14620 VSS.n14619 6.3005
R56439 VSS.n14626 VSS.n14625 6.3005
R56440 VSS.n14632 VSS.n14631 6.3005
R56441 VSS.n14638 VSS.n14637 6.3005
R56442 VSS.n14644 VSS.n14643 6.3005
R56443 VSS.n14650 VSS.n14648 6.3005
R56444 VSS.n14650 VSS.n14649 6.3005
R56445 VSS.n14922 VSS.n14920 6.3005
R56446 VSS.n14914 VSS.n14912 6.3005
R56447 VSS.n14906 VSS.n14904 6.3005
R56448 VSS.n16954 VSS.n16947 6.3005
R56449 VSS.n16959 VSS.n16944 6.3005
R56450 VSS.n16964 VSS.n16941 6.3005
R56451 VSS.n16968 VSS.n14854 6.3005
R56452 VSS.n16974 VSS.n14852 6.3005
R56453 VSS.n16980 VSS.n14850 6.3005
R56454 VSS.n16985 VSS.n14847 6.3005
R56455 VSS.n16995 VSS.n14841 6.3005
R56456 VSS.n17006 VSS.n14836 6.3005
R56457 VSS.n17046 VSS.n17044 6.3005
R56458 VSS.n17052 VSS.n17042 6.3005
R56459 VSS.n17058 VSS.n17040 6.3005
R56460 VSS.n17063 VSS.n17037 6.3005
R56461 VSS.n17098 VSS.n17096 6.3005
R56462 VSS.n17103 VSS.n17093 6.3005
R56463 VSS.n17108 VSS.n17090 6.3005
R56464 VSS.n17113 VSS.n17087 6.3005
R56465 VSS.n17145 VSS.n17143 6.3005
R56466 VSS.n17151 VSS.n17141 6.3005
R56467 VSS.n17157 VSS.n17139 6.3005
R56468 VSS.n17151 VSS.n17150 6.3005
R56469 VSS.n14914 VSS.n14913 6.3005
R56470 VSS.n14922 VSS.n14921 6.3005
R56471 VSS.n17157 VSS.n17156 6.3005
R56472 VSS.n17145 VSS.n17144 6.3005
R56473 VSS.n17113 VSS.n17112 6.3005
R56474 VSS.n17108 VSS.n17107 6.3005
R56475 VSS.n17103 VSS.n17102 6.3005
R56476 VSS.n17098 VSS.n17097 6.3005
R56477 VSS.n17063 VSS.n17062 6.3005
R56478 VSS.n17058 VSS.n17057 6.3005
R56479 VSS.n17052 VSS.n17051 6.3005
R56480 VSS.n17046 VSS.n17045 6.3005
R56481 VSS.n17006 VSS.n17005 6.3005
R56482 VSS.n16995 VSS.n16994 6.3005
R56483 VSS.n16985 VSS.n16984 6.3005
R56484 VSS.n16980 VSS.n16979 6.3005
R56485 VSS.n16974 VSS.n16973 6.3005
R56486 VSS.n16968 VSS.n16967 6.3005
R56487 VSS.n16964 VSS.n16963 6.3005
R56488 VSS.n16959 VSS.n16958 6.3005
R56489 VSS.n16954 VSS.n16953 6.3005
R56490 VSS.n14906 VSS.n14905 6.3005
R56491 VSS.n16513 VSS.n14977 6.3005
R56492 VSS.n16415 VSS.n16413 6.3005
R56493 VSS.n16409 VSS.n16407 6.3005
R56494 VSS.n16454 VSS.n16452 6.3005
R56495 VSS.n16461 VSS.n16459 6.3005
R56496 VSS.n16468 VSS.n16466 6.3005
R56497 VSS.n16475 VSS.n16473 6.3005
R56498 VSS.n16482 VSS.n16480 6.3005
R56499 VSS.n16489 VSS.n16487 6.3005
R56500 VSS.n16496 VSS.n16494 6.3005
R56501 VSS.n16503 VSS.n16501 6.3005
R56502 VSS.n16507 VSS.n14979 6.3005
R56503 VSS.n16557 VSS.n16555 6.3005
R56504 VSS.n16563 VSS.n16553 6.3005
R56505 VSS.n16568 VSS.n16550 6.3005
R56506 VSS.n16574 VSS.n16548 6.3005
R56507 VSS.n16609 VSS.n16607 6.3005
R56508 VSS.n16615 VSS.n16605 6.3005
R56509 VSS.n16620 VSS.n16602 6.3005
R56510 VSS.n16625 VSS.n16599 6.3005
R56511 VSS.n16651 VSS.n16649 6.3005
R56512 VSS.n16657 VSS.n16647 6.3005
R56513 VSS.n16663 VSS.n16645 6.3005
R56514 VSS.n16676 VSS.n16674 6.3005
R56515 VSS.n16676 VSS.n16675 6.3005
R56516 VSS.n16663 VSS.n16662 6.3005
R56517 VSS.n16563 VSS.n16562 6.3005
R56518 VSS.n16557 VSS.n16556 6.3005
R56519 VSS.n16513 VSS.n16512 6.3005
R56520 VSS.n16507 VSS.n16506 6.3005
R56521 VSS.n16503 VSS.n16502 6.3005
R56522 VSS.n16496 VSS.n16495 6.3005
R56523 VSS.n16489 VSS.n16488 6.3005
R56524 VSS.n16482 VSS.n16481 6.3005
R56525 VSS.n16475 VSS.n16474 6.3005
R56526 VSS.n16468 VSS.n16467 6.3005
R56527 VSS.n16461 VSS.n16460 6.3005
R56528 VSS.n16454 VSS.n16453 6.3005
R56529 VSS.n16409 VSS.n16408 6.3005
R56530 VSS.n16415 VSS.n16414 6.3005
R56531 VSS.n16574 VSS.n16573 6.3005
R56532 VSS.n16568 VSS.n16567 6.3005
R56533 VSS.n16615 VSS.n16614 6.3005
R56534 VSS.n16609 VSS.n16608 6.3005
R56535 VSS.n16657 VSS.n16656 6.3005
R56536 VSS.n16651 VSS.n16650 6.3005
R56537 VSS.n16625 VSS.n16624 6.3005
R56538 VSS.n16620 VSS.n16619 6.3005
R56539 VSS.n15890 VSS.n15888 6.3005
R56540 VSS.n15890 VSS.n15889 6.3005
R56541 VSS.n15716 VSS.n15714 6.3005
R56542 VSS.n15722 VSS.n15720 6.3005
R56543 VSS.n15730 VSS.n15728 6.3005
R56544 VSS.n15736 VSS.n15734 6.3005
R56545 VSS.n15744 VSS.n15742 6.3005
R56546 VSS.n15750 VSS.n15748 6.3005
R56547 VSS.n15758 VSS.n15756 6.3005
R56548 VSS.n15764 VSS.n15762 6.3005
R56549 VSS.n15772 VSS.n15770 6.3005
R56550 VSS.n15778 VSS.n15776 6.3005
R56551 VSS.n15786 VSS.n15784 6.3005
R56552 VSS.n15792 VSS.n15790 6.3005
R56553 VSS.n15806 VSS.n15804 6.3005
R56554 VSS.n15816 VSS.n15814 6.3005
R56555 VSS.n15820 VSS.n15818 6.3005
R56556 VSS.n15828 VSS.n15826 6.3005
R56557 VSS.n15834 VSS.n15832 6.3005
R56558 VSS.n15842 VSS.n15840 6.3005
R56559 VSS.n15848 VSS.n15846 6.3005
R56560 VSS.n15866 VSS.n15864 6.3005
R56561 VSS.n15872 VSS.n15870 6.3005
R56562 VSS.n15878 VSS.n15876 6.3005
R56563 VSS.n15884 VSS.n15882 6.3005
R56564 VSS.n15878 VSS.n15877 6.3005
R56565 VSS.n15716 VSS.n15715 6.3005
R56566 VSS.n15722 VSS.n15721 6.3005
R56567 VSS.n15730 VSS.n15729 6.3005
R56568 VSS.n15736 VSS.n15735 6.3005
R56569 VSS.n15744 VSS.n15743 6.3005
R56570 VSS.n15750 VSS.n15749 6.3005
R56571 VSS.n15758 VSS.n15757 6.3005
R56572 VSS.n15764 VSS.n15763 6.3005
R56573 VSS.n15772 VSS.n15771 6.3005
R56574 VSS.n15778 VSS.n15777 6.3005
R56575 VSS.n15786 VSS.n15785 6.3005
R56576 VSS.n15792 VSS.n15791 6.3005
R56577 VSS.n15806 VSS.n15805 6.3005
R56578 VSS.n15816 VSS.n15815 6.3005
R56579 VSS.n15820 VSS.n15819 6.3005
R56580 VSS.n15828 VSS.n15827 6.3005
R56581 VSS.n15834 VSS.n15833 6.3005
R56582 VSS.n15842 VSS.n15841 6.3005
R56583 VSS.n15848 VSS.n15847 6.3005
R56584 VSS.n15866 VSS.n15865 6.3005
R56585 VSS.n15872 VSS.n15871 6.3005
R56586 VSS.n15884 VSS.n15883 6.3005
R56587 VSS.n14169 VSS.n14168 5.91395
R56588 VSS.n21233 VSS.n21232 5.86071
R56589 VSS.n17396 VSS.n17395 5.84304
R56590 VSS.n11415 VSS.n11414 5.84304
R56591 VSS.n11468 VSS.n11467 5.84304
R56592 VSS.n11638 VSS.n11637 5.84304
R56593 VSS.n17384 VSS.n17383 5.84304
R56594 VSS.n11253 VSS.n11252 5.84304
R56595 VSS.n2518 VSS.n2517 5.84304
R56596 VSS.n15897 VSS.n15896 5.7755
R56597 VSS.n19382 VSS.n19370 5.7755
R56598 VSS.n19382 VSS.n19381 5.7755
R56599 VSS.n18484 VSS.n18483 5.7755
R56600 VSS.n18249 VSS.n18248 5.7755
R56601 VSS.n18249 VSS.n18242 5.7755
R56602 VSS.n14962 VSS.n14961 5.7755
R56603 VSS.n14765 VSS.n14763 5.7755
R56604 VSS.n14657 VSS.n14656 5.7755
R56605 VSS.n14931 VSS.n14930 5.7755
R56606 VSS.n16422 VSS.n16421 5.7755
R56607 VSS.n21936 VSS.n35 5.7217
R56608 VSS.n15709 VSS.n15708 5.70391
R56609 VSS.n19241 VSS.n19240 5.70391
R56610 VSS.n18660 VSS.n18659 5.70391
R56611 VSS.n18430 VSS.n18428 5.70391
R56612 VSS.n18430 VSS.n18429 5.70391
R56613 VSS.n16859 VSS.n16858 5.70391
R56614 VSS.n19775 VSS.n19774 5.70391
R56615 VSS.n14464 VSS.n14463 5.70391
R56616 VSS.n17135 VSS.n17134 5.70391
R56617 VSS.n16670 VSS.n16669 5.70391
R56618 VSS.n13655 VSS.n13653 5.70148
R56619 VSS.n14272 VSS.n14269 5.70148
R56620 VSS.n858 VSS.n857 5.2293
R56621 VSS.n11301 VSS.n11300 5.2293
R56622 VSS.n902 VSS.n901 5.2005
R56623 VSS.n15916 VSS.n15915 5.2005
R56624 VSS.n1418 VSS.n1417 5.2005
R56625 VSS.n1417 VSS.n1416 5.2005
R56626 VSS.n16330 VSS.n16329 5.2005
R56627 VSS.n16329 VSS.n16328 5.2005
R56628 VSS.n1428 VSS.n1427 5.2005
R56629 VSS.n16340 VSS.n16339 5.2005
R56630 VSS.n16258 VSS.n16257 5.2005
R56631 VSS.n16260 VSS.n16259 5.2005
R56632 VSS.n1342 VSS.n1341 5.2005
R56633 VSS.n1344 VSS.n1343 5.2005
R56634 VSS.n5662 VSS.n5661 5.2005
R56635 VSS.n20931 VSS.n20930 5.2005
R56636 VSS.n20973 VSS.n20972 5.2005
R56637 VSS.n5762 VSS.n5761 5.2005
R56638 VSS.n20883 VSS.n20882 5.2005
R56639 VSS.n20882 VSS.n20881 5.2005
R56640 VSS.n5754 VSS.n5753 5.2005
R56641 VSS.n5753 VSS.n5752 5.2005
R56642 VSS.n8959 VSS.n8958 5.2005
R56643 VSS.n8957 VSS.n8956 5.2005
R56644 VSS.n9981 VSS.n9980 5.2005
R56645 VSS.n9989 VSS.n9988 5.2005
R56646 VSS.n9997 VSS.n9996 5.2005
R56647 VSS.n10005 VSS.n10004 5.2005
R56648 VSS.n10012 VSS.n10011 5.2005
R56649 VSS.n10019 VSS.n10018 5.2005
R56650 VSS.n10027 VSS.n10026 5.2005
R56651 VSS.n10035 VSS.n10034 5.2005
R56652 VSS.n10043 VSS.n10042 5.2005
R56653 VSS.n10051 VSS.n10050 5.2005
R56654 VSS.n10059 VSS.n10058 5.2005
R56655 VSS.n10066 VSS.n10065 5.2005
R56656 VSS.n10073 VSS.n10072 5.2005
R56657 VSS.n10081 VSS.n10080 5.2005
R56658 VSS.n10089 VSS.n10088 5.2005
R56659 VSS.n10097 VSS.n10096 5.2005
R56660 VSS.n10105 VSS.n10104 5.2005
R56661 VSS.n10113 VSS.n10112 5.2005
R56662 VSS.n10121 VSS.n10120 5.2005
R56663 VSS.n10128 VSS.n10127 5.2005
R56664 VSS.n10135 VSS.n10134 5.2005
R56665 VSS.n10143 VSS.n10142 5.2005
R56666 VSS.n10151 VSS.n10150 5.2005
R56667 VSS.n10160 VSS.n10159 5.2005
R56668 VSS.n10158 VSS.n10157 5.2005
R56669 VSS.n10336 VSS.n10335 5.2005
R56670 VSS.n10344 VSS.n10343 5.2005
R56671 VSS.n10351 VSS.n10350 5.2005
R56672 VSS.n10358 VSS.n10357 5.2005
R56673 VSS.n10366 VSS.n10365 5.2005
R56674 VSS.n10374 VSS.n10373 5.2005
R56675 VSS.n10382 VSS.n10381 5.2005
R56676 VSS.n10390 VSS.n10389 5.2005
R56677 VSS.n10398 VSS.n10397 5.2005
R56678 VSS.n10406 VSS.n10405 5.2005
R56679 VSS.n10413 VSS.n10412 5.2005
R56680 VSS.n10420 VSS.n10419 5.2005
R56681 VSS.n10428 VSS.n10427 5.2005
R56682 VSS.n10436 VSS.n10435 5.2005
R56683 VSS.n10445 VSS.n10444 5.2005
R56684 VSS.n10443 VSS.n10442 5.2005
R56685 VSS.n10318 VSS.n10317 5.2005
R56686 VSS.n10310 VSS.n10309 5.2005
R56687 VSS.n10302 VSS.n10301 5.2005
R56688 VSS.n10295 VSS.n10294 5.2005
R56689 VSS.n10288 VSS.n10287 5.2005
R56690 VSS.n10280 VSS.n10279 5.2005
R56691 VSS.n9889 VSS.n9888 5.2005
R56692 VSS.n9880 VSS.n9879 5.2005
R56693 VSS.n9872 VSS.n9871 5.2005
R56694 VSS.n10531 VSS.n10530 5.2005
R56695 VSS.n9864 VSS.n9863 5.2005
R56696 VSS.n9862 VSS.n9861 5.2005
R56697 VSS.n9858 VSS.n9857 5.2005
R56698 VSS.n9854 VSS.n9853 5.2005
R56699 VSS.n9852 VSS.n9833 5.2005
R56700 VSS.n9833 VSS.n9832 5.2005
R56701 VSS.n9835 VSS.n9834 5.2005
R56702 VSS.n8860 VSS.n8859 5.2005
R56703 VSS.n8864 VSS.n8861 5.2005
R56704 VSS.n12009 VSS.n12008 5.2005
R56705 VSS.n12010 VSS.n12002 5.2005
R56706 VSS.n8864 VSS.n8855 5.2005
R56707 VSS.n8864 VSS.n8851 5.2005
R56708 VSS.n12667 VSS.n12666 5.2005
R56709 VSS.n12663 VSS.n12662 5.2005
R56710 VSS.n12659 VSS.n12658 5.2005
R56711 VSS.n12656 VSS.n12650 5.2005
R56712 VSS.n12650 VSS.n12649 5.2005
R56713 VSS.n12641 VSS.n12640 5.2005
R56714 VSS.n12016 VSS.n12015 5.2005
R56715 VSS.n12669 VSS.n12668 5.2005
R56716 VSS.n12597 VSS.n12596 5.2005
R56717 VSS.n11773 VSS.n11772 5.2005
R56718 VSS.n11781 VSS.n11780 5.2005
R56719 VSS.n12568 VSS.n12567 5.2005
R56720 VSS.n12334 VSS.n12333 5.2005
R56721 VSS.n12342 VSS.n12341 5.2005
R56722 VSS.n12349 VSS.n12348 5.2005
R56723 VSS.n12356 VSS.n12355 5.2005
R56724 VSS.n12364 VSS.n12363 5.2005
R56725 VSS.n12372 VSS.n12371 5.2005
R56726 VSS.n12497 VSS.n12496 5.2005
R56727 VSS.n12499 VSS.n12498 5.2005
R56728 VSS.n12490 VSS.n12489 5.2005
R56729 VSS.n12482 VSS.n12481 5.2005
R56730 VSS.n12474 VSS.n12473 5.2005
R56731 VSS.n12467 VSS.n12466 5.2005
R56732 VSS.n12460 VSS.n12459 5.2005
R56733 VSS.n12452 VSS.n12451 5.2005
R56734 VSS.n12444 VSS.n12443 5.2005
R56735 VSS.n12436 VSS.n12435 5.2005
R56736 VSS.n12428 VSS.n12427 5.2005
R56737 VSS.n12420 VSS.n12419 5.2005
R56738 VSS.n12412 VSS.n12411 5.2005
R56739 VSS.n12405 VSS.n12404 5.2005
R56740 VSS.n12398 VSS.n12397 5.2005
R56741 VSS.n12390 VSS.n12389 5.2005
R56742 VSS.n12209 VSS.n12208 5.2005
R56743 VSS.n12211 VSS.n12210 5.2005
R56744 VSS.n12202 VSS.n12201 5.2005
R56745 VSS.n12194 VSS.n12193 5.2005
R56746 VSS.n12186 VSS.n12185 5.2005
R56747 VSS.n12179 VSS.n12178 5.2005
R56748 VSS.n12172 VSS.n12171 5.2005
R56749 VSS.n12164 VSS.n12163 5.2005
R56750 VSS.n12156 VSS.n12155 5.2005
R56751 VSS.n12148 VSS.n12147 5.2005
R56752 VSS.n12140 VSS.n12139 5.2005
R56753 VSS.n12132 VSS.n12131 5.2005
R56754 VSS.n12124 VSS.n12123 5.2005
R56755 VSS.n12117 VSS.n12116 5.2005
R56756 VSS.n12110 VSS.n12109 5.2005
R56757 VSS.n12102 VSS.n12101 5.2005
R56758 VSS.n12094 VSS.n12093 5.2005
R56759 VSS.n12086 VSS.n12085 5.2005
R56760 VSS.n12078 VSS.n12077 5.2005
R56761 VSS.n12070 VSS.n12069 5.2005
R56762 VSS.n12063 VSS.n12062 5.2005
R56763 VSS.n12056 VSS.n12055 5.2005
R56764 VSS.n12048 VSS.n12047 5.2005
R56765 VSS.n12040 VSS.n12039 5.2005
R56766 VSS.n12032 VSS.n12031 5.2005
R56767 VSS.n12024 VSS.n12023 5.2005
R56768 VSS.n11255 VSS.n11254 5.2005
R56769 VSS.n11260 VSS.n11259 5.2005
R56770 VSS.n11265 VSS.n11264 5.2005
R56771 VSS.n11270 VSS.n11269 5.2005
R56772 VSS.n11275 VSS.n11274 5.2005
R56773 VSS.n11280 VSS.n11279 5.2005
R56774 VSS.n11284 VSS.n11283 5.2005
R56775 VSS.n11289 VSS.n11288 5.2005
R56776 VSS.n11294 VSS.n11293 5.2005
R56777 VSS.n11299 VSS.n11298 5.2005
R56778 VSS.n11305 VSS.n11304 5.2005
R56779 VSS.n15185 VSS.n15184 5.2005
R56780 VSS.n15190 VSS.n15189 5.2005
R56781 VSS.n15195 VSS.n15194 5.2005
R56782 VSS.n15911 VSS.n15910 5.2005
R56783 VSS.n15907 VSS.n15906 5.2005
R56784 VSS.n15200 VSS.n15199 5.2005
R56785 VSS.n15700 VSS.n15699 5.2005
R56786 VSS.n856 VSS.n855 5.2005
R56787 VSS.n1476 VSS.n1475 5.2005
R56788 VSS.n1471 VSS.n1470 5.2005
R56789 VSS.n878 VSS.n877 5.2005
R56790 VSS.n873 VSS.n872 5.2005
R56791 VSS.n868 VSS.n867 5.2005
R56792 VSS.n863 VSS.n862 5.2005
R56793 VSS.n449 VSS.n448 5.2005
R56794 VSS.n454 VSS.n453 5.2005
R56795 VSS.n459 VSS.n458 5.2005
R56796 VSS.n21197 VSS.n21196 5.2005
R56797 VSS.n21202 VSS.n21201 5.2005
R56798 VSS.n21206 VSS.n21205 5.2005
R56799 VSS.n21211 VSS.n21210 5.2005
R56800 VSS.n21216 VSS.n21215 5.2005
R56801 VSS.n21221 VSS.n21220 5.2005
R56802 VSS.n21226 VSS.n21225 5.2005
R56803 VSS.n21231 VSS.n21230 5.2005
R56804 VSS.n5884 VSS.n5883 5.2005
R56805 VSS.n5891 VSS.n5890 5.2005
R56806 VSS.n5419 VSS.n5418 5.2005
R56807 VSS.n5418 VSS.n5417 5.2005
R56808 VSS.n5468 VSS.n5467 5.2005
R56809 VSS.n5463 VSS.n5462 5.2005
R56810 VSS.n5428 VSS.n5427 5.2005
R56811 VSS.n5423 VSS.n5422 5.2005
R56812 VSS.n4864 VSS.n4863 5.2005
R56813 VSS.n4863 VSS.n4862 5.2005
R56814 VSS.n4913 VSS.n4912 5.2005
R56815 VSS.n4908 VSS.n4907 5.2005
R56816 VSS.n4873 VSS.n4872 5.2005
R56817 VSS.n4868 VSS.n4867 5.2005
R56818 VSS.n4802 VSS.n4801 5.2005
R56819 VSS.n4801 VSS.n4800 5.2005
R56820 VSS.n4849 VSS.n4848 5.2005
R56821 VSS.n4844 VSS.n4843 5.2005
R56822 VSS.n4811 VSS.n4810 5.2005
R56823 VSS.n4806 VSS.n4805 5.2005
R56824 VSS.n14301 VSS.n14300 5.2005
R56825 VSS.n14300 VSS.n14299 5.2005
R56826 VSS.n17301 VSS.n17300 5.2005
R56827 VSS.n17296 VSS.n17295 5.2005
R56828 VSS.n17263 VSS.n17262 5.2005
R56829 VSS.n17258 VSS.n17257 5.2005
R56830 VSS.n17254 VSS.n17253 5.2005
R56831 VSS.n17253 VSS.n17252 5.2005
R56832 VSS.n2419 VSS.n2418 5.2005
R56833 VSS.n2414 VSS.n2413 5.2005
R56834 VSS.n2389 VSS.n2388 5.2005
R56835 VSS.n2384 VSS.n2383 5.2005
R56836 VSS.n2458 VSS.n2457 5.2005
R56837 VSS.n2457 VSS.n2456 5.2005
R56838 VSS.n2505 VSS.n2504 5.2005
R56839 VSS.n2500 VSS.n2499 5.2005
R56840 VSS.n2467 VSS.n2466 5.2005
R56841 VSS.n2462 VSS.n2461 5.2005
R56842 VSS.n2455 VSS.n2454 5.2005
R56843 VSS.n2454 VSS.n2453 5.2005
R56844 VSS.n3931 VSS.n3930 5.2005
R56845 VSS.n3926 VSS.n3925 5.2005
R56846 VSS.n3898 VSS.n3897 5.2005
R56847 VSS.n3893 VSS.n3892 5.2005
R56848 VSS.n188 VSS.n187 5.2005
R56849 VSS.n21933 VSS.n188 5.2005
R56850 VSS.n178 VSS.n177 5.2005
R56851 VSS.n183 VSS.n182 5.2005
R56852 VSS.n379 VSS.n378 5.2005
R56853 VSS.n385 VSS.n381 5.2005
R56854 VSS.n385 VSS.n383 5.2005
R56855 VSS.n17382 VSS.n17381 5.2005
R56856 VSS.n17377 VSS.n17376 5.2005
R56857 VSS.n17372 VSS.n17371 5.2005
R56858 VSS.n17368 VSS.n17367 5.2005
R56859 VSS.n17364 VSS.n17363 5.2005
R56860 VSS.n17360 VSS.n17359 5.2005
R56861 VSS.n17356 VSS.n17355 5.2005
R56862 VSS.n17353 VSS.n17352 5.2005
R56863 VSS.n14392 VSS.n14391 5.2005
R56864 VSS.n14435 VSS.n14434 5.2005
R56865 VSS.n14439 VSS.n14438 5.2005
R56866 VSS.n14443 VSS.n14442 5.2005
R56867 VSS.n14447 VSS.n14446 5.2005
R56868 VSS.n14667 VSS.n14666 5.2005
R56869 VSS.n2135 VSS.n2134 5.2005
R56870 VSS.n13438 VSS.n13437 5.2005
R56871 VSS.n13442 VSS.n13441 5.2005
R56872 VSS.n13446 VSS.n13445 5.2005
R56873 VSS.n13450 VSS.n13449 5.2005
R56874 VSS.n13457 VSS.n13456 5.2005
R56875 VSS.n13452 VSS.n13451 5.2005
R56876 VSS.n13371 VSS.n13370 5.2005
R56877 VSS.n13403 VSS.n13402 5.2005
R56878 VSS.n13399 VSS.n13398 5.2005
R56879 VSS.n13395 VSS.n13394 5.2005
R56880 VSS.n13391 VSS.n13390 5.2005
R56881 VSS.n13387 VSS.n13386 5.2005
R56882 VSS.n13383 VSS.n13382 5.2005
R56883 VSS.n13379 VSS.n13378 5.2005
R56884 VSS.n13374 VSS.n13373 5.2005
R56885 VSS.n385 VSS.n380 5.2005
R56886 VSS.n385 VSS.n384 5.2005
R56887 VSS.n14284 VSS.n14283 5.2005
R56888 VSS.n403 VSS.n399 5.2005
R56889 VSS.n403 VSS.n401 5.2005
R56890 VSS.n11636 VSS.n11635 5.2005
R56891 VSS.n11631 VSS.n11630 5.2005
R56892 VSS.n11626 VSS.n11625 5.2005
R56893 VSS.n11621 VSS.n11620 5.2005
R56894 VSS.n11616 VSS.n11615 5.2005
R56895 VSS.n11612 VSS.n11611 5.2005
R56896 VSS.n11608 VSS.n11607 5.2005
R56897 VSS.n11604 VSS.n11603 5.2005
R56898 VSS.n11600 VSS.n11599 5.2005
R56899 VSS.n11597 VSS.n11596 5.2005
R56900 VSS.n15081 VSS.n15080 5.2005
R56901 VSS.n15095 VSS.n15094 5.2005
R56902 VSS.n15091 VSS.n15090 5.2005
R56903 VSS.n15087 VSS.n15086 5.2005
R56904 VSS.n15083 VSS.n15082 5.2005
R56905 VSS.n14941 VSS.n14940 5.2005
R56906 VSS.n738 VSS.n737 5.2005
R56907 VSS.n20046 VSS.n20045 5.2005
R56908 VSS.n20050 VSS.n20049 5.2005
R56909 VSS.n20054 VSS.n20053 5.2005
R56910 VSS.n20058 VSS.n20057 5.2005
R56911 VSS.n20065 VSS.n20064 5.2005
R56912 VSS.n20060 VSS.n20059 5.2005
R56913 VSS.n20693 VSS.n20692 5.2005
R56914 VSS.n20725 VSS.n20724 5.2005
R56915 VSS.n20721 VSS.n20720 5.2005
R56916 VSS.n20717 VSS.n20716 5.2005
R56917 VSS.n20713 VSS.n20712 5.2005
R56918 VSS.n20709 VSS.n20708 5.2005
R56919 VSS.n20705 VSS.n20704 5.2005
R56920 VSS.n20701 VSS.n20700 5.2005
R56921 VSS.n20696 VSS.n20695 5.2005
R56922 VSS.n403 VSS.n398 5.2005
R56923 VSS.n403 VSS.n402 5.2005
R56924 VSS.n397 VSS.n396 5.2005
R56925 VSS.n420 VSS.n416 5.2005
R56926 VSS.n420 VSS.n418 5.2005
R56927 VSS.n11470 VSS.n11469 5.2005
R56928 VSS.n11475 VSS.n11474 5.2005
R56929 VSS.n11480 VSS.n11479 5.2005
R56930 VSS.n11485 VSS.n11484 5.2005
R56931 VSS.n11490 VSS.n11489 5.2005
R56932 VSS.n11494 VSS.n11493 5.2005
R56933 VSS.n11498 VSS.n11497 5.2005
R56934 VSS.n11502 VSS.n11501 5.2005
R56935 VSS.n11509 VSS.n11508 5.2005
R56936 VSS.n11506 VSS.n11505 5.2005
R56937 VSS.n15114 VSS.n15113 5.2005
R56938 VSS.n15128 VSS.n15127 5.2005
R56939 VSS.n15124 VSS.n15123 5.2005
R56940 VSS.n15120 VSS.n15119 5.2005
R56941 VSS.n15116 VSS.n15115 5.2005
R56942 VSS.n14970 VSS.n14969 5.2005
R56943 VSS.n743 VSS.n742 5.2005
R56944 VSS.n2083 VSS.n2082 5.2005
R56945 VSS.n2079 VSS.n2078 5.2005
R56946 VSS.n2075 VSS.n2074 5.2005
R56947 VSS.n2071 VSS.n2070 5.2005
R56948 VSS.n2067 VSS.n2066 5.2005
R56949 VSS.n2062 VSS.n2061 5.2005
R56950 VSS.n20744 VSS.n20743 5.2005
R56951 VSS.n20776 VSS.n20775 5.2005
R56952 VSS.n20772 VSS.n20771 5.2005
R56953 VSS.n20768 VSS.n20767 5.2005
R56954 VSS.n20764 VSS.n20763 5.2005
R56955 VSS.n20760 VSS.n20759 5.2005
R56956 VSS.n20756 VSS.n20755 5.2005
R56957 VSS.n20752 VSS.n20751 5.2005
R56958 VSS.n20747 VSS.n20746 5.2005
R56959 VSS.n420 VSS.n415 5.2005
R56960 VSS.n420 VSS.n419 5.2005
R56961 VSS.n414 VSS.n413 5.2005
R56962 VSS.n437 VSS.n433 5.2005
R56963 VSS.n437 VSS.n435 5.2005
R56964 VSS.n11413 VSS.n11412 5.2005
R56965 VSS.n11408 VSS.n11407 5.2005
R56966 VSS.n11403 VSS.n11402 5.2005
R56967 VSS.n11398 VSS.n11397 5.2005
R56968 VSS.n11393 VSS.n11392 5.2005
R56969 VSS.n11389 VSS.n11388 5.2005
R56970 VSS.n11385 VSS.n11384 5.2005
R56971 VSS.n11381 VSS.n11380 5.2005
R56972 VSS.n11377 VSS.n11376 5.2005
R56973 VSS.n11374 VSS.n11373 5.2005
R56974 VSS.n14998 VSS.n14997 5.2005
R56975 VSS.n16391 VSS.n16390 5.2005
R56976 VSS.n16395 VSS.n16394 5.2005
R56977 VSS.n16399 VSS.n16398 5.2005
R56978 VSS.n16403 VSS.n16402 5.2005
R56979 VSS.n16430 VSS.n16429 5.2005
R56980 VSS.n748 VSS.n747 5.2005
R56981 VSS.n1973 VSS.n1972 5.2005
R56982 VSS.n1977 VSS.n1976 5.2005
R56983 VSS.n1981 VSS.n1980 5.2005
R56984 VSS.n1985 VSS.n1984 5.2005
R56985 VSS.n1992 VSS.n1991 5.2005
R56986 VSS.n1987 VSS.n1986 5.2005
R56987 VSS.n20836 VSS.n20835 5.2005
R56988 VSS.n20868 VSS.n20867 5.2005
R56989 VSS.n20864 VSS.n20863 5.2005
R56990 VSS.n20860 VSS.n20859 5.2005
R56991 VSS.n20856 VSS.n20855 5.2005
R56992 VSS.n20852 VSS.n20851 5.2005
R56993 VSS.n20848 VSS.n20847 5.2005
R56994 VSS.n20844 VSS.n20843 5.2005
R56995 VSS.n20839 VSS.n20838 5.2005
R56996 VSS.n437 VSS.n432 5.2005
R56997 VSS.n437 VSS.n436 5.2005
R56998 VSS.n431 VSS.n430 5.2005
R56999 VSS.n21240 VSS.n21238 5.2005
R57000 VSS.n21240 VSS.n21236 5.2005
R57001 VSS.n17414 VSS.n17413 5.2005
R57002 VSS.n17409 VSS.n17408 5.2005
R57003 VSS.n21686 VSS.n21685 5.2005
R57004 VSS.n17398 VSS.n17397 5.2005
R57005 VSS.n17405 VSS.n17404 5.2005
R57006 VSS.n371 VSS.n370 5.2005
R57007 VSS.n13287 VSS.n13286 5.2005
R57008 VSS.n13301 VSS.n13300 5.2005
R57009 VSS.n13296 VSS.n13295 5.2005
R57010 VSS.n13291 VSS.n13290 5.2005
R57011 VSS.n13304 VSS.n13303 5.2005
R57012 VSS.n13282 VSS.n13281 5.2005
R57013 VSS.n13312 VSS.n13311 5.2005
R57014 VSS.n13308 VSS.n13307 5.2005
R57015 VSS.n17959 VSS.n17958 5.2005
R57016 VSS.n13465 VSS.n13464 5.2005
R57017 VSS.n13469 VSS.n13468 5.2005
R57018 VSS.n17957 VSS.n17956 5.2005
R57019 VSS.n13461 VSS.n13460 5.2005
R57020 VSS.n18129 VSS.n18128 5.2005
R57021 VSS.n18134 VSS.n18133 5.2005
R57022 VSS.n2144 VSS.n2143 5.2005
R57023 VSS.n2139 VSS.n2138 5.2005
R57024 VSS.n353 VSS.n352 5.2005
R57025 VSS.n359 VSS.n355 5.2005
R57026 VSS.n21692 VSS.n21688 5.2005
R57027 VSS.n2520 VSS.n2519 5.2005
R57028 VSS.n21715 VSS.n21714 5.2005
R57029 VSS.n21719 VSS.n21718 5.2005
R57030 VSS.n21723 VSS.n21722 5.2005
R57031 VSS.n21727 VSS.n21726 5.2005
R57032 VSS.n21731 VSS.n21730 5.2005
R57033 VSS.n349 VSS.n348 5.2005
R57034 VSS.n21739 VSS.n21738 5.2005
R57035 VSS.n17877 VSS.n17876 5.2005
R57036 VSS.n17882 VSS.n17881 5.2005
R57037 VSS.n17875 VSS.n17874 5.2005
R57038 VSS.n19024 VSS.n19023 5.2005
R57039 VSS.n19020 VSS.n19019 5.2005
R57040 VSS.n19016 VSS.n19015 5.2005
R57041 VSS.n19012 VSS.n19011 5.2005
R57042 VSS.n4081 VSS.n4080 5.2005
R57043 VSS.n4089 VSS.n4088 5.2005
R57044 VSS.n4099 VSS.n4098 5.2005
R57045 VSS.n4107 VSS.n4106 5.2005
R57046 VSS.n4116 VSS.n4115 5.2005
R57047 VSS.n4104 VSS.n4103 5.2005
R57048 VSS.n4094 VSS.n4093 5.2005
R57049 VSS.n4085 VSS.n4084 5.2005
R57050 VSS.n4077 VSS.n4076 5.2005
R57051 VSS.n3945 VSS.n3944 5.2005
R57052 VSS.n21912 VSS.n21911 5.2005
R57053 VSS.n21903 VSS.n21902 5.2005
R57054 VSS.n21894 VSS.n21893 5.2005
R57055 VSS.n21885 VSS.n21884 5.2005
R57056 VSS.n21877 VSS.n21876 5.2005
R57057 VSS.n2151 VSS.n2150 5.2005
R57058 VSS.n2160 VSS.n2159 5.2005
R57059 VSS.n19166 VSS.n19165 5.2005
R57060 VSS.n19372 VSS.n19371 5.2005
R57061 VSS.n18848 VSS.n18847 5.2005
R57062 VSS.n2181 VSS.n2180 5.2005
R57063 VSS.n21899 VSS.n21898 5.2005
R57064 VSS.n21889 VSS.n21888 5.2005
R57065 VSS.n21881 VSS.n21880 5.2005
R57066 VSS.n346 VSS.n345 5.2005
R57067 VSS.n2156 VSS.n2155 5.2005
R57068 VSS.n19162 VSS.n19161 5.2005
R57069 VSS.n19170 VSS.n19169 5.2005
R57070 VSS.n18844 VSS.n18843 5.2005
R57071 VSS.n2177 VSS.n2176 5.2005
R57072 VSS.n2173 VSS.n2172 5.2005
R57073 VSS.n66 VSS.n65 5.2005
R57074 VSS.n154 VSS.n153 5.2005
R57075 VSS.n161 VSS.n160 5.2005
R57076 VSS.n327 VSS.n326 5.2005
R57077 VSS.n320 VSS.n319 5.2005
R57078 VSS.n289 VSS.n288 5.2005
R57079 VSS.n257 VSS.n256 5.2005
R57080 VSS.n225 VSS.n224 5.2005
R57081 VSS.n59 VSS.n58 5.2005
R57082 VSS.n53 VSS.n52 5.2005
R57083 VSS.n48 VSS.n47 5.2005
R57084 VSS.n43 VSS.n42 5.2005
R57085 VSS.n295 VSS.n294 5.2005
R57086 VSS.n302 VSS.n301 5.2005
R57087 VSS.n307 VSS.n306 5.2005
R57088 VSS.n314 VSS.n313 5.2005
R57089 VSS.n263 VSS.n262 5.2005
R57090 VSS.n270 VSS.n269 5.2005
R57091 VSS.n275 VSS.n274 5.2005
R57092 VSS.n282 VSS.n281 5.2005
R57093 VSS.n231 VSS.n230 5.2005
R57094 VSS.n238 VSS.n237 5.2005
R57095 VSS.n243 VSS.n242 5.2005
R57096 VSS.n250 VSS.n249 5.2005
R57097 VSS.n208 VSS.n207 5.2005
R57098 VSS.n213 VSS.n212 5.2005
R57099 VSS.n218 VSS.n217 5.2005
R57100 VSS.n148 VSS.n147 5.2005
R57101 VSS.n141 VSS.n140 5.2005
R57102 VSS.n136 VSS.n135 5.2005
R57103 VSS.n129 VSS.n128 5.2005
R57104 VSS.n122 VSS.n121 5.2005
R57105 VSS.n342 VSS.n340 5.2005
R57106 VSS.n342 VSS.n338 5.2005
R57107 VSS.n342 VSS.n341 5.2005
R57108 VSS.n21932 VSS.n21931 5.2005
R57109 VSS.n21933 VSS.n21932 5.2005
R57110 VSS.n21930 VSS.n21926 5.2005
R57111 VSS.n21930 VSS.n21928 5.2005
R57112 VSS.n21930 VSS.n21925 5.2005
R57113 VSS.n21930 VSS.n21929 5.2005
R57114 VSS.n117 VSS.n116 5.2005
R57115 VSS.n110 VSS.n109 5.2005
R57116 VSS.n91 VSS.n90 5.2005
R57117 VSS.n85 VSS.n84 5.2005
R57118 VSS.n78 VSS.n77 5.2005
R57119 VSS.n73 VSS.n72 5.2005
R57120 VSS.n98 VSS.n97 5.2005
R57121 VSS.n105 VSS.n104 5.2005
R57122 VSS.n2169 VSS.n2168 5.2005
R57123 VSS.n21692 VSS.n21690 5.2005
R57124 VSS.n19004 VSS.n19003 5.2005
R57125 VSS.n19000 VSS.n18999 5.2005
R57126 VSS.n18996 VSS.n18995 5.2005
R57127 VSS.n18992 VSS.n18991 5.2005
R57128 VSS.n2164 VSS.n2163 5.2005
R57129 VSS.n18983 VSS.n18982 5.2005
R57130 VSS.n4196 VSS.n4195 5.2005
R57131 VSS.n4192 VSS.n4191 5.2005
R57132 VSS.n4184 VSS.n4183 5.2005
R57133 VSS.n4182 VSS.n4181 5.2005
R57134 VSS.n4178 VSS.n4177 5.2005
R57135 VSS.n4173 VSS.n4172 5.2005
R57136 VSS.n4169 VSS.n4168 5.2005
R57137 VSS.n21711 VSS.n21710 5.2005
R57138 VSS.n21704 VSS.n21703 5.2005
R57139 VSS.n21692 VSS.n21687 5.2005
R57140 VSS.n21692 VSS.n21691 5.2005
R57141 VSS.n18125 VSS.n18124 5.2005
R57142 VSS.n17418 VSS.n17417 5.2005
R57143 VSS.n17422 VSS.n17421 5.2005
R57144 VSS.n17426 VSS.n17425 5.2005
R57145 VSS.n17429 VSS.n17428 5.2005
R57146 VSS.n18113 VSS.n18112 5.2005
R57147 VSS.n18117 VSS.n18116 5.2005
R57148 VSS.n18121 VSS.n18120 5.2005
R57149 VSS.n359 VSS.n357 5.2005
R57150 VSS.n359 VSS.n354 5.2005
R57151 VSS.n359 VSS.n358 5.2005
R57152 VSS.n186 VSS.n185 5.2005
R57153 VSS.n5894 VSS.n5893 5.2005
R57154 VSS.n21240 VSS.n21239 5.2005
R57155 VSS.n22225 VSS.n22224 5.2005
R57156 VSS.n22224 VSS.n22223 5.2005
R57157 VSS.n22221 VSS.n22220 5.2005
R57158 VSS.n22233 VSS.n22232 5.2005
R57159 VSS.n22232 VSS.n22231 5.2005
R57160 VSS.n22180 VSS.n22179 5.2005
R57161 VSS.n22179 VSS.n22178 5.2005
R57162 VSS.n22121 VSS.n22120 5.2005
R57163 VSS.n22125 VSS.n22124 5.2005
R57164 VSS.n22130 VSS.n22129 5.2005
R57165 VSS.n22129 VSS.n22128 5.2005
R57166 VSS.n22136 VSS.n22135 5.2005
R57167 VSS.n22135 VSS.n22134 5.2005
R57168 VSS.n22142 VSS.n22141 5.2005
R57169 VSS.n22141 VSS.n22140 5.2005
R57170 VSS.n22148 VSS.n22147 5.2005
R57171 VSS.n22147 VSS.n22146 5.2005
R57172 VSS.n22154 VSS.n22153 5.2005
R57173 VSS.n22153 VSS.n22152 5.2005
R57174 VSS.n22157 VSS.n22156 5.2005
R57175 VSS.n22156 VSS.n22155 5.2005
R57176 VSS.n22172 VSS.n22171 5.2005
R57177 VSS.n22171 VSS.n22170 5.2005
R57178 VSS.n22242 VSS.n22241 5.2005
R57179 VSS.n22241 VSS.n22240 5.2005
R57180 VSS.n22248 VSS.n22247 5.2005
R57181 VSS.n22247 VSS.n22246 5.2005
R57182 VSS.n22217 VSS.n22216 5.2005
R57183 VSS.n22213 VSS.n22212 5.2005
R57184 VSS.n22209 VSS.n22208 5.2005
R57185 VSS.n22205 VSS.n22204 5.2005
R57186 VSS.n22201 VSS.n22200 5.2005
R57187 VSS.n22197 VSS.n22196 5.2005
R57188 VSS.n22193 VSS.n22192 5.2005
R57189 VSS.n22189 VSS.n22188 5.2005
R57190 VSS.n22185 VSS.n22184 5.2005
R57191 VSS.n13640 VSS.n13639 5.2005
R57192 VSS.n13645 VSS.n13644 5.2005
R57193 VSS.n13653 VSS.n13652 5.2005
R57194 VSS.n13651 VSS.n13650 5.2005
R57195 VSS.n13650 VSS.n13649 5.2005
R57196 VSS.n13647 VSS.n13646 5.2005
R57197 VSS.n14262 VSS.n14258 5.2005
R57198 VSS.n14266 VSS.n14265 5.2005
R57199 VSS.n14265 VSS.n14264 5.2005
R57200 VSS.n14257 VSS.n14256 5.2005
R57201 VSS.n14256 VSS.n14255 5.2005
R57202 VSS.n14279 VSS.n14278 5.2005
R57203 VSS.n14278 VSS.n14277 5.2005
R57204 VSS.n14312 VSS.n14311 5.2005
R57205 VSS.n14311 VSS.n14310 5.2005
R57206 VSS.n14325 VSS.n14324 5.2005
R57207 VSS.n14324 VSS.n14323 5.2005
R57208 VSS.n13554 VSS.n13553 5.2005
R57209 VSS.n13553 VSS.n13552 5.2005
R57210 VSS.n13541 VSS.n13540 5.2005
R57211 VSS.n13540 VSS.n13539 5.2005
R57212 VSS.n13575 VSS.n13574 5.2005
R57213 VSS.n13574 VSS.n13573 5.2005
R57214 VSS.n13581 VSS.n13580 5.2005
R57215 VSS.n13580 VSS.n13579 5.2005
R57216 VSS.n13587 VSS.n13586 5.2005
R57217 VSS.n13586 VSS.n13585 5.2005
R57218 VSS.n13593 VSS.n13592 5.2005
R57219 VSS.n13592 VSS.n13591 5.2005
R57220 VSS.n13599 VSS.n13598 5.2005
R57221 VSS.n13598 VSS.n13597 5.2005
R57222 VSS.n13606 VSS.n13605 5.2005
R57223 VSS.n13605 VSS.n13604 5.2005
R57224 VSS.n21982 VSS.n21981 5.2005
R57225 VSS.n21980 VSS.n21979 5.2005
R57226 VSS.n21957 VSS.n21956 5.2005
R57227 VSS.n21955 VSS.n21954 5.2005
R57228 VSS.n21951 VSS.n21950 5.2005
R57229 VSS.n21974 VSS.n21973 5.2005
R57230 VSS.n21964 VSS.n21963 5.2005
R57231 VSS.n5 VSS.n4 5.2005
R57232 VSS.n9 VSS.n8 5.2005
R57233 VSS.n13 VSS.n12 5.2005
R57234 VSS.n17 VSS.n16 5.2005
R57235 VSS.n21 VSS.n20 5.2005
R57236 VSS.n21941 VSS.n21940 5.2005
R57237 VSS.n21940 VSS.n21939 5.2005
R57238 VSS.n21936 VSS.n21935 5.2005
R57239 VSS.n21935 VSS.n21934 5.2005
R57240 VSS.n14269 VSS.n14268 5.2005
R57241 VSS.n14268 VSS.n14267 5.2005
R57242 VSS.n14262 VSS.n14261 5.07814
R57243 VSS.n22228 VSS.n22225 4.83394
R57244 VSS.n22225 VSS.n22222 4.83394
R57245 VSS.n21984 VSS.n21982 4.83394
R57246 VSS.n14370 VSS.n14368 4.60368
R57247 VSS.n13531 VSS.n13530 4.60313
R57248 VSS.n13427 VSS.n13426 4.59757
R57249 VSS.n14354 VSS.n14352 4.59757
R57250 VSS.n9850 VSS.n9838 4.5005
R57251 VSS.n9850 VSS.n9849 4.5005
R57252 VSS.n8864 VSS.n8862 4.5005
R57253 VSS.n8864 VSS.n8863 4.5005
R57254 VSS.n12647 VSS.n12644 4.5005
R57255 VSS.n12647 VSS.n12646 4.5005
R57256 VSS.n21243 VSS.n21241 4.5005
R57257 VSS.n11257 VSS.n11256 4.5005
R57258 VSS.n11263 VSS.n11262 4.5005
R57259 VSS.n11268 VSS.n11267 4.5005
R57260 VSS.n11273 VSS.n11272 4.5005
R57261 VSS.n11278 VSS.n11277 4.5005
R57262 VSS.n11282 VSS.n11281 4.5005
R57263 VSS.n11287 VSS.n11286 4.5005
R57264 VSS.n11292 VSS.n11291 4.5005
R57265 VSS.n11297 VSS.n11296 4.5005
R57266 VSS.n11308 VSS.n11307 4.5005
R57267 VSS.n11303 VSS.n11302 4.5005
R57268 VSS.n15183 VSS.n15182 4.5005
R57269 VSS.n15188 VSS.n15187 4.5005
R57270 VSS.n15193 VSS.n15192 4.5005
R57271 VSS.n15914 VSS.n15913 4.5005
R57272 VSS.n15909 VSS.n15908 4.5005
R57273 VSS.n15905 VSS.n15904 4.5005
R57274 VSS.n15198 VSS.n15197 4.5005
R57275 VSS.n15696 VSS.n15695 4.5005
R57276 VSS.n1479 VSS.n1478 4.5005
R57277 VSS.n1474 VSS.n1473 4.5005
R57278 VSS.n1469 VSS.n1468 4.5005
R57279 VSS.n876 VSS.n875 4.5005
R57280 VSS.n871 VSS.n870 4.5005
R57281 VSS.n866 VSS.n865 4.5005
R57282 VSS.n861 VSS.n860 4.5005
R57283 VSS.n447 VSS.n446 4.5005
R57284 VSS.n452 VSS.n451 4.5005
R57285 VSS.n457 VSS.n456 4.5005
R57286 VSS.n21195 VSS.n21194 4.5005
R57287 VSS.n21200 VSS.n21199 4.5005
R57288 VSS.n21204 VSS.n21203 4.5005
R57289 VSS.n21209 VSS.n21208 4.5005
R57290 VSS.n21214 VSS.n21213 4.5005
R57291 VSS.n21219 VSS.n21218 4.5005
R57292 VSS.n21224 VSS.n21223 4.5005
R57293 VSS.n21229 VSS.n21228 4.5005
R57294 VSS.n389 VSS.n386 4.5005
R57295 VSS.n389 VSS.n377 4.5005
R57296 VSS.n17380 VSS.n17379 4.5005
R57297 VSS.n17375 VSS.n17374 4.5005
R57298 VSS.n17370 VSS.n17369 4.5005
R57299 VSS.n17366 VSS.n17365 4.5005
R57300 VSS.n17362 VSS.n17361 4.5005
R57301 VSS.n17358 VSS.n17357 4.5005
R57302 VSS.n17354 VSS.n17311 4.5005
R57303 VSS.n14390 VSS.n14389 4.5005
R57304 VSS.n14433 VSS.n14432 4.5005
R57305 VSS.n14437 VSS.n14436 4.5005
R57306 VSS.n14441 VSS.n14440 4.5005
R57307 VSS.n14445 VSS.n14444 4.5005
R57308 VSS.n14669 VSS.n14668 4.5005
R57309 VSS.n14665 VSS.n14664 4.5005
R57310 VSS.n2133 VSS.n2132 4.5005
R57311 VSS.n2137 VSS.n2136 4.5005
R57312 VSS.n13440 VSS.n13439 4.5005
R57313 VSS.n13444 VSS.n13443 4.5005
R57314 VSS.n13448 VSS.n13447 4.5005
R57315 VSS.n13459 VSS.n13458 4.5005
R57316 VSS.n13455 VSS.n13454 4.5005
R57317 VSS.n13369 VSS.n13368 4.5005
R57318 VSS.n13405 VSS.n13404 4.5005
R57319 VSS.n13401 VSS.n13400 4.5005
R57320 VSS.n13397 VSS.n13396 4.5005
R57321 VSS.n13393 VSS.n13392 4.5005
R57322 VSS.n13389 VSS.n13388 4.5005
R57323 VSS.n13385 VSS.n13384 4.5005
R57324 VSS.n13381 VSS.n13380 4.5005
R57325 VSS.n13376 VSS.n13375 4.5005
R57326 VSS.n389 VSS.n387 4.5005
R57327 VSS.n389 VSS.n376 4.5005
R57328 VSS.n389 VSS.n388 4.5005
R57329 VSS.n17181 VSS.n17180 4.5005
R57330 VSS.n14344 VSS.n14343 4.5005
R57331 VSS.n14350 VSS.n14349 4.5005
R57332 VSS.n14360 VSS.n14359 4.5005
R57333 VSS.n14364 VSS.n14363 4.5005
R57334 VSS.n14382 VSS.n14381 4.5005
R57335 VSS.n13526 VSS.n13525 4.5005
R57336 VSS.n13516 VSS.n13515 4.5005
R57337 VSS.n13432 VSS.n13431 4.5005
R57338 VSS.n13422 VSS.n13421 4.5005
R57339 VSS.n13274 VSS.n13273 4.5005
R57340 VSS.n13269 VSS.n13268 4.5005
R57341 VSS.n14290 VSS.n14289 4.5005
R57342 VSS.n407 VSS.n404 4.5005
R57343 VSS.n407 VSS.n395 4.5005
R57344 VSS.n11634 VSS.n11633 4.5005
R57345 VSS.n11629 VSS.n11628 4.5005
R57346 VSS.n11624 VSS.n11623 4.5005
R57347 VSS.n11619 VSS.n11618 4.5005
R57348 VSS.n11614 VSS.n11613 4.5005
R57349 VSS.n11610 VSS.n11609 4.5005
R57350 VSS.n11606 VSS.n11605 4.5005
R57351 VSS.n11602 VSS.n11601 4.5005
R57352 VSS.n11598 VSS.n11594 4.5005
R57353 VSS.n15079 VSS.n15078 4.5005
R57354 VSS.n15097 VSS.n15096 4.5005
R57355 VSS.n15093 VSS.n15092 4.5005
R57356 VSS.n15089 VSS.n15088 4.5005
R57357 VSS.n15085 VSS.n15084 4.5005
R57358 VSS.n14943 VSS.n14942 4.5005
R57359 VSS.n14939 VSS.n14938 4.5005
R57360 VSS.n736 VSS.n735 4.5005
R57361 VSS.n20044 VSS.n20043 4.5005
R57362 VSS.n20048 VSS.n20047 4.5005
R57363 VSS.n20052 VSS.n20051 4.5005
R57364 VSS.n20056 VSS.n20055 4.5005
R57365 VSS.n20067 VSS.n20066 4.5005
R57366 VSS.n20063 VSS.n20062 4.5005
R57367 VSS.n20691 VSS.n20690 4.5005
R57368 VSS.n20727 VSS.n20726 4.5005
R57369 VSS.n20723 VSS.n20722 4.5005
R57370 VSS.n20719 VSS.n20718 4.5005
R57371 VSS.n20715 VSS.n20714 4.5005
R57372 VSS.n20711 VSS.n20710 4.5005
R57373 VSS.n20707 VSS.n20706 4.5005
R57374 VSS.n20703 VSS.n20702 4.5005
R57375 VSS.n20698 VSS.n20697 4.5005
R57376 VSS.n407 VSS.n405 4.5005
R57377 VSS.n407 VSS.n394 4.5005
R57378 VSS.n407 VSS.n406 4.5005
R57379 VSS.n424 VSS.n421 4.5005
R57380 VSS.n424 VSS.n412 4.5005
R57381 VSS.n11472 VSS.n11471 4.5005
R57382 VSS.n11478 VSS.n11477 4.5005
R57383 VSS.n11483 VSS.n11482 4.5005
R57384 VSS.n11488 VSS.n11487 4.5005
R57385 VSS.n11492 VSS.n11491 4.5005
R57386 VSS.n11496 VSS.n11495 4.5005
R57387 VSS.n11500 VSS.n11499 4.5005
R57388 VSS.n11511 VSS.n11510 4.5005
R57389 VSS.n11507 VSS.n11503 4.5005
R57390 VSS.n15112 VSS.n15111 4.5005
R57391 VSS.n15130 VSS.n15129 4.5005
R57392 VSS.n15126 VSS.n15125 4.5005
R57393 VSS.n15122 VSS.n15121 4.5005
R57394 VSS.n15118 VSS.n15117 4.5005
R57395 VSS.n14972 VSS.n14971 4.5005
R57396 VSS.n14968 VSS.n14967 4.5005
R57397 VSS.n741 VSS.n740 4.5005
R57398 VSS.n2085 VSS.n2084 4.5005
R57399 VSS.n2081 VSS.n2080 4.5005
R57400 VSS.n2077 VSS.n2076 4.5005
R57401 VSS.n2073 VSS.n2072 4.5005
R57402 VSS.n2069 VSS.n2068 4.5005
R57403 VSS.n2065 VSS.n2064 4.5005
R57404 VSS.n20742 VSS.n20741 4.5005
R57405 VSS.n20778 VSS.n20777 4.5005
R57406 VSS.n20774 VSS.n20773 4.5005
R57407 VSS.n20770 VSS.n20769 4.5005
R57408 VSS.n20766 VSS.n20765 4.5005
R57409 VSS.n20762 VSS.n20761 4.5005
R57410 VSS.n20758 VSS.n20757 4.5005
R57411 VSS.n20754 VSS.n20753 4.5005
R57412 VSS.n20749 VSS.n20748 4.5005
R57413 VSS.n424 VSS.n422 4.5005
R57414 VSS.n424 VSS.n411 4.5005
R57415 VSS.n424 VSS.n423 4.5005
R57416 VSS.n441 VSS.n438 4.5005
R57417 VSS.n441 VSS.n429 4.5005
R57418 VSS.n11411 VSS.n11410 4.5005
R57419 VSS.n11406 VSS.n11405 4.5005
R57420 VSS.n11401 VSS.n11400 4.5005
R57421 VSS.n11396 VSS.n11395 4.5005
R57422 VSS.n11391 VSS.n11390 4.5005
R57423 VSS.n11387 VSS.n11386 4.5005
R57424 VSS.n11383 VSS.n11382 4.5005
R57425 VSS.n11379 VSS.n11378 4.5005
R57426 VSS.n11375 VSS.n11371 4.5005
R57427 VSS.n14996 VSS.n14995 4.5005
R57428 VSS.n16389 VSS.n16388 4.5005
R57429 VSS.n16393 VSS.n16392 4.5005
R57430 VSS.n16397 VSS.n16396 4.5005
R57431 VSS.n16401 VSS.n16400 4.5005
R57432 VSS.n16432 VSS.n16431 4.5005
R57433 VSS.n16428 VSS.n16427 4.5005
R57434 VSS.n746 VSS.n745 4.5005
R57435 VSS.n1971 VSS.n1970 4.5005
R57436 VSS.n1975 VSS.n1974 4.5005
R57437 VSS.n1979 VSS.n1978 4.5005
R57438 VSS.n1983 VSS.n1982 4.5005
R57439 VSS.n1994 VSS.n1993 4.5005
R57440 VSS.n1990 VSS.n1989 4.5005
R57441 VSS.n20834 VSS.n20833 4.5005
R57442 VSS.n20870 VSS.n20869 4.5005
R57443 VSS.n20866 VSS.n20865 4.5005
R57444 VSS.n20862 VSS.n20861 4.5005
R57445 VSS.n20858 VSS.n20857 4.5005
R57446 VSS.n20854 VSS.n20853 4.5005
R57447 VSS.n20850 VSS.n20849 4.5005
R57448 VSS.n20846 VSS.n20845 4.5005
R57449 VSS.n20841 VSS.n20840 4.5005
R57450 VSS.n441 VSS.n439 4.5005
R57451 VSS.n441 VSS.n428 4.5005
R57452 VSS.n441 VSS.n440 4.5005
R57453 VSS.n21243 VSS.n21235 4.5005
R57454 VSS.n21243 VSS.n21242 4.5005
R57455 VSS.n17416 VSS.n17415 4.5005
R57456 VSS.n17412 VSS.n17411 4.5005
R57457 VSS.n17407 VSS.n17406 4.5005
R57458 VSS.n363 VSS.n360 4.5005
R57459 VSS.n363 VSS.n351 4.5005
R57460 VSS.n375 VSS.n374 4.5005
R57461 VSS.n13289 VSS.n13288 4.5005
R57462 VSS.n13302 VSS.n13283 4.5005
R57463 VSS.n13299 VSS.n13298 4.5005
R57464 VSS.n13294 VSS.n13293 4.5005
R57465 VSS.n13306 VSS.n13305 4.5005
R57466 VSS.n13280 VSS.n13279 4.5005
R57467 VSS.n13314 VSS.n13313 4.5005
R57468 VSS.n13310 VSS.n13309 4.5005
R57469 VSS.n17962 VSS.n17961 4.5005
R57470 VSS.n13463 VSS.n13462 4.5005
R57471 VSS.n13471 VSS.n13470 4.5005
R57472 VSS.n13467 VSS.n13466 4.5005
R57473 VSS.n2149 VSS.n2148 4.5005
R57474 VSS.n18127 VSS.n18126 4.5005
R57475 VSS.n18137 VSS.n18136 4.5005
R57476 VSS.n18132 VSS.n18131 4.5005
R57477 VSS.n2146 VSS.n2145 4.5005
R57478 VSS.n21696 VSS.n21693 4.5005
R57479 VSS.n21696 VSS.n21684 4.5005
R57480 VSS.n21717 VSS.n21716 4.5005
R57481 VSS.n21721 VSS.n21720 4.5005
R57482 VSS.n21725 VSS.n21724 4.5005
R57483 VSS.n21729 VSS.n21728 4.5005
R57484 VSS.n21733 VSS.n21732 4.5005
R57485 VSS.n21741 VSS.n21740 4.5005
R57486 VSS.n21737 VSS.n21736 4.5005
R57487 VSS.n17880 VSS.n17879 4.5005
R57488 VSS.n17884 VSS.n17883 4.5005
R57489 VSS.n19026 VSS.n19025 4.5005
R57490 VSS.n19022 VSS.n19021 4.5005
R57491 VSS.n19018 VSS.n19017 4.5005
R57492 VSS.n19014 VSS.n19013 4.5005
R57493 VSS.n19010 VSS.n19009 4.5005
R57494 VSS.n19006 VSS.n19005 4.5005
R57495 VSS.n4079 VSS.n4078 4.5005
R57496 VSS.n4083 VSS.n4082 4.5005
R57497 VSS.n4087 VSS.n4086 4.5005
R57498 VSS.n4092 VSS.n4091 4.5005
R57499 VSS.n4097 VSS.n4096 4.5005
R57500 VSS.n4102 VSS.n4101 4.5005
R57501 VSS.n4105 VSS.n3942 4.5005
R57502 VSS.n4113 VSS.n4112 4.5005
R57503 VSS.n4118 VSS.n4117 4.5005
R57504 VSS.n4075 VSS.n4074 4.5005
R57505 VSS.n2167 VSS.n2166 4.5005
R57506 VSS.n2171 VSS.n2170 4.5005
R57507 VSS.n21909 VSS.n21908 4.5005
R57508 VSS.n21901 VSS.n21900 4.5005
R57509 VSS.n21897 VSS.n21896 4.5005
R57510 VSS.n21892 VSS.n21891 4.5005
R57511 VSS.n21887 VSS.n21886 4.5005
R57512 VSS.n21883 VSS.n21882 4.5005
R57513 VSS.n21879 VSS.n21878 4.5005
R57514 VSS.n21875 VSS.n21874 4.5005
R57515 VSS.n344 VSS.n343 4.5005
R57516 VSS.n2154 VSS.n2153 4.5005
R57517 VSS.n2158 VSS.n2157 4.5005
R57518 VSS.n19160 VSS.n19159 4.5005
R57519 VSS.n19164 VSS.n19163 4.5005
R57520 VSS.n19168 VSS.n19167 4.5005
R57521 VSS.n19172 VSS.n19171 4.5005
R57522 VSS.n19374 VSS.n19373 4.5005
R57523 VSS.n18846 VSS.n18845 4.5005
R57524 VSS.n18850 VSS.n18849 4.5005
R57525 VSS.n2179 VSS.n2178 4.5005
R57526 VSS.n18842 VSS.n18841 4.5005
R57527 VSS.n2175 VSS.n2174 4.5005
R57528 VSS.n63 VSS.n62 4.5005
R57529 VSS.n70 VSS.n69 4.5005
R57530 VSS.n151 VSS.n150 4.5005
R57531 VSS.n158 VSS.n157 4.5005
R57532 VSS.n324 VSS.n323 4.5005
R57533 VSS.n317 VSS.n316 4.5005
R57534 VSS.n292 VSS.n291 4.5005
R57535 VSS.n286 VSS.n285 4.5005
R57536 VSS.n260 VSS.n259 4.5005
R57537 VSS.n254 VSS.n253 4.5005
R57538 VSS.n228 VSS.n227 4.5005
R57539 VSS.n222 VSS.n221 4.5005
R57540 VSS.n56 VSS.n55 4.5005
R57541 VSS.n51 VSS.n50 4.5005
R57542 VSS.n46 VSS.n45 4.5005
R57543 VSS.n40 VSS.n39 4.5005
R57544 VSS.n299 VSS.n298 4.5005
R57545 VSS.n305 VSS.n304 4.5005
R57546 VSS.n311 VSS.n310 4.5005
R57547 VSS.n267 VSS.n266 4.5005
R57548 VSS.n273 VSS.n272 4.5005
R57549 VSS.n279 VSS.n278 4.5005
R57550 VSS.n235 VSS.n234 4.5005
R57551 VSS.n241 VSS.n240 4.5005
R57552 VSS.n247 VSS.n246 4.5005
R57553 VSS.n205 VSS.n204 4.5005
R57554 VSS.n211 VSS.n210 4.5005
R57555 VSS.n216 VSS.n215 4.5005
R57556 VSS.n145 VSS.n144 4.5005
R57557 VSS.n139 VSS.n138 4.5005
R57558 VSS.n133 VSS.n132 4.5005
R57559 VSS.n126 VSS.n125 4.5005
R57560 VSS.n119 VSS.n36 4.5005
R57561 VSS.n21924 VSS.n21921 4.5005
R57562 VSS.n21924 VSS.n21920 4.5005
R57563 VSS.n337 VSS.n335 4.5005
R57564 VSS.n337 VSS.n334 4.5005
R57565 VSS.n337 VSS.n336 4.5005
R57566 VSS.n21924 VSS.n21922 4.5005
R57567 VSS.n21924 VSS.n21919 4.5005
R57568 VSS.n21924 VSS.n21923 4.5005
R57569 VSS.n114 VSS.n113 4.5005
R57570 VSS.n108 VSS.n107 4.5005
R57571 VSS.n95 VSS.n94 4.5005
R57572 VSS.n88 VSS.n87 4.5005
R57573 VSS.n82 VSS.n81 4.5005
R57574 VSS.n76 VSS.n75 4.5005
R57575 VSS.n102 VSS.n101 4.5005
R57576 VSS.n329 VSS.n328 4.5005
R57577 VSS.n163 VSS.n162 4.5005
R57578 VSS.n21914 VSS.n21913 4.5005
R57579 VSS.n21696 VSS.n21694 4.5005
R57580 VSS.n19002 VSS.n19001 4.5005
R57581 VSS.n18998 VSS.n18997 4.5005
R57582 VSS.n18994 VSS.n18993 4.5005
R57583 VSS.n18990 VSS.n18989 4.5005
R57584 VSS.n18985 VSS.n18984 4.5005
R57585 VSS.n18981 VSS.n18980 4.5005
R57586 VSS.n4197 VSS.n4193 4.5005
R57587 VSS.n4190 VSS.n4189 4.5005
R57588 VSS.n4186 VSS.n4185 4.5005
R57589 VSS.n4180 VSS.n4179 4.5005
R57590 VSS.n4176 VSS.n4175 4.5005
R57591 VSS.n4171 VSS.n4170 4.5005
R57592 VSS.n4165 VSS.n4164 4.5005
R57593 VSS.n21713 VSS.n21712 4.5005
R57594 VSS.n21707 VSS.n21706 4.5005
R57595 VSS.n21702 VSS.n21701 4.5005
R57596 VSS.n21696 VSS.n21683 4.5005
R57597 VSS.n21696 VSS.n21695 4.5005
R57598 VSS.n363 VSS.n361 4.5005
R57599 VSS.n2142 VSS.n2141 4.5005
R57600 VSS.n18123 VSS.n18122 4.5005
R57601 VSS.n17420 VSS.n17419 4.5005
R57602 VSS.n17424 VSS.n17423 4.5005
R57603 VSS.n17431 VSS.n17430 4.5005
R57604 VSS.n18111 VSS.n18110 4.5005
R57605 VSS.n18115 VSS.n18114 4.5005
R57606 VSS.n18119 VSS.n18118 4.5005
R57607 VSS.n369 VSS.n368 4.5005
R57608 VSS.n17401 VSS.n17400 4.5005
R57609 VSS.n363 VSS.n350 4.5005
R57610 VSS.n363 VSS.n362 4.5005
R57611 VSS.n13543 VSS.n13542 4.2005
R57612 VSS.n11751 VSS.n11750 4.2005
R57613 VSS.n14314 VSS.n14313 4.2005
R57614 VSS.n14290 VSS.n14280 4.2005
R57615 VSS.n14339 VSS.n14337 4.19666
R57616 VSS.n14370 VSS.n14369 3.98409
R57617 VSS.n13531 VSS.n13529 3.98362
R57618 VSS.n14354 VSS.n14353 3.9788
R57619 VSS.n13427 VSS.n13425 3.9788
R57620 VSS.n11756 VSS.n11755 3.9386
R57621 VSS.n11768 VSS.n11767 3.92116
R57622 VSS.n14333 VSS.n14331 3.90063
R57623 VSS.n14843 VSS.n14842 3.86641
R57624 VSS.n14845 VSS.n14844 3.86641
R57625 VSS.n5694 VSS.n5693 3.71156
R57626 VSS.n20963 VSS.n20962 3.71156
R57627 VSS.n5762 VSS.n5760 3.71156
R57628 VSS.n1216 VSS.n1215 3.71156
R57629 VSS.n14339 VSS.n14338 3.63186
R57630 VSS.n15692 VSS.n15677 3.62347
R57631 VSS.n12001 VSS.n11999 3.58891
R57632 VSS.n11756 VSS.n11754 3.40854
R57633 VSS.n11768 VSS.n11766 3.39344
R57634 VSS.n14333 VSS.n14332 3.37568
R57635 VSS.n19338 VSS.n19336 3.1505
R57636 VSS.n19338 VSS.n19337 3.1505
R57637 VSS.n18568 VSS.n18566 3.1505
R57638 VSS.n18568 VSS.n18567 3.1505
R57639 VSS.n18306 VSS.n18304 3.1505
R57640 VSS.n18306 VSS.n18305 3.1505
R57641 VSS.n16774 VSS.n16772 3.1505
R57642 VSS.n16774 VSS.n16773 3.1505
R57643 VSS.n19826 VSS.n19824 3.1505
R57644 VSS.n19826 VSS.n19825 3.1505
R57645 VSS.n14557 VSS.n14555 3.1505
R57646 VSS.n14557 VSS.n14556 3.1505
R57647 VSS.n17001 VSS.n14839 3.1505
R57648 VSS.n17001 VSS.n17000 3.1505
R57649 VSS.n16518 VSS.n14975 3.1505
R57650 VSS.n16518 VSS.n14974 3.1505
R57651 VSS.n15800 VSS.n15798 3.1505
R57652 VSS.n15800 VSS.n15799 3.1505
R57653 VSS.n15694 VSS.n15693 3.14395
R57654 VSS.n12001 VSS.n12000 3.10592
R57655 VSS.n8854 VSS.n8852 2.91885
R57656 VSS.n12005 VSS.n12004 2.91885
R57657 VSS.n11998 VSS.n11997 2.73983
R57658 VSS.n18487 VSS.n18481 2.6255
R57659 VSS.n14958 VSS.n14957 2.6255
R57660 VSS.n14769 VSS.n14762 2.6255
R57661 VSS.n14653 VSS.n14651 2.6255
R57662 VSS.n17148 VSS.n17142 2.6255
R57663 VSS.n16956 VSS.n16946 2.6255
R57664 VSS.n16961 VSS.n16943 2.6255
R57665 VSS.n16966 VSS.n16965 2.6255
R57666 VSS.n16971 VSS.n14853 2.6255
R57667 VSS.n16982 VSS.n14849 2.6255
R57668 VSS.n16988 VSS.n14846 2.6255
R57669 VSS.n17003 VSS.n14838 2.6255
R57670 VSS.n17008 VSS.n17007 2.6255
R57671 VSS.n17049 VSS.n17043 2.6255
R57672 VSS.n17060 VSS.n17039 2.6255
R57673 VSS.n17100 VSS.n17095 2.6255
R57674 VSS.n17105 VSS.n17092 2.6255
R57675 VSS.n17159 VSS.n17158 2.6255
R57676 VSS.n14641 VSS.n14640 2.6255
R57677 VSS.n14629 VSS.n14628 2.6255
R57678 VSS.n14617 VSS.n14616 2.6255
R57679 VSS.n14605 VSS.n14604 2.6255
R57680 VSS.n14593 VSS.n14592 2.6255
R57681 VSS.n14560 VSS.n14559 2.6255
R57682 VSS.n14546 VSS.n14545 2.6255
R57683 VSS.n14532 VSS.n14531 2.6255
R57684 VSS.n14518 VSS.n14517 2.6255
R57685 VSS.n14504 VSS.n14503 2.6255
R57686 VSS.n14490 VSS.n14489 2.6255
R57687 VSS.n14476 VSS.n14475 2.6255
R57688 VSS.n14469 VSS.n14468 2.6255
R57689 VSS.n14483 VSS.n14482 2.6255
R57690 VSS.n14497 VSS.n14496 2.6255
R57691 VSS.n14511 VSS.n14510 2.6255
R57692 VSS.n14525 VSS.n14524 2.6255
R57693 VSS.n14539 VSS.n14538 2.6255
R57694 VSS.n14553 VSS.n14552 2.6255
R57695 VSS.n14587 VSS.n14452 2.6255
R57696 VSS.n14599 VSS.n14598 2.6255
R57697 VSS.n14611 VSS.n14610 2.6255
R57698 VSS.n14623 VSS.n14622 2.6255
R57699 VSS.n14635 VSS.n14634 2.6255
R57700 VSS.n14647 VSS.n14646 2.6255
R57701 VSS.n14776 VSS.n14775 2.6255
R57702 VSS.n14783 VSS.n14782 2.6255
R57703 VSS.n14790 VSS.n14789 2.6255
R57704 VSS.n14797 VSS.n14796 2.6255
R57705 VSS.n14804 VSS.n14803 2.6255
R57706 VSS.n19829 VSS.n19828 2.6255
R57707 VSS.n19815 VSS.n19814 2.6255
R57708 VSS.n19807 VSS.n19806 2.6255
R57709 VSS.n14711 VSS.n14710 2.6255
R57710 VSS.n19797 VSS.n19796 2.6255
R57711 VSS.n19789 VSS.n19788 2.6255
R57712 VSS.n14681 VSS.n14680 2.6255
R57713 VSS.n19780 VSS.n19779 2.6255
R57714 VSS.n14688 VSS.n14687 2.6255
R57715 VSS.n14696 VSS.n14695 2.6255
R57716 VSS.n14704 VSS.n14703 2.6255
R57717 VSS.n14718 VSS.n14717 2.6255
R57718 VSS.n14726 VSS.n14725 2.6255
R57719 VSS.n19822 VSS.n19821 2.6255
R57720 VSS.n14807 VSS.n14735 2.6255
R57721 VSS.n14800 VSS.n14740 2.6255
R57722 VSS.n14793 VSS.n14745 2.6255
R57723 VSS.n14786 VSS.n14750 2.6255
R57724 VSS.n14779 VSS.n14755 2.6255
R57725 VSS.n14772 VSS.n14760 2.6255
R57726 VSS.n17115 VSS.n17114 2.6255
R57727 VSS.n17110 VSS.n17089 2.6255
R57728 VSS.n17064 VSS.n17036 2.6255
R57729 VSS.n17055 VSS.n17041 2.6255
R57730 VSS.n16992 VSS.n14845 2.6255
R57731 VSS.n16998 VSS.n14840 2.6255
R57732 VSS.n16977 VSS.n14851 2.6255
R57733 VSS.n14918 VSS.n14916 2.6255
R57734 VSS.n14910 VSS.n14908 2.6255
R57735 VSS.n16951 VSS.n16949 2.6255
R57736 VSS.n17154 VSS.n17140 2.6255
R57737 VSS.n14926 VSS.n14924 2.6255
R57738 VSS.n16660 VSS.n16646 2.6255
R57739 VSS.n16560 VSS.n16554 2.6255
R57740 VSS.n16565 VSS.n16552 2.6255
R57741 VSS.n16576 VSS.n16547 2.6255
R57742 VSS.n16617 VSS.n16604 2.6255
R57743 VSS.n16628 VSS.n16626 2.6255
R57744 VSS.n16707 VSS.n16705 2.6255
R57745 VSS.n16721 VSS.n16719 2.6255
R57746 VSS.n16735 VSS.n16733 2.6255
R57747 VSS.n16749 VSS.n16747 2.6255
R57748 VSS.n16763 VSS.n16761 2.6255
R57749 VSS.n16777 VSS.n16775 2.6255
R57750 VSS.n16791 VSS.n16789 2.6255
R57751 VSS.n16805 VSS.n16803 2.6255
R57752 VSS.n16819 VSS.n16817 2.6255
R57753 VSS.n16833 VSS.n16831 2.6255
R57754 VSS.n16847 VSS.n16845 2.6255
R57755 VSS.n16867 VSS.n16865 2.6255
R57756 VSS.n16854 VSS.n16850 2.6255
R57757 VSS.n16840 VSS.n16836 2.6255
R57758 VSS.n16826 VSS.n16822 2.6255
R57759 VSS.n16812 VSS.n16808 2.6255
R57760 VSS.n16798 VSS.n16794 2.6255
R57761 VSS.n16784 VSS.n16780 2.6255
R57762 VSS.n16770 VSS.n16766 2.6255
R57763 VSS.n16758 VSS.n16754 2.6255
R57764 VSS.n16742 VSS.n16738 2.6255
R57765 VSS.n16728 VSS.n16724 2.6255
R57766 VSS.n16714 VSS.n16710 2.6255
R57767 VSS.n14946 VSS.n14945 2.6255
R57768 VSS.n14952 VSS.n14951 2.6255
R57769 VSS.n16654 VSS.n16648 2.6255
R57770 VSS.n16622 VSS.n16601 2.6255
R57771 VSS.n16612 VSS.n16606 2.6255
R57772 VSS.n16571 VSS.n16549 2.6255
R57773 VSS.n16521 VSS.n16519 2.6255
R57774 VSS.n16418 VSS.n16416 2.6255
R57775 VSS.n16412 VSS.n16411 2.6255
R57776 VSS.n16406 VSS.n16405 2.6255
R57777 VSS.n16456 VSS.n16455 2.6255
R57778 VSS.n16463 VSS.n16462 2.6255
R57779 VSS.n16470 VSS.n16469 2.6255
R57780 VSS.n16477 VSS.n16476 2.6255
R57781 VSS.n16484 VSS.n16483 2.6255
R57782 VSS.n16491 VSS.n16490 2.6255
R57783 VSS.n16498 VSS.n16497 2.6255
R57784 VSS.n16505 VSS.n16504 2.6255
R57785 VSS.n16510 VSS.n14978 2.6255
R57786 VSS.n16665 VSS.n16664 2.6255
R57787 VSS.n16678 VSS.n16677 2.6255
R57788 VSS.n16516 VSS.n14976 2.6255
R57789 VSS.n18269 VSS.n18234 2.6255
R57790 VSS.n18522 VSS.n18521 2.6255
R57791 VSS.n18536 VSS.n18535 2.6255
R57792 VSS.n18550 VSS.n18549 2.6255
R57793 VSS.n18564 VSS.n18563 2.6255
R57794 VSS.n18578 VSS.n18577 2.6255
R57795 VSS.n18592 VSS.n18591 2.6255
R57796 VSS.n18606 VSS.n18605 2.6255
R57797 VSS.n18620 VSS.n18619 2.6255
R57798 VSS.n18634 VSS.n18633 2.6255
R57799 VSS.n18648 VSS.n18647 2.6255
R57800 VSS.n18665 VSS.n18664 2.6255
R57801 VSS.n18655 VSS.n18654 2.6255
R57802 VSS.n18641 VSS.n18640 2.6255
R57803 VSS.n18627 VSS.n18626 2.6255
R57804 VSS.n18613 VSS.n18612 2.6255
R57805 VSS.n18599 VSS.n18598 2.6255
R57806 VSS.n18585 VSS.n18584 2.6255
R57807 VSS.n18571 VSS.n18570 2.6255
R57808 VSS.n18560 VSS.n18559 2.6255
R57809 VSS.n18543 VSS.n18542 2.6255
R57810 VSS.n18529 VSS.n18528 2.6255
R57811 VSS.n18515 VSS.n18514 2.6255
R57812 VSS.n18508 VSS.n18507 2.6255
R57813 VSS.n18501 VSS.n18500 2.6255
R57814 VSS.n18494 VSS.n18492 2.6255
R57815 VSS.n19421 VSS.n19420 2.6255
R57816 VSS.n19425 VSS.n19424 2.6255
R57817 VSS.n19429 VSS.n19428 2.6255
R57818 VSS.n19433 VSS.n19432 2.6255
R57819 VSS.n19437 VSS.n19436 2.6255
R57820 VSS.n19341 VSS.n19340 2.6255
R57821 VSS.n19334 VSS.n19333 2.6255
R57822 VSS.n19327 VSS.n19326 2.6255
R57823 VSS.n19320 VSS.n19319 2.6255
R57824 VSS.n19313 VSS.n19312 2.6255
R57825 VSS.n19306 VSS.n19305 2.6255
R57826 VSS.n19299 VSS.n19298 2.6255
R57827 VSS.n19292 VSS.n19291 2.6255
R57828 VSS.n19285 VSS.n19284 2.6255
R57829 VSS.n19278 VSS.n19277 2.6255
R57830 VSS.n19271 VSS.n19270 2.6255
R57831 VSS.n19263 VSS.n19262 2.6255
R57832 VSS.n19255 VSS.n19254 2.6255
R57833 VSS.n19247 VSS.n19246 2.6255
R57834 VSS.n19417 VSS.n19415 2.6255
R57835 VSS.n19391 VSS.n19367 2.6255
R57836 VSS.n19402 VSS.n19362 2.6255
R57837 VSS.n19396 VSS.n19364 2.6255
R57838 VSS.n19387 VSS.n19369 2.6255
R57839 VSS.n19412 VSS.n19358 2.6255
R57840 VSS.n19408 VSS.n19360 2.6255
R57841 VSS.n18278 VSS.n18277 2.6255
R57842 VSS.n18282 VSS.n18281 2.6255
R57843 VSS.n18286 VSS.n18285 2.6255
R57844 VSS.n18290 VSS.n18289 2.6255
R57845 VSS.n18294 VSS.n18293 2.6255
R57846 VSS.n18298 VSS.n18297 2.6255
R57847 VSS.n18302 VSS.n18301 2.6255
R57848 VSS.n18309 VSS.n18308 2.6255
R57849 VSS.n18316 VSS.n18315 2.6255
R57850 VSS.n18323 VSS.n18322 2.6255
R57851 VSS.n18330 VSS.n18329 2.6255
R57852 VSS.n18337 VSS.n18336 2.6255
R57853 VSS.n18344 VSS.n18343 2.6255
R57854 VSS.n18351 VSS.n18350 2.6255
R57855 VSS.n18358 VSS.n18357 2.6255
R57856 VSS.n18389 VSS.n18388 2.6255
R57857 VSS.n18382 VSS.n18381 2.6255
R57858 VSS.n18374 VSS.n18373 2.6255
R57859 VSS.n18366 VSS.n18365 2.6255
R57860 VSS.n18419 VSS.n18418 2.6255
R57861 VSS.n18435 VSS.n18434 2.6255
R57862 VSS.n18274 VSS.n18273 2.6255
R57863 VSS.n18257 VSS.n18238 2.6255
R57864 VSS.n18263 VSS.n18236 2.6255
R57865 VSS.n18252 VSS.n18241 2.6255
R57866 VSS.n16961 VSS.n16942 2.6255
R57867 VSS.n16966 VSS.n14855 2.6255
R57868 VSS.n16982 VSS.n14848 2.6255
R57869 VSS.n17003 VSS.n14837 2.6255
R57870 VSS.n17008 VSS.n14835 2.6255
R57871 VSS.n17060 VSS.n17038 2.6255
R57872 VSS.n17105 VSS.n17091 2.6255
R57873 VSS.n17159 VSS.n17138 2.6255
R57874 VSS.n14647 VSS.n14645 2.6255
R57875 VSS.n14635 VSS.n14633 2.6255
R57876 VSS.n14623 VSS.n14621 2.6255
R57877 VSS.n14611 VSS.n14609 2.6255
R57878 VSS.n14599 VSS.n14597 2.6255
R57879 VSS.n14587 VSS.n14451 2.6255
R57880 VSS.n14553 VSS.n14551 2.6255
R57881 VSS.n14539 VSS.n14537 2.6255
R57882 VSS.n14525 VSS.n14523 2.6255
R57883 VSS.n14511 VSS.n14509 2.6255
R57884 VSS.n14497 VSS.n14495 2.6255
R57885 VSS.n14483 VSS.n14481 2.6255
R57886 VSS.n14469 VSS.n14467 2.6255
R57887 VSS.n14476 VSS.n14474 2.6255
R57888 VSS.n14490 VSS.n14488 2.6255
R57889 VSS.n14504 VSS.n14502 2.6255
R57890 VSS.n14518 VSS.n14516 2.6255
R57891 VSS.n14532 VSS.n14530 2.6255
R57892 VSS.n14546 VSS.n14544 2.6255
R57893 VSS.n14560 VSS.n14558 2.6255
R57894 VSS.n14593 VSS.n14591 2.6255
R57895 VSS.n14605 VSS.n14603 2.6255
R57896 VSS.n14617 VSS.n14615 2.6255
R57897 VSS.n14629 VSS.n14627 2.6255
R57898 VSS.n14641 VSS.n14639 2.6255
R57899 VSS.n14653 VSS.n14652 2.6255
R57900 VSS.n14772 VSS.n14759 2.6255
R57901 VSS.n14779 VSS.n14754 2.6255
R57902 VSS.n14786 VSS.n14749 2.6255
R57903 VSS.n14793 VSS.n14744 2.6255
R57904 VSS.n14800 VSS.n14739 2.6255
R57905 VSS.n14807 VSS.n14734 2.6255
R57906 VSS.n19822 VSS.n19820 2.6255
R57907 VSS.n14726 VSS.n14724 2.6255
R57908 VSS.n14718 VSS.n14716 2.6255
R57909 VSS.n14704 VSS.n14702 2.6255
R57910 VSS.n14696 VSS.n14694 2.6255
R57911 VSS.n14688 VSS.n14686 2.6255
R57912 VSS.n19780 VSS.n19778 2.6255
R57913 VSS.n14681 VSS.n14679 2.6255
R57914 VSS.n19789 VSS.n19787 2.6255
R57915 VSS.n19797 VSS.n19795 2.6255
R57916 VSS.n14711 VSS.n14709 2.6255
R57917 VSS.n19807 VSS.n19805 2.6255
R57918 VSS.n19815 VSS.n19813 2.6255
R57919 VSS.n19829 VSS.n19827 2.6255
R57920 VSS.n14804 VSS.n14737 2.6255
R57921 VSS.n14797 VSS.n14742 2.6255
R57922 VSS.n14790 VSS.n14747 2.6255
R57923 VSS.n14783 VSS.n14752 2.6255
R57924 VSS.n14776 VSS.n14757 2.6255
R57925 VSS.n14769 VSS.n14768 2.6255
R57926 VSS.n17154 VSS.n17153 2.6255
R57927 VSS.n17148 VSS.n17147 2.6255
R57928 VSS.n17115 VSS.n17086 2.6255
R57929 VSS.n17110 VSS.n17088 2.6255
R57930 VSS.n17100 VSS.n17094 2.6255
R57931 VSS.n17064 VSS.n17035 2.6255
R57932 VSS.n17055 VSS.n17054 2.6255
R57933 VSS.n17049 VSS.n17048 2.6255
R57934 VSS.n16992 VSS.n14843 2.6255
R57935 VSS.n16998 VSS.n16997 2.6255
R57936 VSS.n16988 VSS.n16987 2.6255
R57937 VSS.n16977 VSS.n16976 2.6255
R57938 VSS.n16971 VSS.n16970 2.6255
R57939 VSS.n16956 VSS.n16945 2.6255
R57940 VSS.n16951 VSS.n16948 2.6255
R57941 VSS.n14910 VSS.n14909 2.6255
R57942 VSS.n14926 VSS.n14925 2.6255
R57943 VSS.n14918 VSS.n14917 2.6255
R57944 VSS.n16418 VSS.n16417 2.6255
R57945 VSS.n16412 VSS.n16410 2.6255
R57946 VSS.n16406 VSS.n16404 2.6255
R57947 VSS.n16456 VSS.n16451 2.6255
R57948 VSS.n16463 VSS.n16458 2.6255
R57949 VSS.n16470 VSS.n16465 2.6255
R57950 VSS.n16477 VSS.n16472 2.6255
R57951 VSS.n16484 VSS.n16479 2.6255
R57952 VSS.n16491 VSS.n16486 2.6255
R57953 VSS.n16498 VSS.n16493 2.6255
R57954 VSS.n16505 VSS.n14980 2.6255
R57955 VSS.n16565 VSS.n16551 2.6255
R57956 VSS.n16576 VSS.n16575 2.6255
R57957 VSS.n16622 VSS.n16600 2.6255
R57958 VSS.n16628 VSS.n16627 2.6255
R57959 VSS.n16665 VSS.n16644 2.6255
R57960 VSS.n16678 VSS.n16673 2.6255
R57961 VSS.n14952 VSS.n14950 2.6255
R57962 VSS.n14946 VSS.n14944 2.6255
R57963 VSS.n16707 VSS.n16706 2.6255
R57964 VSS.n16714 VSS.n16709 2.6255
R57965 VSS.n16721 VSS.n16720 2.6255
R57966 VSS.n16728 VSS.n16723 2.6255
R57967 VSS.n16735 VSS.n16734 2.6255
R57968 VSS.n16742 VSS.n16737 2.6255
R57969 VSS.n16749 VSS.n16748 2.6255
R57970 VSS.n16758 VSS.n16753 2.6255
R57971 VSS.n16763 VSS.n16762 2.6255
R57972 VSS.n16770 VSS.n16765 2.6255
R57973 VSS.n16777 VSS.n16776 2.6255
R57974 VSS.n16784 VSS.n16779 2.6255
R57975 VSS.n16791 VSS.n16790 2.6255
R57976 VSS.n16798 VSS.n16793 2.6255
R57977 VSS.n16805 VSS.n16804 2.6255
R57978 VSS.n16812 VSS.n16807 2.6255
R57979 VSS.n16819 VSS.n16818 2.6255
R57980 VSS.n16826 VSS.n16821 2.6255
R57981 VSS.n16833 VSS.n16832 2.6255
R57982 VSS.n16840 VSS.n16835 2.6255
R57983 VSS.n16847 VSS.n16846 2.6255
R57984 VSS.n16854 VSS.n16849 2.6255
R57985 VSS.n16867 VSS.n16866 2.6255
R57986 VSS.n14958 VSS.n14956 2.6255
R57987 VSS.n16660 VSS.n16659 2.6255
R57988 VSS.n16654 VSS.n16653 2.6255
R57989 VSS.n16617 VSS.n16603 2.6255
R57990 VSS.n16612 VSS.n16611 2.6255
R57991 VSS.n16571 VSS.n16570 2.6255
R57992 VSS.n16521 VSS.n16520 2.6255
R57993 VSS.n16516 VSS.n16515 2.6255
R57994 VSS.n16510 VSS.n16509 2.6255
R57995 VSS.n16560 VSS.n16559 2.6255
R57996 VSS.n18515 VSS.n18513 2.6255
R57997 VSS.n18529 VSS.n18527 2.6255
R57998 VSS.n18543 VSS.n18541 2.6255
R57999 VSS.n18560 VSS.n18558 2.6255
R58000 VSS.n18571 VSS.n18569 2.6255
R58001 VSS.n18585 VSS.n18583 2.6255
R58002 VSS.n18599 VSS.n18597 2.6255
R58003 VSS.n18613 VSS.n18611 2.6255
R58004 VSS.n18627 VSS.n18625 2.6255
R58005 VSS.n18641 VSS.n18639 2.6255
R58006 VSS.n18655 VSS.n18653 2.6255
R58007 VSS.n18665 VSS.n18663 2.6255
R58008 VSS.n18648 VSS.n18646 2.6255
R58009 VSS.n18634 VSS.n18632 2.6255
R58010 VSS.n18620 VSS.n18618 2.6255
R58011 VSS.n18606 VSS.n18604 2.6255
R58012 VSS.n18592 VSS.n18590 2.6255
R58013 VSS.n18578 VSS.n18576 2.6255
R58014 VSS.n18564 VSS.n18556 2.6255
R58015 VSS.n18550 VSS.n18548 2.6255
R58016 VSS.n18536 VSS.n18534 2.6255
R58017 VSS.n18522 VSS.n18520 2.6255
R58018 VSS.n18508 VSS.n18506 2.6255
R58019 VSS.n18501 VSS.n18499 2.6255
R58020 VSS.n18494 VSS.n18493 2.6255
R58021 VSS.n18487 VSS.n18480 2.6255
R58022 VSS.n19247 VSS.n19245 2.6255
R58023 VSS.n19255 VSS.n19253 2.6255
R58024 VSS.n19263 VSS.n19261 2.6255
R58025 VSS.n19271 VSS.n19269 2.6255
R58026 VSS.n19278 VSS.n19276 2.6255
R58027 VSS.n19285 VSS.n19283 2.6255
R58028 VSS.n19292 VSS.n19290 2.6255
R58029 VSS.n19299 VSS.n19297 2.6255
R58030 VSS.n19306 VSS.n19304 2.6255
R58031 VSS.n19313 VSS.n19311 2.6255
R58032 VSS.n19320 VSS.n19318 2.6255
R58033 VSS.n19327 VSS.n19325 2.6255
R58034 VSS.n19334 VSS.n19332 2.6255
R58035 VSS.n19341 VSS.n19339 2.6255
R58036 VSS.n19437 VSS.n19346 2.6255
R58037 VSS.n19433 VSS.n19348 2.6255
R58038 VSS.n19429 VSS.n19350 2.6255
R58039 VSS.n19425 VSS.n19352 2.6255
R58040 VSS.n19421 VSS.n19354 2.6255
R58041 VSS.n19417 VSS.n19416 2.6255
R58042 VSS.n19396 VSS.n19395 2.6255
R58043 VSS.n19391 VSS.n19366 2.6255
R58044 VSS.n19387 VSS.n19386 2.6255
R58045 VSS.n19402 VSS.n19401 2.6255
R58046 VSS.n19408 VSS.n19407 2.6255
R58047 VSS.n19412 VSS.n19357 2.6255
R58048 VSS.n18435 VSS.n18433 2.6255
R58049 VSS.n18419 VSS.n18417 2.6255
R58050 VSS.n18366 VSS.n18364 2.6255
R58051 VSS.n18374 VSS.n18372 2.6255
R58052 VSS.n18382 VSS.n18380 2.6255
R58053 VSS.n18389 VSS.n18387 2.6255
R58054 VSS.n18358 VSS.n18356 2.6255
R58055 VSS.n18351 VSS.n18349 2.6255
R58056 VSS.n18344 VSS.n18342 2.6255
R58057 VSS.n18337 VSS.n18335 2.6255
R58058 VSS.n18330 VSS.n18328 2.6255
R58059 VSS.n18323 VSS.n18321 2.6255
R58060 VSS.n18316 VSS.n18314 2.6255
R58061 VSS.n18309 VSS.n18307 2.6255
R58062 VSS.n18302 VSS.n18218 2.6255
R58063 VSS.n18298 VSS.n18220 2.6255
R58064 VSS.n18294 VSS.n18222 2.6255
R58065 VSS.n18290 VSS.n18224 2.6255
R58066 VSS.n18286 VSS.n18226 2.6255
R58067 VSS.n18282 VSS.n18228 2.6255
R58068 VSS.n18278 VSS.n18230 2.6255
R58069 VSS.n18274 VSS.n18232 2.6255
R58070 VSS.n18263 VSS.n18262 2.6255
R58071 VSS.n18269 VSS.n18268 2.6255
R58072 VSS.n18257 VSS.n18256 2.6255
R58073 VSS.n18252 VSS.n18240 2.6255
R58074 VSS.n15869 VSS.n15867 2.6255
R58075 VSS.n15854 VSS.n15853 2.6255
R58076 VSS.n15850 VSS.n15845 2.6255
R58077 VSS.n15843 VSS.n15839 2.6255
R58078 VSS.n15836 VSS.n15831 2.6255
R58079 VSS.n15829 VSS.n15825 2.6255
R58080 VSS.n15822 VSS.n15817 2.6255
R58081 VSS.n15813 VSS.n15812 2.6255
R58082 VSS.n15808 VSS.n15803 2.6255
R58083 VSS.n15801 VSS.n15797 2.6255
R58084 VSS.n15794 VSS.n15789 2.6255
R58085 VSS.n15787 VSS.n15783 2.6255
R58086 VSS.n15780 VSS.n15775 2.6255
R58087 VSS.n15773 VSS.n15769 2.6255
R58088 VSS.n15766 VSS.n15761 2.6255
R58089 VSS.n15759 VSS.n15755 2.6255
R58090 VSS.n15752 VSS.n15747 2.6255
R58091 VSS.n15745 VSS.n15741 2.6255
R58092 VSS.n15738 VSS.n15733 2.6255
R58093 VSS.n15731 VSS.n15727 2.6255
R58094 VSS.n15724 VSS.n15719 2.6255
R58095 VSS.n15717 VSS.n15713 2.6255
R58096 VSS.n15717 VSS.n15712 2.6255
R58097 VSS.n15724 VSS.n15723 2.6255
R58098 VSS.n15731 VSS.n15726 2.6255
R58099 VSS.n15738 VSS.n15737 2.6255
R58100 VSS.n15745 VSS.n15740 2.6255
R58101 VSS.n15752 VSS.n15751 2.6255
R58102 VSS.n15759 VSS.n15754 2.6255
R58103 VSS.n15766 VSS.n15765 2.6255
R58104 VSS.n15773 VSS.n15768 2.6255
R58105 VSS.n15780 VSS.n15779 2.6255
R58106 VSS.n15787 VSS.n15782 2.6255
R58107 VSS.n15794 VSS.n15793 2.6255
R58108 VSS.n15801 VSS.n15796 2.6255
R58109 VSS.n15808 VSS.n15807 2.6255
R58110 VSS.n15813 VSS.n15811 2.6255
R58111 VSS.n15822 VSS.n15821 2.6255
R58112 VSS.n15829 VSS.n15824 2.6255
R58113 VSS.n15836 VSS.n15835 2.6255
R58114 VSS.n15843 VSS.n15838 2.6255
R58115 VSS.n15850 VSS.n15849 2.6255
R58116 VSS.n15854 VSS.n15852 2.6255
R58117 VSS.n15869 VSS.n15868 2.6255
R58118 VSS.n15875 VSS.n15874 2.6255
R58119 VSS.n15875 VSS.n15873 2.6255
R58120 VSS.n15881 VSS.n15879 2.6255
R58121 VSS.n15881 VSS.n15880 2.6255
R58122 VSS.n15887 VSS.n15885 2.6255
R58123 VSS.n15887 VSS.n15886 2.6255
R58124 VSS.n15893 VSS.n15891 2.6255
R58125 VSS.n15893 VSS.n15892 2.6255
R58126 VSS.n16298 VSS.n16294 2.61893
R58127 VSS.n1381 VSS.n1380 2.61893
R58128 VSS.n5701 VSS.n5641 2.61893
R58129 VSS.n20970 VSS.n20905 2.61893
R58130 VSS.n1422 VSS.n1421 2.6005
R58131 VSS.n1421 VSS.n1420 2.6005
R58132 VSS.n906 VSS.n905 2.6005
R58133 VSS.n899 VSS.n898 2.6005
R58134 VSS.n896 VSS.n895 2.6005
R58135 VSS.n891 VSS.n890 2.6005
R58136 VSS.n1492 VSS.n1491 2.6005
R58137 VSS.n1489 VSS.n1488 2.6005
R58138 VSS.n1486 VSS.n1485 2.6005
R58139 VSS.n1483 VSS.n1482 2.6005
R58140 VSS.n15209 VSS.n15208 2.6005
R58141 VSS.n15202 VSS.n15201 2.6005
R58142 VSS.n15215 VSS.n15214 2.6005
R58143 VSS.n15212 VSS.n15211 2.6005
R58144 VSS.n15931 VSS.n15930 2.6005
R58145 VSS.n15928 VSS.n15927 2.6005
R58146 VSS.n15925 VSS.n15924 2.6005
R58147 VSS.n15920 VSS.n15919 2.6005
R58148 VSS.n16333 VSS.n16332 2.6005
R58149 VSS.n16336 VSS.n16335 2.6005
R58150 VSS.n16335 VSS.n16334 2.6005
R58151 VSS.n1431 VSS.n1430 2.6005
R58152 VSS.n1430 VSS.n1429 2.6005
R58153 VSS.n16343 VSS.n16342 2.6005
R58154 VSS.n16342 VSS.n16341 2.6005
R58155 VSS.n1424 VSS.n1423 2.6005
R58156 VSS.n1378 VSS.n1377 2.6005
R58157 VSS.n1385 VSS.n1384 2.6005
R58158 VSS.n16302 VSS.n16301 2.6005
R58159 VSS.n16297 VSS.n16296 2.6005
R58160 VSS.n16262 VSS.n16261 2.6005
R58161 VSS.n1351 VSS.n1350 2.6005
R58162 VSS.n16267 VSS.n16266 2.6005
R58163 VSS.n1346 VSS.n1345 2.6005
R58164 VSS.n15971 VSS.n15970 2.6005
R58165 VSS.n15975 VSS.n15974 2.6005
R58166 VSS.n15979 VSS.n15978 2.6005
R58167 VSS.n15983 VSS.n15982 2.6005
R58168 VSS.n15576 VSS.n15575 2.6005
R58169 VSS.n15581 VSS.n15580 2.6005
R58170 VSS.n15262 VSS.n15261 2.6005
R58171 VSS.n15266 VSS.n15265 2.6005
R58172 VSS.n1553 VSS.n1552 2.6005
R58173 VSS.n957 VSS.n956 2.6005
R58174 VSS.n949 VSS.n948 2.6005
R58175 VSS.n1555 VSS.n1554 2.6005
R58176 VSS.n1559 VSS.n1558 2.6005
R58177 VSS.n1561 VSS.n1560 2.6005
R58178 VSS.n944 VSS.n943 2.6005
R58179 VSS.n952 VSS.n951 2.6005
R58180 VSS.n20923 VSS.n20922 2.6005
R58181 VSS.n20913 VSS.n20912 2.6005
R58182 VSS.n1013 VSS.n1012 2.6005
R58183 VSS.n1009 VSS.n1008 2.6005
R58184 VSS.n1045 VSS.n1044 2.6005
R58185 VSS.n1621 VSS.n1620 2.6005
R58186 VSS.n1627 VSS.n1626 2.6005
R58187 VSS.n15303 VSS.n15302 2.6005
R58188 VSS.n15301 VSS.n15300 2.6005
R58189 VSS.n15308 VSS.n15307 2.6005
R58190 VSS.n16040 VSS.n16039 2.6005
R58191 VSS.n16031 VSS.n16030 2.6005
R58192 VSS.n5529 VSS.n5528 2.6005
R58193 VSS.n5647 VSS.n5646 2.6005
R58194 VSS.n5656 VSS.n5655 2.6005
R58195 VSS.n5650 VSS.n5649 2.6005
R58196 VSS.n5535 VSS.n5534 2.6005
R58197 VSS.n16076 VSS.n16075 2.6005
R58198 VSS.n16045 VSS.n16044 2.6005
R58199 VSS.n16034 VSS.n16033 2.6005
R58200 VSS.n1614 VSS.n1613 2.6005
R58201 VSS.n1041 VSS.n1040 2.6005
R58202 VSS.n1006 VSS.n1005 2.6005
R58203 VSS.n1019 VSS.n1018 2.6005
R58204 VSS.n20907 VSS.n20906 2.6005
R58205 VSS.n20917 VSS.n20916 2.6005
R58206 VSS.n20933 VSS.n20932 2.6005
R58207 VSS.n5700 VSS.n5699 2.6005
R58208 VSS.n5664 VSS.n5663 2.6005
R58209 VSS.n5696 VSS.n5695 2.6005
R58210 VSS.n20965 VSS.n20964 2.6005
R58211 VSS.n20969 VSS.n20968 2.6005
R58212 VSS.n5705 VSS.n5704 2.6005
R58213 VSS.n20976 VSS.n20975 2.6005
R58214 VSS.n20975 VSS.n20974 2.6005
R58215 VSS.n5751 VSS.n5750 2.6005
R58216 VSS.n1212 VSS.n1211 2.6005
R58217 VSS.n20903 VSS.n20902 2.6005
R58218 VSS.n20902 VSS.n20901 2.6005
R58219 VSS.n5765 VSS.n5764 2.6005
R58220 VSS.n5764 VSS.n5763 2.6005
R58221 VSS.n1218 VSS.n1217 2.6005
R58222 VSS.n5757 VSS.n5756 2.6005
R58223 VSS.n5756 VSS.n5755 2.6005
R58224 VSS.n1306 VSS.n1305 2.6005
R58225 VSS.n968 VSS.n967 2.6005
R58226 VSS.n960 VSS.n959 2.6005
R58227 VSS.n1579 VSS.n1578 2.6005
R58228 VSS.n1572 VSS.n1571 2.6005
R58229 VSS.n15272 VSS.n15271 2.6005
R58230 VSS.n15559 VSS.n15558 2.6005
R58231 VSS.n16000 VSS.n15999 2.6005
R58232 VSS.n15997 VSS.n15996 2.6005
R58233 VSS.n15994 VSS.n15993 2.6005
R58234 VSS.n15989 VSS.n15988 2.6005
R58235 VSS.n5485 VSS.n5484 2.6005
R58236 VSS.n5488 VSS.n5487 2.6005
R58237 VSS.n5481 VSS.n5480 2.6005
R58238 VSS.n5498 VSS.n5497 2.6005
R58239 VSS.n5495 VSS.n5494 2.6005
R58240 VSS.n1303 VSS.n1302 2.6005
R58241 VSS.n964 VSS.n963 2.6005
R58242 VSS.n1576 VSS.n1575 2.6005
R58243 VSS.n1570 VSS.n1569 2.6005
R58244 VSS.n15276 VSS.n15275 2.6005
R58245 VSS.n15270 VSS.n15269 2.6005
R58246 VSS.n21178 VSS.n21177 2.6005
R58247 VSS.n20891 VSS.n20890 2.6005
R58248 VSS.n20877 VSS.n20876 2.6005
R58249 VSS.n20887 VSS.n20886 2.6005
R58250 VSS.n10329 VSS.n10328 2.6005
R58251 VSS.n12383 VSS.n12382 2.6005
R58252 VSS.n14663 VSS.n14662 2.6005
R58253 VSS.n17172 VSS.n17171 2.6005
R58254 VSS.n14937 VSS.n14936 2.6005
R58255 VSS.n14966 VSS.n14965 2.6005
R58256 VSS.n16426 VSS.n16425 2.6005
R58257 VSS.n19378 VSS.n19377 2.6005
R58258 VSS.n19008 VSS.n19007 2.6005
R58259 VSS.n18245 VSS.n18244 2.6005
R58260 VSS.n14298 VSS.n14297 2.6005
R58261 VSS.n14297 VSS.n14296 2.6005
R58262 VSS.n14286 VSS.n14285 2.6005
R58263 VSS.n35 VSS.n34 2.6005
R58264 VSS.n14261 VSS.n14260 2.6005
R58265 VSS.n14260 VSS.n14259 2.6005
R58266 VSS.n14662 VSS.n14660 2.54004
R58267 VSS.n14662 VSS.n14661 2.54004
R58268 VSS.n17174 VSS.n17172 2.54004
R58269 VSS.n14936 VSS.n14934 2.54004
R58270 VSS.n14936 VSS.n14935 2.54004
R58271 VSS.n19377 VSS.n19375 2.54004
R58272 VSS.n19377 VSS.n19376 2.54004
R58273 VSS.n12005 VSS.n12003 2.52606
R58274 VSS.n8854 VSS.n8853 2.52606
R58275 VSS.n5886 VSS.n5885 2.41287
R58276 VSS.n14247 VSS.n14243 2.41287
R58277 VSS.n13547 VSS.n13543 2.41287
R58278 VSS.n17178 VSS.n11751 2.41287
R58279 VSS.n14318 VSS.n14314 2.41287
R58280 VSS.n14305 VSS.n14290 2.41287
R58281 VSS.n2417 VSS.n2416 2.41287
R58282 VSS.n2382 VSS.n2381 2.41287
R58283 VSS.n2460 VSS.n2459 2.41287
R58284 VSS.n2387 VSS.n2386 2.41287
R58285 VSS.n2412 VSS.n2411 2.41287
R58286 VSS.n2452 VSS.n2451 2.41287
R58287 VSS.n2465 VSS.n2464 2.41287
R58288 VSS.n3896 VSS.n3895 2.41287
R58289 VSS.n176 VSS.n175 2.41287
R58290 VSS.n173 VSS.n172 2.41287
R58291 VSS.n3891 VSS.n3890 2.41287
R58292 VSS.n3924 VSS.n3923 2.41287
R58293 VSS.n3929 VSS.n3928 2.41287
R58294 VSS.n2498 VSS.n2497 2.41287
R58295 VSS.n2503 VSS.n2502 2.41287
R58296 VSS.n3889 VSS.n3888 2.41287
R58297 VSS.n5896 VSS.n5895 2.41287
R58298 VSS.n5889 VSS.n5888 2.41287
R58299 VSS.n5416 VSS.n5415 2.41287
R58300 VSS.n5466 VSS.n5465 2.41287
R58301 VSS.n5461 VSS.n5460 2.41287
R58302 VSS.n5426 VSS.n5425 2.41287
R58303 VSS.n5421 VSS.n5420 2.41287
R58304 VSS.n4861 VSS.n4860 2.41287
R58305 VSS.n4911 VSS.n4910 2.41287
R58306 VSS.n4906 VSS.n4905 2.41287
R58307 VSS.n4871 VSS.n4870 2.41287
R58308 VSS.n4866 VSS.n4865 2.41287
R58309 VSS.n4799 VSS.n4798 2.41287
R58310 VSS.n4847 VSS.n4846 2.41287
R58311 VSS.n4842 VSS.n4841 2.41287
R58312 VSS.n4809 VSS.n4808 2.41287
R58313 VSS.n4804 VSS.n4803 2.41287
R58314 VSS.n14305 VSS.n14304 2.41287
R58315 VSS.n14318 VSS.n14317 2.41287
R58316 VSS.n17178 VSS.n17177 2.41287
R58317 VSS.n13547 VSS.n13546 2.41287
R58318 VSS.n14247 VSS.n14246 2.41287
R58319 VSS.n17251 VSS.n17250 2.41287
R58320 VSS.n17299 VSS.n17298 2.41287
R58321 VSS.n17294 VSS.n17293 2.41287
R58322 VSS.n17261 VSS.n17260 2.41287
R58323 VSS.n17256 VSS.n17255 2.41287
R58324 VSS.n2380 VSS.n2379 2.41287
R58325 VSS.n181 VSS.n180 2.41287
R58326 VSS.n13655 VSS.n13654 2.41287
R58327 VSS.n22228 VSS.n22227 2.41287
R58328 VSS.n22227 VSS.n22226 2.41287
R58329 VSS.n22169 VSS.n22168 2.41287
R58330 VSS.n22168 VSS.n22167 2.41287
R58331 VSS.n22160 VSS.n22159 2.41287
R58332 VSS.n22159 VSS.n22158 2.41287
R58333 VSS.n22145 VSS.n22144 2.41287
R58334 VSS.n22144 VSS.n22143 2.41287
R58335 VSS.n22133 VSS.n22132 2.41287
R58336 VSS.n22132 VSS.n22131 2.41287
R58337 VSS.n22123 VSS.n22122 2.41287
R58338 VSS.n22127 VSS.n22126 2.41287
R58339 VSS.n22139 VSS.n22138 2.41287
R58340 VSS.n22138 VSS.n22137 2.41287
R58341 VSS.n22151 VSS.n22150 2.41287
R58342 VSS.n22150 VSS.n22149 2.41287
R58343 VSS.n22173 VSS.n22166 2.41287
R58344 VSS.n22166 VSS.n22165 2.41287
R58345 VSS.n22245 VSS.n22244 2.41287
R58346 VSS.n22244 VSS.n22243 2.41287
R58347 VSS.n22251 VSS.n22250 2.41287
R58348 VSS.n22250 VSS.n22249 2.41287
R58349 VSS.n22236 VSS.n22235 2.41287
R58350 VSS.n22235 VSS.n22234 2.41287
R58351 VSS.n22219 VSS.n22218 2.41287
R58352 VSS.n22215 VSS.n22214 2.41287
R58353 VSS.n22211 VSS.n22210 2.41287
R58354 VSS.n22207 VSS.n22206 2.41287
R58355 VSS.n22203 VSS.n22202 2.41287
R58356 VSS.n22199 VSS.n22198 2.41287
R58357 VSS.n22195 VSS.n22194 2.41287
R58358 VSS.n22191 VSS.n22190 2.41287
R58359 VSS.n22187 VSS.n22186 2.41287
R58360 VSS.n22183 VSS.n22182 2.41287
R58361 VSS.n13642 VSS.n13641 2.41287
R58362 VSS.n22222 VSS.n22181 2.41287
R58363 VSS.n14272 VSS.n14271 2.41287
R58364 VSS.n14271 VSS.n14270 2.41287
R58365 VSS.n21942 VSS.n21938 2.41287
R58366 VSS.n13609 VSS.n13608 2.41287
R58367 VSS.n13608 VSS.n13607 2.41287
R58368 VSS.n14276 VSS.n13556 2.41287
R58369 VSS.n13556 VSS.n13555 2.41287
R58370 VSS.n14308 VSS.n14307 2.41287
R58371 VSS.n14307 VSS.n14306 2.41287
R58372 VSS.n14321 VSS.n14320 2.41287
R58373 VSS.n14320 VSS.n14319 2.41287
R58374 VSS.n14327 VSS.n14326 2.41287
R58375 VSS.n14328 VSS.n14327 2.41287
R58376 VSS.n13550 VSS.n13549 2.41287
R58377 VSS.n13549 VSS.n13548 2.41287
R58378 VSS.n14250 VSS.n14249 2.41287
R58379 VSS.n14249 VSS.n14248 2.41287
R58380 VSS.n13578 VSS.n13577 2.41287
R58381 VSS.n13577 VSS.n13576 2.41287
R58382 VSS.n13584 VSS.n13583 2.41287
R58383 VSS.n13583 VSS.n13582 2.41287
R58384 VSS.n13590 VSS.n13589 2.41287
R58385 VSS.n13589 VSS.n13588 2.41287
R58386 VSS.n13596 VSS.n13595 2.41287
R58387 VSS.n13595 VSS.n13594 2.41287
R58388 VSS.n13602 VSS.n13601 2.41287
R58389 VSS.n13601 VSS.n13600 2.41287
R58390 VSS.n21984 VSS.n21983 2.41287
R58391 VSS.n21946 VSS.n21945 2.41287
R58392 VSS.n21959 VSS.n21958 2.41287
R58393 VSS.n21953 VSS.n21952 2.41287
R58394 VSS.n21972 VSS.n21971 2.41287
R58395 VSS.n21976 VSS.n21975 2.41287
R58396 VSS.n21966 VSS.n21965 2.41287
R58397 VSS.n7 VSS.n6 2.41287
R58398 VSS.n11 VSS.n10 2.41287
R58399 VSS.n15 VSS.n14 2.41287
R58400 VSS.n19 VSS.n18 2.41287
R58401 VSS.n24 VSS.n23 2.41287
R58402 VSS.n23 VSS.n22 2.41287
R58403 VSS.n21938 VSS.n21937 2.41287
R58404 VSS.n5471 VSS.n5416 2.41258
R58405 VSS.n4916 VSS.n4861 2.41258
R58406 VSS.n4852 VSS.n4799 2.41258
R58407 VSS.n14304 VSS.n14303 2.41258
R58408 VSS.n17304 VSS.n17251 2.41258
R58409 VSS.n2422 VSS.n2380 2.41258
R58410 VSS.n2508 VSS.n2452 2.41258
R58411 VSS.n3934 VSS.n3889 2.41258
R58412 VSS.n5897 VSS.n5896 2.41193
R58413 VSS.n174 VSS.n173 2.41193
R58414 VSS.n8881 VSS.n8879 2.41108
R58415 VSS.n8877 VSS.n8876 2.41079
R58416 VSS.n11992 VSS.n11991 2.41079
R58417 VSS.n8869 VSS.n8867 2.40893
R58418 VSS.n11984 VSS.n11982 2.40888
R58419 VSS.n11998 VSS.n11996 2.37114
R58420 VSS.n20926 VSS.n20925 2.35296
R58421 VSS.n20880 VSS.n20879 2.35296
R58422 VSS.n5643 VSS.n5642 2.32427
R58423 VSS.n5492 VSS.n5491 2.32427
R58424 VSS.n201 VSS.n200 2.3132
R58425 VSS.n15691 VSS.n15680 2.3132
R58426 VSS.n16145 VSS.n16144 2.25091
R58427 VSS.n1125 VSS.n1124 2.25091
R58428 VSS.n15399 VSS.n15286 2.25089
R58429 VSS.n1715 VSS.n1599 2.25089
R58430 VSS.n16133 VSS.n16019 2.25087
R58431 VSS.n1113 VSS.n1000 2.25087
R58432 VSS.n15393 VSS.n15297 2.25084
R58433 VSS.n1709 VSS.n1610 2.25084
R58434 VSS.n5563 VSS.n5538 2.25082
R58435 VSS.n16079 VSS.n16078 2.25082
R58436 VSS.n1058 VSS.n1022 2.25082
R58437 VSS.n15336 VSS.n15311 2.25079
R58438 VSS.n1652 VSS.n1629 2.25079
R58439 VSS.n8919 VSS.n8914 2.25078
R58440 VSS.n8919 VSS.n8904 2.25073
R58441 VSS.n8992 VSS.n8985 2.25073
R58442 VSS.n8919 VSS.n8912 2.25069
R58443 VSS.n17394 VSS.n17393 2.25065
R58444 VSS.n8992 VSS.n8973 2.25065
R58445 VSS.n8919 VSS.n8918 2.25051
R58446 VSS.n8841 VSS.n8840 2.25051
R58447 VSS.n15582 VSS.n15577 2.2505
R58448 VSS.n15579 VSS.n15578 2.2505
R58449 VSS.n15268 VSS.n15267 2.2505
R58450 VSS.n15264 VSS.n15263 2.2505
R58451 VSS.n15207 VSS.n15204 2.2505
R58452 VSS.n15210 VSS.n15203 2.2505
R58453 VSS.n15218 VSS.n15217 2.2505
R58454 VSS.n15216 VSS.n15213 2.2505
R58455 VSS.n15305 VSS.n15304 2.2505
R58456 VSS.n15299 VSS.n15298 2.2505
R58457 VSS.n5658 VSS.n5643 2.2505
R58458 VSS.n5653 VSS.n5652 2.2505
R58459 VSS.n5648 VSS.n5644 2.2505
R58460 VSS.n5538 VSS.n5537 2.2505
R58461 VSS.n5532 VSS.n5531 2.2505
R58462 VSS.n15311 VSS.n15310 2.2505
R58463 VSS.n15315 VSS.n15314 2.2505
R58464 VSS.n16243 VSS.n16242 2.2505
R58465 VSS.n15977 VSS.n15976 2.2505
R58466 VSS.n15973 VSS.n15972 2.2505
R58467 VSS.n15985 VSS.n15984 2.2505
R58468 VSS.n15981 VSS.n15980 2.2505
R58469 VSS.n15934 VSS.n15933 2.2505
R58470 VSS.n15932 VSS.n15929 2.2505
R58471 VSS.n15923 VSS.n15922 2.2505
R58472 VSS.n15926 VSS.n15921 2.2505
R58473 VSS.n15918 VSS.n15917 2.2505
R58474 VSS.n16078 VSS.n16074 2.2505
R58475 VSS.n16028 VSS.n16027 2.2505
R58476 VSS.n16047 VSS.n16046 2.2505
R58477 VSS.n16042 VSS.n16032 2.2505
R58478 VSS.n16037 VSS.n16036 2.2505
R58479 VSS.n15391 VSS.n15390 2.2505
R58480 VSS.n15278 VSS.n15277 2.2505
R58481 VSS.n15280 VSS.n15279 2.2505
R58482 VSS.n15274 VSS.n15273 2.2505
R58483 VSS.n15561 VSS.n15560 2.2505
R58484 VSS.n16003 VSS.n16002 2.2505
R58485 VSS.n16001 VSS.n15998 2.2505
R58486 VSS.n15992 VSS.n15991 2.2505
R58487 VSS.n15995 VSS.n15990 2.2505
R58488 VSS.n15987 VSS.n15986 2.2505
R58489 VSS.n5486 VSS.n5483 2.2505
R58490 VSS.n5489 VSS.n5482 2.2505
R58491 VSS.n5479 VSS.n5478 2.2505
R58492 VSS.n5499 VSS.n5496 2.2505
R58493 VSS.n5493 VSS.n5492 2.2505
R58494 VSS.n21180 VSS.n21179 2.2505
R58495 VSS.n20892 VSS.n20889 2.2505
R58496 VSS.n20875 VSS.n20874 2.2505
R58497 VSS.n20888 VSS.n20878 2.2505
R58498 VSS.n20885 VSS.n20880 2.2505
R58499 VSS.n21001 VSS.n21000 2.2505
R58500 VSS.n20910 VSS.n20909 2.2505
R58501 VSS.n20915 VSS.n20914 2.2505
R58502 VSS.n20920 VSS.n20919 2.2505
R58503 VSS.n20927 VSS.n20926 2.2505
R58504 VSS.n1307 VSS.n1304 2.2505
R58505 VSS.n970 VSS.n969 2.2505
R58506 VSS.n962 VSS.n961 2.2505
R58507 VSS.n966 VSS.n965 2.2505
R58508 VSS.n1313 VSS.n1312 2.2505
R58509 VSS.n904 VSS.n903 2.2505
R58510 VSS.n907 VSS.n900 2.2505
R58511 VSS.n894 VSS.n893 2.2505
R58512 VSS.n897 VSS.n892 2.2505
R58513 VSS.n1455 VSS.n1454 2.2505
R58514 VSS.n1320 VSS.n1319 2.2505
R58515 VSS.n950 VSS.n945 2.2505
R58516 VSS.n947 VSS.n946 2.2505
R58517 VSS.n958 VSS.n953 2.2505
R58518 VSS.n955 VSS.n954 2.2505
R58519 VSS.n1047 VSS.n1043 2.2505
R58520 VSS.n1003 VSS.n1002 2.2505
R58521 VSS.n1010 VSS.n1007 2.2505
R58522 VSS.n1022 VSS.n1021 2.2505
R58523 VSS.n1016 VSS.n1015 2.2505
R58524 VSS.n1707 VSS.n1706 2.2505
R58525 VSS.n1580 VSS.n1577 2.2505
R58526 VSS.n1582 VSS.n1581 2.2505
R58527 VSS.n1574 VSS.n1573 2.2505
R58528 VSS.n1849 VSS.n1848 2.2505
R58529 VSS.n1493 VSS.n1490 2.2505
R58530 VSS.n1495 VSS.n1494 2.2505
R58531 VSS.n1487 VSS.n1484 2.2505
R58532 VSS.n1481 VSS.n1480 2.2505
R58533 VSS.n1557 VSS.n1556 2.2505
R58534 VSS.n1565 VSS.n1564 2.2505
R58535 VSS.n1563 VSS.n1562 2.2505
R58536 VSS.n1568 VSS.n1567 2.2505
R58537 VSS.n1629 VSS.n1625 2.2505
R58538 VSS.n1612 VSS.n1611 2.2505
R58539 VSS.n1622 VSS.n1615 2.2505
R58540 VSS.n1618 VSS.n1617 2.2505
R58541 VSS.n9005 VSS.n9004 2.2505
R58542 VSS.n21002 VSS.n21001 2.25047
R58543 VSS.n1048 VSS.n1047 2.25047
R58544 VSS.n8919 VSS.n8916 2.25047
R58545 VSS.n16081 VSS.n16047 2.25042
R58546 VSS.n16375 VSS.n15926 2.25042
R58547 VSS.n16248 VSS.n15977 2.25042
R58548 VSS.n16246 VSS.n15985 2.25042
R58549 VSS.n16373 VSS.n15932 2.25042
R58550 VSS.n16235 VSS.n15995 2.25042
R58551 VSS.n5874 VSS.n5489 2.25042
R58552 VSS.n5872 VSS.n5499 2.25042
R58553 VSS.n16233 VSS.n16001 2.25042
R58554 VSS.n21183 VSS.n20888 2.25042
R58555 VSS.n21181 VSS.n21180 2.25042
R58556 VSS.n1300 VSS.n970 2.25042
R58557 VSS.n1060 VSS.n1010 2.25042
R58558 VSS.n1308 VSS.n1307 2.25042
R58559 VSS.n1327 VSS.n958 2.25042
R58560 VSS.n1329 VSS.n950 2.25042
R58561 VSS.n1450 VSS.n907 2.25042
R58562 VSS.n1456 VSS.n1455 2.25042
R58563 VSS.n1458 VSS.n897 2.25042
R58564 VSS.n1321 VSS.n1320 2.25042
R58565 VSS.n1314 VSS.n1313 2.25042
R58566 VSS.n1316 VSS.n966 2.25042
R58567 VSS.n8992 VSS.n8969 2.25038
R58568 VSS.n8992 VSS.n8951 2.25038
R58569 VSS.n15326 VSS.n15315 2.25037
R58570 VSS.n15667 VSS.n15210 2.25031
R58571 VSS.n15573 VSS.n15268 2.25031
R58572 VSS.n15583 VSS.n15582 2.25031
R58573 VSS.n15665 VSS.n15216 2.25031
R58574 VSS.n15338 VSS.n15305 2.25031
R58575 VSS.n15552 VSS.n15280 2.25031
R58576 VSS.n15554 VSS.n15278 2.25031
R58577 VSS.n15562 VSS.n15561 2.25031
R58578 VSS.n15564 VSS.n15274 2.25031
R58579 VSS.n1840 VSS.n1582 2.25031
R58580 VSS.n1654 VSS.n1622 2.25031
R58581 VSS.n1842 VSS.n1580 2.25031
R58582 VSS.n1925 VSS.n1487 2.25031
R58583 VSS.n1863 VSS.n1557 2.25031
R58584 VSS.n1861 VSS.n1563 2.25031
R58585 VSS.n1923 VSS.n1493 2.25031
R58586 VSS.n1857 VSS.n1568 2.25031
R58587 VSS.n1850 VSS.n1849 2.25031
R58588 VSS.n1852 VSS.n1574 2.25031
R58589 VSS.n8992 VSS.n8979 2.25029
R58590 VSS.n8992 VSS.n8991 2.25029
R58591 VSS.n4120 VSS.n4119 2.2502
R58592 VSS.n8841 VSS.n8797 2.25016
R58593 VSS.n8841 VSS.n8792 2.25016
R58594 VSS.n16131 VSS.n16025 2.25007
R58595 VSS.n8992 VSS.n8936 2.24994
R58596 VSS.n16135 VSS.n16009 2.24839
R58597 VSS.n1115 VSS.n990 2.24839
R58598 VSS.n15395 VSS.n15290 2.24789
R58599 VSS.n1711 VSS.n1607 2.24789
R58600 VSS.n16244 VSS.n16243 2.24737
R58601 VSS.n16371 VSS.n15934 2.24737
R58602 VSS.n16231 VSS.n16003 2.24737
R58603 VSS.n21175 VSS.n20892 2.24737
R58604 VSS.n15663 VSS.n15218 2.24668
R58605 VSS.n1859 VSS.n1565 2.24668
R58606 VSS.n1921 VSS.n1495 2.24668
R58607 VSS.n21931 VSS.n342 2.20947
R58608 VSS.n187 VSS.n186 2.20947
R58609 VSS.n14378 VSS.n14377 2.19825
R58610 VSS.n17174 VSS.n17173 2.19825
R58611 VSS.n359 VSS.n353 2.18432
R58612 VSS.n21692 VSS.n21686 2.18432
R58613 VSS.n420 VSS.n414 2.18432
R58614 VSS.n403 VSS.n397 2.18432
R58615 VSS.n14288 VSS.n14284 2.18432
R58616 VSS.n14288 VSS.n14286 2.18432
R58617 VSS.n385 VSS.n379 2.18432
R58618 VSS.n2507 VSS.n2455 2.18432
R58619 VSS.n2507 VSS.n2458 2.18432
R58620 VSS.n17303 VSS.n17254 2.18432
R58621 VSS.n14302 VSS.n14298 2.18432
R58622 VSS.n14302 VSS.n14301 2.18432
R58623 VSS.n4851 VSS.n4802 2.18432
R58624 VSS.n4915 VSS.n4864 2.18432
R58625 VSS.n437 VSS.n431 2.1605
R58626 VSS.n5470 VSS.n5419 2.1605
R58627 VSS.n21931 VSS.n21930 2.15918
R58628 VSS.n15691 VSS.n15690 2.0485
R58629 VSS.n201 VSS.n198 2.0485
R58630 VSS.n5894 VSS.n5887 1.85305
R58631 VSS.n5894 VSS.n5892 1.85305
R58632 VSS.n5470 VSS.n5469 1.85305
R58633 VSS.n5470 VSS.n5464 1.85305
R58634 VSS.n5470 VSS.n5429 1.85305
R58635 VSS.n5470 VSS.n5424 1.85305
R58636 VSS.n4915 VSS.n4914 1.85305
R58637 VSS.n4915 VSS.n4909 1.85305
R58638 VSS.n4915 VSS.n4874 1.85305
R58639 VSS.n4915 VSS.n4869 1.85305
R58640 VSS.n4851 VSS.n4850 1.85305
R58641 VSS.n4851 VSS.n4845 1.85305
R58642 VSS.n4851 VSS.n4812 1.85305
R58643 VSS.n4851 VSS.n4807 1.85305
R58644 VSS.n17303 VSS.n17302 1.85305
R58645 VSS.n17303 VSS.n17297 1.85305
R58646 VSS.n17303 VSS.n17264 1.85305
R58647 VSS.n17303 VSS.n17259 1.85305
R58648 VSS.n2421 VSS.n2420 1.85305
R58649 VSS.n2421 VSS.n2415 1.85305
R58650 VSS.n2421 VSS.n2390 1.85305
R58651 VSS.n2421 VSS.n2385 1.85305
R58652 VSS.n2507 VSS.n2506 1.85305
R58653 VSS.n2507 VSS.n2501 1.85305
R58654 VSS.n2507 VSS.n2468 1.85305
R58655 VSS.n2507 VSS.n2463 1.85305
R58656 VSS.n3933 VSS.n3932 1.85305
R58657 VSS.n3933 VSS.n3927 1.85305
R58658 VSS.n3933 VSS.n3899 1.85305
R58659 VSS.n3933 VSS.n3894 1.85305
R58660 VSS.n186 VSS.n179 1.85305
R58661 VSS.n186 VSS.n184 1.85305
R58662 VSS.n22123 VSS.n22121 1.83517
R58663 VSS.n21942 VSS.n21936 1.83517
R58664 VSS.n1435 VSS.n1434 1.73383
R58665 VSS.n1434 VSS.n1433 1.73383
R58666 VSS.n1411 VSS.n1410 1.73383
R58667 VSS.n1410 VSS.n1409 1.73383
R58668 VSS.n921 VSS.n920 1.73383
R58669 VSS.n920 VSS.n919 1.73383
R58670 VSS.n913 VSS.n912 1.73383
R58671 VSS.n912 VSS.n911 1.73383
R58672 VSS.n1518 VSS.n1517 1.73383
R58673 VSS.n1517 VSS.n1516 1.73383
R58674 VSS.n1513 VSS.n1512 1.73383
R58675 VSS.n1512 VSS.n1511 1.73383
R58676 VSS.n1509 VSS.n1508 1.73383
R58677 VSS.n1508 VSS.n1507 1.73383
R58678 VSS.n1501 VSS.n1500 1.73383
R58679 VSS.n1500 VSS.n1499 1.73383
R58680 VSS.n15640 VSS.n15639 1.73383
R58681 VSS.n15639 VSS.n15638 1.73383
R58682 VSS.n15235 VSS.n15234 1.73383
R58683 VSS.n15234 VSS.n15233 1.73383
R58684 VSS.n15227 VSS.n15226 1.73383
R58685 VSS.n15226 VSS.n15225 1.73383
R58686 VSS.n15221 VSS.n15220 1.73383
R58687 VSS.n15220 VSS.n15219 1.73383
R58688 VSS.n15948 VSS.n15947 1.73383
R58689 VSS.n15947 VSS.n15946 1.73383
R58690 VSS.n15940 VSS.n15939 1.73383
R58691 VSS.n15939 VSS.n15938 1.73383
R58692 VSS.n16354 VSS.n16353 1.73383
R58693 VSS.n16353 VSS.n16352 1.73383
R58694 VSS.n16349 VSS.n16348 1.73383
R58695 VSS.n16348 VSS.n16347 1.73383
R58696 VSS.n1389 VSS.n1388 1.73383
R58697 VSS.n1375 VSS.n1374 1.73383
R58698 VSS.n930 VSS.n929 1.73383
R58699 VSS.n926 VSS.n925 1.73383
R58700 VSS.n1533 VSS.n1532 1.73383
R58701 VSS.n1531 VSS.n1530 1.73383
R58702 VSS.n1527 VSS.n1526 1.73383
R58703 VSS.n1523 VSS.n1522 1.73383
R58704 VSS.n15616 VSS.n15615 1.73383
R58705 VSS.n15246 VSS.n15245 1.73383
R58706 VSS.n15242 VSS.n15241 1.73383
R58707 VSS.n15238 VSS.n15237 1.73383
R58708 VSS.n15957 VSS.n15956 1.73383
R58709 VSS.n15953 VSS.n15952 1.73383
R58710 VSS.n16308 VSS.n16307 1.73383
R58711 VSS.n16306 VSS.n16305 1.73383
R58712 VSS.n16271 VSS.n16270 1.73383
R58713 VSS.n16274 VSS.n16273 1.73383
R58714 VSS.n15963 VSS.n15962 1.73383
R58715 VSS.n15968 VSS.n15967 1.73383
R58716 VSS.n15250 VSS.n15249 1.73383
R58717 VSS.n15254 VSS.n15253 1.73383
R58718 VSS.n15259 VSS.n15258 1.73383
R58719 VSS.n15593 VSS.n15592 1.73383
R58720 VSS.n1539 VSS.n1538 1.73383
R58721 VSS.n1544 VSS.n1543 1.73383
R58722 VSS.n1547 VSS.n1546 1.73383
R58723 VSS.n1550 VSS.n1549 1.73383
R58724 VSS.n936 VSS.n935 1.73383
R58725 VSS.n941 VSS.n940 1.73383
R58726 VSS.n1339 VSS.n1338 1.73383
R58727 VSS.n1355 VSS.n1354 1.73383
R58728 VSS.n20941 VSS.n20940 1.73383
R58729 VSS.n15284 VSS.n15283 1.73383
R58730 VSS.n16022 VSS.n16021 1.73383
R58731 VSS.n16006 VSS.n16005 1.73383
R58732 VSS.n16142 VSS.n16141 1.73383
R58733 VSS.n16140 VSS.n16139 1.73383
R58734 VSS.n16015 VSS.n16014 1.73383
R58735 VSS.n5666 VSS.n5665 1.73383
R58736 VSS.n5672 VSS.n5671 1.73383
R58737 VSS.n5678 VSS.n5677 1.73383
R58738 VSS.n5682 VSS.n5681 1.73383
R58739 VSS.n5688 VSS.n5687 1.73383
R58740 VSS.n20957 VSS.n20956 1.73383
R58741 VSS.n996 VSS.n995 1.73383
R58742 VSS.n15292 VSS.n15291 1.73383
R58743 VSS.n15282 VSS.n15281 1.73383
R58744 VSS.n20951 VSS.n20950 1.73383
R58745 VSS.n20947 VSS.n20946 1.73383
R58746 VSS.n20935 VSS.n20934 1.73383
R58747 VSS.n1120 VSS.n1119 1.73383
R58748 VSS.n1122 VSS.n1121 1.73383
R58749 VSS.n987 VSS.n986 1.73383
R58750 VSS.n1604 VSS.n1603 1.73383
R58751 VSS.n1601 VSS.n1600 1.73383
R58752 VSS.n1598 VSS.n1597 1.73383
R58753 VSS.n1595 VSS.n1594 1.73383
R58754 VSS.n20982 VSS.n20981 1.73383
R58755 VSS.n20981 VSS.n20980 1.73383
R58756 VSS.n20898 VSS.n20897 1.73383
R58757 VSS.n20897 VSS.n20896 1.73383
R58758 VSS.n21100 VSS.n21099 1.73383
R58759 VSS.n21099 VSS.n21098 1.73383
R58760 VSS.n21095 VSS.n21094 1.73383
R58761 VSS.n21094 VSS.n21093 1.73383
R58762 VSS.n1147 VSS.n1146 1.73383
R58763 VSS.n1150 VSS.n1149 1.73383
R58764 VSS.n1143 VSS.n1142 1.73383
R58765 VSS.n979 VSS.n978 1.73383
R58766 VSS.n974 VSS.n973 1.73383
R58767 VSS.n1590 VSS.n1589 1.73383
R58768 VSS.n1584 VSS.n1583 1.73383
R58769 VSS.n15430 VSS.n15429 1.73383
R58770 VSS.n15420 VSS.n15419 1.73383
R58771 VSS.n5505 VSS.n5504 1.73383
R58772 VSS.n5509 VSS.n5508 1.73383
R58773 VSS.n5513 VSS.n5512 1.73383
R58774 VSS.n5517 VSS.n5516 1.73383
R58775 VSS.n5521 VSS.n5520 1.73383
R58776 VSS.n1588 VSS.n1587 1.73383
R58777 VSS.n1737 VSS.n1736 1.73383
R58778 VSS.n15434 VSS.n15433 1.73383
R58779 VSS.n15424 VSS.n15423 1.73383
R58780 VSS.n5525 VSS.n5524 1.73383
R58781 VSS.n5503 VSS.n5502 1.73383
R58782 VSS.n5711 VSS.n5710 1.73383
R58783 VSS.n5709 VSS.n5708 1.73383
R58784 VSS.n1256 VSS.n1255 1.73383
R58785 VSS.n1255 VSS.n1254 1.73383
R58786 VSS.n1265 VSS.n1264 1.73383
R58787 VSS.n1264 VSS.n1263 1.73383
R58788 VSS.n1207 VSS.n1206 1.73383
R58789 VSS.n1206 VSS.n1205 1.73383
R58790 VSS.n1198 VSS.n1197 1.73383
R58791 VSS.n1197 VSS.n1196 1.73383
R58792 VSS.n1791 VSS.n1790 1.73383
R58793 VSS.n1790 VSS.n1789 1.73383
R58794 VSS.n1804 VSS.n1803 1.73383
R58795 VSS.n1803 VSS.n1802 1.73383
R58796 VSS.n15502 VSS.n15501 1.73383
R58797 VSS.n15501 VSS.n15500 1.73383
R58798 VSS.n15487 VSS.n15486 1.73383
R58799 VSS.n15486 VSS.n15485 1.73383
R58800 VSS.n15478 VSS.n15477 1.73383
R58801 VSS.n15477 VSS.n15476 1.73383
R58802 VSS.n5799 VSS.n5798 1.73383
R58803 VSS.n5798 VSS.n5797 1.73383
R58804 VSS.n5803 VSS.n5802 1.73383
R58805 VSS.n5802 VSS.n5801 1.73383
R58806 VSS.n5810 VSS.n5809 1.73383
R58807 VSS.n5809 VSS.n5808 1.73383
R58808 VSS.n5817 VSS.n5816 1.73383
R58809 VSS.n5816 VSS.n5815 1.73383
R58810 VSS.n5826 VSS.n5825 1.73383
R58811 VSS.n5825 VSS.n5824 1.73383
R58812 VSS.n5833 VSS.n5832 1.73383
R58813 VSS.n5832 VSS.n5831 1.73383
R58814 VSS.n5783 VSS.n5782 1.73383
R58815 VSS.n5782 VSS.n5781 1.73383
R58816 VSS.n5774 VSS.n5773 1.73383
R58817 VSS.n5773 VSS.n5772 1.73383
R58818 VSS.n1798 VSS.n1797 1.73383
R58819 VSS.n1797 VSS.n1796 1.73383
R58820 VSS.n1786 VSS.n1785 1.73383
R58821 VSS.n1785 VSS.n1784 1.73383
R58822 VSS.n15516 VSS.n15515 1.73383
R58823 VSS.n15515 VSS.n15514 1.73383
R58824 VSS.n1235 VSS.n1234 1.73383
R58825 VSS.n1225 VSS.n1224 1.73383
R58826 VSS.n1232 VSS.n1231 1.73383
R58827 VSS.n1241 VSS.n1240 1.73383
R58828 VSS.n1249 VSS.n1248 1.73383
R58829 VSS.n1248 VSS.n1247 1.73383
R58830 VSS.n15496 VSS.n15495 1.73383
R58831 VSS.n15495 VSS.n15494 1.73383
R58832 VSS.n202 VSS.n201 1.73383
R58833 VSS.n13537 VSS.n13536 1.7277
R58834 VSS.n13534 VSS.n13533 1.7277
R58835 VSS.n13528 VSS.n13527 1.7277
R58836 VSS.n13518 VSS.n13517 1.7277
R58837 VSS.n13434 VSS.n13433 1.7277
R58838 VSS.n13424 VSS.n13423 1.7277
R58839 VSS.n13276 VSS.n13275 1.7277
R58840 VSS.n13271 VSS.n13270 1.7277
R58841 VSS.n11765 VSS.n11764 1.7277
R58842 VSS.n11762 VSS.n11761 1.7277
R58843 VSS.n11759 VSS.n11758 1.7277
R58844 VSS.n14336 VSS.n14334 1.7277
R58845 VSS.n17179 VSS.n11749 1.7277
R58846 VSS.n14345 VSS.n14340 1.7277
R58847 VSS.n14351 VSS.n14346 1.7277
R58848 VSS.n14361 VSS.n14355 1.7277
R58849 VSS.n14365 VSS.n14362 1.7277
R58850 VSS.n14367 VSS.n14366 1.7277
R58851 VSS.n14373 VSS.n14371 1.7277
R58852 VSS.n14376 VSS.n14374 1.7277
R58853 VSS.n17178 VSS.n14330 1.69393
R58854 VSS.n15696 VSS.n15676 1.68445
R58855 VSS.n15696 VSS.n15694 1.68445
R58856 VSS.n17293 VSS.n17265 1.68445
R58857 VSS.n17178 VSS.n11753 1.68445
R58858 VSS.n4841 VSS.n4813 1.68445
R58859 VSS.n4905 VSS.n4875 1.68445
R58860 VSS.n5460 VSS.n5430 1.68445
R58861 VSS.n2497 VSS.n2496 1.68445
R58862 VSS.n17293 VSS.n17283 1.61232
R58863 VSS.n17293 VSS.n17284 1.61232
R58864 VSS.n17293 VSS.n17285 1.61232
R58865 VSS.n17293 VSS.n17287 1.61232
R58866 VSS.n17293 VSS.n17288 1.61232
R58867 VSS.n17293 VSS.n17289 1.61232
R58868 VSS.n17293 VSS.n17291 1.61232
R58869 VSS.n17293 VSS.n17292 1.61232
R58870 VSS.n17293 VSS.n17280 1.61232
R58871 VSS.n17293 VSS.n17279 1.61232
R58872 VSS.n17293 VSS.n17277 1.61232
R58873 VSS.n17293 VSS.n17276 1.61232
R58874 VSS.n17293 VSS.n17275 1.61232
R58875 VSS.n17293 VSS.n17273 1.61232
R58876 VSS.n17293 VSS.n17272 1.61232
R58877 VSS.n17293 VSS.n17271 1.61232
R58878 VSS.n17293 VSS.n17269 1.61232
R58879 VSS.n17293 VSS.n17268 1.61232
R58880 VSS.n17293 VSS.n17267 1.61232
R58881 VSS.n17178 VSS.n14336 1.61232
R58882 VSS.n17179 VSS.n17178 1.61232
R58883 VSS.n17178 VSS.n14345 1.61232
R58884 VSS.n17178 VSS.n14351 1.61232
R58885 VSS.n17178 VSS.n14361 1.61232
R58886 VSS.n17178 VSS.n14365 1.61232
R58887 VSS.n17178 VSS.n14367 1.61232
R58888 VSS.n17178 VSS.n14373 1.61232
R58889 VSS.n17178 VSS.n14376 1.61232
R58890 VSS.n17178 VSS.n13537 1.61232
R58891 VSS.n17178 VSS.n13534 1.61232
R58892 VSS.n17178 VSS.n13528 1.61232
R58893 VSS.n17178 VSS.n13518 1.61232
R58894 VSS.n17178 VSS.n13434 1.61232
R58895 VSS.n17178 VSS.n13424 1.61232
R58896 VSS.n17178 VSS.n13276 1.61232
R58897 VSS.n17178 VSS.n13271 1.61232
R58898 VSS.n17178 VSS.n11765 1.61232
R58899 VSS.n17178 VSS.n11762 1.61232
R58900 VSS.n17178 VSS.n11759 1.61232
R58901 VSS.n4841 VSS.n4831 1.61232
R58902 VSS.n4841 VSS.n4832 1.61232
R58903 VSS.n4841 VSS.n4833 1.61232
R58904 VSS.n4841 VSS.n4835 1.61232
R58905 VSS.n4841 VSS.n4836 1.61232
R58906 VSS.n4841 VSS.n4837 1.61232
R58907 VSS.n4841 VSS.n4839 1.61232
R58908 VSS.n4841 VSS.n4840 1.61232
R58909 VSS.n4841 VSS.n4828 1.61232
R58910 VSS.n4841 VSS.n4827 1.61232
R58911 VSS.n4841 VSS.n4825 1.61232
R58912 VSS.n4841 VSS.n4824 1.61232
R58913 VSS.n4841 VSS.n4823 1.61232
R58914 VSS.n4841 VSS.n4821 1.61232
R58915 VSS.n4841 VSS.n4820 1.61232
R58916 VSS.n4841 VSS.n4819 1.61232
R58917 VSS.n4841 VSS.n4817 1.61232
R58918 VSS.n4841 VSS.n4816 1.61232
R58919 VSS.n4841 VSS.n4815 1.61232
R58920 VSS.n4905 VSS.n4893 1.61232
R58921 VSS.n4905 VSS.n4894 1.61232
R58922 VSS.n4905 VSS.n4895 1.61232
R58923 VSS.n4905 VSS.n4897 1.61232
R58924 VSS.n4905 VSS.n4898 1.61232
R58925 VSS.n4905 VSS.n4899 1.61232
R58926 VSS.n4905 VSS.n4901 1.61232
R58927 VSS.n4905 VSS.n4902 1.61232
R58928 VSS.n4905 VSS.n4890 1.61232
R58929 VSS.n4905 VSS.n4889 1.61232
R58930 VSS.n4905 VSS.n4887 1.61232
R58931 VSS.n4905 VSS.n4886 1.61232
R58932 VSS.n4905 VSS.n4885 1.61232
R58933 VSS.n4905 VSS.n4883 1.61232
R58934 VSS.n4905 VSS.n4882 1.61232
R58935 VSS.n4905 VSS.n4881 1.61232
R58936 VSS.n4905 VSS.n4879 1.61232
R58937 VSS.n4905 VSS.n4878 1.61232
R58938 VSS.n4905 VSS.n4877 1.61232
R58939 VSS.n5460 VSS.n5448 1.61232
R58940 VSS.n5460 VSS.n5449 1.61232
R58941 VSS.n5460 VSS.n5450 1.61232
R58942 VSS.n5460 VSS.n5452 1.61232
R58943 VSS.n5460 VSS.n5453 1.61232
R58944 VSS.n5460 VSS.n5454 1.61232
R58945 VSS.n5460 VSS.n5456 1.61232
R58946 VSS.n5460 VSS.n5457 1.61232
R58947 VSS.n5460 VSS.n5445 1.61232
R58948 VSS.n5460 VSS.n5444 1.61232
R58949 VSS.n5460 VSS.n5442 1.61232
R58950 VSS.n5460 VSS.n5441 1.61232
R58951 VSS.n5460 VSS.n5440 1.61232
R58952 VSS.n5460 VSS.n5438 1.61232
R58953 VSS.n5460 VSS.n5437 1.61232
R58954 VSS.n5460 VSS.n5436 1.61232
R58955 VSS.n5460 VSS.n5434 1.61232
R58956 VSS.n5460 VSS.n5433 1.61232
R58957 VSS.n5460 VSS.n5432 1.61232
R58958 VSS.n2411 VSS.n2397 1.61232
R58959 VSS.n2411 VSS.n2396 1.61232
R58960 VSS.n2411 VSS.n2395 1.61232
R58961 VSS.n2411 VSS.n2394 1.61232
R58962 VSS.n2411 VSS.n2393 1.61232
R58963 VSS.n2411 VSS.n2392 1.61232
R58964 VSS.n2497 VSS.n2481 1.61232
R58965 VSS.n2497 VSS.n2482 1.61232
R58966 VSS.n2497 VSS.n2483 1.61232
R58967 VSS.n2497 VSS.n2485 1.61232
R58968 VSS.n2497 VSS.n2486 1.61232
R58969 VSS.n2497 VSS.n2487 1.61232
R58970 VSS.n2497 VSS.n2489 1.61232
R58971 VSS.n2497 VSS.n2490 1.61232
R58972 VSS.n2497 VSS.n2491 1.61232
R58973 VSS.n2497 VSS.n2493 1.61232
R58974 VSS.n2497 VSS.n2494 1.61232
R58975 VSS.n2497 VSS.n2480 1.61232
R58976 VSS.n3923 VSS.n3914 1.61232
R58977 VSS.n3923 VSS.n3915 1.61232
R58978 VSS.n3923 VSS.n3911 1.61232
R58979 VSS.n3923 VSS.n3909 1.61232
R58980 VSS.n3923 VSS.n3907 1.61232
R58981 VSS.n3923 VSS.n3917 1.61232
R58982 VSS.n3923 VSS.n3918 1.61232
R58983 VSS.n3923 VSS.n3905 1.61232
R58984 VSS.n3923 VSS.n3919 1.61232
R58985 VSS.n3923 VSS.n3920 1.61232
R58986 VSS.n3923 VSS.n3903 1.61232
R58987 VSS.n3923 VSS.n3921 1.61232
R58988 VSS.n3923 VSS.n3901 1.61232
R58989 VSS.n3923 VSS.n3922 1.61232
R58990 VSS.n3923 VSS.n3900 1.61232
R58991 VSS.n2497 VSS.n2479 1.61232
R58992 VSS.n2497 VSS.n2477 1.61232
R58993 VSS.n2497 VSS.n2476 1.61232
R58994 VSS.n2497 VSS.n2475 1.61232
R58995 VSS.n2497 VSS.n2473 1.61232
R58996 VSS.n2497 VSS.n2472 1.61232
R58997 VSS.n2497 VSS.n2471 1.61232
R58998 VSS.n2411 VSS.n2391 1.61232
R58999 VSS.n2411 VSS.n2405 1.61232
R59000 VSS.n2411 VSS.n2406 1.61232
R59001 VSS.n2411 VSS.n2407 1.61232
R59002 VSS.n2411 VSS.n2409 1.61232
R59003 VSS.n2411 VSS.n2410 1.61232
R59004 VSS.n11753 VSS.n11752 1.57222
R59005 VSS.n17227 VSS.n17226 1.5539
R59006 VSS.n14330 VSS.n14329 1.5518
R59007 VSS.n17218 VSS.n17217 1.5296
R59008 VSS.n13659 VSS.n13622 1.50371
R59009 VSS.n16966 VSS.n16940 1.5005
R59010 VSS.n17009 VSS.n17008 1.5005
R59011 VSS.n17160 VSS.n17159 1.5005
R59012 VSS.n14561 VSS.n14560 1.5005
R59013 VSS.n14547 VSS.n14546 1.5005
R59014 VSS.n14533 VSS.n14532 1.5005
R59015 VSS.n14519 VSS.n14518 1.5005
R59016 VSS.n14505 VSS.n14504 1.5005
R59017 VSS.n14491 VSS.n14490 1.5005
R59018 VSS.n14477 VSS.n14476 1.5005
R59019 VSS.n14470 VSS.n14469 1.5005
R59020 VSS.n14484 VSS.n14483 1.5005
R59021 VSS.n14498 VSS.n14497 1.5005
R59022 VSS.n14512 VSS.n14511 1.5005
R59023 VSS.n14526 VSS.n14525 1.5005
R59024 VSS.n14540 VSS.n14539 1.5005
R59025 VSS.n14554 VSS.n14553 1.5005
R59026 VSS.n14587 VSS.n14586 1.5005
R59027 VSS.n14712 VSS.n14711 1.5005
R59028 VSS.n14682 VSS.n14681 1.5005
R59029 VSS.n14689 VSS.n14688 1.5005
R59030 VSS.n14697 VSS.n14696 1.5005
R59031 VSS.n14705 VSS.n14704 1.5005
R59032 VSS.n14719 VSS.n14718 1.5005
R59033 VSS.n14727 VSS.n14726 1.5005
R59034 VSS.n14808 VSS.n14807 1.5005
R59035 VSS.n17116 VSS.n17115 1.5005
R59036 VSS.n17065 VSS.n17064 1.5005
R59037 VSS.n15647 VSS.n15642 1.5005
R59038 VSS.n15642 VSS.n15641 1.5005
R59039 VSS.n15232 VSS.n15231 1.5005
R59040 VSS.n15231 VSS.n15230 1.5005
R59041 VSS.n15236 VSS.n15229 1.5005
R59042 VSS.n15229 VSS.n15228 1.5005
R59043 VSS.n15224 VSS.n15223 1.5005
R59044 VSS.n15223 VSS.n15222 1.5005
R59045 VSS.n15620 VSS.n15619 1.5005
R59046 VSS.n15244 VSS.n15243 1.5005
R59047 VSS.n15248 VSS.n15247 1.5005
R59048 VSS.n15240 VSS.n15239 1.5005
R59049 VSS.n15252 VSS.n15251 1.5005
R59050 VSS.n15260 VSS.n15255 1.5005
R59051 VSS.n15257 VSS.n15256 1.5005
R59052 VSS.n15597 VSS.n15594 1.5005
R59053 VSS.n16577 VSS.n16576 1.5005
R59054 VSS.n16629 VSS.n16628 1.5005
R59055 VSS.n16708 VSS.n16707 1.5005
R59056 VSS.n16722 VSS.n16721 1.5005
R59057 VSS.n16736 VSS.n16735 1.5005
R59058 VSS.n16750 VSS.n16749 1.5005
R59059 VSS.n16764 VSS.n16763 1.5005
R59060 VSS.n16778 VSS.n16777 1.5005
R59061 VSS.n16792 VSS.n16791 1.5005
R59062 VSS.n16806 VSS.n16805 1.5005
R59063 VSS.n16820 VSS.n16819 1.5005
R59064 VSS.n16834 VSS.n16833 1.5005
R59065 VSS.n16848 VSS.n16847 1.5005
R59066 VSS.n16868 VSS.n16867 1.5005
R59067 VSS.n16855 VSS.n16854 1.5005
R59068 VSS.n16841 VSS.n16840 1.5005
R59069 VSS.n16827 VSS.n16826 1.5005
R59070 VSS.n16813 VSS.n16812 1.5005
R59071 VSS.n16799 VSS.n16798 1.5005
R59072 VSS.n16785 VSS.n16784 1.5005
R59073 VSS.n16771 VSS.n16770 1.5005
R59074 VSS.n16758 VSS.n16751 1.5005
R59075 VSS.n16743 VSS.n16742 1.5005
R59076 VSS.n16729 VSS.n16728 1.5005
R59077 VSS.n16715 VSS.n16714 1.5005
R59078 VSS.n16522 VSS.n16521 1.5005
R59079 VSS.n16457 VSS.n16456 1.5005
R59080 VSS.n16464 VSS.n16463 1.5005
R59081 VSS.n16471 VSS.n16470 1.5005
R59082 VSS.n16478 VSS.n16477 1.5005
R59083 VSS.n16485 VSS.n16484 1.5005
R59084 VSS.n16492 VSS.n16491 1.5005
R59085 VSS.n16499 VSS.n16498 1.5005
R59086 VSS.n16505 VSS.n16500 1.5005
R59087 VSS.n16666 VSS.n16665 1.5005
R59088 VSS.n16679 VSS.n16678 1.5005
R59089 VSS.n18523 VSS.n18522 1.5005
R59090 VSS.n18537 VSS.n18536 1.5005
R59091 VSS.n18551 VSS.n18550 1.5005
R59092 VSS.n18565 VSS.n18564 1.5005
R59093 VSS.n18579 VSS.n18578 1.5005
R59094 VSS.n18593 VSS.n18592 1.5005
R59095 VSS.n18607 VSS.n18606 1.5005
R59096 VSS.n18621 VSS.n18620 1.5005
R59097 VSS.n18635 VSS.n18634 1.5005
R59098 VSS.n18649 VSS.n18648 1.5005
R59099 VSS.n18666 VSS.n18665 1.5005
R59100 VSS.n18656 VSS.n18655 1.5005
R59101 VSS.n18642 VSS.n18641 1.5005
R59102 VSS.n18628 VSS.n18627 1.5005
R59103 VSS.n18614 VSS.n18613 1.5005
R59104 VSS.n18600 VSS.n18599 1.5005
R59105 VSS.n18586 VSS.n18585 1.5005
R59106 VSS.n18572 VSS.n18571 1.5005
R59107 VSS.n18560 VSS.n18552 1.5005
R59108 VSS.n18544 VSS.n18543 1.5005
R59109 VSS.n18530 VSS.n18529 1.5005
R59110 VSS.n18516 VSS.n18515 1.5005
R59111 VSS.n18509 VSS.n18508 1.5005
R59112 VSS.n18502 VSS.n18501 1.5005
R59113 VSS.n18495 VSS.n18494 1.5005
R59114 VSS.n18488 VSS.n18487 1.5005
R59115 VSS.n18303 VSS.n18302 1.5005
R59116 VSS.n18310 VSS.n18309 1.5005
R59117 VSS.n18317 VSS.n18316 1.5005
R59118 VSS.n18324 VSS.n18323 1.5005
R59119 VSS.n18331 VSS.n18330 1.5005
R59120 VSS.n18338 VSS.n18337 1.5005
R59121 VSS.n18345 VSS.n18344 1.5005
R59122 VSS.n18352 VSS.n18351 1.5005
R59123 VSS.n18359 VSS.n18358 1.5005
R59124 VSS.n18390 VSS.n18389 1.5005
R59125 VSS.n18420 VSS.n18419 1.5005
R59126 VSS.n18436 VSS.n18435 1.5005
R59127 VSS.n15945 VSS.n15944 1.5005
R59128 VSS.n15944 VSS.n15943 1.5005
R59129 VSS.n15949 VSS.n15942 1.5005
R59130 VSS.n15942 VSS.n15941 1.5005
R59131 VSS.n15937 VSS.n15936 1.5005
R59132 VSS.n15936 VSS.n15935 1.5005
R59133 VSS.n16355 VSS.n16351 1.5005
R59134 VSS.n16351 VSS.n16350 1.5005
R59135 VSS.n15955 VSS.n15954 1.5005
R59136 VSS.n15959 VSS.n15958 1.5005
R59137 VSS.n15951 VSS.n15950 1.5005
R59138 VSS.n16310 VSS.n16309 1.5005
R59139 VSS.n16304 VSS.n16303 1.5005
R59140 VSS.n16269 VSS.n16268 1.5005
R59141 VSS.n16275 VSS.n16272 1.5005
R59142 VSS.n15961 VSS.n15960 1.5005
R59143 VSS.n15969 VSS.n15964 1.5005
R59144 VSS.n15966 VSS.n15965 1.5005
R59145 VSS.n16346 VSS.n16345 1.5005
R59146 VSS.n16345 VSS.n16344 1.5005
R59147 VSS.n15297 VSS.n15296 1.5005
R59148 VSS.n15390 VSS.n15389 1.5005
R59149 VSS.n15290 VSS.n15289 1.5005
R59150 VSS.n16025 VSS.n16024 1.5005
R59151 VSS.n16009 VSS.n16008 1.5005
R59152 VSS.n16144 VSS.n16143 1.5005
R59153 VSS.n16019 VSS.n16018 1.5005
R59154 VSS.n16012 VSS.n16011 1.5005
R59155 VSS.n5669 VSS.n5668 1.5005
R59156 VSS.n5675 VSS.n5674 1.5005
R59157 VSS.n5680 VSS.n5679 1.5005
R59158 VSS.n5685 VSS.n5684 1.5005
R59159 VSS.n5691 VSS.n5690 1.5005
R59160 VSS.n15286 VSS.n15285 1.5005
R59161 VSS.n15438 VSS.n15437 1.5005
R59162 VSS.n15432 VSS.n15431 1.5005
R59163 VSS.n15422 VSS.n15421 1.5005
R59164 VSS.n15426 VSS.n15425 1.5005
R59165 VSS.n15418 VSS.n15417 1.5005
R59166 VSS.n5507 VSS.n5506 1.5005
R59167 VSS.n5511 VSS.n5510 1.5005
R59168 VSS.n5515 VSS.n5514 1.5005
R59169 VSS.n5519 VSS.n5518 1.5005
R59170 VSS.n5523 VSS.n5522 1.5005
R59171 VSS.n5527 VSS.n5526 1.5005
R59172 VSS.n5501 VSS.n5500 1.5005
R59173 VSS.n5713 VSS.n5712 1.5005
R59174 VSS.n5707 VSS.n5706 1.5005
R59175 VSS.n15511 VSS.n15504 1.5005
R59176 VSS.n15504 VSS.n15503 1.5005
R59177 VSS.n15519 VSS.n15518 1.5005
R59178 VSS.n15518 VSS.n15517 1.5005
R59179 VSS.n15482 VSS.n15481 1.5005
R59180 VSS.n15481 VSS.n15480 1.5005
R59181 VSS.n5795 VSS.n5793 1.5005
R59182 VSS.n5793 VSS.n5792 1.5005
R59183 VSS.n5800 VSS.n5791 1.5005
R59184 VSS.n5791 VSS.n5790 1.5005
R59185 VSS.n5805 VSS.n5789 1.5005
R59186 VSS.n5789 VSS.n5788 1.5005
R59187 VSS.n5812 VSS.n5787 1.5005
R59188 VSS.n5787 VSS.n5786 1.5005
R59189 VSS.n5822 VSS.n5821 1.5005
R59190 VSS.n5821 VSS.n5820 1.5005
R59191 VSS.n5829 VSS.n5785 1.5005
R59192 VSS.n5785 VSS.n5784 1.5005
R59193 VSS.n5779 VSS.n5778 1.5005
R59194 VSS.n5778 VSS.n5777 1.5005
R59195 VSS.n5770 VSS.n5769 1.5005
R59196 VSS.n5769 VSS.n5768 1.5005
R59197 VSS.n5836 VSS.n5835 1.5005
R59198 VSS.n5835 VSS.n5834 1.5005
R59199 VSS.n15492 VSS.n15491 1.5005
R59200 VSS.n15491 VSS.n15490 1.5005
R59201 VSS.n15499 VSS.n15498 1.5005
R59202 VSS.n15498 VSS.n15497 1.5005
R59203 VSS.n1222 VSS.n1221 1.5005
R59204 VSS.n1228 VSS.n1227 1.5005
R59205 VSS.n1233 VSS.n1210 1.5005
R59206 VSS.n1238 VSS.n1237 1.5005
R59207 VSS.n1245 VSS.n1244 1.5005
R59208 VSS.n20983 VSS.n20900 1.5005
R59209 VSS.n20900 VSS.n20899 1.5005
R59210 VSS.n20895 VSS.n20894 1.5005
R59211 VSS.n20894 VSS.n20893 1.5005
R59212 VSS.n21101 VSS.n21097 1.5005
R59213 VSS.n21097 VSS.n21096 1.5005
R59214 VSS.n21092 VSS.n21091 1.5005
R59215 VSS.n21091 VSS.n21090 1.5005
R59216 VSS.n20979 VSS.n20978 1.5005
R59217 VSS.n20978 VSS.n20977 1.5005
R59218 VSS.n20954 VSS.n20953 1.5005
R59219 VSS.n20949 VSS.n20948 1.5005
R59220 VSS.n20944 VSS.n20943 1.5005
R59221 VSS.n20938 VSS.n20937 1.5005
R59222 VSS.n20960 VSS.n20959 1.5005
R59223 VSS.n1252 VSS.n1209 1.5005
R59224 VSS.n1209 VSS.n1208 1.5005
R59225 VSS.n1261 VSS.n1260 1.5005
R59226 VSS.n1260 VSS.n1259 1.5005
R59227 VSS.n1268 VSS.n1267 1.5005
R59228 VSS.n1267 VSS.n1266 1.5005
R59229 VSS.n1203 VSS.n1202 1.5005
R59230 VSS.n1202 VSS.n1201 1.5005
R59231 VSS.n1194 VSS.n1193 1.5005
R59232 VSS.n1193 VSS.n1192 1.5005
R59233 VSS.n1432 VSS.n1415 1.5005
R59234 VSS.n1415 VSS.n1414 1.5005
R59235 VSS.n1436 VSS.n1413 1.5005
R59236 VSS.n1413 VSS.n1412 1.5005
R59237 VSS.n918 VSS.n917 1.5005
R59238 VSS.n917 VSS.n916 1.5005
R59239 VSS.n922 VSS.n915 1.5005
R59240 VSS.n915 VSS.n914 1.5005
R59241 VSS.n910 VSS.n909 1.5005
R59242 VSS.n909 VSS.n908 1.5005
R59243 VSS.n1387 VSS.n1386 1.5005
R59244 VSS.n1391 VSS.n1390 1.5005
R59245 VSS.n928 VSS.n927 1.5005
R59246 VSS.n932 VSS.n931 1.5005
R59247 VSS.n924 VSS.n923 1.5005
R59248 VSS.n934 VSS.n933 1.5005
R59249 VSS.n942 VSS.n937 1.5005
R59250 VSS.n939 VSS.n938 1.5005
R59251 VSS.n1356 VSS.n1340 1.5005
R59252 VSS.n1353 VSS.n1352 1.5005
R59253 VSS.n1148 VSS.n1145 1.5005
R59254 VSS.n1151 VSS.n1144 1.5005
R59255 VSS.n977 VSS.n976 1.5005
R59256 VSS.n980 VSS.n975 1.5005
R59257 VSS.n972 VSS.n971 1.5005
R59258 VSS.n1000 VSS.n999 1.5005
R59259 VSS.n1124 VSS.n1123 1.5005
R59260 VSS.n990 VSS.n989 1.5005
R59261 VSS.n984 VSS.n983 1.5005
R59262 VSS.n993 VSS.n992 1.5005
R59263 VSS.n1794 VSS.n1788 1.5005
R59264 VSS.n1788 VSS.n1787 1.5005
R59265 VSS.n1801 VSS.n1800 1.5005
R59266 VSS.n1800 VSS.n1799 1.5005
R59267 VSS.n1807 VSS.n1806 1.5005
R59268 VSS.n1806 VSS.n1805 1.5005
R59269 VSS.n19823 VSS.n19822 1.5005
R59270 VSS.n19781 VSS.n19780 1.5005
R59271 VSS.n19790 VSS.n19789 1.5005
R59272 VSS.n19798 VSS.n19797 1.5005
R59273 VSS.n19808 VSS.n19807 1.5005
R59274 VSS.n19816 VSS.n19815 1.5005
R59275 VSS.n19830 VSS.n19829 1.5005
R59276 VSS.n1519 VSS.n1515 1.5005
R59277 VSS.n1515 VSS.n1514 1.5005
R59278 VSS.n1506 VSS.n1505 1.5005
R59279 VSS.n1505 VSS.n1504 1.5005
R59280 VSS.n1510 VSS.n1503 1.5005
R59281 VSS.n1503 VSS.n1502 1.5005
R59282 VSS.n1498 VSS.n1497 1.5005
R59283 VSS.n1497 VSS.n1496 1.5005
R59284 VSS.n1535 VSS.n1534 1.5005
R59285 VSS.n1525 VSS.n1524 1.5005
R59286 VSS.n1529 VSS.n1528 1.5005
R59287 VSS.n1521 VSS.n1520 1.5005
R59288 VSS.n1537 VSS.n1536 1.5005
R59289 VSS.n1545 VSS.n1540 1.5005
R59290 VSS.n1542 VSS.n1541 1.5005
R59291 VSS.n1551 VSS.n1548 1.5005
R59292 VSS.n19279 VSS.n19278 1.5005
R59293 VSS.n19286 VSS.n19285 1.5005
R59294 VSS.n19293 VSS.n19292 1.5005
R59295 VSS.n19300 VSS.n19299 1.5005
R59296 VSS.n19307 VSS.n19306 1.5005
R59297 VSS.n19314 VSS.n19313 1.5005
R59298 VSS.n19321 VSS.n19320 1.5005
R59299 VSS.n19328 VSS.n19327 1.5005
R59300 VSS.n19335 VSS.n19334 1.5005
R59301 VSS.n19342 VSS.n19341 1.5005
R59302 VSS.n19438 VSS.n19437 1.5005
R59303 VSS.n1592 VSS.n1591 1.5005
R59304 VSS.n1586 VSS.n1585 1.5005
R59305 VSS.n1735 VSS.n1734 1.5005
R59306 VSS.n1738 VSS.n1733 1.5005
R59307 VSS.n1781 VSS.n1780 1.5005
R59308 VSS.n1780 VSS.n1779 1.5005
R59309 VSS.n1607 VSS.n1606 1.5005
R59310 VSS.n1706 VSS.n1705 1.5005
R59311 VSS.n1610 VSS.n1609 1.5005
R59312 VSS.n1599 VSS.n1596 1.5005
R59313 VSS.n15855 VSS.n15854 1.5005
R59314 VSS.n15844 VSS.n15843 1.5005
R59315 VSS.n15830 VSS.n15829 1.5005
R59316 VSS.n15813 VSS.n15810 1.5005
R59317 VSS.n15802 VSS.n15801 1.5005
R59318 VSS.n15788 VSS.n15787 1.5005
R59319 VSS.n15774 VSS.n15773 1.5005
R59320 VSS.n15760 VSS.n15759 1.5005
R59321 VSS.n15746 VSS.n15745 1.5005
R59322 VSS.n15732 VSS.n15731 1.5005
R59323 VSS.n15718 VSS.n15717 1.5005
R59324 VSS.n15725 VSS.n15724 1.5005
R59325 VSS.n15739 VSS.n15738 1.5005
R59326 VSS.n15753 VSS.n15752 1.5005
R59327 VSS.n15767 VSS.n15766 1.5005
R59328 VSS.n15781 VSS.n15780 1.5005
R59329 VSS.n15795 VSS.n15794 1.5005
R59330 VSS.n15809 VSS.n15808 1.5005
R59331 VSS.n15823 VSS.n15822 1.5005
R59332 VSS.n15837 VSS.n15836 1.5005
R59333 VSS.n15851 VSS.n15850 1.5005
R59334 VSS.n13656 VSS.n13655 1.5005
R59335 VSS.n22229 VSS.n22228 1.5005
R59336 VSS.n13643 VSS.n13642 1.5005
R59337 VSS.n14273 VSS.n14272 1.5005
R59338 VSS.n14276 VSS.n14275 1.5005
R59339 VSS.n14251 VSS.n14250 1.5005
R59340 VSS.n13603 VSS.n13602 1.5005
R59341 VSS.n13610 VSS.n13609 1.5005
R59342 VSS.n21943 VSS.n21942 1.5005
R59343 VSS.n21985 VSS.n21984 1.5005
R59344 VSS.n22174 VSS.n22173 1.5005
R59345 VSS.n22161 VSS.n22160 1.5005
R59346 VSS.n22252 VSS.n22251 1.5005
R59347 VSS.n22237 VSS.n22236 1.5005
R59348 VSS.n21947 VSS.n21946 1.5005
R59349 VSS.n21960 VSS.n21959 1.5005
R59350 VSS.n21977 VSS.n21976 1.5005
R59351 VSS.n21967 VSS.n21966 1.5005
R59352 VSS.n33 VSS.n24 1.5005
R59353 VSS.n4187 VSS.n4186 1.50017
R59354 VSS.n16358 VSS.n15949 1.50017
R59355 VSS.n16313 VSS.n15959 1.50017
R59356 VSS.n16278 VSS.n15969 1.50017
R59357 VSS.n18986 VSS.n18985 1.50017
R59358 VSS.n5716 VSS.n5527 1.50017
R59359 VSS.n21742 VSS.n21741 1.50017
R59360 VSS.n21104 VSS.n20983 1.50017
R59361 VSS.n19027 VSS.n19026 1.50017
R59362 VSS.n4165 VSS.n4163 1.50017
R59363 VSS.n18990 VSS.n18988 1.50013
R59364 VSS.n5714 VSS.n5713 1.50013
R59365 VSS.n21734 VSS.n21733 1.50013
R59366 VSS.n21102 VSS.n21101 1.50013
R59367 VSS.n17885 VSS.n17884 1.50013
R59368 VSS.n21707 VSS.n21682 1.50013
R59369 VSS.n21455 VSS.n375 1.50013
R59370 VSS.n18111 VSS.n18109 1.50009
R59371 VSS.n17963 VSS.n17962 1.50009
R59372 VSS.n1154 VSS.n980 1.50006
R59373 VSS.n1359 VSS.n942 1.50006
R59374 VSS.n1394 VSS.n932 1.50006
R59375 VSS.n1439 VSS.n922 1.50006
R59376 VSS.n18944 VSS.n18850 1.50006
R59377 VSS.n4075 VSS.n4073 1.50006
R59378 VSS.n21875 VSS.n21873 1.50006
R59379 VSS.n19160 VSS.n19158 1.50006
R59380 VSS.n4198 VSS.n4197 1.50002
R59381 VSS.n16356 VSS.n16355 1.50002
R59382 VSS.n16311 VSS.n16310 1.50002
R59383 VSS.n16276 VSS.n16275 1.50002
R59384 VSS.n5837 VSS.n5836 1.50002
R59385 VSS.n1152 VSS.n1151 1.50002
R59386 VSS.n1269 VSS.n1268 1.50002
R59387 VSS.n1357 VSS.n1356 1.50002
R59388 VSS.n1392 VSS.n1391 1.50002
R59389 VSS.n1437 VSS.n1436 1.50002
R59390 VSS.n1741 VSS.n1592 1.49999
R59391 VSS.n15439 VSS.n15438 1.49999
R59392 VSS.n17479 VSS.n17431 1.49998
R59393 VSS.n13350 VSS.n13314 1.49998
R59394 VSS.n13493 VSS.n13471 1.49998
R59395 VSS.n15427 VSS.n15426 1.49994
R59396 VSS.n18138 VSS.n18137 1.49989
R59397 VSS.n19709 VSS.n2149 1.49989
R59398 VSS.n15600 VSS.n15260 1.49987
R59399 VSS.n15623 VSS.n15248 1.49987
R59400 VSS.n15650 VSS.n15236 1.49987
R59401 VSS.n1908 VSS.n1510 1.49987
R59402 VSS.n1891 VSS.n1529 1.49987
R59403 VSS.n1874 VSS.n1545 1.49987
R59404 VSS.n19512 VSS.n19172 1.49987
R59405 VSS.n18842 VSS.n18840 1.49987
R59406 VSS.n15598 VSS.n15597 1.49983
R59407 VSS.n15621 VSS.n15620 1.49983
R59408 VSS.n15648 VSS.n15647 1.49983
R59409 VSS.n15520 VSS.n15519 1.49983
R59410 VSS.n1808 VSS.n1807 1.49983
R59411 VSS.n1906 VSS.n1519 1.49983
R59412 VSS.n1889 VSS.n1535 1.49983
R59413 VSS.n1872 VSS.n1551 1.49983
R59414 VSS.n1739 VSS.n1738 1.49983
R59415 VSS.n19717 VSS.n2146 1.49978
R59416 VSS.n184 VSS.n183 1.49689
R59417 VSS.n179 VSS.n178 1.49689
R59418 VSS.n3894 VSS.n3893 1.49689
R59419 VSS.n3899 VSS.n3898 1.49689
R59420 VSS.n3927 VSS.n3926 1.49689
R59421 VSS.n3932 VSS.n3931 1.49689
R59422 VSS.n2463 VSS.n2462 1.49689
R59423 VSS.n2468 VSS.n2467 1.49689
R59424 VSS.n2501 VSS.n2500 1.49689
R59425 VSS.n2506 VSS.n2505 1.49689
R59426 VSS.n2385 VSS.n2384 1.49689
R59427 VSS.n2390 VSS.n2389 1.49689
R59428 VSS.n2415 VSS.n2414 1.49689
R59429 VSS.n2420 VSS.n2419 1.49689
R59430 VSS.n17259 VSS.n17258 1.49689
R59431 VSS.n17264 VSS.n17263 1.49689
R59432 VSS.n17297 VSS.n17296 1.49689
R59433 VSS.n17302 VSS.n17301 1.49689
R59434 VSS.n14245 VSS.n14244 1.49689
R59435 VSS.n13545 VSS.n13544 1.49689
R59436 VSS.n17176 VSS.n17175 1.49689
R59437 VSS.n14316 VSS.n14315 1.49689
R59438 VSS.n4807 VSS.n4806 1.49689
R59439 VSS.n4812 VSS.n4811 1.49689
R59440 VSS.n4845 VSS.n4844 1.49689
R59441 VSS.n4850 VSS.n4849 1.49689
R59442 VSS.n4869 VSS.n4868 1.49689
R59443 VSS.n4874 VSS.n4873 1.49689
R59444 VSS.n4909 VSS.n4908 1.49689
R59445 VSS.n4914 VSS.n4913 1.49689
R59446 VSS.n5424 VSS.n5423 1.49689
R59447 VSS.n5429 VSS.n5428 1.49689
R59448 VSS.n5464 VSS.n5463 1.49689
R59449 VSS.n5469 VSS.n5468 1.49689
R59450 VSS.n5892 VSS.n5891 1.49689
R59451 VSS.n5887 VSS.n5886 1.49689
R59452 VSS.n5887 VSS.n5884 1.49689
R59453 VSS.n5892 VSS.n5889 1.49689
R59454 VSS.n5469 VSS.n5466 1.49689
R59455 VSS.n5464 VSS.n5461 1.49689
R59456 VSS.n5429 VSS.n5426 1.49689
R59457 VSS.n5424 VSS.n5421 1.49689
R59458 VSS.n4914 VSS.n4911 1.49689
R59459 VSS.n4909 VSS.n4906 1.49689
R59460 VSS.n4874 VSS.n4871 1.49689
R59461 VSS.n4869 VSS.n4866 1.49689
R59462 VSS.n4850 VSS.n4847 1.49689
R59463 VSS.n4845 VSS.n4842 1.49689
R59464 VSS.n4812 VSS.n4809 1.49689
R59465 VSS.n4807 VSS.n4804 1.49689
R59466 VSS.n14317 VSS.n14316 1.49689
R59467 VSS.n17177 VSS.n17176 1.49689
R59468 VSS.n13546 VSS.n13545 1.49689
R59469 VSS.n14246 VSS.n14245 1.49689
R59470 VSS.n17302 VSS.n17299 1.49689
R59471 VSS.n17297 VSS.n17294 1.49689
R59472 VSS.n17264 VSS.n17261 1.49689
R59473 VSS.n17259 VSS.n17256 1.49689
R59474 VSS.n2420 VSS.n2417 1.49689
R59475 VSS.n2415 VSS.n2412 1.49689
R59476 VSS.n2390 VSS.n2387 1.49689
R59477 VSS.n2385 VSS.n2382 1.49689
R59478 VSS.n2506 VSS.n2503 1.49689
R59479 VSS.n2501 VSS.n2498 1.49689
R59480 VSS.n2468 VSS.n2465 1.49689
R59481 VSS.n2463 VSS.n2460 1.49689
R59482 VSS.n3932 VSS.n3929 1.49689
R59483 VSS.n3927 VSS.n3924 1.49689
R59484 VSS.n3899 VSS.n3896 1.49689
R59485 VSS.n3894 VSS.n3891 1.49689
R59486 VSS.n179 VSS.n176 1.49689
R59487 VSS.n184 VSS.n181 1.49689
R59488 VSS.n9081 VSS.n9063 1.49632
R59489 VSS.n2663 VSS.n2662 1.49617
R59490 VSS.n9079 VSS.n9078 1.49613
R59491 VSS.n8158 VSS.n8146 1.49541
R59492 VSS.n4101 VSS.n4100 1.49526
R59493 VSS.n4096 VSS.n4095 1.49526
R59494 VSS.n4091 VSS.n4090 1.49526
R59495 VSS.n21891 VSS.n21890 1.49526
R59496 VSS.n21896 VSS.n21895 1.49526
R59497 VSS.n4175 VSS.n4174 1.49526
R59498 VSS.n17411 VSS.n17410 1.49526
R59499 VSS.n2148 VSS.n2147 1.49526
R59500 VSS.n11405 VSS.n11404 1.49526
R59501 VSS.n11400 VSS.n11399 1.49526
R59502 VSS.n11395 VSS.n11394 1.49526
R59503 VSS.n11477 VSS.n11476 1.49526
R59504 VSS.n11482 VSS.n11481 1.49526
R59505 VSS.n11487 VSS.n11486 1.49526
R59506 VSS.n11628 VSS.n11627 1.49526
R59507 VSS.n11623 VSS.n11622 1.49526
R59508 VSS.n11618 VSS.n11617 1.49526
R59509 VSS.n14336 VSS.n14335 1.49526
R59510 VSS.n17180 VSS.n17179 1.49526
R59511 VSS.n14345 VSS.n14344 1.49526
R59512 VSS.n14351 VSS.n14350 1.49526
R59513 VSS.n14361 VSS.n14360 1.49526
R59514 VSS.n14365 VSS.n14364 1.49526
R59515 VSS.n14381 VSS.n14367 1.49526
R59516 VSS.n14373 VSS.n14372 1.49526
R59517 VSS.n14376 VSS.n14375 1.49526
R59518 VSS.n17374 VSS.n17373 1.49526
R59519 VSS.n13537 VSS.n13535 1.49526
R59520 VSS.n13534 VSS.n13532 1.49526
R59521 VSS.n13528 VSS.n13526 1.49526
R59522 VSS.n13518 VSS.n13516 1.49526
R59523 VSS.n13434 VSS.n13432 1.49526
R59524 VSS.n13424 VSS.n13422 1.49526
R59525 VSS.n13276 VSS.n13274 1.49526
R59526 VSS.n13271 VSS.n13269 1.49526
R59527 VSS.n11765 VSS.n11763 1.49526
R59528 VSS.n11762 VSS.n11760 1.49526
R59529 VSS.n11759 VSS.n11757 1.49526
R59530 VSS.n13298 VSS.n13297 1.49526
R59531 VSS.n13293 VSS.n13292 1.49526
R59532 VSS.n18136 VSS.n18135 1.49526
R59533 VSS.n18131 VSS.n18130 1.49526
R59534 VSS.n2141 VSS.n2140 1.49526
R59535 VSS.n8156 VSS.n8155 1.4952
R59536 VSS.n22254 VSS.n22230 1.49219
R59537 VSS.n21987 VSS.n21986 1.49219
R59538 VSS.n14254 VSS.n14253 1.48921
R59539 VSS.n13658 VSS.n13631 1.48921
R59540 VSS.n21987 VSS.n21978 1.48921
R59541 VSS.n22254 VSS.n22175 1.48921
R59542 VSS.n22254 VSS.n22253 1.47742
R59543 VSS.n21987 VSS.n21961 1.47742
R59544 VSS.n18244 VSS.n18243 1.47246
R59545 VSS.n15690 VSS.n15689 1.4635
R59546 VSS.n198 VSS.n197 1.4635
R59547 VSS.n157 VSS.n156 1.36071
R59548 VSS.n94 VSS.n93 1.36071
R59549 VSS.n69 VSS.n68 1.36071
R59550 VSS.n62 VSS.n61 1.36071
R59551 VSS.n221 VSS.n220 1.36071
R59552 VSS.n253 VSS.n252 1.36071
R59553 VSS.n285 VSS.n284 1.36071
R59554 VSS.n4112 VSS.n4111 1.36071
R59555 VSS.n11262 VSS.n11261 1.36071
R59556 VSS.n11267 VSS.n11266 1.36071
R59557 VSS.n11272 VSS.n11271 1.36071
R59558 VSS.n11277 VSS.n11276 1.36071
R59559 VSS.n11286 VSS.n11285 1.36071
R59560 VSS.n11291 VSS.n11290 1.36071
R59561 VSS.n11296 VSS.n11295 1.36071
R59562 VSS.n11307 VSS.n11306 1.36071
R59563 VSS.n15182 VSS.n15181 1.36071
R59564 VSS.n15187 VSS.n15186 1.36071
R59565 VSS.n15192 VSS.n15191 1.36071
R59566 VSS.n15913 VSS.n15912 1.36071
R59567 VSS.n15904 VSS.n15903 1.36071
R59568 VSS.n15197 VSS.n15196 1.36071
R59569 VSS.n15676 VSS.n15675 1.36071
R59570 VSS.n1478 VSS.n1477 1.36071
R59571 VSS.n1473 VSS.n1472 1.36071
R59572 VSS.n875 VSS.n874 1.36071
R59573 VSS.n870 VSS.n869 1.36071
R59574 VSS.n865 VSS.n864 1.36071
R59575 VSS.n860 VSS.n859 1.36071
R59576 VSS.n451 VSS.n450 1.36071
R59577 VSS.n456 VSS.n455 1.36071
R59578 VSS.n21194 VSS.n21193 1.36071
R59579 VSS.n21199 VSS.n21198 1.36071
R59580 VSS.n21208 VSS.n21207 1.36071
R59581 VSS.n21213 VSS.n21212 1.36071
R59582 VSS.n21218 VSS.n21217 1.36071
R59583 VSS.n21223 VSS.n21222 1.36071
R59584 VSS.n374 VSS.n373 1.36071
R59585 VSS.n21908 VSS.n21907 1.36071
R59586 VSS.n323 VSS.n322 1.36071
R59587 VSS.n50 VSS.n49 1.36071
R59588 VSS.n45 VSS.n44 1.36071
R59589 VSS.n39 VSS.n38 1.36071
R59590 VSS.n298 VSS.n297 1.36071
R59591 VSS.n304 VSS.n303 1.36071
R59592 VSS.n310 VSS.n309 1.36071
R59593 VSS.n266 VSS.n265 1.36071
R59594 VSS.n272 VSS.n271 1.36071
R59595 VSS.n278 VSS.n277 1.36071
R59596 VSS.n234 VSS.n233 1.36071
R59597 VSS.n240 VSS.n239 1.36071
R59598 VSS.n246 VSS.n245 1.36071
R59599 VSS.n210 VSS.n209 1.36071
R59600 VSS.n215 VSS.n214 1.36071
R59601 VSS.n144 VSS.n143 1.36071
R59602 VSS.n138 VSS.n137 1.36071
R59603 VSS.n132 VSS.n131 1.36071
R59604 VSS.n125 VSS.n124 1.36071
R59605 VSS.n113 VSS.n112 1.36071
R59606 VSS.n107 VSS.n106 1.36071
R59607 VSS.n81 VSS.n80 1.36071
R59608 VSS.n75 VSS.n74 1.36071
R59609 VSS.n101 VSS.n100 1.36071
R59610 VSS.n16294 VSS.n16293 1.35477
R59611 VSS.n1380 VSS.n1379 1.35477
R59612 VSS.n5641 VSS.n5640 1.35477
R59613 VSS.n20905 VSS.n20904 1.35477
R59614 VSS.n12816 VSS.n12815 1.30851
R59615 VSS.n7546 VSS.n7545 1.30851
R59616 VSS.n11235 VSS.n11234 1.30851
R59617 VSS.n515 VSS.n514 1.30851
R59618 VSS.n12615 VSS.n12614 1.3005
R59619 VSS.n12614 VSS.n12613 1.3005
R59620 VSS.n12627 VSS.n12626 1.3005
R59621 VSS.n12626 VSS.n12625 1.3005
R59622 VSS.n6824 VSS.n6823 1.3005
R59623 VSS.n6823 VSS.n6822 1.3005
R59624 VSS.n6818 VSS.n6817 1.3005
R59625 VSS.n6817 VSS.n6816 1.3005
R59626 VSS.n8653 VSS.n8652 1.3005
R59627 VSS.n8652 VSS.n8651 1.3005
R59628 VSS.n8502 VSS.n8501 1.3005
R59629 VSS.n8501 VSS.n8500 1.3005
R59630 VSS.n9643 VSS.n9642 1.3005
R59631 VSS.n9642 VSS.n9641 1.3005
R59632 VSS.n9628 VSS.n9627 1.3005
R59633 VSS.n9627 VSS.n9626 1.3005
R59634 VSS.n9526 VSS.n9525 1.3005
R59635 VSS.n9525 VSS.n9524 1.3005
R59636 VSS.n9511 VSS.n9510 1.3005
R59637 VSS.n9510 VSS.n9509 1.3005
R59638 VSS.n9517 VSS.n9516 1.3005
R59639 VSS.n9516 VSS.n9515 1.3005
R59640 VSS.n9520 VSS.n9519 1.3005
R59641 VSS.n9519 VSS.n9518 1.3005
R59642 VSS.n9634 VSS.n9633 1.3005
R59643 VSS.n9633 VSS.n9632 1.3005
R59644 VSS.n9637 VSS.n9636 1.3005
R59645 VSS.n9636 VSS.n9635 1.3005
R59646 VSS.n8493 VSS.n8492 1.3005
R59647 VSS.n8492 VSS.n8491 1.3005
R59648 VSS.n8644 VSS.n8643 1.3005
R59649 VSS.n8643 VSS.n8642 1.3005
R59650 VSS.n8647 VSS.n8646 1.3005
R59651 VSS.n8646 VSS.n8645 1.3005
R59652 VSS.n6830 VSS.n6829 1.3005
R59653 VSS.n6829 VSS.n6828 1.3005
R59654 VSS.n12609 VSS.n12608 1.3005
R59655 VSS.n12608 VSS.n12607 1.3005
R59656 VSS.n12621 VSS.n12620 1.3005
R59657 VSS.n12620 VSS.n12619 1.3005
R59658 VSS.n12633 VSS.n12632 1.3005
R59659 VSS.n12632 VSS.n12631 1.3005
R59660 VSS.n9841 VSS.n9840 1.3005
R59661 VSS.n9840 VSS.n9839 1.3005
R59662 VSS.n9054 VSS.n9053 1.3005
R59663 VSS.n9053 VSS.n9052 1.3005
R59664 VSS.n8143 VSS.n8142 1.3005
R59665 VSS.n8142 VSS.n8141 1.3005
R59666 VSS.n6541 VSS.n6540 1.3005
R59667 VSS.n6540 VSS.n6539 1.3005
R59668 VSS.n9236 VSS.n9235 1.3005
R59669 VSS.n9235 VSS.n9234 1.3005
R59670 VSS.n9210 VSS.n9209 1.3005
R59671 VSS.n9209 VSS.n9208 1.3005
R59672 VSS.n6392 VSS.n6391 1.3005
R59673 VSS.n6391 VSS.n6390 1.3005
R59674 VSS.n6551 VSS.n6550 1.3005
R59675 VSS.n6550 VSS.n6549 1.3005
R59676 VSS.n6544 VSS.n6543 1.3005
R59677 VSS.n6543 VSS.n6542 1.3005
R59678 VSS.n6557 VSS.n6556 1.3005
R59679 VSS.n6556 VSS.n6555 1.3005
R59680 VSS.n6409 VSS.n6408 1.3005
R59681 VSS.n6408 VSS.n6407 1.3005
R59682 VSS.n6397 VSS.n6396 1.3005
R59683 VSS.n6396 VSS.n6395 1.3005
R59684 VSS.n6406 VSS.n6405 1.3005
R59685 VSS.n6405 VSS.n6404 1.3005
R59686 VSS.n6386 VSS.n6385 1.3005
R59687 VSS.n6385 VSS.n6384 1.3005
R59688 VSS.n8152 VSS.n8151 1.3005
R59689 VSS.n8151 VSS.n8150 1.3005
R59690 VSS.n9204 VSS.n9203 1.3005
R59691 VSS.n9203 VSS.n9202 1.3005
R59692 VSS.n9216 VSS.n9215 1.3005
R59693 VSS.n9215 VSS.n9214 1.3005
R59694 VSS.n9239 VSS.n9238 1.3005
R59695 VSS.n9238 VSS.n9237 1.3005
R59696 VSS.n9222 VSS.n9221 1.3005
R59697 VSS.n9221 VSS.n9220 1.3005
R59698 VSS.n9230 VSS.n9229 1.3005
R59699 VSS.n9229 VSS.n9228 1.3005
R59700 VSS.n9075 VSS.n9074 1.3005
R59701 VSS.n9074 VSS.n9073 1.3005
R59702 VSS.n9069 VSS.n9068 1.3005
R59703 VSS.n9068 VSS.n9067 1.3005
R59704 VSS.n9060 VSS.n9059 1.3005
R59705 VSS.n9059 VSS.n9058 1.3005
R59706 VSS.n16266 VSS.n16265 1.24924
R59707 VSS.n16301 VSS.n16300 1.24924
R59708 VSS.n16342 VSS.n16340 1.24924
R59709 VSS.n5695 VSS.n5694 1.24924
R59710 VSS.n5704 VSS.n5703 1.24924
R59711 VSS.n5764 VSS.n5762 1.24924
R59712 VSS.n17178 VSS.n14378 1.23547
R59713 VSS.n17178 VSS.n17174 1.23547
R59714 VSS.n4905 VSS.n4903 1.23547
R59715 VSS.n4905 VSS.n4904 1.23547
R59716 VSS.n5460 VSS.n5458 1.23547
R59717 VSS.n5460 VSS.n5459 1.23547
R59718 VSS.n1350 VSS.n1349 1.23166
R59719 VSS.n1384 VSS.n1383 1.23166
R59720 VSS.n1430 VSS.n1428 1.23166
R59721 VSS.n20964 VSS.n20963 1.23166
R59722 VSS.n20975 VSS.n20973 1.23166
R59723 VSS.n1217 VSS.n1216 1.23166
R59724 VSS.n5876 VSS.n5875 1.17298
R59725 VSS.n21185 VSS.n21184 1.17298
R59726 VSS.n12010 VSS.n11998 1.14278
R59727 VSS.n8876 VSS.n8875 1.13013
R59728 VSS.n15702 VSS.n15701 1.1255
R59729 VSS.n15901 VSS.n15900 1.1255
R59730 VSS.n9514 VSS.n9513 1.1255
R59731 VSS.n9513 VSS.n9512 1.1255
R59732 VSS.n9529 VSS.n9528 1.1255
R59733 VSS.n9528 VSS.n9527 1.1255
R59734 VSS.n9523 VSS.n9522 1.1255
R59735 VSS.n9522 VSS.n9521 1.1255
R59736 VSS.n9625 VSS.n9624 1.1255
R59737 VSS.n9624 VSS.n9623 1.1255
R59738 VSS.n9631 VSS.n9630 1.1255
R59739 VSS.n9630 VSS.n9629 1.1255
R59740 VSS.n9646 VSS.n9645 1.1255
R59741 VSS.n9645 VSS.n9644 1.1255
R59742 VSS.n9640 VSS.n9639 1.1255
R59743 VSS.n9639 VSS.n9638 1.1255
R59744 VSS.n8490 VSS.n8489 1.1255
R59745 VSS.n8489 VSS.n8488 1.1255
R59746 VSS.n8505 VSS.n8504 1.1255
R59747 VSS.n8504 VSS.n8503 1.1255
R59748 VSS.n8499 VSS.n8498 1.1255
R59749 VSS.n8498 VSS.n8497 1.1255
R59750 VSS.n8641 VSS.n8640 1.1255
R59751 VSS.n8640 VSS.n8639 1.1255
R59752 VSS.n8656 VSS.n8655 1.1255
R59753 VSS.n8655 VSS.n8654 1.1255
R59754 VSS.n8650 VSS.n8649 1.1255
R59755 VSS.n8649 VSS.n8648 1.1255
R59756 VSS.n6815 VSS.n6814 1.1255
R59757 VSS.n6814 VSS.n6813 1.1255
R59758 VSS.n6833 VSS.n6832 1.1255
R59759 VSS.n6832 VSS.n6831 1.1255
R59760 VSS.n6827 VSS.n6826 1.1255
R59761 VSS.n6826 VSS.n6825 1.1255
R59762 VSS.n6821 VSS.n6820 1.1255
R59763 VSS.n6820 VSS.n6819 1.1255
R59764 VSS.n12612 VSS.n12611 1.1255
R59765 VSS.n12611 VSS.n12610 1.1255
R59766 VSS.n12618 VSS.n12617 1.1255
R59767 VSS.n12617 VSS.n12616 1.1255
R59768 VSS.n12624 VSS.n12623 1.1255
R59769 VSS.n12623 VSS.n12622 1.1255
R59770 VSS.n12630 VSS.n12629 1.1255
R59771 VSS.n12629 VSS.n12628 1.1255
R59772 VSS.n9508 VSS.n9507 1.1255
R59773 VSS.n9507 VSS.n9506 1.1255
R59774 VSS.n6560 VSS.n6559 1.1255
R59775 VSS.n6559 VSS.n6558 1.1255
R59776 VSS.n6554 VSS.n6553 1.1255
R59777 VSS.n6553 VSS.n6552 1.1255
R59778 VSS.n6538 VSS.n6537 1.1255
R59779 VSS.n6537 VSS.n6536 1.1255
R59780 VSS.n6398 VSS.n6394 1.1255
R59781 VSS.n6394 VSS.n6393 1.1255
R59782 VSS.n6403 VSS.n6402 1.1255
R59783 VSS.n6402 VSS.n6401 1.1255
R59784 VSS.n6412 VSS.n6411 1.1255
R59785 VSS.n6411 VSS.n6410 1.1255
R59786 VSS.n6389 VSS.n6388 1.1255
R59787 VSS.n6388 VSS.n6387 1.1255
R59788 VSS.n8155 VSS.n8154 1.1255
R59789 VSS.n8154 VSS.n8153 1.1255
R59790 VSS.n6383 VSS.n6382 1.1255
R59791 VSS.n6382 VSS.n6381 1.1255
R59792 VSS.n8146 VSS.n8145 1.1255
R59793 VSS.n8145 VSS.n8144 1.1255
R59794 VSS.n9207 VSS.n9206 1.1255
R59795 VSS.n9206 VSS.n9205 1.1255
R59796 VSS.n9201 VSS.n9200 1.1255
R59797 VSS.n9200 VSS.n9199 1.1255
R59798 VSS.n9213 VSS.n9212 1.1255
R59799 VSS.n9212 VSS.n9211 1.1255
R59800 VSS.n9242 VSS.n9241 1.1255
R59801 VSS.n9241 VSS.n9240 1.1255
R59802 VSS.n9225 VSS.n9224 1.1255
R59803 VSS.n9224 VSS.n9223 1.1255
R59804 VSS.n9219 VSS.n9218 1.1255
R59805 VSS.n9218 VSS.n9217 1.1255
R59806 VSS.n9233 VSS.n9232 1.1255
R59807 VSS.n9232 VSS.n9231 1.1255
R59808 VSS.n9072 VSS.n9071 1.1255
R59809 VSS.n9071 VSS.n9070 1.1255
R59810 VSS.n9078 VSS.n9077 1.1255
R59811 VSS.n9077 VSS.n9076 1.1255
R59812 VSS.n9057 VSS.n9056 1.1255
R59813 VSS.n9056 VSS.n9055 1.1255
R59814 VSS.n9063 VSS.n9062 1.1255
R59815 VSS.n9062 VSS.n9061 1.1255
R59816 VSS.n6547 VSS.n6546 1.1255
R59817 VSS.n6546 VSS.n6545 1.1255
R59818 VSS.n1469 VSS.n1467 1.12142
R59819 VSS.n21195 VSS.n21192 1.12142
R59820 VSS.n16384 VSS.n15914 1.12142
R59821 VSS.n11309 VSS.n11308 1.12142
R59822 VSS.n21246 VSS.n21245 1.12124
R59823 VSS.n17386 VSS.n17385 1.12124
R59824 VSS.n17239 VSS.n17238 1.12124
R59825 VSS.n11640 VSS.n11639 1.12124
R59826 VSS.n11466 VSS.n11465 1.12124
R59827 VSS.n11417 VSS.n11416 1.12124
R59828 VSS.n11251 VSS.n11250 1.12124
R59829 VSS.n11602 VSS.n11593 1.12072
R59830 VSS.n11512 VSS.n11511 1.12072
R59831 VSS.n11379 VSS.n11370 1.12072
R59832 VSS.n13262 VSS.n13254 1.12072
R59833 VSS.n13262 VSS.n12999 1.12072
R59834 VSS.n17539 VSS.n17482 1.12072
R59835 VSS.n14433 VSS.n14431 1.12072
R59836 VSS.n15098 VSS.n15097 1.12072
R59837 VSS.n15131 VSS.n15130 1.12072
R59838 VSS.n16389 VSS.n16387 1.12072
R59839 VSS.n18106 VSS.n18105 1.12072
R59840 VSS.n20297 VSS.n682 1.12072
R59841 VSS.n13406 VSS.n13405 1.12072
R59842 VSS.n13421 VSS.n13420 1.12072
R59843 VSS.n20728 VSS.n20727 1.12072
R59844 VSS.n20779 VSS.n20778 1.12072
R59845 VSS.n20871 VSS.n20870 1.12072
R59846 VSS.n20604 VSS.n20590 1.12072
R59847 VSS.n17813 VSS.n2337 1.12072
R59848 VSS.n9243 VSS.n9242 1.12072
R59849 VSS.n6563 VSS.n6547 1.12072
R59850 VSS.n6561 VSS.n6560 1.12072
R59851 VSS.n9226 VSS.n9225 1.12072
R59852 VSS.n13511 VSS.n13459 1.12072
R59853 VSS.n13515 VSS.n13514 1.12072
R59854 VSS.n20068 VSS.n20067 1.12072
R59855 VSS.n2069 VSS.n2060 1.12072
R59856 VSS.n1995 VSS.n1994 1.12072
R59857 VSS.n20167 VSS.n20166 1.12072
R59858 VSS.n17967 VSS.n17966 1.12072
R59859 VSS.n6413 VSS.n6412 1.12072
R59860 VSS.n7564 VSS.n7541 1.12072
R59861 VSS.n9342 VSS.n9320 1.12072
R59862 VSS.n7851 VSS.n7850 1.12072
R59863 VSS.n9396 VSS.n9157 1.12072
R59864 VSS.n6699 VSS.n6685 1.12072
R59865 VSS.n6759 VSS.n6535 1.12072
R59866 VSS.n8075 VSS.n6904 1.12072
R59867 VSS.n8024 VSS.n7006 1.12072
R59868 VSS.n9778 VSS.n9594 1.12072
R59869 VSS.n9724 VSS.n9711 1.12072
R59870 VSS.n3847 VSS.n3184 1.12072
R59871 VSS.n4695 VSS.n4694 1.12072
R59872 VSS.n4755 VSS.n4754 1.12072
R59873 VSS.n11218 VSS.n5923 1.12072
R59874 VSS.n11721 VSS.n11720 1.12072
R59875 VSS.n11439 VSS.n5413 1.12072
R59876 VSS.n3810 VSS.n3779 1.12072
R59877 VSS.n11184 VSS.n11183 1.12072
R59878 VSS.n3289 VSS.n3288 1.12072
R59879 VSS.n20374 VSS.n680 1.12072
R59880 VSS.n10626 VSS.n10625 1.12072
R59881 VSS.n9530 VSS.n9529 1.12072
R59882 VSS.n9647 VSS.n9646 1.12072
R59883 VSS.n6834 VSS.n6833 1.12072
R59884 VSS.n17354 VSS.n17350 1.12053
R59885 VSS.n4636 VSS.n4211 1.12053
R59886 VSS.n20351 VSS.n681 1.12053
R59887 VSS.n6399 VSS.n6398 1.12053
R59888 VSS.n1934 VSS.n1479 1.12051
R59889 VSS.n15905 VSS.n15902 1.12051
R59890 VSS.n14670 VSS.n14669 1.11968
R59891 VSS.n17166 VSS.n17165 1.11968
R59892 VSS.n16873 VSS.n14943 1.11968
R59893 VSS.n16684 VSS.n14972 1.11968
R59894 VSS.n16433 VSS.n16432 1.11968
R59895 VSS.n8431 VSS.n8430 1.11968
R59896 VSS.n8763 VSS.n8575 1.11968
R59897 VSS.n8727 VSS.n8726 1.11968
R59898 VSS.n8270 VSS.n8238 1.11968
R59899 VSS.n19767 VSS.n2137 1.11968
R59900 VSS.n19857 VSS.n2131 1.11968
R59901 VSS.n20044 VSS.n20042 1.11968
R59902 VSS.n2086 VSS.n2085 1.11968
R59903 VSS.n1971 VSS.n1969 1.11968
R59904 VSS.n8506 VSS.n8505 1.11968
R59905 VSS.n8657 VSS.n8656 1.11968
R59906 VSS.n14208 VSS.n14207 1.11241
R59907 VSS.n17232 VSS.n17231 1.11241
R59908 VSS.n17232 VSS.n11748 1.11241
R59909 VSS.n17587 VSS.n17585 1.11241
R59910 VSS.n17587 VSS.n17586 1.11241
R59911 VSS.n17579 VSS.n2341 1.11241
R59912 VSS.n4666 VSS.n4651 1.11241
R59913 VSS.n4671 VSS.n2448 1.11241
R59914 VSS.n4666 VSS.n4665 1.11241
R59915 VSS.n4666 VSS.n2449 1.11241
R59916 VSS.n4671 VSS.n4670 1.11241
R59917 VSS.n4671 VSS.n2447 1.11241
R59918 VSS.n17579 VSS.n2342 1.11241
R59919 VSS.n17579 VSS.n2339 1.11241
R59920 VSS.n14148 VSS.n14131 1.11241
R59921 VSS.n14274 VSS.n14254 1.10465
R59922 VSS.n13658 VSS.n13657 1.10465
R59923 VSS.n14254 VSS.n13611 1.10458
R59924 VSS.n21987 VSS.n21944 1.10458
R59925 VSS.n8876 VSS.n8873 1.05973
R59926 VSS.n8876 VSS.n8872 1.05973
R59927 VSS.n11991 VSS.n11989 1.05973
R59928 VSS.n11991 VSS.n11988 1.05973
R59929 VSS.n12010 VSS.n12005 1.05973
R59930 VSS.n8864 VSS.n8854 1.05973
R59931 VSS.n21426 VSS.n392 0.897595
R59932 VSS.n21415 VSS.n393 0.897595
R59933 VSS.n21316 VSS.n410 0.897595
R59934 VSS.n21305 VSS.n427 0.897595
R59935 VSS.n21253 VSS.n444 0.897595
R59936 VSS.n15692 VSS.n15691 0.87334
R59937 VSS.n15206 VSS.n15205 0.867167
R59938 VSS.n15644 VSS.n15643 0.867167
R59939 VSS.n15507 VSS.n15506 0.867167
R59940 VSS.n1847 VSS.n1846 0.867167
R59941 VSS.n12661 VSS.n12659 0.771929
R59942 VSS.n12663 VSS.n12661 0.771929
R59943 VSS.n12665 VSS.n12663 0.771929
R59944 VSS.n12667 VSS.n12665 0.771929
R59945 VSS.n12671 VSS.n12667 0.771929
R59946 VSS.n12671 VSS.n12669 0.771929
R59947 VSS.n12599 VSS.n12597 0.771929
R59948 VSS.n11775 VSS.n11773 0.771929
R59949 VSS.n11783 VSS.n11781 0.771929
R59950 VSS.n12570 VSS.n12568 0.771929
R59951 VSS.n12336 VSS.n12334 0.771929
R59952 VSS.n12344 VSS.n12342 0.771929
R59953 VSS.n12351 VSS.n12349 0.771929
R59954 VSS.n12358 VSS.n12356 0.771929
R59955 VSS.n12366 VSS.n12364 0.771929
R59956 VSS.n12374 VSS.n12372 0.771929
R59957 VSS.n12501 VSS.n12497 0.771929
R59958 VSS.n12501 VSS.n12499 0.771929
R59959 VSS.n12492 VSS.n12490 0.771929
R59960 VSS.n12484 VSS.n12482 0.771929
R59961 VSS.n12476 VSS.n12474 0.771929
R59962 VSS.n12469 VSS.n12467 0.771929
R59963 VSS.n12462 VSS.n12460 0.771929
R59964 VSS.n12454 VSS.n12452 0.771929
R59965 VSS.n12446 VSS.n12444 0.771929
R59966 VSS.n12438 VSS.n12436 0.771929
R59967 VSS.n12430 VSS.n12428 0.771929
R59968 VSS.n12422 VSS.n12420 0.771929
R59969 VSS.n12414 VSS.n12412 0.771929
R59970 VSS.n12407 VSS.n12405 0.771929
R59971 VSS.n12400 VSS.n12398 0.771929
R59972 VSS.n12392 VSS.n12390 0.771929
R59973 VSS.n12385 VSS.n12383 0.771929
R59974 VSS.n12213 VSS.n12209 0.771929
R59975 VSS.n12213 VSS.n12211 0.771929
R59976 VSS.n12204 VSS.n12202 0.771929
R59977 VSS.n12196 VSS.n12194 0.771929
R59978 VSS.n12188 VSS.n12186 0.771929
R59979 VSS.n12181 VSS.n12179 0.771929
R59980 VSS.n12174 VSS.n12172 0.771929
R59981 VSS.n12166 VSS.n12164 0.771929
R59982 VSS.n12158 VSS.n12156 0.771929
R59983 VSS.n12150 VSS.n12148 0.771929
R59984 VSS.n12142 VSS.n12140 0.771929
R59985 VSS.n12134 VSS.n12132 0.771929
R59986 VSS.n12126 VSS.n12124 0.771929
R59987 VSS.n12119 VSS.n12117 0.771929
R59988 VSS.n12112 VSS.n12110 0.771929
R59989 VSS.n12104 VSS.n12102 0.771929
R59990 VSS.n12096 VSS.n12094 0.771929
R59991 VSS.n12088 VSS.n12086 0.771929
R59992 VSS.n12080 VSS.n12078 0.771929
R59993 VSS.n12072 VSS.n12070 0.771929
R59994 VSS.n12065 VSS.n12063 0.771929
R59995 VSS.n12058 VSS.n12056 0.771929
R59996 VSS.n12050 VSS.n12048 0.771929
R59997 VSS.n12042 VSS.n12040 0.771929
R59998 VSS.n12034 VSS.n12032 0.771929
R59999 VSS.n12026 VSS.n12024 0.771929
R60000 VSS.n12018 VSS.n12016 0.771929
R60001 VSS.n12010 VSS.n12009 0.771929
R60002 VSS.n12009 VSS.n12007 0.771929
R60003 VSS.n12007 VSS.n12006 0.771929
R60004 VSS.n11982 VSS.n11981 0.771929
R60005 VSS.n11987 VSS.n11986 0.771929
R60006 VSS.n11991 VSS.n11987 0.771929
R60007 VSS.n9856 VSS.n9854 0.771929
R60008 VSS.n9858 VSS.n9856 0.771929
R60009 VSS.n9860 VSS.n9858 0.771929
R60010 VSS.n9862 VSS.n9860 0.771929
R60011 VSS.n9866 VSS.n9862 0.771929
R60012 VSS.n9866 VSS.n9864 0.771929
R60013 VSS.n10533 VSS.n10531 0.771929
R60014 VSS.n9874 VSS.n9872 0.771929
R60015 VSS.n9882 VSS.n9880 0.771929
R60016 VSS.n9891 VSS.n9889 0.771929
R60017 VSS.n10282 VSS.n10280 0.771929
R60018 VSS.n10290 VSS.n10288 0.771929
R60019 VSS.n10297 VSS.n10295 0.771929
R60020 VSS.n10304 VSS.n10302 0.771929
R60021 VSS.n10312 VSS.n10310 0.771929
R60022 VSS.n10320 VSS.n10318 0.771929
R60023 VSS.n10447 VSS.n10443 0.771929
R60024 VSS.n10447 VSS.n10445 0.771929
R60025 VSS.n10438 VSS.n10436 0.771929
R60026 VSS.n10430 VSS.n10428 0.771929
R60027 VSS.n10422 VSS.n10420 0.771929
R60028 VSS.n10415 VSS.n10413 0.771929
R60029 VSS.n10408 VSS.n10406 0.771929
R60030 VSS.n10400 VSS.n10398 0.771929
R60031 VSS.n10392 VSS.n10390 0.771929
R60032 VSS.n10384 VSS.n10382 0.771929
R60033 VSS.n10376 VSS.n10374 0.771929
R60034 VSS.n10368 VSS.n10366 0.771929
R60035 VSS.n10360 VSS.n10358 0.771929
R60036 VSS.n10353 VSS.n10351 0.771929
R60037 VSS.n10346 VSS.n10344 0.771929
R60038 VSS.n10338 VSS.n10336 0.771929
R60039 VSS.n10331 VSS.n10329 0.771929
R60040 VSS.n10162 VSS.n10158 0.771929
R60041 VSS.n10162 VSS.n10160 0.771929
R60042 VSS.n10153 VSS.n10151 0.771929
R60043 VSS.n10145 VSS.n10143 0.771929
R60044 VSS.n10137 VSS.n10135 0.771929
R60045 VSS.n10130 VSS.n10128 0.771929
R60046 VSS.n10123 VSS.n10121 0.771929
R60047 VSS.n10115 VSS.n10113 0.771929
R60048 VSS.n10107 VSS.n10105 0.771929
R60049 VSS.n10099 VSS.n10097 0.771929
R60050 VSS.n10091 VSS.n10089 0.771929
R60051 VSS.n10083 VSS.n10081 0.771929
R60052 VSS.n10075 VSS.n10073 0.771929
R60053 VSS.n10068 VSS.n10066 0.771929
R60054 VSS.n10061 VSS.n10059 0.771929
R60055 VSS.n10053 VSS.n10051 0.771929
R60056 VSS.n10045 VSS.n10043 0.771929
R60057 VSS.n10037 VSS.n10035 0.771929
R60058 VSS.n10029 VSS.n10027 0.771929
R60059 VSS.n10021 VSS.n10019 0.771929
R60060 VSS.n10014 VSS.n10012 0.771929
R60061 VSS.n10007 VSS.n10005 0.771929
R60062 VSS.n9999 VSS.n9997 0.771929
R60063 VSS.n9991 VSS.n9989 0.771929
R60064 VSS.n9983 VSS.n9981 0.771929
R60065 VSS.n8961 VSS.n8957 0.771929
R60066 VSS.n8961 VSS.n8959 0.771929
R60067 VSS.n8864 VSS.n8860 0.771929
R60068 VSS.n8860 VSS.n8858 0.771929
R60069 VSS.n8858 VSS.n8856 0.771929
R60070 VSS.n8867 VSS.n8866 0.771929
R60071 VSS.n8876 VSS.n8871 0.771929
R60072 VSS.n8858 VSS.n8857 0.754407
R60073 VSS.n12579 VSS.n11785 0.7505
R60074 VSS.n12602 VSS.n12601 0.7505
R60075 VSS.n12573 VSS.n12572 0.7505
R60076 VSS.n12586 VSS.n11777 0.7505
R60077 VSS.n10541 VSS.n9868 0.7505
R60078 VSS.n8838 VSS.n8837 0.7505
R60079 VSS.n10514 VSS.n9884 0.7505
R60080 VSS.n10521 VSS.n9876 0.7505
R60081 VSS.n10536 VSS.n10535 0.7505
R60082 VSS.n10508 VSS.n9893 0.7505
R60083 VSS.n8965 VSS.n8964 0.7505
R60084 VSS.n8899 VSS.n8888 0.7505
R60085 VSS.n12673 VSS.n12672 0.7505
R60086 VSS.n12010 VSS.n12001 0.748877
R60087 VSS.n11991 VSS.n11990 0.7005
R60088 VSS.n8876 VSS.n8874 0.7005
R60089 VSS.n9849 VSS.n9848 0.696929
R60090 VSS.n9856 VSS.n9855 0.696929
R60091 VSS.n10283 VSS.n10282 0.696929
R60092 VSS.n10282 VSS.n10281 0.696929
R60093 VSS.n10291 VSS.n10290 0.696929
R60094 VSS.n10290 VSS.n10289 0.696929
R60095 VSS.n10423 VSS.n10422 0.696929
R60096 VSS.n10422 VSS.n10421 0.696929
R60097 VSS.n10385 VSS.n10384 0.696929
R60098 VSS.n10384 VSS.n10383 0.696929
R60099 VSS.n10377 VSS.n10376 0.696929
R60100 VSS.n10376 VSS.n10375 0.696929
R60101 VSS.n10361 VSS.n10360 0.696929
R60102 VSS.n10360 VSS.n10359 0.696929
R60103 VSS.n10146 VSS.n10145 0.696929
R60104 VSS.n10145 VSS.n10144 0.696929
R60105 VSS.n10138 VSS.n10137 0.696929
R60106 VSS.n10137 VSS.n10136 0.696929
R60107 VSS.n10100 VSS.n10099 0.696929
R60108 VSS.n10099 VSS.n10098 0.696929
R60109 VSS.n10084 VSS.n10083 0.696929
R60110 VSS.n10083 VSS.n10082 0.696929
R60111 VSS.n10076 VSS.n10075 0.696929
R60112 VSS.n10075 VSS.n10074 0.696929
R60113 VSS.n10030 VSS.n10029 0.696929
R60114 VSS.n10029 VSS.n10028 0.696929
R60115 VSS.n10022 VSS.n10021 0.696929
R60116 VSS.n10021 VSS.n10020 0.696929
R60117 VSS.n8836 VSS.n8835 0.696929
R60118 VSS.n8835 VSS.n8834 0.696929
R60119 VSS.n10275 VSS.n10274 0.696929
R60120 VSS.n10274 VSS.n10273 0.696929
R60121 VSS.n10305 VSS.n10304 0.696929
R60122 VSS.n10304 VSS.n10303 0.696929
R60123 VSS.n10313 VSS.n10312 0.696929
R60124 VSS.n10312 VSS.n10311 0.696929
R60125 VSS.n10321 VSS.n10320 0.696929
R60126 VSS.n10320 VSS.n10319 0.696929
R60127 VSS.n10439 VSS.n10438 0.696929
R60128 VSS.n10438 VSS.n10437 0.696929
R60129 VSS.n10431 VSS.n10430 0.696929
R60130 VSS.n10430 VSS.n10429 0.696929
R60131 VSS.n10409 VSS.n10408 0.696929
R60132 VSS.n10408 VSS.n10407 0.696929
R60133 VSS.n10401 VSS.n10400 0.696929
R60134 VSS.n10400 VSS.n10399 0.696929
R60135 VSS.n10393 VSS.n10392 0.696929
R60136 VSS.n10392 VSS.n10391 0.696929
R60137 VSS.n10369 VSS.n10368 0.696929
R60138 VSS.n10368 VSS.n10367 0.696929
R60139 VSS.n10347 VSS.n10346 0.696929
R60140 VSS.n10346 VSS.n10345 0.696929
R60141 VSS.n10339 VSS.n10338 0.696929
R60142 VSS.n10338 VSS.n10337 0.696929
R60143 VSS.n10163 VSS.n10162 0.696929
R60144 VSS.n10162 VSS.n10161 0.696929
R60145 VSS.n10154 VSS.n10153 0.696929
R60146 VSS.n10153 VSS.n10152 0.696929
R60147 VSS.n10124 VSS.n10123 0.696929
R60148 VSS.n10123 VSS.n10122 0.696929
R60149 VSS.n10116 VSS.n10115 0.696929
R60150 VSS.n10115 VSS.n10114 0.696929
R60151 VSS.n10108 VSS.n10107 0.696929
R60152 VSS.n10107 VSS.n10106 0.696929
R60153 VSS.n10092 VSS.n10091 0.696929
R60154 VSS.n10091 VSS.n10090 0.696929
R60155 VSS.n10062 VSS.n10061 0.696929
R60156 VSS.n10061 VSS.n10060 0.696929
R60157 VSS.n10054 VSS.n10053 0.696929
R60158 VSS.n10053 VSS.n10052 0.696929
R60159 VSS.n10046 VSS.n10045 0.696929
R60160 VSS.n10045 VSS.n10044 0.696929
R60161 VSS.n10038 VSS.n10037 0.696929
R60162 VSS.n10037 VSS.n10036 0.696929
R60163 VSS.n10008 VSS.n10007 0.696929
R60164 VSS.n10007 VSS.n10006 0.696929
R60165 VSS.n10000 VSS.n9999 0.696929
R60166 VSS.n9999 VSS.n9998 0.696929
R60167 VSS.n9992 VSS.n9991 0.696929
R60168 VSS.n9991 VSS.n9990 0.696929
R60169 VSS.n9883 VSS.n9882 0.696929
R60170 VSS.n9882 VSS.n9881 0.696929
R60171 VSS.n9875 VSS.n9874 0.696929
R60172 VSS.n9874 VSS.n9873 0.696929
R60173 VSS.n10534 VSS.n10533 0.696929
R60174 VSS.n10533 VSS.n10532 0.696929
R60175 VSS.n9892 VSS.n9891 0.696929
R60176 VSS.n9891 VSS.n9890 0.696929
R60177 VSS.n9984 VSS.n9983 0.696929
R60178 VSS.n9983 VSS.n9982 0.696929
R60179 VSS.n9860 VSS.n9859 0.696929
R60180 VSS.n8962 VSS.n8961 0.696929
R60181 VSS.n8961 VSS.n8960 0.696929
R60182 VSS.n9838 VSS.n9837 0.696929
R60183 VSS.n12011 VSS.n12010 0.696929
R60184 VSS.n8865 VSS.n8864 0.696929
R60185 VSS.n12073 VSS.n12072 0.696929
R60186 VSS.n12072 VSS.n12071 0.696929
R60187 VSS.n12081 VSS.n12080 0.696929
R60188 VSS.n12080 VSS.n12079 0.696929
R60189 VSS.n12127 VSS.n12126 0.696929
R60190 VSS.n12126 VSS.n12125 0.696929
R60191 VSS.n12135 VSS.n12134 0.696929
R60192 VSS.n12134 VSS.n12133 0.696929
R60193 VSS.n12151 VSS.n12150 0.696929
R60194 VSS.n12150 VSS.n12149 0.696929
R60195 VSS.n12189 VSS.n12188 0.696929
R60196 VSS.n12188 VSS.n12187 0.696929
R60197 VSS.n12197 VSS.n12196 0.696929
R60198 VSS.n12196 VSS.n12195 0.696929
R60199 VSS.n12415 VSS.n12414 0.696929
R60200 VSS.n12414 VSS.n12413 0.696929
R60201 VSS.n12431 VSS.n12430 0.696929
R60202 VSS.n12430 VSS.n12429 0.696929
R60203 VSS.n12439 VSS.n12438 0.696929
R60204 VSS.n12438 VSS.n12437 0.696929
R60205 VSS.n12477 VSS.n12476 0.696929
R60206 VSS.n12476 VSS.n12475 0.696929
R60207 VSS.n12345 VSS.n12344 0.696929
R60208 VSS.n12344 VSS.n12343 0.696929
R60209 VSS.n12337 VSS.n12336 0.696929
R60210 VSS.n12336 VSS.n12335 0.696929
R60211 VSS.n12043 VSS.n12042 0.696929
R60212 VSS.n12042 VSS.n12041 0.696929
R60213 VSS.n12359 VSS.n12358 0.696929
R60214 VSS.n12358 VSS.n12357 0.696929
R60215 VSS.n12367 VSS.n12366 0.696929
R60216 VSS.n12366 VSS.n12365 0.696929
R60217 VSS.n12375 VSS.n12374 0.696929
R60218 VSS.n12374 VSS.n12373 0.696929
R60219 VSS.n12493 VSS.n12492 0.696929
R60220 VSS.n12492 VSS.n12491 0.696929
R60221 VSS.n12485 VSS.n12484 0.696929
R60222 VSS.n12484 VSS.n12483 0.696929
R60223 VSS.n12463 VSS.n12462 0.696929
R60224 VSS.n12462 VSS.n12461 0.696929
R60225 VSS.n12455 VSS.n12454 0.696929
R60226 VSS.n12454 VSS.n12453 0.696929
R60227 VSS.n12447 VSS.n12446 0.696929
R60228 VSS.n12446 VSS.n12445 0.696929
R60229 VSS.n12423 VSS.n12422 0.696929
R60230 VSS.n12422 VSS.n12421 0.696929
R60231 VSS.n12401 VSS.n12400 0.696929
R60232 VSS.n12400 VSS.n12399 0.696929
R60233 VSS.n12393 VSS.n12392 0.696929
R60234 VSS.n12392 VSS.n12391 0.696929
R60235 VSS.n12214 VSS.n12213 0.696929
R60236 VSS.n12213 VSS.n12212 0.696929
R60237 VSS.n12205 VSS.n12204 0.696929
R60238 VSS.n12204 VSS.n12203 0.696929
R60239 VSS.n12175 VSS.n12174 0.696929
R60240 VSS.n12174 VSS.n12173 0.696929
R60241 VSS.n12167 VSS.n12166 0.696929
R60242 VSS.n12166 VSS.n12165 0.696929
R60243 VSS.n12159 VSS.n12158 0.696929
R60244 VSS.n12158 VSS.n12157 0.696929
R60245 VSS.n12143 VSS.n12142 0.696929
R60246 VSS.n12142 VSS.n12141 0.696929
R60247 VSS.n12113 VSS.n12112 0.696929
R60248 VSS.n12112 VSS.n12111 0.696929
R60249 VSS.n12105 VSS.n12104 0.696929
R60250 VSS.n12104 VSS.n12103 0.696929
R60251 VSS.n12097 VSS.n12096 0.696929
R60252 VSS.n12096 VSS.n12095 0.696929
R60253 VSS.n12089 VSS.n12088 0.696929
R60254 VSS.n12088 VSS.n12087 0.696929
R60255 VSS.n12059 VSS.n12058 0.696929
R60256 VSS.n12058 VSS.n12057 0.696929
R60257 VSS.n12051 VSS.n12050 0.696929
R60258 VSS.n12050 VSS.n12049 0.696929
R60259 VSS.n12665 VSS.n12664 0.696929
R60260 VSS.n12035 VSS.n12034 0.696929
R60261 VSS.n12034 VSS.n12033 0.696929
R60262 VSS.n12027 VSS.n12026 0.696929
R60263 VSS.n12026 VSS.n12025 0.696929
R60264 VSS.n9868 VSS.n9866 0.696929
R60265 VSS.n9866 VSS.n9865 0.696929
R60266 VSS.n10298 VSS.n10297 0.696929
R60267 VSS.n10297 VSS.n10296 0.696929
R60268 VSS.n10448 VSS.n10447 0.696929
R60269 VSS.n10447 VSS.n10446 0.696929
R60270 VSS.n10416 VSS.n10415 0.696929
R60271 VSS.n10415 VSS.n10414 0.696929
R60272 VSS.n10354 VSS.n10353 0.696929
R60273 VSS.n10353 VSS.n10352 0.696929
R60274 VSS.n10332 VSS.n10331 0.696929
R60275 VSS.n10331 VSS.n10330 0.696929
R60276 VSS.n10326 VSS.n10325 0.696929
R60277 VSS.n10325 VSS.n10324 0.696929
R60278 VSS.n10131 VSS.n10130 0.696929
R60279 VSS.n10130 VSS.n10129 0.696929
R60280 VSS.n10069 VSS.n10068 0.696929
R60281 VSS.n10068 VSS.n10067 0.696929
R60282 VSS.n10015 VSS.n10014 0.696929
R60283 VSS.n10014 VSS.n10013 0.696929
R60284 VSS.n12644 VSS.n12643 0.696929
R60285 VSS.n12646 VSS.n12645 0.696929
R60286 VSS.n12661 VSS.n12660 0.696929
R60287 VSS.n12066 VSS.n12065 0.696929
R60288 VSS.n12065 VSS.n12064 0.696929
R60289 VSS.n12120 VSS.n12119 0.696929
R60290 VSS.n12119 VSS.n12118 0.696929
R60291 VSS.n12182 VSS.n12181 0.696929
R60292 VSS.n12181 VSS.n12180 0.696929
R60293 VSS.n12380 VSS.n12379 0.696929
R60294 VSS.n12379 VSS.n12378 0.696929
R60295 VSS.n12386 VSS.n12385 0.696929
R60296 VSS.n12385 VSS.n12384 0.696929
R60297 VSS.n12408 VSS.n12407 0.696929
R60298 VSS.n12407 VSS.n12406 0.696929
R60299 VSS.n12470 VSS.n12469 0.696929
R60300 VSS.n12469 VSS.n12468 0.696929
R60301 VSS.n12502 VSS.n12501 0.696929
R60302 VSS.n12501 VSS.n12500 0.696929
R60303 VSS.n12352 VSS.n12351 0.696929
R60304 VSS.n12351 VSS.n12350 0.696929
R60305 VSS.n12329 VSS.n12328 0.696929
R60306 VSS.n12328 VSS.n12327 0.696929
R60307 VSS.n12571 VSS.n12570 0.696929
R60308 VSS.n12570 VSS.n12569 0.696929
R60309 VSS.n11784 VSS.n11783 0.696929
R60310 VSS.n11783 VSS.n11782 0.696929
R60311 VSS.n11776 VSS.n11775 0.696929
R60312 VSS.n11775 VSS.n11774 0.696929
R60313 VSS.n12600 VSS.n12599 0.696929
R60314 VSS.n12599 VSS.n12598 0.696929
R60315 VSS.n12672 VSS.n12671 0.696929
R60316 VSS.n12671 VSS.n12670 0.696929
R60317 VSS.n12019 VSS.n12018 0.696929
R60318 VSS.n12018 VSS.n12017 0.696929
R60319 VSS.n12644 VSS.n12641 0.686214
R60320 VSS.n9838 VSS.n9835 0.686214
R60321 VSS.n13651 VSS.n13647 0.685697
R60322 VSS.n14266 VSS.n14262 0.685697
R60323 VSS.n4167 DVSS 0.66425
R60324 VSS.n21709 DVSS 0.66425
R60325 VSS.n11409 DVSS 0.66425
R60326 VSS.n20842 DVSS 0.66425
R60327 VSS.n11473 DVSS 0.66425
R60328 VSS.n20750 DVSS 0.66425
R60329 VSS.n11632 DVSS 0.66425
R60330 VSS.n20699 DVSS 0.66425
R60331 VSS.n17234 DVSS 0.66425
R60332 VSS.n13258 DVSS 0.66425
R60333 VSS.n17378 DVSS 0.66425
R60334 VSS.n13377 DVSS 0.66425
R60335 VSS.n17403 DVSS 0.66425
R60336 VSS.n13285 DVSS 0.66425
R60337 VSS.n21227 DVSS 0.66425
R60338 VSS.n11258 DVSS 0.66425
R60339 VSS.n4108 DVSS 0.66425
R60340 VSS.n21904 DVSS 0.66425
R60341 VSS.n15646 VSS.n15645 0.6505
R60342 VSS.n15645 VSS.n15644 0.6505
R60343 VSS.n15618 VSS.n15617 0.6505
R60344 VSS.n15596 VSS.n15595 0.6505
R60345 VSS.n15507 VSS.n15505 0.6505
R60346 VSS.n15436 VSS.n15435 0.6505
R60347 VSS.n15508 VSS.n15507 0.6505
R60348 VSS.n15509 VSS.n15508 0.6505
R60349 VSS.n21934 VSS.n21933 0.647738
R60350 VSS.n15689 VSS.n15686 0.632106
R60351 VSS.n15689 VSS.n15682 0.632106
R60352 VSS.n197 VSS.n191 0.632106
R60353 VSS.n197 VSS.n196 0.632106
R60354 VSS.n15696 VSS.n15692 0.624161
R60355 VSS.n21421 VSS.n21420 0.623413
R60356 VSS.n21311 VSS.n21310 0.623413
R60357 VSS.n17241 VSS.n17240 0.623413
R60358 VSS.n4931 VSS.n4930 0.623413
R60359 VSS.n21661 VSS.n21660 0.617744
R60360 VSS.n4122 VSS.n4121 0.617744
R60361 VSS.n21248 VSS.n21247 0.616858
R60362 VSS.n11249 VSS.n11248 0.616858
R60363 VSS.n17338 VSS.n17337 0.612075
R60364 VSS.n11514 VSS.n11513 0.612075
R60365 VSS.n13253 VSS.n13252 0.612075
R60366 VSS.n12892 VSS.n12891 0.612075
R60367 VSS.n14430 VSS.n14429 0.612075
R60368 VSS.n15100 VSS.n15099 0.612075
R60369 VSS.n13408 VSS.n13407 0.612075
R60370 VSS.n20730 VSS.n20729 0.612075
R60371 VSS.n13513 VSS.n13512 0.612075
R60372 VSS.n2059 VSS.n2058 0.612075
R60373 VSS.n587 VSS.n586 0.612075
R60374 VSS.n3956 VSS.n3955 0.61172
R60375 VSS.n13124 VSS.n13123 0.61172
R60376 VSS.n18969 VSS.n18968 0.61172
R60377 VSS.n21754 VSS.n21753 0.61172
R60378 VSS.n19039 VSS.n19038 0.61172
R60379 VSS.n11311 VSS.n11310 0.611189
R60380 VSS.n12825 VSS.n12824 0.611189
R60381 VSS.n16386 VSS.n16385 0.611189
R60382 VSS.n20873 VSS.n20872 0.611189
R60383 VSS.n889 VSS.n888 0.611189
R60384 VSS.n524 VSS.n523 0.611189
R60385 VSS.n21432 VSS.n21431 0.606228
R60386 VSS.n17388 VSS.n17387 0.606228
R60387 VSS.n15689 VSS.n15685 0.604265
R60388 VSS.n15689 VSS.n15681 0.604265
R60389 VSS.n17293 VSS.n17281 0.604265
R60390 VSS.n17178 VSS.n14333 0.604265
R60391 VSS.n2411 VSS.n2399 0.604265
R60392 VSS.n197 VSS.n193 0.604265
R60393 VSS.n197 VSS.n192 0.604265
R60394 VSS.n2497 VSS.n2469 0.604265
R60395 VSS.n13240 VSS.n13239 0.600559
R60396 VSS.n13357 VSS.n13356 0.600559
R60397 VSS.n13500 VSS.n13499 0.600559
R60398 VSS.n17293 VSS.n17270 0.594741
R60399 VSS.n17178 VSS.n11768 0.594741
R60400 VSS.n4841 VSS.n4830 0.594741
R60401 VSS.n4841 VSS.n4818 0.594741
R60402 VSS.n4905 VSS.n4892 0.594741
R60403 VSS.n4905 VSS.n4880 0.594741
R60404 VSS.n5460 VSS.n5447 0.594741
R60405 VSS.n5460 VSS.n5435 0.594741
R60406 VSS.n2411 VSS.n2401 0.594741
R60407 VSS.n2497 VSS.n2484 0.594741
R60408 VSS.n3923 VSS.n3913 0.594741
R60409 VSS.n3923 VSS.n3908 0.594741
R60410 VSS.n17293 VSS.n17266 0.586651
R60411 VSS.n17178 VSS.n11756 0.586651
R60412 VSS.n4841 VSS.n4829 0.586651
R60413 VSS.n4841 VSS.n4814 0.586651
R60414 VSS.n4905 VSS.n4891 0.586651
R60415 VSS.n4905 VSS.n4876 0.586651
R60416 VSS.n5460 VSS.n5446 0.586651
R60417 VSS.n5460 VSS.n5431 0.586651
R60418 VSS.n2411 VSS.n2400 0.586651
R60419 VSS.n3923 VSS.n3912 0.586651
R60420 VSS.n3923 VSS.n3916 0.586651
R60421 VSS.n2497 VSS.n2495 0.586651
R60422 VSS.n200 VSS.n199 0.576595
R60423 VSS.n15680 VSS.n15679 0.576595
R60424 VSS.n8496 VSS.n8495 0.5205
R60425 VSS.n8495 VSS.n8494 0.5205
R60426 VSS.n9198 VSS.n9197 0.5205
R60427 VSS.n9197 VSS.n9196 0.5205
R60428 VSS.n10449 VSS.n10448 0.5005
R60429 VSS.n10164 VSS.n10163 0.5005
R60430 VSS.n12503 VSS.n12502 0.5005
R60431 VSS.n12215 VSS.n12214 0.5005
R60432 VSS.n17293 VSS.n17282 0.466929
R60433 VSS.n17178 VSS.n14339 0.466929
R60434 VSS.n2411 VSS.n2398 0.466929
R60435 VSS.n2497 VSS.n2470 0.466929
R60436 VSS.n1422 VSS.n1418 0.403878
R60437 VSS.n16333 VSS.n16330 0.403878
R60438 VSS.n16262 VSS.n16260 0.403878
R60439 VSS.n1346 VSS.n1344 0.403878
R60440 VSS.n15566 VSS.n15565 0.394514
R60441 VSS.n1854 VSS.n1853 0.394514
R60442 VSS.n1493 VSS.n1492 0.376311
R60443 VSS.n1563 VSS.n1561 0.376311
R60444 VSS.n1580 VSS.n1579 0.376311
R60445 VSS.n15216 VSS.n15212 0.375905
R60446 VSS.n15582 VSS.n15576 0.375905
R60447 VSS.n15561 VSS.n15559 0.375905
R60448 VSS.n5486 VSS.n5485 0.373473
R60449 VSS.n1307 VSS.n1306 0.373473
R60450 VSS.n858 DVSS 0.37265
R60451 VSS.n11301 DVSS 0.37265
R60452 VSS.n16035 VSS.n16034 0.371446
R60453 VSS.n1042 VSS.n1041 0.371041
R60454 VSS.n5530 VSS.n5529 0.368608
R60455 VSS.n1014 VSS.n1013 0.368608
R60456 VSS.n4025 VSS.n4024 0.345264
R60457 VSS.n13052 VSS.n13051 0.345264
R60458 VSS.n18896 VSS.n18895 0.345264
R60459 VSS.n21825 VSS.n21824 0.345264
R60460 VSS.n19110 VSS.n19109 0.345264
R60461 VSS.n21596 VSS.n21595 0.345264
R60462 VSS.n3827 VSS.n3826 0.345264
R60463 VSS.n2363 VSS.n2362 0.344378
R60464 VSS.n13173 VSS.n13172 0.344378
R60465 VSS.n2262 VSS.n2261 0.344378
R60466 VSS.n2313 VSS.n2312 0.344378
R60467 VSS.n17921 VSS.n17920 0.344378
R60468 VSS.n21500 VSS.n21499 0.344378
R60469 VSS.n4716 VSS.n4715 0.344378
R60470 VSS.n12775 VSS.n12774 0.340835
R60471 VSS.n7587 VSS.n7586 0.340835
R60472 VSS.n11198 VSS.n11197 0.340835
R60473 VSS.n478 VSS.n477 0.340835
R60474 VSS.n4194 DVSS 0.332375
R60475 VSS.n17878 DVSS 0.332375
R60476 VSS.n11372 DVSS 0.332375
R60477 VSS.n1988 DVSS 0.332375
R60478 VSS.n11504 DVSS 0.332375
R60479 VSS.n2063 DVSS 0.332375
R60480 VSS.n11595 DVSS 0.332375
R60481 VSS.n20061 DVSS 0.332375
R60482 VSS.n14357 DVSS 0.332375
R60483 VSS.n13430 DVSS 0.332375
R60484 VSS.n17351 DVSS 0.332375
R60485 VSS.n13453 DVSS 0.332375
R60486 VSS.n17427 DVSS 0.332375
R60487 VSS.n17960 DVSS 0.332375
R60488 VSS.n3943 DVSS 0.332375
R60489 VSS.n2152 DVSS 0.332375
R60490 VSS.n16237 VSS.n16236 0.330913
R60491 VSS.n1318 VSS.n1317 0.330913
R60492 VSS.n15689 VSS.n15687 0.28898
R60493 VSS.n15689 VSS.n15683 0.28898
R60494 VSS.n197 VSS.n194 0.28898
R60495 VSS.n197 VSS.n189 0.28898
R60496 VSS.n15689 VSS.n15684 0.287336
R60497 VSS.n197 VSS.n190 0.287336
R60498 VSS.n197 VSS.n195 0.287336
R60499 VSS.n15689 VSS.n15688 0.287064
R60500 VSS.n21259 VSS.n21258 0.285913
R60501 VSS.n11419 VSS.n11418 0.285913
R60502 VSS.n904 VSS.n902 0.284689
R60503 VSS.n15918 VSS.n15916 0.284284
R60504 VSS.n17293 VSS.n17286 0.280941
R60505 VSS.n17293 VSS.n17274 0.280941
R60506 VSS.n17178 VSS.n14354 0.280941
R60507 VSS.n17178 VSS.n13427 0.280941
R60508 VSS.n4841 VSS.n4834 0.280941
R60509 VSS.n4841 VSS.n4822 0.280941
R60510 VSS.n4905 VSS.n4896 0.280941
R60511 VSS.n4905 VSS.n4884 0.280941
R60512 VSS.n5460 VSS.n5451 0.280941
R60513 VSS.n5460 VSS.n5439 0.280941
R60514 VSS.n2411 VSS.n2402 0.280941
R60515 VSS.n2497 VSS.n2488 0.280941
R60516 VSS.n3923 VSS.n3910 0.280941
R60517 VSS.n3923 VSS.n3906 0.280941
R60518 VSS.n2497 VSS.n2474 0.280941
R60519 VSS.n2411 VSS.n2408 0.280941
R60520 VSS.n11369 VSS.n11368 0.280244
R60521 VSS.n12838 VSS.n12837 0.280244
R60522 VSS.n15170 VSS.n15169 0.280244
R60523 VSS.n20822 VSS.n20821 0.280244
R60524 VSS.n1997 VSS.n1996 0.280244
R60525 VSS.n537 VSS.n536 0.280244
R60526 VSS.n17293 VSS.n17278 0.278361
R60527 VSS.n17178 VSS.n13531 0.278361
R60528 VSS.n4841 VSS.n4826 0.278361
R60529 VSS.n4905 VSS.n4888 0.278361
R60530 VSS.n5460 VSS.n5443 0.278361
R60531 VSS.n2411 VSS.n2403 0.278361
R60532 VSS.n2411 VSS.n2404 0.278361
R60533 VSS.n3923 VSS.n3904 0.278361
R60534 VSS.n3923 VSS.n3902 0.278361
R60535 VSS.n2497 VSS.n2478 0.278361
R60536 VSS.n17293 VSS.n17290 0.278105
R60537 VSS.n17178 VSS.n14370 0.278105
R60538 VSS.n4841 VSS.n4838 0.278105
R60539 VSS.n4905 VSS.n4900 0.278105
R60540 VSS.n5460 VSS.n5455 0.278105
R60541 VSS.n2497 VSS.n2492 0.278105
R60542 VSS.n15669 VSS.n15668 0.268599
R60543 VSS.n1927 VSS.n1926 0.268599
R60544 VSS.n5664 VSS.n5662 0.266041
R60545 VSS.n5757 VSS.n5754 0.266041
R60546 VSS.n20933 VSS.n20931 0.265635
R60547 VSS.n3186 VSS.n3185 0.257472
R60548 VSS.n3211 VSS.n3210 0.2505
R60549 VSS.n3677 VSS.n3676 0.2505
R60550 VSS.n3676 VSS.n3675 0.2505
R60551 VSS.n3652 VSS.n3651 0.2505
R60552 VSS.n3650 VSS.n3649 0.2505
R60553 VSS.n3648 VSS.n3647 0.2505
R60554 VSS.n3646 VSS.n3645 0.2505
R60555 VSS.n3639 VSS.n3638 0.2505
R60556 VSS.n3629 VSS.n3628 0.2505
R60557 VSS.n3620 VSS.n3619 0.2505
R60558 VSS.n3612 VSS.n3611 0.2505
R60559 VSS.n3609 VSS.n3608 0.2505
R60560 VSS.n3607 VSS.n3606 0.2505
R60561 VSS.n3604 VSS.n3603 0.2505
R60562 VSS.n3596 VSS.n3595 0.2505
R60563 VSS.n3586 VSS.n3585 0.2505
R60564 VSS.n3577 VSS.n3576 0.2505
R60565 VSS.n3569 VSS.n3568 0.2505
R60566 VSS.n3566 VSS.n3565 0.2505
R60567 VSS.n3564 VSS.n3563 0.2505
R60568 VSS.n3562 VSS.n3561 0.2505
R60569 VSS.n3560 VSS.n3559 0.2505
R60570 VSS.n3558 VSS.n3557 0.2505
R60571 VSS.n3556 VSS.n3555 0.2505
R60572 VSS.n3554 VSS.n3553 0.2505
R60573 VSS.n3552 VSS.n3551 0.2505
R60574 VSS.n3550 VSS.n3549 0.2505
R60575 VSS.n3547 VSS.n3546 0.2505
R60576 VSS.n3544 VSS.n3543 0.2505
R60577 VSS.n3537 VSS.n3536 0.2505
R60578 VSS.n3527 VSS.n3526 0.2505
R60579 VSS.n3518 VSS.n3517 0.2505
R60580 VSS.n3509 VSS.n3508 0.2505
R60581 VSS.n3502 VSS.n3501 0.2505
R60582 VSS.n3497 VSS.n3496 0.2505
R60583 VSS.n3495 VSS.n3494 0.2505
R60584 VSS.n3493 VSS.n3492 0.2505
R60585 VSS.n3490 VSS.n3489 0.2505
R60586 VSS.n3487 VSS.n3486 0.2505
R60587 VSS.n3485 VSS.n3484 0.2505
R60588 VSS.n3478 VSS.n3477 0.2505
R60589 VSS.n3471 VSS.n3470 0.2505
R60590 VSS.n3457 VSS.n3456 0.2505
R60591 VSS.n3452 VSS.n3451 0.2505
R60592 VSS.n3439 VSS.n3438 0.2505
R60593 VSS.n3430 VSS.n3429 0.2505
R60594 VSS.n3421 VSS.n3420 0.2505
R60595 VSS.n3418 VSS.n3417 0.2505
R60596 VSS.n3414 VSS.n3413 0.2505
R60597 VSS.n3411 VSS.n3410 0.2505
R60598 VSS.n3406 VSS.n3405 0.2505
R60599 VSS.n3401 VSS.n3400 0.2505
R60600 VSS.n3399 VSS.n3398 0.2505
R60601 VSS.n3397 VSS.n3396 0.2505
R60602 VSS.n3392 VSS.n3391 0.2505
R60603 VSS.n3386 VSS.n3385 0.2505
R60604 VSS.n3377 VSS.n3376 0.2505
R60605 VSS.n3367 VSS.n3366 0.2505
R60606 VSS.n3363 VSS.n3362 0.2505
R60607 VSS.n3361 VSS.n3360 0.2505
R60608 VSS.n3359 VSS.n3358 0.2505
R60609 VSS.n3357 VSS.n3356 0.2505
R60610 VSS.n3355 VSS.n3354 0.2505
R60611 VSS.n3353 VSS.n3352 0.2505
R60612 VSS.n3351 VSS.n3350 0.2505
R60613 VSS.n3349 VSS.n3348 0.2505
R60614 VSS.n3347 VSS.n3346 0.2505
R60615 VSS.n3345 VSS.n3344 0.2505
R60616 VSS.n3343 VSS.n3342 0.2505
R60617 VSS.n3338 VSS.n3337 0.2505
R60618 VSS.n3332 VSS.n3331 0.2505
R60619 VSS.n3323 VSS.n3322 0.2505
R60620 VSS.n3314 VSS.n3313 0.2505
R60621 VSS.n3311 VSS.n3310 0.2505
R60622 VSS.n3309 VSS.n3308 0.2505
R60623 VSS.n3307 VSS.n3306 0.2505
R60624 VSS.n3305 VSS.n3304 0.2505
R60625 VSS.n3300 VSS.n3299 0.2505
R60626 VSS.n3294 VSS.n3293 0.2505
R60627 VSS.n3192 VSS.n3190 0.2505
R60628 VSS.n3193 VSS.n3192 0.2505
R60629 VSS.n3775 VSS.n3774 0.2505
R60630 VSS.n3776 VSS.n3775 0.2505
R60631 VSS.n3217 VSS.n3216 0.2505
R60632 VSS.n3222 VSS.n3221 0.2505
R60633 VSS.n3224 VSS.n3223 0.2505
R60634 VSS.n3226 VSS.n3225 0.2505
R60635 VSS.n3228 VSS.n3227 0.2505
R60636 VSS.n3231 VSS.n3230 0.2505
R60637 VSS.n3240 VSS.n3239 0.2505
R60638 VSS.n1474 VSS.n1471 0.233545
R60639 VSS.n15907 VSS.n15905 0.233293
R60640 VSS.n2523 VSS.n2522 0.231864
R60641 VSS.n4933 VSS.n4932 0.231864
R60642 VSS.n5905 VSS.n5904 0.231864
R60643 VSS.n2432 VSS.n2431 0.231864
R60644 VSS.n4733 VSS.n4732 0.231864
R60645 VSS.n225 VSS.n223 0.231534
R60646 VSS.n59 VSS.n57 0.231282
R60647 VSS.n22008 VSS.n21989 0.23125
R60648 VSS.n60 VSS.n59 0.230528
R60649 VSS.n13664 VSS.n13661 0.230514
R60650 VSS.n226 VSS.n225 0.230277
R60651 VSS.n92 VSS.n91 0.228768
R60652 VSS.n91 VSS.n89 0.228768
R60653 VSS.n257 VSS.n255 0.228768
R60654 VSS.n258 VSS.n257 0.228768
R60655 VSS.n13676 VSS.n13675 0.2255
R60656 VSS.n13679 VSS.n13678 0.2255
R60657 VSS.n13681 VSS.n13680 0.2255
R60658 VSS.n13683 VSS.n13682 0.2255
R60659 VSS.n13685 VSS.n13684 0.2255
R60660 VSS.n13687 VSS.n13686 0.2255
R60661 VSS.n13689 VSS.n13688 0.2255
R60662 VSS.n13691 VSS.n13690 0.2255
R60663 VSS.n13693 VSS.n13692 0.2255
R60664 VSS.n13695 VSS.n13694 0.2255
R60665 VSS.n13697 VSS.n13696 0.2255
R60666 VSS.n13699 VSS.n13698 0.2255
R60667 VSS.n13701 VSS.n13700 0.2255
R60668 VSS.n13703 VSS.n13702 0.2255
R60669 VSS.n13705 VSS.n13704 0.2255
R60670 VSS.n13707 VSS.n13706 0.2255
R60671 VSS.n13709 VSS.n13708 0.2255
R60672 VSS.n13711 VSS.n13710 0.2255
R60673 VSS.n13713 VSS.n13712 0.2255
R60674 VSS.n13715 VSS.n13714 0.2255
R60675 VSS.n13717 VSS.n13716 0.2255
R60676 VSS.n13719 VSS.n13718 0.2255
R60677 VSS.n13721 VSS.n13720 0.2255
R60678 VSS.n13723 VSS.n13722 0.2255
R60679 VSS.n13725 VSS.n13724 0.2255
R60680 VSS.n13727 VSS.n13726 0.2255
R60681 VSS.n13729 VSS.n13728 0.2255
R60682 VSS.n13731 VSS.n13730 0.2255
R60683 VSS.n13733 VSS.n13732 0.2255
R60684 VSS.n13735 VSS.n13734 0.2255
R60685 VSS.n13737 VSS.n13736 0.2255
R60686 VSS.n13739 VSS.n13738 0.2255
R60687 VSS.n13741 VSS.n13740 0.2255
R60688 VSS.n13743 VSS.n13742 0.2255
R60689 VSS.n13746 VSS.n13745 0.2255
R60690 VSS.n13749 VSS.n13748 0.2255
R60691 VSS.n13752 VSS.n13751 0.2255
R60692 VSS.n13755 VSS.n13754 0.2255
R60693 VSS.n13757 VSS.n13756 0.2255
R60694 VSS.n13759 VSS.n13758 0.2255
R60695 VSS.n13761 VSS.n13760 0.2255
R60696 VSS.n13763 VSS.n13762 0.2255
R60697 VSS.n13765 VSS.n13764 0.2255
R60698 VSS.n13767 VSS.n13766 0.2255
R60699 VSS.n13770 VSS.n13769 0.2255
R60700 VSS.n13773 VSS.n13772 0.2255
R60701 VSS.n13775 VSS.n13774 0.2255
R60702 VSS.n13777 VSS.n13776 0.2255
R60703 VSS.n13779 VSS.n13778 0.2255
R60704 VSS.n13781 VSS.n13780 0.2255
R60705 VSS.n13783 VSS.n13782 0.2255
R60706 VSS.n13785 VSS.n13784 0.2255
R60707 VSS.n13787 VSS.n13786 0.2255
R60708 VSS.n13789 VSS.n13788 0.2255
R60709 VSS.n13791 VSS.n13790 0.2255
R60710 VSS.n13794 VSS.n13793 0.2255
R60711 VSS.n13797 VSS.n13796 0.2255
R60712 VSS.n13799 VSS.n13798 0.2255
R60713 VSS.n13801 VSS.n13800 0.2255
R60714 VSS.n13803 VSS.n13802 0.2255
R60715 VSS.n13805 VSS.n13804 0.2255
R60716 VSS.n13807 VSS.n13806 0.2255
R60717 VSS.n13809 VSS.n13808 0.2255
R60718 VSS.n13811 VSS.n13810 0.2255
R60719 VSS.n13813 VSS.n13812 0.2255
R60720 VSS.n13815 VSS.n13814 0.2255
R60721 VSS.n13817 VSS.n13816 0.2255
R60722 VSS.n13819 VSS.n13818 0.2255
R60723 VSS.n13821 VSS.n13820 0.2255
R60724 VSS.n13823 VSS.n13822 0.2255
R60725 VSS.n13825 VSS.n13824 0.2255
R60726 VSS.n13827 VSS.n13826 0.2255
R60727 VSS.n13829 VSS.n13828 0.2255
R60728 VSS.n13831 VSS.n13830 0.2255
R60729 VSS.n13833 VSS.n13832 0.2255
R60730 VSS.n13836 VSS.n13835 0.2255
R60731 VSS.n13840 VSS.n13839 0.2255
R60732 VSS.n13845 VSS.n13844 0.2255
R60733 VSS.n13849 VSS.n13848 0.2255
R60734 VSS.n13852 VSS.n13851 0.2255
R60735 VSS.n13851 VSS.n13850 0.2255
R60736 VSS.n13670 VSS.n13669 0.2255
R60737 VSS.n13668 VSS.n13667 0.2255
R60738 VSS.n13666 VSS.n13665 0.2255
R60739 VSS.n14239 VSS.n14238 0.2255
R60740 VSS.n14230 VSS.n14229 0.2255
R60741 VSS.n14228 VSS.n14227 0.2255
R60742 VSS.n14226 VSS.n14225 0.2255
R60743 VSS.n14224 VSS.n14223 0.2255
R60744 VSS.n14222 VSS.n14221 0.2255
R60745 VSS.n14220 VSS.n14219 0.2255
R60746 VSS.n14218 VSS.n14217 0.2255
R60747 VSS.n14216 VSS.n14215 0.2255
R60748 VSS.n14213 VSS.n14212 0.2255
R60749 VSS.n14214 VSS.n14213 0.2255
R60750 VSS.n13941 VSS.n13940 0.2255
R60751 VSS.n13942 VSS.n13941 0.2255
R60752 VSS.n2553 VSS.n2552 0.2255
R60753 VSS.n2575 VSS.n2574 0.2255
R60754 VSS.n2574 VSS.n2573 0.2255
R60755 VSS.n2876 VSS.n2875 0.2255
R60756 VSS.n2888 VSS.n2887 0.2255
R60757 VSS.n2898 VSS.n2897 0.2255
R60758 VSS.n2903 VSS.n2902 0.2255
R60759 VSS.n2906 VSS.n2905 0.2255
R60760 VSS.n2909 VSS.n2908 0.2255
R60761 VSS.n2911 VSS.n2910 0.2255
R60762 VSS.n2913 VSS.n2912 0.2255
R60763 VSS.n2915 VSS.n2914 0.2255
R60764 VSS.n2917 VSS.n2916 0.2255
R60765 VSS.n2920 VSS.n2919 0.2255
R60766 VSS.n2930 VSS.n2929 0.2255
R60767 VSS.n2940 VSS.n2939 0.2255
R60768 VSS.n2951 VSS.n2950 0.2255
R60769 VSS.n2959 VSS.n2958 0.2255
R60770 VSS.n2961 VSS.n2960 0.2255
R60771 VSS.n2963 VSS.n2962 0.2255
R60772 VSS.n2965 VSS.n2964 0.2255
R60773 VSS.n2967 VSS.n2966 0.2255
R60774 VSS.n2969 VSS.n2968 0.2255
R60775 VSS.n2971 VSS.n2970 0.2255
R60776 VSS.n2973 VSS.n2972 0.2255
R60777 VSS.n2976 VSS.n2975 0.2255
R60778 VSS.n2979 VSS.n2978 0.2255
R60779 VSS.n2981 VSS.n2980 0.2255
R60780 VSS.n2984 VSS.n2983 0.2255
R60781 VSS.n2994 VSS.n2993 0.2255
R60782 VSS.n3005 VSS.n3004 0.2255
R60783 VSS.n3015 VSS.n3014 0.2255
R60784 VSS.n3023 VSS.n3022 0.2255
R60785 VSS.n3025 VSS.n3024 0.2255
R60786 VSS.n3027 VSS.n3026 0.2255
R60787 VSS.n3029 VSS.n3028 0.2255
R60788 VSS.n3032 VSS.n3031 0.2255
R60789 VSS.n3042 VSS.n3041 0.2255
R60790 VSS.n3053 VSS.n3052 0.2255
R60791 VSS.n3063 VSS.n3062 0.2255
R60792 VSS.n3072 VSS.n3071 0.2255
R60793 VSS.n3075 VSS.n3074 0.2255
R60794 VSS.n3077 VSS.n3076 0.2255
R60795 VSS.n3084 VSS.n3083 0.2255
R60796 VSS.n3083 VSS.n3082 0.2255
R60797 VSS.n2864 VSS.n2863 0.2255
R60798 VSS.n2802 VSS.n2801 0.2255
R60799 VSS.n2806 VSS.n2805 0.2255
R60800 VSS.n2808 VSS.n2807 0.2255
R60801 VSS.n2810 VSS.n2809 0.2255
R60802 VSS.n2812 VSS.n2811 0.2255
R60803 VSS.n2814 VSS.n2813 0.2255
R60804 VSS.n2816 VSS.n2815 0.2255
R60805 VSS.n2818 VSS.n2817 0.2255
R60806 VSS.n2820 VSS.n2819 0.2255
R60807 VSS.n2822 VSS.n2821 0.2255
R60808 VSS.n2824 VSS.n2823 0.2255
R60809 VSS.n2833 VSS.n2832 0.2255
R60810 VSS.n2845 VSS.n2844 0.2255
R60811 VSS.n2859 VSS.n2858 0.2255
R60812 VSS.n2699 VSS.n2698 0.2255
R60813 VSS.n2704 VSS.n2703 0.2255
R60814 VSS.n2715 VSS.n2714 0.2255
R60815 VSS.n2726 VSS.n2725 0.2255
R60816 VSS.n2752 VSS.n2751 0.2255
R60817 VSS.n2775 VSS.n2774 0.2255
R60818 VSS.n2786 VSS.n2785 0.2255
R60819 VSS.n2529 VSS.n2528 0.2255
R60820 VSS.n2540 VSS.n2539 0.2255
R60821 VSS.n2541 VSS.n2540 0.2255
R60822 VSS.n3181 VSS.n3180 0.2255
R60823 VSS.n3182 VSS.n3181 0.2255
R60824 VSS.n2579 VSS.n2578 0.2255
R60825 VSS.n2581 VSS.n2580 0.2255
R60826 VSS.n2584 VSS.n2583 0.2255
R60827 VSS.n2587 VSS.n2586 0.2255
R60828 VSS.n2671 VSS.n2670 0.2255
R60829 VSS.n2681 VSS.n2680 0.2255
R60830 VSS.n2689 VSS.n2688 0.2255
R60831 VSS.n4964 VSS.n4954 0.2255
R60832 VSS.n4964 VSS.n4963 0.2255
R60833 VSS.n4973 VSS.n4972 0.2255
R60834 VSS.n4972 VSS.n4971 0.2255
R60835 VSS.n5312 VSS.n5311 0.2255
R60836 VSS.n5311 VSS.n5310 0.2255
R60837 VSS.n5307 VSS.n5306 0.2255
R60838 VSS.n5305 VSS.n5304 0.2255
R60839 VSS.n5303 VSS.n5302 0.2255
R60840 VSS.n5301 VSS.n5300 0.2255
R60841 VSS.n5296 VSS.n5295 0.2255
R60842 VSS.n5288 VSS.n5287 0.2255
R60843 VSS.n5281 VSS.n5280 0.2255
R60844 VSS.n5275 VSS.n5274 0.2255
R60845 VSS.n5272 VSS.n5271 0.2255
R60846 VSS.n5270 VSS.n5269 0.2255
R60847 VSS.n5268 VSS.n5267 0.2255
R60848 VSS.n5266 VSS.n5265 0.2255
R60849 VSS.n5261 VSS.n5260 0.2255
R60850 VSS.n5253 VSS.n5252 0.2255
R60851 VSS.n5247 VSS.n5246 0.2255
R60852 VSS.n5240 VSS.n5239 0.2255
R60853 VSS.n5237 VSS.n5236 0.2255
R60854 VSS.n5235 VSS.n5234 0.2255
R60855 VSS.n5233 VSS.n5232 0.2255
R60856 VSS.n5231 VSS.n5230 0.2255
R60857 VSS.n5229 VSS.n5228 0.2255
R60858 VSS.n5227 VSS.n5226 0.2255
R60859 VSS.n5225 VSS.n5224 0.2255
R60860 VSS.n5223 VSS.n5222 0.2255
R60861 VSS.n5221 VSS.n5220 0.2255
R60862 VSS.n5219 VSS.n5218 0.2255
R60863 VSS.n5217 VSS.n5216 0.2255
R60864 VSS.n5215 VSS.n5214 0.2255
R60865 VSS.n5210 VSS.n5209 0.2255
R60866 VSS.n5202 VSS.n5201 0.2255
R60867 VSS.n5196 VSS.n5195 0.2255
R60868 VSS.n5189 VSS.n5188 0.2255
R60869 VSS.n5186 VSS.n5185 0.2255
R60870 VSS.n5184 VSS.n5183 0.2255
R60871 VSS.n5182 VSS.n5181 0.2255
R60872 VSS.n5180 VSS.n5179 0.2255
R60873 VSS.n5178 VSS.n5177 0.2255
R60874 VSS.n5176 VSS.n5175 0.2255
R60875 VSS.n5174 VSS.n5173 0.2255
R60876 VSS.n5172 VSS.n5171 0.2255
R60877 VSS.n5170 VSS.n5169 0.2255
R60878 VSS.n5168 VSS.n5167 0.2255
R60879 VSS.n5166 VSS.n5165 0.2255
R60880 VSS.n5164 VSS.n5163 0.2255
R60881 VSS.n5159 VSS.n5158 0.2255
R60882 VSS.n5152 VSS.n5151 0.2255
R60883 VSS.n5140 VSS.n5139 0.2255
R60884 VSS.n4939 VSS.n4937 0.2255
R60885 VSS.n4940 VSS.n4939 0.2255
R60886 VSS.n5410 VSS.n5409 0.2255
R60887 VSS.n5411 VSS.n5410 0.2255
R60888 VSS.n4981 VSS.n4980 0.2255
R60889 VSS.n4986 VSS.n4985 0.2255
R60890 VSS.n4994 VSS.n4993 0.2255
R60891 VSS.n5001 VSS.n5000 0.2255
R60892 VSS.n5005 VSS.n5004 0.2255
R60893 VSS.n5008 VSS.n5007 0.2255
R60894 VSS.n5010 VSS.n5009 0.2255
R60895 VSS.n5012 VSS.n5011 0.2255
R60896 VSS.n5014 VSS.n5013 0.2255
R60897 VSS.n5016 VSS.n5015 0.2255
R60898 VSS.n5024 VSS.n5023 0.2255
R60899 VSS.n5031 VSS.n5030 0.2255
R60900 VSS.n5035 VSS.n5034 0.2255
R60901 VSS.n5038 VSS.n5037 0.2255
R60902 VSS.n5040 VSS.n5039 0.2255
R60903 VSS.n5042 VSS.n5041 0.2255
R60904 VSS.n5045 VSS.n5044 0.2255
R60905 VSS.n5048 VSS.n5047 0.2255
R60906 VSS.n5050 VSS.n5049 0.2255
R60907 VSS.n5053 VSS.n5052 0.2255
R60908 VSS.n5056 VSS.n5055 0.2255
R60909 VSS.n5060 VSS.n5059 0.2255
R60910 VSS.n5070 VSS.n5069 0.2255
R60911 VSS.n5077 VSS.n5076 0.2255
R60912 VSS.n5081 VSS.n5080 0.2255
R60913 VSS.n5084 VSS.n5083 0.2255
R60914 VSS.n5086 VSS.n5085 0.2255
R60915 VSS.n5088 VSS.n5087 0.2255
R60916 VSS.n5090 VSS.n5089 0.2255
R60917 VSS.n5093 VSS.n5092 0.2255
R60918 VSS.n5096 VSS.n5095 0.2255
R60919 VSS.n5098 VSS.n5097 0.2255
R60920 VSS.n5100 VSS.n5099 0.2255
R60921 VSS.n5102 VSS.n5101 0.2255
R60922 VSS.n5104 VSS.n5103 0.2255
R60923 VSS.n5106 VSS.n5105 0.2255
R60924 VSS.n5109 VSS.n5108 0.2255
R60925 VSS.n5115 VSS.n5114 0.2255
R60926 VSS.n5124 VSS.n5123 0.2255
R60927 VSS.n5135 VSS.n5134 0.2255
R60928 VSS.n5920 VSS.n5918 0.2255
R60929 VSS.n7529 VSS.n7528 0.2255
R60930 VSS.n7538 VSS.n7537 0.2255
R60931 VSS.n7539 VSS.n7538 0.2255
R60932 VSS.n5921 VSS.n5920 0.2255
R60933 VSS.n7421 VSS.n7420 0.2255
R60934 VSS.n7420 VSS.n7419 0.2255
R60935 VSS.n7417 VSS.n7416 0.2255
R60936 VSS.n7415 VSS.n7414 0.2255
R60937 VSS.n7413 VSS.n7412 0.2255
R60938 VSS.n7411 VSS.n7410 0.2255
R60939 VSS.n7404 VSS.n7403 0.2255
R60940 VSS.n7395 VSS.n7394 0.2255
R60941 VSS.n7390 VSS.n7389 0.2255
R60942 VSS.n7387 VSS.n7386 0.2255
R60943 VSS.n7385 VSS.n7384 0.2255
R60944 VSS.n7383 VSS.n7382 0.2255
R60945 VSS.n7381 VSS.n7380 0.2255
R60946 VSS.n7379 VSS.n7378 0.2255
R60947 VSS.n7372 VSS.n7371 0.2255
R60948 VSS.n7361 VSS.n7360 0.2255
R60949 VSS.n7354 VSS.n7353 0.2255
R60950 VSS.n7349 VSS.n7348 0.2255
R60951 VSS.n7345 VSS.n7344 0.2255
R60952 VSS.n7343 VSS.n7342 0.2255
R60953 VSS.n7341 VSS.n7340 0.2255
R60954 VSS.n7339 VSS.n7338 0.2255
R60955 VSS.n7337 VSS.n7336 0.2255
R60956 VSS.n7333 VSS.n7332 0.2255
R60957 VSS.n7331 VSS.n7330 0.2255
R60958 VSS.n7318 VSS.n7317 0.2255
R60959 VSS.n7307 VSS.n7306 0.2255
R60960 VSS.n7300 VSS.n7299 0.2255
R60961 VSS.n7295 VSS.n7294 0.2255
R60962 VSS.n7291 VSS.n7290 0.2255
R60963 VSS.n7289 VSS.n7288 0.2255
R60964 VSS.n7287 VSS.n7286 0.2255
R60965 VSS.n7285 VSS.n7284 0.2255
R60966 VSS.n7283 VSS.n7282 0.2255
R60967 VSS.n7281 VSS.n7280 0.2255
R60968 VSS.n7279 VSS.n7278 0.2255
R60969 VSS.n7277 VSS.n7276 0.2255
R60970 VSS.n7275 VSS.n7274 0.2255
R60971 VSS.n7273 VSS.n7272 0.2255
R60972 VSS.n7271 VSS.n7270 0.2255
R60973 VSS.n7263 VSS.n7262 0.2255
R60974 VSS.n7256 VSS.n7255 0.2255
R60975 VSS.n7245 VSS.n7244 0.2255
R60976 VSS.n7239 VSS.n7238 0.2255
R60977 VSS.n7230 VSS.n7229 0.2255
R60978 VSS.n7221 VSS.n7220 0.2255
R60979 VSS.n7213 VSS.n7212 0.2255
R60980 VSS.n7211 VSS.n7210 0.2255
R60981 VSS.n7209 VSS.n7208 0.2255
R60982 VSS.n7207 VSS.n7206 0.2255
R60983 VSS.n7205 VSS.n7204 0.2255
R60984 VSS.n7203 VSS.n7202 0.2255
R60985 VSS.n7201 VSS.n7200 0.2255
R60986 VSS.n7199 VSS.n7198 0.2255
R60987 VSS.n7197 VSS.n7196 0.2255
R60988 VSS.n7191 VSS.n7190 0.2255
R60989 VSS.n7189 VSS.n7188 0.2255
R60990 VSS.n7182 VSS.n7181 0.2255
R60991 VSS.n7173 VSS.n7172 0.2255
R60992 VSS.n7163 VSS.n7162 0.2255
R60993 VSS.n7154 VSS.n7153 0.2255
R60994 VSS.n7152 VSS.n7151 0.2255
R60995 VSS.n7138 VSS.n7137 0.2255
R60996 VSS.n7123 VSS.n7122 0.2255
R60997 VSS.n7114 VSS.n7113 0.2255
R60998 VSS.n7104 VSS.n7103 0.2255
R60999 VSS.n7095 VSS.n7094 0.2255
R61000 VSS.n7089 VSS.n7088 0.2255
R61001 VSS.n7081 VSS.n7080 0.2255
R61002 VSS.n7074 VSS.n7073 0.2255
R61003 VSS.n7067 VSS.n7066 0.2255
R61004 VSS.n7058 VSS.n7057 0.2255
R61005 VSS.n7054 VSS.n7053 0.2255
R61006 VSS.n7519 VSS.n7518 0.2255
R61007 VSS.n7520 VSS.n7519 0.2255
R61008 VSS.n5911 VSS.n5910 0.2255
R61009 VSS.n4213 VSS.n2445 0.2255
R61010 VSS.n4691 VSS.n2445 0.2255
R61011 VSS.n4686 VSS.n4685 0.2255
R61012 VSS.n4681 VSS.n4680 0.2255
R61013 VSS.n4679 VSS.n4678 0.2255
R61014 VSS.n4677 VSS.n4676 0.2255
R61015 VSS.n4675 VSS.n4674 0.2255
R61016 VSS.n4673 VSS.n4672 0.2255
R61017 VSS.n4669 VSS.n4668 0.2255
R61018 VSS.n4649 VSS.n4648 0.2255
R61019 VSS.n4647 VSS.n4646 0.2255
R61020 VSS.n4645 VSS.n4644 0.2255
R61021 VSS.n4643 VSS.n4642 0.2255
R61022 VSS.n4641 VSS.n4640 0.2255
R61023 VSS.n4639 VSS.n4638 0.2255
R61024 VSS.n4634 VSS.n4633 0.2255
R61025 VSS.n4625 VSS.n4624 0.2255
R61026 VSS.n4620 VSS.n4619 0.2255
R61027 VSS.n4617 VSS.n4616 0.2255
R61028 VSS.n4615 VSS.n4614 0.2255
R61029 VSS.n4613 VSS.n4612 0.2255
R61030 VSS.n4611 VSS.n4610 0.2255
R61031 VSS.n4609 VSS.n4608 0.2255
R61032 VSS.n4607 VSS.n4606 0.2255
R61033 VSS.n4605 VSS.n4604 0.2255
R61034 VSS.n4603 VSS.n4602 0.2255
R61035 VSS.n4601 VSS.n4600 0.2255
R61036 VSS.n4599 VSS.n4598 0.2255
R61037 VSS.n4597 VSS.n4596 0.2255
R61038 VSS.n4595 VSS.n4594 0.2255
R61039 VSS.n4593 VSS.n4592 0.2255
R61040 VSS.n4588 VSS.n4587 0.2255
R61041 VSS.n4579 VSS.n4578 0.2255
R61042 VSS.n4574 VSS.n4573 0.2255
R61043 VSS.n4571 VSS.n4570 0.2255
R61044 VSS.n4569 VSS.n4568 0.2255
R61045 VSS.n4567 VSS.n4566 0.2255
R61046 VSS.n4565 VSS.n4564 0.2255
R61047 VSS.n4563 VSS.n4562 0.2255
R61048 VSS.n4561 VSS.n4560 0.2255
R61049 VSS.n4559 VSS.n4558 0.2255
R61050 VSS.n4557 VSS.n4556 0.2255
R61051 VSS.n4555 VSS.n4554 0.2255
R61052 VSS.n4553 VSS.n4552 0.2255
R61053 VSS.n4551 VSS.n4550 0.2255
R61054 VSS.n4549 VSS.n4548 0.2255
R61055 VSS.n4547 VSS.n4546 0.2255
R61056 VSS.n4541 VSS.n4540 0.2255
R61057 VSS.n4534 VSS.n4533 0.2255
R61058 VSS.n4522 VSS.n4521 0.2255
R61059 VSS.n4516 VSS.n4515 0.2255
R61060 VSS.n4506 VSS.n4505 0.2255
R61061 VSS.n4497 VSS.n4496 0.2255
R61062 VSS.n4491 VSS.n4490 0.2255
R61063 VSS.n4489 VSS.n4488 0.2255
R61064 VSS.n4487 VSS.n4486 0.2255
R61065 VSS.n4485 VSS.n4484 0.2255
R61066 VSS.n4483 VSS.n4482 0.2255
R61067 VSS.n4481 VSS.n4480 0.2255
R61068 VSS.n4479 VSS.n4478 0.2255
R61069 VSS.n4477 VSS.n4476 0.2255
R61070 VSS.n4475 VSS.n4474 0.2255
R61071 VSS.n4473 VSS.n4472 0.2255
R61072 VSS.n4471 VSS.n4470 0.2255
R61073 VSS.n4467 VSS.n4466 0.2255
R61074 VSS.n4461 VSS.n4460 0.2255
R61075 VSS.n4454 VSS.n4453 0.2255
R61076 VSS.n4447 VSS.n4446 0.2255
R61077 VSS.n4440 VSS.n4439 0.2255
R61078 VSS.n4438 VSS.n4437 0.2255
R61079 VSS.n4436 VSS.n4435 0.2255
R61080 VSS.n4434 VSS.n4433 0.2255
R61081 VSS.n4432 VSS.n4431 0.2255
R61082 VSS.n4430 VSS.n4429 0.2255
R61083 VSS.n4428 VSS.n4427 0.2255
R61084 VSS.n4426 VSS.n4425 0.2255
R61085 VSS.n4424 VSS.n4423 0.2255
R61086 VSS.n4422 VSS.n4421 0.2255
R61087 VSS.n4420 VSS.n4419 0.2255
R61088 VSS.n4418 VSS.n4417 0.2255
R61089 VSS.n4416 VSS.n4415 0.2255
R61090 VSS.n4410 VSS.n4409 0.2255
R61091 VSS.n4403 VSS.n4402 0.2255
R61092 VSS.n4396 VSS.n4395 0.2255
R61093 VSS.n4389 VSS.n4388 0.2255
R61094 VSS.n4387 VSS.n4386 0.2255
R61095 VSS.n4385 VSS.n4384 0.2255
R61096 VSS.n4383 VSS.n4382 0.2255
R61097 VSS.n4381 VSS.n4380 0.2255
R61098 VSS.n4375 VSS.n4374 0.2255
R61099 VSS.n4368 VSS.n4367 0.2255
R61100 VSS.n4361 VSS.n4360 0.2255
R61101 VSS.n4354 VSS.n4353 0.2255
R61102 VSS.n4352 VSS.n4351 0.2255
R61103 VSS.n4350 VSS.n4349 0.2255
R61104 VSS.n4348 VSS.n4347 0.2255
R61105 VSS.n4346 VSS.n4322 0.2255
R61106 VSS.n4346 VSS.n4345 0.2255
R61107 VSS.n4321 VSS.n4320 0.2255
R61108 VSS.n2438 VSS.n2437 0.2255
R61109 VSS.n2439 VSS.n2438 0.2255
R61110 VSS.n17713 VSS.n17712 0.2255
R61111 VSS.n4739 VSS.n4737 0.2255
R61112 VSS.n4740 VSS.n4739 0.2255
R61113 VSS.n4751 VSS.n4750 0.2255
R61114 VSS.n4750 VSS.n4749 0.2255
R61115 VSS.n17605 VSS.n17604 0.2255
R61116 VSS.n17604 VSS.n17603 0.2255
R61117 VSS.n17599 VSS.n17598 0.2255
R61118 VSS.n17597 VSS.n17596 0.2255
R61119 VSS.n17595 VSS.n17594 0.2255
R61120 VSS.n17593 VSS.n17592 0.2255
R61121 VSS.n17591 VSS.n17590 0.2255
R61122 VSS.n17582 VSS.n17581 0.2255
R61123 VSS.n17576 VSS.n17575 0.2255
R61124 VSS.n17574 VSS.n17573 0.2255
R61125 VSS.n17557 VSS.n17556 0.2255
R61126 VSS.n17546 VSS.n17545 0.2255
R61127 VSS.n17530 VSS.n17529 0.2255
R61128 VSS.n17499 VSS.n17498 0.2255
R61129 VSS.n17488 VSS.n17487 0.2255
R61130 VSS.n18096 VSS.n18095 0.2255
R61131 VSS.n18090 VSS.n18089 0.2255
R61132 VSS.n18088 VSS.n18087 0.2255
R61133 VSS.n18086 VSS.n18085 0.2255
R61134 VSS.n18084 VSS.n18083 0.2255
R61135 VSS.n18082 VSS.n18081 0.2255
R61136 VSS.n18080 VSS.n18079 0.2255
R61137 VSS.n18078 VSS.n18077 0.2255
R61138 VSS.n18076 VSS.n18075 0.2255
R61139 VSS.n18074 VSS.n18073 0.2255
R61140 VSS.n18072 VSS.n18071 0.2255
R61141 VSS.n18066 VSS.n18065 0.2255
R61142 VSS.n18055 VSS.n18054 0.2255
R61143 VSS.n18041 VSS.n18040 0.2255
R61144 VSS.n18035 VSS.n18034 0.2255
R61145 VSS.n18025 VSS.n18024 0.2255
R61146 VSS.n18014 VSS.n18013 0.2255
R61147 VSS.n18006 VSS.n18005 0.2255
R61148 VSS.n18004 VSS.n18003 0.2255
R61149 VSS.n18000 VSS.n17999 0.2255
R61150 VSS.n17998 VSS.n17997 0.2255
R61151 VSS.n17994 VSS.n17993 0.2255
R61152 VSS.n17992 VSS.n17991 0.2255
R61153 VSS.n17990 VSS.n17989 0.2255
R61154 VSS.n17988 VSS.n17987 0.2255
R61155 VSS.n17986 VSS.n17985 0.2255
R61156 VSS.n17984 VSS.n17983 0.2255
R61157 VSS.n17982 VSS.n17981 0.2255
R61158 VSS.n17974 VSS.n17973 0.2255
R61159 VSS.n17870 VSS.n17869 0.2255
R61160 VSS.n17861 VSS.n17860 0.2255
R61161 VSS.n17852 VSS.n17851 0.2255
R61162 VSS.n17850 VSS.n17849 0.2255
R61163 VSS.n17848 VSS.n17847 0.2255
R61164 VSS.n17846 VSS.n17845 0.2255
R61165 VSS.n17844 VSS.n17843 0.2255
R61166 VSS.n17842 VSS.n17841 0.2255
R61167 VSS.n17838 VSS.n17837 0.2255
R61168 VSS.n17836 VSS.n17835 0.2255
R61169 VSS.n17834 VSS.n17833 0.2255
R61170 VSS.n17832 VSS.n17831 0.2255
R61171 VSS.n17830 VSS.n17829 0.2255
R61172 VSS.n17828 VSS.n17827 0.2255
R61173 VSS.n17820 VSS.n17819 0.2255
R61174 VSS.n17809 VSS.n17808 0.2255
R61175 VSS.n17800 VSS.n17799 0.2255
R61176 VSS.n17791 VSS.n17790 0.2255
R61177 VSS.n17789 VSS.n17788 0.2255
R61178 VSS.n17787 VSS.n17786 0.2255
R61179 VSS.n17783 VSS.n17782 0.2255
R61180 VSS.n17775 VSS.n17774 0.2255
R61181 VSS.n17764 VSS.n17763 0.2255
R61182 VSS.n17755 VSS.n17754 0.2255
R61183 VSS.n17746 VSS.n17745 0.2255
R61184 VSS.n17744 VSS.n17743 0.2255
R61185 VSS.n17742 VSS.n17741 0.2255
R61186 VSS.n17740 VSS.n17739 0.2255
R61187 VSS.n17738 VSS.n17701 0.2255
R61188 VSS.n17738 VSS.n17737 0.2255
R61189 VSS.n14125 VSS.n14124 0.2255
R61190 VSS.n22007 VSS.n22006 0.2255
R61191 VSS.n22005 VSS.n21990 0.2255
R61192 VSS.n22004 VSS.n22003 0.2255
R61193 VSS.n22000 VSS.n21999 0.2255
R61194 VSS.n21998 VSS.n21992 0.2255
R61195 VSS.n21996 VSS.n21994 0.2255
R61196 VSS.n14129 VSS.n14128 0.2255
R61197 VSS.n14117 VSS.n13950 0.2255
R61198 VSS.n14116 VSS.n14115 0.2255
R61199 VSS.n14114 VSS.n13951 0.2255
R61200 VSS.n14113 VSS.n14112 0.2255
R61201 VSS.n14111 VSS.n13952 0.2255
R61202 VSS.n14107 VSS.n13956 0.2255
R61203 VSS.n14106 VSS.n14105 0.2255
R61204 VSS.n14103 VSS.n14102 0.2255
R61205 VSS.n14099 VSS.n14098 0.2255
R61206 VSS.n14095 VSS.n14094 0.2255
R61207 VSS.n14090 VSS.n13959 0.2255
R61208 VSS.n14089 VSS.n14088 0.2255
R61209 VSS.n14087 VSS.n13960 0.2255
R61210 VSS.n14086 VSS.n14085 0.2255
R61211 VSS.n14084 VSS.n13961 0.2255
R61212 VSS.n14083 VSS.n14082 0.2255
R61213 VSS.n14081 VSS.n13962 0.2255
R61214 VSS.n14080 VSS.n14079 0.2255
R61215 VSS.n14078 VSS.n13963 0.2255
R61216 VSS.n14077 VSS.n14076 0.2255
R61217 VSS.n14075 VSS.n13964 0.2255
R61218 VSS.n14074 VSS.n14073 0.2255
R61219 VSS.n14072 VSS.n13965 0.2255
R61220 VSS.n14070 VSS.n13967 0.2255
R61221 VSS.n14069 VSS.n14068 0.2255
R61222 VSS.n14067 VSS.n13968 0.2255
R61223 VSS.n14066 VSS.n14065 0.2255
R61224 VSS.n14064 VSS.n13969 0.2255
R61225 VSS.n14063 VSS.n14062 0.2255
R61226 VSS.n14061 VSS.n13970 0.2255
R61227 VSS.n14060 VSS.n14059 0.2255
R61228 VSS.n14058 VSS.n13971 0.2255
R61229 VSS.n14057 VSS.n14056 0.2255
R61230 VSS.n14055 VSS.n13972 0.2255
R61231 VSS.n14054 VSS.n14053 0.2255
R61232 VSS.n14052 VSS.n13973 0.2255
R61233 VSS.n14051 VSS.n14050 0.2255
R61234 VSS.n14049 VSS.n13974 0.2255
R61235 VSS.n14048 VSS.n14047 0.2255
R61236 VSS.n14046 VSS.n13975 0.2255
R61237 VSS.n14045 VSS.n14044 0.2255
R61238 VSS.n14043 VSS.n13976 0.2255
R61239 VSS.n14042 VSS.n14041 0.2255
R61240 VSS.n14039 VSS.n14038 0.2255
R61241 VSS.n14034 VSS.n13979 0.2255
R61242 VSS.n14033 VSS.n14032 0.2255
R61243 VSS.n14030 VSS.n14029 0.2255
R61244 VSS.n14027 VSS.n13980 0.2255
R61245 VSS.n14026 VSS.n14025 0.2255
R61246 VSS.n14021 VSS.n14020 0.2255
R61247 VSS.n14015 VSS.n14014 0.2255
R61248 VSS.n14012 VSS.n13981 0.2255
R61249 VSS.n14011 VSS.n14010 0.2255
R61250 VSS.n14009 VSS.n13982 0.2255
R61251 VSS.n14008 VSS.n14007 0.2255
R61252 VSS.n14006 VSS.n13983 0.2255
R61253 VSS.n14004 VSS.n13985 0.2255
R61254 VSS.n14001 VSS.n14000 0.2255
R61255 VSS.n13997 VSS.n13986 0.2255
R61256 VSS.n13996 VSS.n13995 0.2255
R61257 VSS.n13994 VSS.n13987 0.2255
R61258 VSS.n13993 VSS.n13992 0.2255
R61259 VSS.n13991 VSS.n13988 0.2255
R61260 VSS.n13990 VSS.n13989 0.2255
R61261 VSS.n22263 VSS.n0 0.2255
R61262 VSS.n22265 VSS.n22262 0.2255
R61263 VSS.n22265 VSS.n22264 0.2255
R61264 VSS.n2 VSS.n1 0.2255
R61265 VSS.n22107 VSS.n22106 0.2255
R61266 VSS.n22258 VSS.n22257 0.2255
R61267 VSS.n16377 VSS.n16376 0.225323
R61268 VSS.n1460 VSS.n1459 0.225323
R61269 VSS.n11303 VSS.n11301 0.225249
R61270 VSS.n1519 VSS.n1518 0.222388
R61271 VSS.n1535 VSS.n1533 0.222388
R61272 VSS.n1551 VSS.n1550 0.222388
R61273 VSS.n15420 VSS.n15418 0.222388
R61274 VSS.n1592 VSS.n1590 0.222388
R61275 VSS.n15224 VSS.n15221 0.222149
R61276 VSS.n15240 VSS.n15238 0.222149
R61277 VSS.n15252 VSS.n15250 0.222149
R61278 VSS.n15426 VSS.n15420 0.222149
R61279 VSS.n5523 VSS.n5521 0.220713
R61280 VSS.n5521 VSS.n5519 0.220713
R61281 VSS.n1148 VSS.n1147 0.220713
R61282 VSS.n1605 VSS.n1604 0.220473
R61283 VSS.n1792 VSS.n1791 0.220473
R61284 VSS.n15488 VSS.n15487 0.220234
R61285 VSS.n16023 VSS.n16022 0.219516
R61286 VSS.n15487 VSS.n15484 0.219516
R61287 VSS.n5667 VSS.n5666 0.21784
R61288 VSS.n20936 VSS.n20935 0.21784
R61289 VSS.n5818 VSS.n5817 0.21784
R61290 VSS.n5817 VSS.n5814 0.21784
R61291 VSS.n1250 VSS.n1249 0.21784
R61292 VSS.n1249 VSS.n1246 0.21784
R61293 VSS.n14248 VSS.n14247 0.216246
R61294 VSS.n13539 VSS.n13538 0.216246
R61295 VSS.n13548 VSS.n13547 0.216246
R61296 VSS.n13552 VSS.n13551 0.216246
R61297 VSS.n17178 VSS.n14328 0.216246
R61298 VSS.n14323 VSS.n14322 0.216246
R61299 VSS.n14319 VSS.n14318 0.216246
R61300 VSS.n14310 VSS.n14309 0.216246
R61301 VSS.n14306 VSS.n14305 0.216246
R61302 VSS.n15410 VSS.n15409 0.214725
R61303 VSS.n1726 VSS.n1725 0.214725
R61304 VSS.n5758 VSS.n5751 0.208878
R61305 VSS.n5698 VSS.n5664 0.208878
R61306 VSS.n20970 VSS.n20969 0.208878
R61307 VSS.n20969 VSS.n20967 0.208878
R61308 VSS.n20967 VSS.n20933 0.208878
R61309 VSS.n5701 VSS.n5700 0.208878
R61310 VSS.n5700 VSS.n5698 0.208878
R61311 VSS.n1213 VSS.n1212 0.208878
R61312 VSS.n20970 VSS.n20903 0.208878
R61313 VSS.n5758 VSS.n5757 0.208878
R61314 VSS.n16338 VSS.n16337 0.199888
R61315 VSS.n1426 VSS.n1425 0.199888
R61316 VSS.n16299 VSS.n16298 0.199888
R61317 VSS.n1382 VSS.n1381 0.199888
R61318 VSS.n16264 VSS.n16263 0.199888
R61319 VSS.n1348 VSS.n1347 0.199888
R61320 VSS.n9219 VSS.n9216 0.185308
R61321 VSS.n6386 VSS.n6383 0.185308
R61322 VSS.n9640 VSS.n9637 0.185308
R61323 VSS.n8650 VSS.n8647 0.185308
R61324 VSS.n9216 VSS.n9213 0.185115
R61325 VSS.n6389 VSS.n6386 0.185115
R61326 VSS.n9233 VSS.n9230 0.183192
R61327 VSS.n6412 VSS.n6409 0.183192
R61328 VSS.n9523 VSS.n9520 0.183192
R61329 VSS.n12612 VSS.n12609 0.183192
R61330 VSS.n5633 VSS.n5632 0.180146
R61331 VSS.n16155 VSS.n16154 0.180146
R61332 VSS.n21083 VSS.n21082 0.180146
R61333 VSS.n1135 VSS.n1134 0.180146
R61334 VSS.n1432 VSS.n1431 0.168293
R61335 VSS.n1387 VSS.n1385 0.168293
R61336 VSS.n1353 VSS.n1351 0.168293
R61337 VSS.n16346 VSS.n16343 0.168053
R61338 VSS.n16304 VSS.n16302 0.168053
R61339 VSS.n16269 VSS.n16267 0.168053
R61340 VSS.n861 VSS.n858 0.137763
R61341 DVSS VSS.n1469 0.136254
R61342 VSS.n15909 DVSS 0.136254
R61343 VSS.n15447 VSS.n15446 0.136134
R61344 VSS.n1749 VSS.n1748 0.136134
R61345 VSS.n19020 VSS.n19018 0.133972
R61346 VSS.n1977 VSS.n1975 0.133972
R61347 VSS.n2081 VSS.n2079 0.133972
R61348 VSS.n20050 VSS.n20048 0.133972
R61349 VSS.n13521 VSS.n13520 0.133972
R61350 VSS.n13442 VSS.n13440 0.133972
R61351 VSS.n13461 VSS.n2149 0.133972
R61352 VSS.n19168 VSS.n19166 0.133972
R61353 VSS.n18998 VSS.n18996 0.133833
R61354 VSS.n16401 VSS.n16399 0.133833
R61355 VSS.n15120 VSS.n15118 0.133833
R61356 VSS.n15087 VSS.n15085 0.133833
R61357 VSS.n14386 VSS.n14385 0.133833
R61358 VSS.n14445 VSS.n14443 0.133833
R61359 VSS.n18127 VSS.n18125 0.133833
R61360 VSS.n18848 VSS.n18846 0.133833
R61361 VSS.n15551 VSS.n15550 0.13381
R61362 VSS.n1839 VSS.n1838 0.13381
R61363 VSS.n4197 VSS.n4196 0.132444
R61364 VSS.n11375 VSS.n11374 0.132444
R61365 VSS.n11507 VSS.n11506 0.132444
R61366 VSS.n11598 VSS.n11597 0.132444
R61367 VSS.n17354 VSS.n17353 0.132444
R61368 VSS.n17431 VSS.n17429 0.132444
R61369 VSS.n4075 VSS.n3945 0.132444
R61370 VSS.n15631 VSS.n15630 0.128739
R61371 VSS.n15608 VSS.n15607 0.128739
R61372 VSS.n1899 VSS.n1898 0.128739
R61373 VSS.n1882 VSS.n1881 0.128739
R61374 VSS.n15658 VSS.n15657 0.128106
R61375 VSS.n1916 VSS.n1915 0.128106
R61376 VSS.n15585 VSS.n15584 0.127894
R61377 VSS.n1865 VSS.n1864 0.127894
R61378 VSS.n14237 VSS.n14236 0.120204
R61379 VSS.n22009 VSS.n22008 0.116341
R61380 VSS.n13664 VSS.n13663 0.116325
R61381 VSS VSS.n22259 0.115811
R61382 VSS.n21300 VSS.n21299 0.114949
R61383 VSS.n11456 VSS.n11455 0.114949
R61384 VSS.n5724 VSS.n5723 0.11424
R61385 VSS.n16172 VSS.n16171 0.11424
R61386 VSS.n21112 VSS.n21111 0.11424
R61387 VSS.n1162 VSS.n1161 0.11424
R61388 VSS.n5865 VSS.n5864 0.112291
R61389 VSS.n16226 VSS.n16225 0.112291
R61390 VSS.n21170 VSS.n21169 0.112291
R61391 VSS.n1299 VSS.n1298 0.112291
R61392 VSS.n8799 VSS.n8798 0.110613
R61393 VSS.n9412 VSS.n9411 0.110613
R61394 VSS.n6154 VSS.n6153 0.110613
R61395 VSS.n7027 VSS.n7026 0.110523
R61396 VSS.n7930 VSS.n7920 0.109536
R61397 VSS.n6359 VSS.n6349 0.109536
R61398 VSS.n11332 VSS.n11331 0.10928
R61399 VSS.n12879 VSS.n12878 0.10928
R61400 VSS.n15133 VSS.n15132 0.10928
R61401 VSS.n20781 VSS.n20780 0.10928
R61402 VSS.n2038 VSS.n2037 0.10928
R61403 VSS.n574 VSS.n573 0.10928
R61404 VSS.n17880 VSS.n17878 0.108278
R61405 VSS.n1990 VSS.n1988 0.108278
R61406 VSS.n2065 VSS.n2063 0.108278
R61407 VSS.n20063 VSS.n20061 0.108278
R61408 VSS.n14359 VSS.n14357 0.108278
R61409 VSS.n13431 VSS.n13430 0.108278
R61410 VSS.n13455 VSS.n13453 0.108278
R61411 VSS.n17962 VSS.n17960 0.108278
R61412 VSS.n2154 VSS.n2152 0.108278
R61413 VSS.n16321 VSS.n16320 0.108039
R61414 VSS.n16286 VSS.n16285 0.108039
R61415 VSS.n1402 VSS.n1401 0.108039
R61416 VSS.n1367 VSS.n1366 0.108039
R61417 VSS.n11717 VSS.n11716 0.107643
R61418 VSS.n20537 VSS.n20526 0.107643
R61419 VSS.n20537 VSS.n20536 0.107643
R61420 VSS.n20363 VSS.n20362 0.107643
R61421 VSS.n20349 VSS.n20348 0.107643
R61422 VSS.n20341 VSS.n20340 0.107643
R61423 VSS.n20335 VSS.n20334 0.107643
R61424 VSS.n20332 VSS.n20331 0.107643
R61425 VSS.n20330 VSS.n20329 0.107643
R61426 VSS.n20326 VSS.n20325 0.107643
R61427 VSS.n20324 VSS.n20323 0.107643
R61428 VSS.n20322 VSS.n20321 0.107643
R61429 VSS.n20320 VSS.n20319 0.107643
R61430 VSS.n20318 VSS.n20317 0.107643
R61431 VSS.n20316 VSS.n20315 0.107643
R61432 VSS.n20314 VSS.n20313 0.107643
R61433 VSS.n20312 VSS.n20311 0.107643
R61434 VSS.n20310 VSS.n20309 0.107643
R61435 VSS.n20308 VSS.n20307 0.107643
R61436 VSS.n20303 VSS.n20302 0.107643
R61437 VSS.n20295 VSS.n20294 0.107643
R61438 VSS.n20289 VSS.n20288 0.107643
R61439 VSS.n20286 VSS.n20285 0.107643
R61440 VSS.n20284 VSS.n20283 0.107643
R61441 VSS.n20282 VSS.n20281 0.107643
R61442 VSS.n20256 VSS.n20255 0.107643
R61443 VSS.n20247 VSS.n20246 0.107643
R61444 VSS.n20236 VSS.n20235 0.107643
R61445 VSS.n20219 VSS.n20218 0.107643
R61446 VSS.n20210 VSS.n20209 0.107643
R61447 VSS.n20202 VSS.n20201 0.107643
R61448 VSS.n20194 VSS.n20193 0.107643
R61449 VSS.n20192 VSS.n20191 0.107643
R61450 VSS.n20188 VSS.n20187 0.107643
R61451 VSS.n20186 VSS.n20185 0.107643
R61452 VSS.n20182 VSS.n20181 0.107643
R61453 VSS.n20180 VSS.n20179 0.107643
R61454 VSS.n20178 VSS.n20177 0.107643
R61455 VSS.n20173 VSS.n20172 0.107643
R61456 VSS.n732 VSS.n731 0.107643
R61457 VSS.n725 VSS.n724 0.107643
R61458 VSS.n717 VSS.n716 0.107643
R61459 VSS.n715 VSS.n714 0.107643
R61460 VSS.n713 VSS.n712 0.107643
R61461 VSS.n711 VSS.n710 0.107643
R61462 VSS.n709 VSS.n708 0.107643
R61463 VSS.n707 VSS.n706 0.107643
R61464 VSS.n705 VSS.n704 0.107643
R61465 VSS.n703 VSS.n702 0.107643
R61466 VSS.n701 VSS.n700 0.107643
R61467 VSS.n699 VSS.n698 0.107643
R61468 VSS.n697 VSS.n696 0.107643
R61469 VSS.n693 VSS.n692 0.107643
R61470 VSS.n687 VSS.n686 0.107643
R61471 VSS.n20588 VSS.n20587 0.107643
R61472 VSS.n20488 VSS.n20487 0.107643
R61473 VSS.n20490 VSS.n20489 0.107643
R61474 VSS.n20492 VSS.n20491 0.107643
R61475 VSS.n20494 VSS.n20493 0.107643
R61476 VSS.n20496 VSS.n20495 0.107643
R61477 VSS.n20498 VSS.n20497 0.107643
R61478 VSS.n20502 VSS.n20501 0.107643
R61479 VSS.n20506 VSS.n20505 0.107643
R61480 VSS.n20510 VSS.n20509 0.107643
R61481 VSS.n20512 VSS.n20511 0.107643
R61482 VSS.n20514 VSS.n20513 0.107643
R61483 VSS.n20516 VSS.n20515 0.107643
R61484 VSS.n20518 VSS.n20517 0.107643
R61485 VSS.n20550 VSS.n20549 0.107643
R61486 VSS.n20551 VSS.n20550 0.107643
R61487 VSS.n20548 VSS.n20547 0.107643
R61488 VSS.n20547 VSS.n20546 0.107643
R61489 VSS.n20401 VSS.n20400 0.107643
R61490 VSS.n20400 VSS.n20399 0.107643
R61491 VSS.n20396 VSS.n20395 0.107643
R61492 VSS.n20393 VSS.n20392 0.107643
R61493 VSS.n20391 VSS.n20390 0.107643
R61494 VSS.n20389 VSS.n20388 0.107643
R61495 VSS.n20387 VSS.n20386 0.107643
R61496 VSS.n20385 VSS.n20384 0.107643
R61497 VSS.n20380 VSS.n20379 0.107643
R61498 VSS.n20372 VSS.n20371 0.107643
R61499 VSS.n7034 VSS.n7033 0.107643
R61500 VSS.n8813 VSS.n8812 0.107643
R61501 VSS.n8817 VSS.n8816 0.107643
R61502 VSS.n8820 VSS.n8819 0.107643
R61503 VSS.n8822 VSS.n8821 0.107643
R61504 VSS.n8824 VSS.n8823 0.107643
R61505 VSS.n8826 VSS.n8825 0.107643
R61506 VSS.n8828 VSS.n8827 0.107643
R61507 VSS.n8846 VSS.n8845 0.107643
R61508 VSS.n8925 VSS.n8924 0.107643
R61509 VSS.n8995 VSS.n8994 0.107643
R61510 VSS.n9008 VSS.n9007 0.107643
R61511 VSS.n9012 VSS.n9011 0.107643
R61512 VSS.n9014 VSS.n9013 0.107643
R61513 VSS.n9403 VSS.n9402 0.107643
R61514 VSS.n9393 VSS.n9392 0.107643
R61515 VSS.n9385 VSS.n9384 0.107643
R61516 VSS.n9380 VSS.n9379 0.107643
R61517 VSS.n9378 VSS.n9377 0.107643
R61518 VSS.n9376 VSS.n9375 0.107643
R61519 VSS.n9374 VSS.n9373 0.107643
R61520 VSS.n9372 VSS.n9371 0.107643
R61521 VSS.n9370 VSS.n9369 0.107643
R61522 VSS.n9368 VSS.n9367 0.107643
R61523 VSS.n9366 VSS.n9365 0.107643
R61524 VSS.n9364 VSS.n9363 0.107643
R61525 VSS.n9362 VSS.n9361 0.107643
R61526 VSS.n9360 VSS.n9359 0.107643
R61527 VSS.n9358 VSS.n9357 0.107643
R61528 VSS.n9356 VSS.n9355 0.107643
R61529 VSS.n9349 VSS.n9348 0.107643
R61530 VSS.n9339 VSS.n9338 0.107643
R61531 VSS.n9331 VSS.n9330 0.107643
R61532 VSS.n9326 VSS.n9325 0.107643
R61533 VSS.n8439 VSS.n8438 0.107643
R61534 VSS.n8303 VSS.n8302 0.107643
R61535 VSS.n8292 VSS.n8291 0.107643
R61536 VSS.n8276 VSS.n8275 0.107643
R61537 VSS.n8265 VSS.n8264 0.107643
R61538 VSS.n8256 VSS.n8255 0.107643
R61539 VSS.n8242 VSS.n8241 0.107643
R61540 VSS.n6774 VSS.n6773 0.107643
R61541 VSS.n6765 VSS.n6764 0.107643
R61542 VSS.n6755 VSS.n6754 0.107643
R61543 VSS.n6745 VSS.n6744 0.107643
R61544 VSS.n6737 VSS.n6736 0.107643
R61545 VSS.n6735 VSS.n6734 0.107643
R61546 VSS.n6729 VSS.n6728 0.107643
R61547 VSS.n6727 VSS.n6726 0.107643
R61548 VSS.n6725 VSS.n6724 0.107643
R61549 VSS.n6723 VSS.n6722 0.107643
R61550 VSS.n6721 VSS.n6720 0.107643
R61551 VSS.n6714 VSS.n6713 0.107643
R61552 VSS.n6705 VSS.n6704 0.107643
R61553 VSS.n6695 VSS.n6694 0.107643
R61554 VSS.n7905 VSS.n7904 0.107643
R61555 VSS.n7901 VSS.n7900 0.107643
R61556 VSS.n7899 VSS.n7898 0.107643
R61557 VSS.n7892 VSS.n7891 0.107643
R61558 VSS.n7883 VSS.n7882 0.107643
R61559 VSS.n7873 VSS.n7872 0.107643
R61560 VSS.n7865 VSS.n7864 0.107643
R61561 VSS.n7019 VSS.n7018 0.107643
R61562 VSS.n7021 VSS.n7020 0.107643
R61563 VSS.n7858 VSS.n7857 0.107643
R61564 VSS.n7860 VSS.n7859 0.107643
R61565 VSS.n7855 VSS.n7854 0.107643
R61566 VSS.n7854 VSS.n7853 0.107643
R61567 VSS.n7043 VSS.n7042 0.107643
R61568 VSS.n7044 VSS.n7043 0.107643
R61569 VSS.n8805 VSS.n8804 0.107643
R61570 VSS.n8733 VSS.n8732 0.107643
R61571 VSS.n8602 VSS.n8601 0.107643
R61572 VSS.n8593 VSS.n8592 0.107643
R61573 VSS.n8090 VSS.n8089 0.107643
R61574 VSS.n8081 VSS.n8080 0.107643
R61575 VSS.n8071 VSS.n8070 0.107643
R61576 VSS.n8061 VSS.n8060 0.107643
R61577 VSS.n8059 VSS.n8058 0.107643
R61578 VSS.n8041 VSS.n8040 0.107643
R61579 VSS.n8037 VSS.n8036 0.107643
R61580 VSS.n8030 VSS.n8029 0.107643
R61581 VSS.n8021 VSS.n8020 0.107643
R61582 VSS.n8011 VSS.n8010 0.107643
R61583 VSS.n8001 VSS.n8000 0.107643
R61584 VSS.n7998 VSS.n7997 0.107643
R61585 VSS.n7994 VSS.n7993 0.107643
R61586 VSS.n7992 VSS.n7991 0.107643
R61587 VSS.n7985 VSS.n7984 0.107643
R61588 VSS.n7976 VSS.n7975 0.107643
R61589 VSS.n7966 VSS.n7965 0.107643
R61590 VSS.n7958 VSS.n7957 0.107643
R61591 VSS.n7954 VSS.n7918 0.107643
R61592 VSS.n7951 VSS.n7940 0.107643
R61593 VSS.n7951 VSS.n7950 0.107643
R61594 VSS.n7939 VSS.n7938 0.107643
R61595 VSS.n7938 VSS.n7937 0.107643
R61596 VSS.n7930 VSS.n7929 0.107643
R61597 VSS.n7929 VSS.n7928 0.107643
R61598 VSS.n9717 VSS.n9716 0.107643
R61599 VSS.n9715 VSS.n9714 0.107643
R61600 VSS.n8771 VSS.n8770 0.107643
R61601 VSS.n8760 VSS.n8759 0.107643
R61602 VSS.n8749 VSS.n8748 0.107643
R61603 VSS.n9418 VSS.n9417 0.107643
R61604 VSS.n9425 VSS.n9424 0.107643
R61605 VSS.n9430 VSS.n9429 0.107643
R61606 VSS.n9433 VSS.n9432 0.107643
R61607 VSS.n9435 VSS.n9434 0.107643
R61608 VSS.n9437 VSS.n9436 0.107643
R61609 VSS.n9439 VSS.n9438 0.107643
R61610 VSS.n9441 VSS.n9440 0.107643
R61611 VSS.n9449 VSS.n9448 0.107643
R61612 VSS.n9459 VSS.n9458 0.107643
R61613 VSS.n9465 VSS.n9464 0.107643
R61614 VSS.n9470 VSS.n9469 0.107643
R61615 VSS.n9472 VSS.n9471 0.107643
R61616 VSS.n9474 VSS.n9473 0.107643
R61617 VSS.n9476 VSS.n9475 0.107643
R61618 VSS.n9801 VSS.n9800 0.107643
R61619 VSS.n9794 VSS.n9793 0.107643
R61620 VSS.n9784 VSS.n9783 0.107643
R61621 VSS.n9776 VSS.n9775 0.107643
R61622 VSS.n9771 VSS.n9770 0.107643
R61623 VSS.n9767 VSS.n9766 0.107643
R61624 VSS.n9765 VSS.n9764 0.107643
R61625 VSS.n9763 VSS.n9762 0.107643
R61626 VSS.n9761 VSS.n9760 0.107643
R61627 VSS.n9759 VSS.n9758 0.107643
R61628 VSS.n9757 VSS.n9756 0.107643
R61629 VSS.n9755 VSS.n9754 0.107643
R61630 VSS.n9753 VSS.n9752 0.107643
R61631 VSS.n9751 VSS.n9750 0.107643
R61632 VSS.n9749 VSS.n9748 0.107643
R61633 VSS.n9747 VSS.n9746 0.107643
R61634 VSS.n9740 VSS.n9739 0.107643
R61635 VSS.n9730 VSS.n9729 0.107643
R61636 VSS.n9722 VSS.n9721 0.107643
R61637 VSS.n6359 VSS.n6358 0.107643
R61638 VSS.n6358 VSS.n6357 0.107643
R61639 VSS.n11071 VSS.n11070 0.107643
R61640 VSS.n11072 VSS.n6348 0.107643
R61641 VSS.n11079 VSS.n11078 0.107643
R61642 VSS.n11076 VSS.n6379 0.107643
R61643 VSS.n11076 VSS.n11075 0.107643
R61644 VSS.n6378 VSS.n6377 0.107643
R61645 VSS.n6377 VSS.n6376 0.107643
R61646 VSS.n6368 VSS.n6367 0.107643
R61647 VSS.n6367 VSS.n6366 0.107643
R61648 VSS.n11065 VSS.n11064 0.107643
R61649 VSS.n11054 VSS.n11053 0.107643
R61650 VSS.n11045 VSS.n11044 0.107643
R61651 VSS.n11036 VSS.n11035 0.107643
R61652 VSS.n11034 VSS.n11033 0.107643
R61653 VSS.n11032 VSS.n11031 0.107643
R61654 VSS.n11030 VSS.n11029 0.107643
R61655 VSS.n11027 VSS.n11026 0.107643
R61656 VSS.n10923 VSS.n10922 0.107643
R61657 VSS.n10934 VSS.n10933 0.107643
R61658 VSS.n10946 VSS.n10945 0.107643
R61659 VSS.n11001 VSS.n11000 0.107643
R61660 VSS.n11014 VSS.n11013 0.107643
R61661 VSS.n10910 VSS.n10909 0.107643
R61662 VSS.n10896 VSS.n10895 0.107643
R61663 VSS.n10868 VSS.n10867 0.107643
R61664 VSS.n10957 VSS.n10956 0.107643
R61665 VSS.n10960 VSS.n10959 0.107643
R61666 VSS.n10963 VSS.n10962 0.107643
R61667 VSS.n10968 VSS.n10967 0.107643
R61668 VSS.n10976 VSS.n10975 0.107643
R61669 VSS.n10990 VSS.n10989 0.107643
R61670 VSS.n10857 VSS.n10856 0.107643
R61671 VSS.n10842 VSS.n10841 0.107643
R61672 VSS.n10826 VSS.n10825 0.107643
R61673 VSS.n10814 VSS.n10813 0.107643
R61674 VSS.n10800 VSS.n10799 0.107643
R61675 VSS.n10789 VSS.n10788 0.107643
R61676 VSS.n10760 VSS.n10759 0.107643
R61677 VSS.n10757 VSS.n10756 0.107643
R61678 VSS.n10749 VSS.n10748 0.107643
R61679 VSS.n10729 VSS.n10728 0.107643
R61680 VSS.n10741 VSS.n10740 0.107643
R61681 VSS.n10718 VSS.n10717 0.107643
R61682 VSS.n10716 VSS.n10715 0.107643
R61683 VSS.n10714 VSS.n10713 0.107643
R61684 VSS.n10712 VSS.n10711 0.107643
R61685 VSS.n10710 VSS.n10709 0.107643
R61686 VSS.n10708 VSS.n10707 0.107643
R61687 VSS.n10706 VSS.n10705 0.107643
R61688 VSS.n10704 VSS.n10703 0.107643
R61689 VSS.n10702 VSS.n10701 0.107643
R61690 VSS.n10699 VSS.n10698 0.107643
R61691 VSS.n10696 VSS.n10695 0.107643
R61692 VSS.n10694 VSS.n10693 0.107643
R61693 VSS.n10687 VSS.n10686 0.107643
R61694 VSS.n10679 VSS.n10678 0.107643
R61695 VSS.n10638 VSS.n10637 0.107643
R61696 VSS.n10643 VSS.n10642 0.107643
R61697 VSS.n10645 VSS.n10644 0.107643
R61698 VSS.n10647 VSS.n10646 0.107643
R61699 VSS.n10653 VSS.n10652 0.107643
R61700 VSS.n10656 VSS.n10655 0.107643
R61701 VSS.n10667 VSS.n10666 0.107643
R61702 VSS.n6160 VSS.n6159 0.107643
R61703 VSS.n11180 VSS.n11178 0.107643
R61704 VSS.n11181 VSS.n11180 0.107643
R61705 VSS.n9805 VSS.n9804 0.107643
R61706 VSS.n9808 VSS.n9807 0.107643
R61707 VSS.n9810 VSS.n9809 0.107643
R61708 VSS.n9812 VSS.n9811 0.107643
R61709 VSS.n9814 VSS.n9813 0.107643
R61710 VSS.n9816 VSS.n9815 0.107643
R61711 VSS.n9823 VSS.n9822 0.107643
R61712 VSS.n10632 VSS.n10631 0.107643
R61713 VSS.n16366 VSS.n16365 0.107508
R61714 VSS.n1447 VSS.n1446 0.107508
R61715 VSS.n16250 VSS.n16249 0.107331
R61716 VSS.n1331 VSS.n1330 0.107331
R61717 VSS.n1425 VSS.n1422 0.101041
R61718 VSS.n16337 VSS.n16333 0.101041
R61719 VSS.n16337 VSS.n16336 0.101041
R61720 VSS.n1425 VSS.n1424 0.101041
R61721 VSS.n1381 VSS.n1378 0.101041
R61722 VSS.n16298 VSS.n16297 0.101041
R61723 VSS.n16263 VSS.n16262 0.101041
R61724 VSS.n1347 VSS.n1346 0.101041
R61725 DVSS VSS.n15907 0.0977905
R61726 VSS.n1471 DVSS 0.0975391
R61727 VSS.n21226 VSS.n21224 0.0945223
R61728 VSS.n11263 VSS.n11260 0.0945223
R61729 VSS.n155 VSS.n154 0.093014
R61730 VSS.n321 VSS.n320 0.093014
R61731 VSS.n21410 VSS.n21409 0.0929803
R61732 VSS.n11735 VSS.n11734 0.0929803
R61733 VSS.n154 VSS.n152 0.0915056
R61734 VSS.n320 VSS.n318 0.0915056
R61735 VSS.n13631 VSS.n13630 0.0913803
R61736 VSS.n14253 VSS.n14252 0.0913803
R61737 VSS.n22175 VSS.n22174 0.0913803
R61738 VSS.n21978 VSS.n21977 0.0913803
R61739 VSS.n21204 VSS.n21202 0.0889916
R61740 VSS.n11284 VSS.n11282 0.0889916
R61741 VSS.n17325 VSS.n17324 0.087311
R61742 VSS.n12993 VSS.n12992 0.087311
R61743 VSS.n14417 VSS.n14416 0.087311
R61744 VSS.n20153 VSS.n20152 0.087311
R61745 VSS.n123 VSS.n122 0.0859749
R61746 VSS.n122 VSS.n120 0.0859749
R61747 VSS.n289 VSS.n287 0.0859749
R61748 VSS.n290 VSS.n289 0.0859749
R61749 VSS.n22110 VSS.n22109 0.081839
R61750 VSS.n22112 VSS.n22111 0.081839
R61751 VSS.n22114 VSS.n22113 0.081839
R61752 VSS.n22116 VSS.n22115 0.081839
R61753 VSS.n22118 VSS.n22117 0.081839
R61754 VSS.n22161 VSS.n22119 0.081839
R61755 VSS.n22164 VSS.n22163 0.081839
R61756 VSS.n22252 VSS.n22239 0.081839
R61757 VSS.n13570 VSS.n13569 0.081839
R61758 VSS.n13568 VSS.n13567 0.081839
R61759 VSS.n13566 VSS.n13565 0.081839
R61760 VSS.n14251 VSS.n14242 0.081839
R61761 VSS.n13558 VSS.n13557 0.081839
R61762 VSS.n13560 VSS.n13559 0.081839
R61763 VSS.n13562 VSS.n13561 0.081839
R61764 VSS.n14275 VSS.n13563 0.081839
R61765 VSS.n13619 VSS.n13618 0.081839
R61766 VSS.n13617 VSS.n13616 0.081839
R61767 VSS.n13625 VSS.n13624 0.081839
R61768 VSS.n13627 VSS.n13626 0.081839
R61769 VSS.n13629 VSS.n13628 0.081839
R61770 VSS.n13633 VSS.n13632 0.081839
R61771 VSS.n13635 VSS.n13634 0.081839
R61772 VSS.n13637 VSS.n13636 0.081839
R61773 VSS.n13643 VSS.n13638 0.081839
R61774 VSS.n30 VSS.n29 0.081839
R61775 VSS.n28 VSS.n27 0.081839
R61776 VSS.n26 VSS.n25 0.081839
R61777 VSS.n21967 VSS.n21962 0.081839
R61778 VSS.n21970 VSS.n21969 0.081839
R61779 VSS.n21960 VSS.n21949 0.081839
R61780 VSS.n9842 VSS.n9841 0.0797308
R61781 VSS.n12634 VSS.n12633 0.0797308
R61782 DVSS VSS.n18994 0.0796667
R61783 VSS.n19022 DVSS 0.0796667
R61784 DVSS VSS.n16397 0.0796667
R61785 VSS.n1979 DVSS 0.0796667
R61786 VSS.n15122 DVSS 0.0796667
R61787 DVSS VSS.n2077 0.0796667
R61788 VSS.n15089 DVSS 0.0796667
R61789 VSS.n20052 DVSS 0.0796667
R61790 DVSS VSS.n14384 0.0796667
R61791 VSS.n13522 DVSS 0.0796667
R61792 DVSS VSS.n14441 0.0796667
R61793 VSS.n13444 DVSS 0.0796667
R61794 DVSS VSS.n18123 0.0796667
R61795 VSS.n13463 DVSS 0.0796667
R61796 VSS.n18850 DVSS 0.0796667
R61797 DVSS VSS.n19164 0.0796667
R61798 VSS.n21227 VSS.n21226 0.075919
R61799 VSS.n11260 VSS.n11258 0.075919
R61800 VSS.n4178 VSS.n4176 0.0728611
R61801 VSS.n17183 VSS.n17182 0.0728611
R61802 VSS.n17370 VSS.n17368 0.0728611
R61803 VSS.n17414 VSS.n17412 0.0728611
R61804 VSS.n8332 VSS.n8331 0.0693732
R61805 VSS.n8128 VSS.n8127 0.0693732
R61806 VSS.n13657 VSS.n13643 0.0687349
R61807 VSS.n14275 VSS.n14274 0.0687349
R61808 VSS.n13611 VSS.n13603 0.0682096
R61809 VSS.n21944 VSS.n33 0.0682096
R61810 VSS.n16260 VSS.n16258 0.0673919
R61811 VSS.n1344 VSS.n1342 0.0669865
R61812 VSS.n6554 VSS.n6551 0.0599231
R61813 VSS.n12633 VSS.n12630 0.0599231
R61814 VSS.n9063 VSS.n9054 0.0597308
R61815 VSS.n9039 VSS.n9038 0.0582559
R61816 VSS.n9182 VSS.n9181 0.0582559
R61817 VSS.n6672 VSS.n6671 0.0582559
R61818 VSS.n6522 VSS.n6521 0.0582559
R61819 VSS.n7675 VSS.n7674 0.0582559
R61820 VSS.n7763 VSS.n7762 0.0582559
R61821 VSS.n6086 VSS.n6085 0.0582559
R61822 VSS.n6005 VSS.n6004 0.0582559
R61823 VSS.n5662 VSS.n5660 0.0576622
R61824 VSS.n20931 VSS.n20929 0.0576622
R61825 VSS.n20884 VSS.n20883 0.0576622
R61826 VSS.n15900 VSS.n15899 0.056075
R61827 VSS.n22253 VSS.n22252 0.0550258
R61828 VSS.n21961 VSS.n21960 0.0550258
R61829 VSS.n18996 DVSS 0.0548056
R61830 VSS.n16399 DVSS 0.0548056
R61831 DVSS VSS.n15120 0.0548056
R61832 DVSS VSS.n15087 0.0548056
R61833 VSS.n14385 DVSS 0.0548056
R61834 VSS.n14443 DVSS 0.0548056
R61835 VSS.n18125 DVSS 0.0548056
R61836 DVSS VSS.n18848 0.0548056
R61837 VSS.n22253 VSS.n22237 0.0546818
R61838 VSS.n21961 VSS.n21947 0.0546818
R61839 DVSS VSS.n19020 0.0546667
R61840 DVSS VSS.n1977 0.0546667
R61841 VSS.n2079 DVSS 0.0546667
R61842 DVSS VSS.n20050 0.0546667
R61843 DVSS VSS.n13521 0.0546667
R61844 DVSS VSS.n13442 0.0546667
R61845 DVSS VSS.n13461 0.0546667
R61846 VSS.n19166 DVSS 0.0546667
R61847 VSS.n21713 VSS.n21711 0.0545278
R61848 VSS.n11408 VSS.n11406 0.0545278
R61849 VSS.n20846 VSS.n20844 0.0545278
R61850 VSS.n11478 VSS.n11475 0.0545278
R61851 VSS.n20754 VSS.n20752 0.0545278
R61852 VSS.n11631 VSS.n11629 0.0545278
R61853 VSS.n20703 VSS.n20701 0.0545278
R61854 VSS.n13260 VSS.n13259 0.0545278
R61855 VSS.n13381 VSS.n13379 0.0545278
R61856 VSS.n13289 VSS.n13287 0.0545278
R61857 VSS.n4107 VSS.n4105 0.0545278
R61858 VSS.n21903 VSS.n21901 0.0545278
R61859 VSS.n13603 VSS.n13572 0.0545
R61860 VSS.n13572 VSS.n13571 0.0545
R61861 VSS.n13622 VSS.n13621 0.0545
R61862 VSS.n13621 VSS.n13620 0.0545
R61863 VSS.n33 VSS.n32 0.0545
R61864 VSS.n32 VSS.n31 0.0545
R61865 VSS.n14672 VSS.n14671 0.0539507
R61866 VSS.n17164 VSS.n17163 0.0539507
R61867 VSS.n16872 VSS.n16871 0.0539507
R61868 VSS.n16683 VSS.n16682 0.0539507
R61869 VSS.n15703 VSS.n14994 0.0539507
R61870 VSS.n19769 VSS.n19768 0.0539507
R61871 VSS.n19859 VSS.n19858 0.0539507
R61872 VSS.n2130 VSS.n2129 0.0539507
R61873 VSS.n749 VSS.n739 0.0539507
R61874 VSS.n1968 VSS.n1967 0.0539507
R61875 VSS.n18474 VSS.n18473 0.0537394
R61876 VSS.n14572 VSS.n14571 0.0537394
R61877 VSS.n14823 VSS.n14822 0.0537394
R61878 VSS.n16696 VSS.n16695 0.0537394
R61879 VSS.n16445 VSS.n16444 0.0537394
R61880 VSS.n19565 VSS.n19564 0.0537394
R61881 VSS.n19756 VSS.n19755 0.0537394
R61882 VSS.n19846 VSS.n19845 0.0537394
R61883 VSS.n2098 VSS.n2097 0.0537394
R61884 VSS.n844 VSS.n843 0.0537394
R61885 VSS.n21727 VSS.n21725 0.0535556
R61886 VSS.n11391 VSS.n11389 0.0535556
R61887 VSS.n20860 VSS.n20858 0.0535556
R61888 VSS.n11494 VSS.n11492 0.0535556
R61889 VSS.n20768 VSS.n20766 0.0535556
R61890 VSS.n11614 VSS.n11612 0.0535556
R61891 VSS.n20717 VSS.n20715 0.0535556
R61892 VSS.n13267 VSS.n13266 0.0535556
R61893 VSS.n13395 VSS.n13393 0.0535556
R61894 VSS.n13304 VSS.n13302 0.0535556
R61895 VSS.n4092 VSS.n4089 0.0535556
R61896 VSS.n21887 VSS.n21885 0.0535556
R61897 VSS.n18670 VSS.n18669 0.0535282
R61898 VSS.n19533 VSS.n19532 0.0535282
R61899 VSS.n15901 VSS.n15863 0.0526831
R61900 VSS.n1936 VSS.n1935 0.0526831
R61901 VSS.n4171 VSS.n4169 0.0524444
R61902 VSS.n17233 VSS.n17232 0.0524444
R61903 VSS.n17377 VSS.n17375 0.0524444
R61904 VSS.n17407 VSS.n17405 0.0524444
R61905 VSS.n5702 VSS.n5701 0.0510053
R61906 VSS.n20971 VSS.n20970 0.0510053
R61907 VSS.n5698 VSS.n5697 0.0510053
R61908 VSS.n20967 VSS.n20966 0.0510053
R61909 VSS.n5759 VSS.n5758 0.0510053
R61910 VSS.n1214 VSS.n1213 0.0510053
R61911 DVSS VSS.n21200 0.0487682
R61912 VSS.n11287 DVSS 0.0487682
R61913 VSS.n14139 VSS.n14138 0.04775
R61914 VSS.n14143 VSS.n14142 0.04775
R61915 VSS.n14154 VSS.n14153 0.04775
R61916 VSS.n14158 VSS.n14157 0.04775
R61917 VSS.n14177 VSS.n14176 0.04775
R61918 VSS.n14181 VSS.n14180 0.04775
R61919 VSS.n14202 VSS.n14201 0.04775
R61920 VSS.n14198 VSS.n14197 0.04775
R61921 VSS.n14150 VSS.n14149 0.0455
R61922 VSS.n14207 VSS.n14185 0.0451759
R61923 VSS.n14148 VSS.n14147 0.0449197
R61924 VSS.n17231 VSS.n17230 0.0449145
R61925 VSS.n17220 VSS.n17219 0.0449145
R61926 VSS.n11748 VSS.n11747 0.0445103
R61927 VSS.n17225 VSS.n17224 0.0445103
R61928 VSS.n14207 VSS.n14206 0.0443278
R61929 VSS.n21711 VSS.n21709 0.04425
R61930 VSS.n11409 VSS.n11408 0.04425
R61931 VSS.n20844 VSS.n20842 0.04425
R61932 VSS.n11475 VSS.n11473 0.04425
R61933 VSS.n20752 VSS.n20750 0.04425
R61934 VSS.n11632 VSS.n11631 0.04425
R61935 VSS.n20701 VSS.n20699 0.04425
R61936 VSS.n13259 VSS.n13258 0.04425
R61937 VSS.n13379 VSS.n13377 0.04425
R61938 VSS.n13287 VSS.n13285 0.04425
R61939 VSS.n4108 VSS.n4107 0.04425
R61940 VSS.n21904 VSS.n21903 0.04425
R61941 VSS.n4169 VSS.n4167 0.0421667
R61942 VSS.n17234 VSS.n17233 0.0421667
R61943 VSS.n17378 VSS.n17377 0.0421667
R61944 VSS.n17405 VSS.n17403 0.0421667
R61945 DVSS VSS.n4178 0.0420278
R61946 VSS.n17182 DVSS 0.0420278
R61947 VSS.n17368 DVSS 0.0420278
R61948 DVSS VSS.n17414 0.0420278
R61949 VSS.n13611 VSS.n13610 0.0420015
R61950 VSS.n21944 VSS.n21943 0.0420015
R61951 VSS.n14274 VSS.n14273 0.0414881
R61952 VSS.n13657 VSS.n13656 0.0414881
R61953 VSS.n21202 DVSS 0.0407235
R61954 DVSS VSS.n11284 0.0407235
R61955 VSS.n22125 VSS.n22123 0.0403361
R61956 VSS.n22127 VSS.n22125 0.0403361
R61957 VSS.n22130 VSS.n22127 0.0403361
R61958 VSS.n22133 VSS.n22130 0.0403361
R61959 VSS.n22136 VSS.n22133 0.0403361
R61960 VSS.n22139 VSS.n22136 0.0403361
R61961 VSS.n22142 VSS.n22139 0.0403361
R61962 VSS.n22145 VSS.n22142 0.0403361
R61963 VSS.n22148 VSS.n22145 0.0403361
R61964 VSS.n22151 VSS.n22148 0.0403361
R61965 VSS.n22154 VSS.n22151 0.0403361
R61966 VSS.n22160 VSS.n22154 0.0403361
R61967 VSS.n22160 VSS.n22157 0.0403361
R61968 VSS.n22173 VSS.n22172 0.0403361
R61969 VSS.n22172 VSS.n22169 0.0403361
R61970 VSS.n22245 VSS.n22242 0.0403361
R61971 VSS.n22248 VSS.n22245 0.0403361
R61972 VSS.n22251 VSS.n22248 0.0403361
R61973 VSS.n22236 VSS.n22233 0.0403361
R61974 VSS.n22228 VSS.n22180 0.0403361
R61975 VSS.n22222 VSS.n22221 0.0403361
R61976 VSS.n22221 VSS.n22219 0.0403361
R61977 VSS.n22219 VSS.n22217 0.0403361
R61978 VSS.n22217 VSS.n22215 0.0403361
R61979 VSS.n22215 VSS.n22213 0.0403361
R61980 VSS.n22213 VSS.n22211 0.0403361
R61981 VSS.n22211 VSS.n22209 0.0403361
R61982 VSS.n22209 VSS.n22207 0.0403361
R61983 VSS.n22207 VSS.n22205 0.0403361
R61984 VSS.n22205 VSS.n22203 0.0403361
R61985 VSS.n22203 VSS.n22201 0.0403361
R61986 VSS.n22201 VSS.n22199 0.0403361
R61987 VSS.n22199 VSS.n22197 0.0403361
R61988 VSS.n22197 VSS.n22195 0.0403361
R61989 VSS.n22195 VSS.n22193 0.0403361
R61990 VSS.n22193 VSS.n22191 0.0403361
R61991 VSS.n22191 VSS.n22189 0.0403361
R61992 VSS.n22189 VSS.n22187 0.0403361
R61993 VSS.n22187 VSS.n22185 0.0403361
R61994 VSS.n22185 VSS.n22183 0.0403361
R61995 VSS.n13642 VSS.n13640 0.0403361
R61996 VSS.n13655 VSS.n13645 0.0403361
R61997 VSS.n21942 VSS.n21941 0.0403361
R61998 VSS.n24 VSS.n21 0.0403361
R61999 VSS.n21 VSS.n19 0.0403361
R62000 VSS.n19 VSS.n17 0.0403361
R62001 VSS.n17 VSS.n15 0.0403361
R62002 VSS.n15 VSS.n13 0.0403361
R62003 VSS.n13 VSS.n11 0.0403361
R62004 VSS.n11 VSS.n9 0.0403361
R62005 VSS.n9 VSS.n7 0.0403361
R62006 VSS.n7 VSS.n5 0.0403361
R62007 VSS.n21966 VSS.n21964 0.0403361
R62008 VSS.n21976 VSS.n21974 0.0403361
R62009 VSS.n21974 VSS.n21972 0.0403361
R62010 VSS.n21953 VSS.n21951 0.0403361
R62011 VSS.n21955 VSS.n21953 0.0403361
R62012 VSS.n21959 VSS.n21955 0.0403361
R62013 VSS.n21959 VSS.n21957 0.0403361
R62014 VSS.n21984 VSS.n21980 0.0403361
R62015 VSS.n13609 VSS.n13606 0.0403361
R62016 VSS.n13602 VSS.n13599 0.0403361
R62017 VSS.n13599 VSS.n13596 0.0403361
R62018 VSS.n13596 VSS.n13593 0.0403361
R62019 VSS.n13593 VSS.n13590 0.0403361
R62020 VSS.n13590 VSS.n13587 0.0403361
R62021 VSS.n13587 VSS.n13584 0.0403361
R62022 VSS.n13584 VSS.n13581 0.0403361
R62023 VSS.n13581 VSS.n13578 0.0403361
R62024 VSS.n13578 VSS.n13575 0.0403361
R62025 VSS.n13550 VSS.n13541 0.0403361
R62026 VSS.n13554 VSS.n13550 0.0403361
R62027 VSS.n14326 VSS.n13554 0.0403361
R62028 VSS.n14326 VSS.n14325 0.0403361
R62029 VSS.n14325 VSS.n14321 0.0403361
R62030 VSS.n14321 VSS.n14312 0.0403361
R62031 VSS.n14312 VSS.n14308 0.0403361
R62032 VSS.n14308 VSS.n14279 0.0403361
R62033 VSS.n14279 VSS.n14276 0.0403361
R62034 VSS.n14272 VSS.n14257 0.0403361
R62035 VSS.n14458 VSS.n14457 0.0402183
R62036 VSS.n19724 VSS.n19723 0.0402183
R62037 VSS.n19379 VSS.n19378 0.0401
R62038 VSS.n19008 VSS.n2162 0.0401
R62039 VSS.n18246 VSS.n18245 0.0401
R62040 VSS.n14966 VSS.n14964 0.0401
R62041 VSS.n17171 VSS.n14379 0.0401
R62042 VSS.n14663 VSS.n14659 0.0401
R62043 VSS.n14937 VSS.n14933 0.0401
R62044 VSS.n16426 VSS.n16424 0.0401
R62045 VSS.n17221 VSS.n17220 0.037361
R62046 VSS.n17230 VSS.n17229 0.037361
R62047 VSS.n17224 VSS.n17223 0.0372894
R62048 VSS.n11747 VSS.n11746 0.0372894
R62049 VSS.n14173 VSS.n14172 0.03515
R62050 VSS.n14194 VSS.n14193 0.03515
R62051 VSS.n20885 VSS.n20884 0.0337432
R62052 VSS.n15207 VSS.n15206 0.0333378
R62053 VSS.n1568 VSS.n1566 0.0333378
R62054 VSS.n5493 VSS.n5490 0.0333378
R62055 VSS.n1849 VSS.n1847 0.0333378
R62056 VSS.n17186 VSS.n17185 0.03245
R62057 VSS.n17192 VSS.n17191 0.032
R62058 VSS.n17206 VSS.n17205 0.032
R62059 VSS.n17212 VSS.n17211 0.032
R62060 VSS.n14185 VSS.n14184 0.0319852
R62061 VSS.n14147 VSS.n14146 0.0319852
R62062 VSS.n4180 DVSS 0.0313333
R62063 VSS.n21729 DVSS 0.0313333
R62064 DVSS VSS.n11387 0.0313333
R62065 VSS.n20862 DVSS 0.0313333
R62066 VSS.n11496 DVSS 0.0313333
R62067 VSS.n20770 DVSS 0.0313333
R62068 DVSS VSS.n11610 0.0313333
R62069 VSS.n20719 DVSS 0.0313333
R62070 DVSS VSS.n17181 0.0313333
R62071 VSS.n13268 DVSS 0.0313333
R62072 DVSS VSS.n17366 0.0313333
R62073 VSS.n13397 DVSS 0.0313333
R62074 VSS.n17416 DVSS 0.0313333
R62075 VSS.n13306 DVSS 0.0313333
R62076 DVSS VSS.n4087 0.0313333
R62077 DVSS VSS.n21883 0.0313333
R62078 VSS.n14206 VSS.n14205 0.0308013
R62079 VSS.n4654 VSS.n4653 0.03065
R62080 VSS.n4661 VSS.n4660 0.03065
R62081 VSS.n4663 VSS.n4662 0.03065
R62082 VSS.n1624 VSS.n1623 0.0300946
R62083 VSS.n17226 VSS.n17225 0.0291833
R62084 VSS.n11748 VSS.n11745 0.0291833
R62085 VSS.n4665 VSS.n4664 0.0291833
R62086 VSS.n14149 VSS.n14148 0.0291833
R62087 VSS.n17219 VSS.n17218 0.0289271
R62088 VSS.n17231 VSS.n17227 0.0289271
R62089 VSS.n2447 VSS.n2446 0.0289271
R62090 VSS.n2341 VSS.n2340 0.0289271
R62091 VSS.n20929 VSS.n20928 0.0288784
R62092 VSS.n14166 VSS.n14165 0.0285987
R62093 VSS.n14189 VSS.n14188 0.0285987
R62094 VSS.n5660 VSS.n5659 0.028473
R62095 VSS.n13620 VSS.n13619 0.027839
R62096 VSS.n13618 VSS.n13617 0.027839
R62097 VSS.n13626 VSS.n13625 0.027839
R62098 VSS.n13628 VSS.n13627 0.027839
R62099 VSS.n13634 VSS.n13633 0.027839
R62100 VSS.n13636 VSS.n13635 0.027839
R62101 VSS.n13638 VSS.n13637 0.027839
R62102 VSS.n13563 VSS.n13562 0.027839
R62103 VSS.n13561 VSS.n13560 0.027839
R62104 VSS.n13559 VSS.n13558 0.027839
R62105 VSS.n13567 VSS.n13566 0.027839
R62106 VSS.n13569 VSS.n13568 0.027839
R62107 VSS.n13571 VSS.n13570 0.027839
R62108 VSS.n22174 VSS.n22164 0.027839
R62109 VSS.n22119 VSS.n22118 0.027839
R62110 VSS.n22115 VSS.n22114 0.027839
R62111 VSS.n22111 VSS.n22110 0.027839
R62112 VSS.n22109 VSS.n22108 0.027839
R62113 VSS.n22113 VSS.n22112 0.027839
R62114 VSS.n22117 VSS.n22116 0.027839
R62115 VSS.n22163 VSS.n22162 0.027839
R62116 VSS.n22239 VSS.n22238 0.027839
R62117 VSS.n21949 VSS.n21948 0.027839
R62118 VSS.n21969 VSS.n21968 0.027839
R62119 VSS.n21977 VSS.n21970 0.027839
R62120 VSS.n27 VSS.n26 0.027839
R62121 VSS.n29 VSS.n28 0.027839
R62122 VSS.n31 VSS.n30 0.027839
R62123 VSS.n4653 VSS.n4652 0.02615
R62124 VSS.n4655 VSS.n4654 0.02615
R62125 VSS.n4662 VSS.n4661 0.02615
R62126 VSS.n4664 VSS.n4663 0.02615
R62127 VSS.n21245 VSS.n21234 0.0248803
R62128 VSS.n4196 VSS.n4194 0.0246667
R62129 VSS.n17878 VSS.n17877 0.0246667
R62130 VSS.n11374 VSS.n11372 0.0246667
R62131 VSS.n1988 VSS.n1987 0.0246667
R62132 VSS.n11506 VSS.n11504 0.0246667
R62133 VSS.n2063 VSS.n2062 0.0246667
R62134 VSS.n11597 VSS.n11595 0.0246667
R62135 VSS.n20061 VSS.n20060 0.0246667
R62136 VSS.n14357 VSS.n14356 0.0246667
R62137 VSS.n13430 VSS.n13429 0.0246667
R62138 VSS.n17353 VSS.n17351 0.0246667
R62139 VSS.n13453 VSS.n13452 0.0246667
R62140 VSS.n17429 VSS.n17427 0.0246667
R62141 VSS.n17960 VSS.n17959 0.0246667
R62142 VSS.n3945 VSS.n3943 0.0246667
R62143 VSS.n2152 VSS.n2151 0.0246667
R62144 VSS.n14136 VSS.n14135 0.024601
R62145 VSS.n14190 VSS.n14189 0.0245016
R62146 VSS.n14165 VSS.n14164 0.0245016
R62147 VSS.n14162 VSS.n14161 0.0243765
R62148 VSS.n14161 VSS.n14160 0.0237031
R62149 VSS.n14135 VSS.n14134 0.0234786
R62150 VSS.n15701 VSS.n15698 0.02345
R62151 VSS.n9201 VSS.n9198 0.0233846
R62152 VSS.n8499 VSS.n8496 0.0233846
R62153 VSS.n18757 VSS.n18756 0.0233169
R62154 VSS.n18758 VSS.n18757 0.0233169
R62155 VSS.n18759 VSS.n18758 0.0233169
R62156 VSS.n18760 VSS.n18759 0.0233169
R62157 VSS.n18761 VSS.n18760 0.0233169
R62158 VSS.n18762 VSS.n18761 0.0233169
R62159 VSS.n18763 VSS.n18762 0.0233169
R62160 VSS.n18764 VSS.n18763 0.0233169
R62161 VSS.n18765 VSS.n18764 0.0233169
R62162 VSS.n18766 VSS.n18765 0.0233169
R62163 VSS.n18767 VSS.n18766 0.0233169
R62164 VSS.n18768 VSS.n18767 0.0233169
R62165 VSS.n18769 VSS.n18768 0.0233169
R62166 VSS.n18770 VSS.n18769 0.0233169
R62167 VSS.n18771 VSS.n18770 0.0233169
R62168 VSS.n18772 VSS.n18771 0.0233169
R62169 VSS.n18666 VSS.n18656 0.0233169
R62170 VSS.n18656 VSS.n18649 0.0233169
R62171 VSS.n18649 VSS.n18642 0.0233169
R62172 VSS.n18642 VSS.n18635 0.0233169
R62173 VSS.n18635 VSS.n18628 0.0233169
R62174 VSS.n18628 VSS.n18621 0.0233169
R62175 VSS.n18621 VSS.n18614 0.0233169
R62176 VSS.n18614 VSS.n18607 0.0233169
R62177 VSS.n18607 VSS.n18600 0.0233169
R62178 VSS.n18600 VSS.n18593 0.0233169
R62179 VSS.n18593 VSS.n18586 0.0233169
R62180 VSS.n18586 VSS.n18579 0.0233169
R62181 VSS.n18579 VSS.n18572 0.0233169
R62182 VSS.n18572 VSS.n18565 0.0233169
R62183 VSS.n18565 VSS.n18552 0.0233169
R62184 VSS.n18552 VSS.n18551 0.0233169
R62185 VSS.n18551 VSS.n18544 0.0233169
R62186 VSS.n18544 VSS.n18537 0.0233169
R62187 VSS.n18537 VSS.n18530 0.0233169
R62188 VSS.n18530 VSS.n18523 0.0233169
R62189 VSS.n18523 VSS.n18516 0.0233169
R62190 VSS.n18516 VSS.n18509 0.0233169
R62191 VSS.n18509 VSS.n18502 0.0233169
R62192 VSS.n18502 VSS.n18495 0.0233169
R62193 VSS.n18495 VSS.n18488 0.0233169
R62194 VSS.n18390 VSS.n18359 0.0233169
R62195 VSS.n18359 VSS.n18352 0.0233169
R62196 VSS.n18352 VSS.n18345 0.0233169
R62197 VSS.n18345 VSS.n18338 0.0233169
R62198 VSS.n18338 VSS.n18331 0.0233169
R62199 VSS.n18331 VSS.n18324 0.0233169
R62200 VSS.n18324 VSS.n18317 0.0233169
R62201 VSS.n18317 VSS.n18310 0.0233169
R62202 VSS.n18310 VSS.n18303 0.0233169
R62203 VSS.n18303 VSS.n18214 0.0233169
R62204 VSS.n18214 VSS.n18213 0.0233169
R62205 VSS.n18213 VSS.n18212 0.0233169
R62206 VSS.n18212 VSS.n18211 0.0233169
R62207 VSS.n18211 VSS.n18210 0.0233169
R62208 VSS.n18210 VSS.n18209 0.0233169
R62209 VSS.n18209 VSS.n18208 0.0233169
R62210 VSS.n14477 VSS.n14470 0.0233169
R62211 VSS.n14484 VSS.n14477 0.0233169
R62212 VSS.n14491 VSS.n14484 0.0233169
R62213 VSS.n14498 VSS.n14491 0.0233169
R62214 VSS.n14505 VSS.n14498 0.0233169
R62215 VSS.n14512 VSS.n14505 0.0233169
R62216 VSS.n14519 VSS.n14512 0.0233169
R62217 VSS.n14526 VSS.n14519 0.0233169
R62218 VSS.n14533 VSS.n14526 0.0233169
R62219 VSS.n14540 VSS.n14533 0.0233169
R62220 VSS.n14547 VSS.n14540 0.0233169
R62221 VSS.n14554 VSS.n14547 0.0233169
R62222 VSS.n14561 VSS.n14554 0.0233169
R62223 VSS.n14586 VSS.n14561 0.0233169
R62224 VSS.n14586 VSS.n14585 0.0233169
R62225 VSS.n14585 VSS.n14584 0.0233169
R62226 VSS.n14584 VSS.n14583 0.0233169
R62227 VSS.n14583 VSS.n14582 0.0233169
R62228 VSS.n14582 VSS.n14581 0.0233169
R62229 VSS.n14581 VSS.n14580 0.0233169
R62230 VSS.n14580 VSS.n14579 0.0233169
R62231 VSS.n14579 VSS.n14578 0.0233169
R62232 VSS.n14578 VSS.n14577 0.0233169
R62233 VSS.n14577 VSS.n14576 0.0233169
R62234 VSS.n14576 VSS.n14575 0.0233169
R62235 VSS.n14682 VSS.n14675 0.0233169
R62236 VSS.n14689 VSS.n14682 0.0233169
R62237 VSS.n14690 VSS.n14689 0.0233169
R62238 VSS.n14697 VSS.n14690 0.0233169
R62239 VSS.n14698 VSS.n14697 0.0233169
R62240 VSS.n14705 VSS.n14698 0.0233169
R62241 VSS.n14712 VSS.n14705 0.0233169
R62242 VSS.n14719 VSS.n14712 0.0233169
R62243 VSS.n14720 VSS.n14719 0.0233169
R62244 VSS.n14727 VSS.n14720 0.0233169
R62245 VSS.n14728 VSS.n14727 0.0233169
R62246 VSS.n14729 VSS.n14728 0.0233169
R62247 VSS.n14730 VSS.n14729 0.0233169
R62248 VSS.n14808 VSS.n14730 0.0233169
R62249 VSS.n14809 VSS.n14808 0.0233169
R62250 VSS.n14810 VSS.n14809 0.0233169
R62251 VSS.n14811 VSS.n14810 0.0233169
R62252 VSS.n14812 VSS.n14811 0.0233169
R62253 VSS.n14813 VSS.n14812 0.0233169
R62254 VSS.n14814 VSS.n14813 0.0233169
R62255 VSS.n14815 VSS.n14814 0.0233169
R62256 VSS.n14816 VSS.n14815 0.0233169
R62257 VSS.n14817 VSS.n14816 0.0233169
R62258 VSS.n14818 VSS.n14817 0.0233169
R62259 VSS.n14819 VSS.n14818 0.0233169
R62260 VSS.n16868 VSS.n16855 0.0233169
R62261 VSS.n16855 VSS.n16848 0.0233169
R62262 VSS.n16848 VSS.n16841 0.0233169
R62263 VSS.n16841 VSS.n16834 0.0233169
R62264 VSS.n16834 VSS.n16827 0.0233169
R62265 VSS.n16827 VSS.n16820 0.0233169
R62266 VSS.n16820 VSS.n16813 0.0233169
R62267 VSS.n16813 VSS.n16806 0.0233169
R62268 VSS.n16806 VSS.n16799 0.0233169
R62269 VSS.n16799 VSS.n16792 0.0233169
R62270 VSS.n16792 VSS.n16785 0.0233169
R62271 VSS.n16785 VSS.n16778 0.0233169
R62272 VSS.n16778 VSS.n16771 0.0233169
R62273 VSS.n16771 VSS.n16764 0.0233169
R62274 VSS.n16764 VSS.n16751 0.0233169
R62275 VSS.n16751 VSS.n16750 0.0233169
R62276 VSS.n16750 VSS.n16743 0.0233169
R62277 VSS.n16743 VSS.n16736 0.0233169
R62278 VSS.n16736 VSS.n16729 0.0233169
R62279 VSS.n16729 VSS.n16722 0.0233169
R62280 VSS.n16722 VSS.n16715 0.0233169
R62281 VSS.n16715 VSS.n16708 0.0233169
R62282 VSS.n16708 VSS.n16701 0.0233169
R62283 VSS.n16701 VSS.n16700 0.0233169
R62284 VSS.n16700 VSS.n16699 0.0233169
R62285 VSS.n16679 VSS.n16666 0.0233169
R62286 VSS.n16500 VSS.n16499 0.0233169
R62287 VSS.n16499 VSS.n16492 0.0233169
R62288 VSS.n16492 VSS.n16485 0.0233169
R62289 VSS.n16485 VSS.n16478 0.0233169
R62290 VSS.n16478 VSS.n16471 0.0233169
R62291 VSS.n16471 VSS.n16464 0.0233169
R62292 VSS.n16464 VSS.n16457 0.0233169
R62293 VSS.n16457 VSS.n16450 0.0233169
R62294 VSS.n16450 VSS.n16449 0.0233169
R62295 VSS.n16449 VSS.n16448 0.0233169
R62296 VSS.n15725 VSS.n15718 0.0233169
R62297 VSS.n15732 VSS.n15725 0.0233169
R62298 VSS.n15739 VSS.n15732 0.0233169
R62299 VSS.n15746 VSS.n15739 0.0233169
R62300 VSS.n15753 VSS.n15746 0.0233169
R62301 VSS.n15760 VSS.n15753 0.0233169
R62302 VSS.n15767 VSS.n15760 0.0233169
R62303 VSS.n15774 VSS.n15767 0.0233169
R62304 VSS.n15781 VSS.n15774 0.0233169
R62305 VSS.n15788 VSS.n15781 0.0233169
R62306 VSS.n15795 VSS.n15788 0.0233169
R62307 VSS.n15802 VSS.n15795 0.0233169
R62308 VSS.n15809 VSS.n15802 0.0233169
R62309 VSS.n15810 VSS.n15809 0.0233169
R62310 VSS.n15823 VSS.n15810 0.0233169
R62311 VSS.n15830 VSS.n15823 0.0233169
R62312 VSS.n15837 VSS.n15830 0.0233169
R62313 VSS.n15844 VSS.n15837 0.0233169
R62314 VSS.n15851 VSS.n15844 0.0233169
R62315 VSS.n15855 VSS.n15851 0.0233169
R62316 VSS.n15856 VSS.n15855 0.0233169
R62317 VSS.n15857 VSS.n15856 0.0233169
R62318 VSS.n15858 VSS.n15857 0.0233169
R62319 VSS.n15859 VSS.n15858 0.0233169
R62320 VSS.n15860 VSS.n15859 0.0233169
R62321 VSS.n19286 VSS.n19279 0.0233169
R62322 VSS.n19293 VSS.n19286 0.0233169
R62323 VSS.n19300 VSS.n19293 0.0233169
R62324 VSS.n19307 VSS.n19300 0.0233169
R62325 VSS.n19314 VSS.n19307 0.0233169
R62326 VSS.n19321 VSS.n19314 0.0233169
R62327 VSS.n19328 VSS.n19321 0.0233169
R62328 VSS.n19335 VSS.n19328 0.0233169
R62329 VSS.n19342 VSS.n19335 0.0233169
R62330 VSS.n19438 VSS.n19342 0.0233169
R62331 VSS.n19439 VSS.n19438 0.0233169
R62332 VSS.n19440 VSS.n19439 0.0233169
R62333 VSS.n19441 VSS.n19440 0.0233169
R62334 VSS.n19442 VSS.n19441 0.0233169
R62335 VSS.n19443 VSS.n19442 0.0233169
R62336 VSS.n19444 VSS.n19443 0.0233169
R62337 VSS.n19537 VSS.n19536 0.0233169
R62338 VSS.n19538 VSS.n19537 0.0233169
R62339 VSS.n19539 VSS.n19538 0.0233169
R62340 VSS.n19540 VSS.n19539 0.0233169
R62341 VSS.n19541 VSS.n19540 0.0233169
R62342 VSS.n19542 VSS.n19541 0.0233169
R62343 VSS.n19543 VSS.n19542 0.0233169
R62344 VSS.n19544 VSS.n19543 0.0233169
R62345 VSS.n19545 VSS.n19544 0.0233169
R62346 VSS.n19546 VSS.n19545 0.0233169
R62347 VSS.n19547 VSS.n19546 0.0233169
R62348 VSS.n19548 VSS.n19547 0.0233169
R62349 VSS.n19549 VSS.n19548 0.0233169
R62350 VSS.n19550 VSS.n19549 0.0233169
R62351 VSS.n19551 VSS.n19550 0.0233169
R62352 VSS.n19552 VSS.n19551 0.0233169
R62353 VSS.n19553 VSS.n19552 0.0233169
R62354 VSS.n19554 VSS.n19553 0.0233169
R62355 VSS.n19555 VSS.n19554 0.0233169
R62356 VSS.n19556 VSS.n19555 0.0233169
R62357 VSS.n19557 VSS.n19556 0.0233169
R62358 VSS.n19558 VSS.n19557 0.0233169
R62359 VSS.n19559 VSS.n19558 0.0233169
R62360 VSS.n19560 VSS.n19559 0.0233169
R62361 VSS.n19561 VSS.n19560 0.0233169
R62362 VSS.n19632 VSS.n19631 0.0233169
R62363 VSS.n19633 VSS.n19632 0.0233169
R62364 VSS.n19634 VSS.n19633 0.0233169
R62365 VSS.n19635 VSS.n19634 0.0233169
R62366 VSS.n19636 VSS.n19635 0.0233169
R62367 VSS.n19637 VSS.n19636 0.0233169
R62368 VSS.n19638 VSS.n19637 0.0233169
R62369 VSS.n19639 VSS.n19638 0.0233169
R62370 VSS.n19640 VSS.n19639 0.0233169
R62371 VSS.n19641 VSS.n19640 0.0233169
R62372 VSS.n19642 VSS.n19641 0.0233169
R62373 VSS.n19643 VSS.n19642 0.0233169
R62374 VSS.n19644 VSS.n19643 0.0233169
R62375 VSS.n19645 VSS.n19644 0.0233169
R62376 VSS.n19646 VSS.n19645 0.0233169
R62377 VSS.n19647 VSS.n19646 0.0233169
R62378 VSS.n19728 VSS.n19727 0.0233169
R62379 VSS.n19729 VSS.n19728 0.0233169
R62380 VSS.n19730 VSS.n19729 0.0233169
R62381 VSS.n19731 VSS.n19730 0.0233169
R62382 VSS.n19732 VSS.n19731 0.0233169
R62383 VSS.n19733 VSS.n19732 0.0233169
R62384 VSS.n19734 VSS.n19733 0.0233169
R62385 VSS.n19735 VSS.n19734 0.0233169
R62386 VSS.n19736 VSS.n19735 0.0233169
R62387 VSS.n19737 VSS.n19736 0.0233169
R62388 VSS.n19738 VSS.n19737 0.0233169
R62389 VSS.n19739 VSS.n19738 0.0233169
R62390 VSS.n19740 VSS.n19739 0.0233169
R62391 VSS.n19741 VSS.n19740 0.0233169
R62392 VSS.n19742 VSS.n19741 0.0233169
R62393 VSS.n19743 VSS.n19742 0.0233169
R62394 VSS.n19744 VSS.n19743 0.0233169
R62395 VSS.n19745 VSS.n19744 0.0233169
R62396 VSS.n19746 VSS.n19745 0.0233169
R62397 VSS.n19747 VSS.n19746 0.0233169
R62398 VSS.n19748 VSS.n19747 0.0233169
R62399 VSS.n19749 VSS.n19748 0.0233169
R62400 VSS.n19750 VSS.n19749 0.0233169
R62401 VSS.n19751 VSS.n19750 0.0233169
R62402 VSS.n19752 VSS.n19751 0.0233169
R62403 VSS.n19782 VSS.n19781 0.0233169
R62404 VSS.n19783 VSS.n19782 0.0233169
R62405 VSS.n19790 VSS.n19783 0.0233169
R62406 VSS.n19791 VSS.n19790 0.0233169
R62407 VSS.n19798 VSS.n19791 0.0233169
R62408 VSS.n19799 VSS.n19798 0.0233169
R62409 VSS.n19800 VSS.n19799 0.0233169
R62410 VSS.n19801 VSS.n19800 0.0233169
R62411 VSS.n19808 VSS.n19801 0.0233169
R62412 VSS.n19809 VSS.n19808 0.0233169
R62413 VSS.n19816 VSS.n19809 0.0233169
R62414 VSS.n19823 VSS.n19816 0.0233169
R62415 VSS.n19830 VSS.n19823 0.0233169
R62416 VSS.n19831 VSS.n19830 0.0233169
R62417 VSS.n19832 VSS.n19831 0.0233169
R62418 VSS.n19833 VSS.n19832 0.0233169
R62419 VSS.n19834 VSS.n19833 0.0233169
R62420 VSS.n19835 VSS.n19834 0.0233169
R62421 VSS.n19836 VSS.n19835 0.0233169
R62422 VSS.n19837 VSS.n19836 0.0233169
R62423 VSS.n19838 VSS.n19837 0.0233169
R62424 VSS.n19839 VSS.n19838 0.0233169
R62425 VSS.n19840 VSS.n19839 0.0233169
R62426 VSS.n19841 VSS.n19840 0.0233169
R62427 VSS.n19842 VSS.n19841 0.0233169
R62428 VSS.n2126 VSS.n2125 0.0233169
R62429 VSS.n2125 VSS.n2124 0.0233169
R62430 VSS.n2124 VSS.n2123 0.0233169
R62431 VSS.n2123 VSS.n2122 0.0233169
R62432 VSS.n2122 VSS.n2121 0.0233169
R62433 VSS.n2121 VSS.n2120 0.0233169
R62434 VSS.n2120 VSS.n2119 0.0233169
R62435 VSS.n2119 VSS.n2118 0.0233169
R62436 VSS.n2118 VSS.n2117 0.0233169
R62437 VSS.n2117 VSS.n2116 0.0233169
R62438 VSS.n2116 VSS.n2115 0.0233169
R62439 VSS.n2115 VSS.n2114 0.0233169
R62440 VSS.n2114 VSS.n2113 0.0233169
R62441 VSS.n2113 VSS.n2112 0.0233169
R62442 VSS.n2112 VSS.n2111 0.0233169
R62443 VSS.n2111 VSS.n2110 0.0233169
R62444 VSS.n2110 VSS.n2109 0.0233169
R62445 VSS.n2109 VSS.n2108 0.0233169
R62446 VSS.n2108 VSS.n2107 0.0233169
R62447 VSS.n2107 VSS.n2106 0.0233169
R62448 VSS.n2106 VSS.n2105 0.0233169
R62449 VSS.n2105 VSS.n2104 0.0233169
R62450 VSS.n2104 VSS.n2103 0.0233169
R62451 VSS.n2103 VSS.n2102 0.0233169
R62452 VSS.n2102 VSS.n2101 0.0233169
R62453 VSS.n753 VSS.n752 0.0233169
R62454 VSS.n831 VSS.n830 0.0233169
R62455 VSS.n832 VSS.n831 0.0233169
R62456 VSS.n833 VSS.n832 0.0233169
R62457 VSS.n834 VSS.n833 0.0233169
R62458 VSS.n835 VSS.n834 0.0233169
R62459 VSS.n836 VSS.n835 0.0233169
R62460 VSS.n837 VSS.n836 0.0233169
R62461 VSS.n838 VSS.n837 0.0233169
R62462 VSS.n839 VSS.n838 0.0233169
R62463 VSS.n840 VSS.n839 0.0233169
R62464 VSS.n1964 VSS.n1963 0.0233169
R62465 VSS.n1963 VSS.n1962 0.0233169
R62466 VSS.n1962 VSS.n1961 0.0233169
R62467 VSS.n1961 VSS.n1960 0.0233169
R62468 VSS.n1960 VSS.n1959 0.0233169
R62469 VSS.n1959 VSS.n1958 0.0233169
R62470 VSS.n1958 VSS.n1957 0.0233169
R62471 VSS.n1957 VSS.n1956 0.0233169
R62472 VSS.n1956 VSS.n1955 0.0233169
R62473 VSS.n1955 VSS.n1954 0.0233169
R62474 VSS.n1954 VSS.n1953 0.0233169
R62475 VSS.n1953 VSS.n1952 0.0233169
R62476 VSS.n1952 VSS.n1951 0.0233169
R62477 VSS.n1951 VSS.n1950 0.0233169
R62478 VSS.n1950 VSS.n1949 0.0233169
R62479 VSS.n1949 VSS.n1948 0.0233169
R62480 VSS.n1948 VSS.n1947 0.0233169
R62481 VSS.n1947 VSS.n1946 0.0233169
R62482 VSS.n1946 VSS.n1945 0.0233169
R62483 VSS.n1945 VSS.n1944 0.0233169
R62484 VSS.n1944 VSS.n1943 0.0233169
R62485 VSS.n1943 VSS.n1942 0.0233169
R62486 VSS.n1942 VSS.n1941 0.0233169
R62487 VSS.n1941 VSS.n1940 0.0233169
R62488 VSS.n1940 VSS.n1939 0.0233169
R62489 DVSS VSS.n21727 0.0227222
R62490 VSS.n11389 DVSS 0.0227222
R62491 DVSS VSS.n20860 0.0227222
R62492 DVSS VSS.n11494 0.0227222
R62493 DVSS VSS.n20768 0.0227222
R62494 VSS.n11612 DVSS 0.0227222
R62495 DVSS VSS.n20717 0.0227222
R62496 DVSS VSS.n13267 0.0227222
R62497 DVSS VSS.n13395 0.0227222
R62498 DVSS VSS.n13304 0.0227222
R62499 VSS.n4089 DVSS 0.0227222
R62500 VSS.n21885 DVSS 0.0227222
R62501 VSS.n15542 VSS.n15541 0.0226831
R62502 VSS.n15538 VSS.n15537 0.0226831
R62503 VSS.n15460 VSS.n15459 0.0226831
R62504 VSS.n15451 VSS.n15450 0.0226831
R62505 VSS.n15372 VSS.n15371 0.0226831
R62506 VSS.n15368 VSS.n15367 0.0226831
R62507 VSS.n15364 VSS.n15363 0.0226831
R62508 VSS.n15355 VSS.n15354 0.0226831
R62509 VSS.n15351 VSS.n15350 0.0226831
R62510 VSS.n8458 VSS.n8457 0.0226831
R62511 VSS.n8462 VSS.n8461 0.0226831
R62512 VSS.n8471 VSS.n8470 0.0226831
R62513 VSS.n8475 VSS.n8474 0.0226831
R62514 VSS.n8522 VSS.n8521 0.0226831
R62515 VSS.n8574 VSS.n8573 0.0226831
R62516 VSS.n8570 VSS.n8569 0.0226831
R62517 VSS.n8566 VSS.n8565 0.0226831
R62518 VSS.n8557 VSS.n8556 0.0226831
R62519 VSS.n8553 VSS.n8552 0.0226831
R62520 VSS.n8544 VSS.n8543 0.0226831
R62521 VSS.n8540 VSS.n8539 0.0226831
R62522 VSS.n8310 VSS.n8309 0.0226831
R62523 VSS.n8319 VSS.n8318 0.0226831
R62524 VSS.n8323 VSS.n8322 0.0226831
R62525 VSS.n8336 VSS.n8335 0.0226831
R62526 VSS.n8340 VSS.n8339 0.0226831
R62527 VSS.n8429 VSS.n8428 0.0226831
R62528 VSS.n8425 VSS.n8424 0.0226831
R62529 VSS.n8421 VSS.n8420 0.0226831
R62530 VSS.n8412 VSS.n8411 0.0226831
R62531 VSS.n8408 VSS.n8407 0.0226831
R62532 VSS.n8399 VSS.n8398 0.0226831
R62533 VSS.n8395 VSS.n8394 0.0226831
R62534 VSS.n8382 VSS.n8381 0.0226831
R62535 VSS.n8378 VSS.n8377 0.0226831
R62536 VSS.n8369 VSS.n8368 0.0226831
R62537 VSS.n8365 VSS.n8364 0.0226831
R62538 VSS.n1830 VSS.n1829 0.0226831
R62539 VSS.n1826 VSS.n1825 0.0226831
R62540 VSS.n1762 VSS.n1761 0.0226831
R62541 VSS.n1753 VSS.n1752 0.0226831
R62542 VSS.n1688 VSS.n1687 0.0226831
R62543 VSS.n1684 VSS.n1683 0.0226831
R62544 VSS.n1680 VSS.n1679 0.0226831
R62545 VSS.n1671 VSS.n1670 0.0226831
R62546 VSS.n1667 VSS.n1666 0.0226831
R62547 VSS.n8609 VSS.n8608 0.0226831
R62548 VSS.n8613 VSS.n8612 0.0226831
R62549 VSS.n8622 VSS.n8621 0.0226831
R62550 VSS.n8626 VSS.n8625 0.0226831
R62551 VSS.n8673 VSS.n8672 0.0226831
R62552 VSS.n8725 VSS.n8724 0.0226831
R62553 VSS.n8721 VSS.n8720 0.0226831
R62554 VSS.n8717 VSS.n8716 0.0226831
R62555 VSS.n8708 VSS.n8707 0.0226831
R62556 VSS.n8704 VSS.n8703 0.0226831
R62557 VSS.n8695 VSS.n8694 0.0226831
R62558 VSS.n8691 VSS.n8690 0.0226831
R62559 VSS.n8106 VSS.n8105 0.0226831
R62560 VSS.n8115 VSS.n8114 0.0226831
R62561 VSS.n8119 VSS.n8118 0.0226831
R62562 VSS.n8132 VSS.n8131 0.0226831
R62563 VSS.n8136 VSS.n8135 0.0226831
R62564 VSS.n8237 VSS.n8236 0.0226831
R62565 VSS.n8233 VSS.n8232 0.0226831
R62566 VSS.n8229 VSS.n8228 0.0226831
R62567 VSS.n8220 VSS.n8219 0.0226831
R62568 VSS.n8216 VSS.n8215 0.0226831
R62569 VSS.n8207 VSS.n8206 0.0226831
R62570 VSS.n8203 VSS.n8202 0.0226831
R62571 VSS.n8190 VSS.n8189 0.0226831
R62572 VSS.n8186 VSS.n8185 0.0226831
R62573 VSS.n8177 VSS.n8176 0.0226831
R62574 VSS.n8173 VSS.n8172 0.0226831
R62575 VSS.n15920 VSS.n15918 0.0223919
R62576 VSS.n15926 VSS.n15920 0.0223919
R62577 VSS.n15926 VSS.n15925 0.0223919
R62578 VSS.n15925 VSS.n15923 0.0223919
R62579 VSS.n15932 VSS.n15928 0.0223919
R62580 VSS.n15932 VSS.n15931 0.0223919
R62581 VSS.n15216 VSS.n15215 0.0223919
R62582 VSS.n15210 VSS.n15202 0.0223919
R62583 VSS.n15210 VSS.n15209 0.0223919
R62584 VSS.n15209 VSS.n15207 0.0223919
R62585 VSS.n1483 VSS.n1481 0.0223919
R62586 VSS.n1487 VSS.n1483 0.0223919
R62587 VSS.n1487 VSS.n1486 0.0223919
R62588 VSS.n1493 VSS.n1489 0.0223919
R62589 VSS.n897 VSS.n891 0.0223919
R62590 VSS.n897 VSS.n896 0.0223919
R62591 VSS.n896 VSS.n894 0.0223919
R62592 VSS.n907 VSS.n899 0.0223919
R62593 VSS.n907 VSS.n906 0.0223919
R62594 VSS.n906 VSS.n904 0.0223919
R62595 VSS.n15977 VSS.n15971 0.0223919
R62596 VSS.n15977 VSS.n15975 0.0223919
R62597 VSS.n15975 VSS.n15973 0.0223919
R62598 VSS.n15985 VSS.n15979 0.0223919
R62599 VSS.n15985 VSS.n15983 0.0223919
R62600 VSS.n15983 VSS.n15981 0.0223919
R62601 VSS.n15582 VSS.n15581 0.0223919
R62602 VSS.n15581 VSS.n15579 0.0223919
R62603 VSS.n15268 VSS.n15262 0.0223919
R62604 VSS.n15268 VSS.n15266 0.0223919
R62605 VSS.n15266 VSS.n15264 0.0223919
R62606 VSS.n1557 VSS.n1553 0.0223919
R62607 VSS.n1557 VSS.n1555 0.0223919
R62608 VSS.n1563 VSS.n1559 0.0223919
R62609 VSS.n950 VSS.n944 0.0223919
R62610 VSS.n950 VSS.n949 0.0223919
R62611 VSS.n949 VSS.n947 0.0223919
R62612 VSS.n958 VSS.n952 0.0223919
R62613 VSS.n958 VSS.n957 0.0223919
R62614 VSS.n957 VSS.n955 0.0223919
R62615 VSS.n5650 VSS.n5648 0.0223919
R62616 VSS.n5648 VSS.n5647 0.0223919
R62617 VSS.n16047 VSS.n16031 0.0223919
R62618 VSS.n16047 VSS.n16045 0.0223919
R62619 VSS.n15301 VSS.n15299 0.0223919
R62620 VSS.n15305 VSS.n15301 0.0223919
R62621 VSS.n15305 VSS.n15303 0.0223919
R62622 VSS.n1614 VSS.n1612 0.0223919
R62623 VSS.n1622 VSS.n1614 0.0223919
R62624 VSS.n1622 VSS.n1621 0.0223919
R62625 VSS.n1010 VSS.n1006 0.0223919
R62626 VSS.n1010 VSS.n1009 0.0223919
R62627 VSS.n20915 VSS.n20913 0.0223919
R62628 VSS.n20917 VSS.n20915 0.0223919
R62629 VSS.n5495 VSS.n5493 0.0223919
R62630 VSS.n5499 VSS.n5495 0.0223919
R62631 VSS.n5499 VSS.n5498 0.0223919
R62632 VSS.n5481 VSS.n5479 0.0223919
R62633 VSS.n5489 VSS.n5481 0.0223919
R62634 VSS.n5489 VSS.n5488 0.0223919
R62635 VSS.n5488 VSS.n5486 0.0223919
R62636 VSS.n15989 VSS.n15987 0.0223919
R62637 VSS.n15995 VSS.n15989 0.0223919
R62638 VSS.n15995 VSS.n15994 0.0223919
R62639 VSS.n15994 VSS.n15992 0.0223919
R62640 VSS.n16001 VSS.n15997 0.0223919
R62641 VSS.n16001 VSS.n16000 0.0223919
R62642 VSS.n15274 VSS.n15270 0.0223919
R62643 VSS.n15274 VSS.n15272 0.0223919
R62644 VSS.n15278 VSS.n15276 0.0223919
R62645 VSS.n1574 VSS.n1570 0.0223919
R62646 VSS.n1574 VSS.n1572 0.0223919
R62647 VSS.n1580 VSS.n1576 0.0223919
R62648 VSS.n966 VSS.n960 0.0223919
R62649 VSS.n966 VSS.n964 0.0223919
R62650 VSS.n964 VSS.n962 0.0223919
R62651 VSS.n970 VSS.n968 0.0223919
R62652 VSS.n1307 VSS.n1303 0.0223919
R62653 VSS.n21180 VSS.n21178 0.0223919
R62654 VSS.n20892 VSS.n20891 0.0223919
R62655 VSS.n20877 VSS.n20875 0.0223919
R62656 VSS.n20888 VSS.n20877 0.0223919
R62657 VSS.n20888 VSS.n20887 0.0223919
R62658 VSS.n20887 VSS.n20885 0.0223919
R62659 VSS.n21322 VSS.n21321 0.0217598
R62660 VSS.n11642 VSS.n11641 0.0217598
R62661 VSS.n8526 VSS.n8525 0.0214155
R62662 VSS.n8344 VSS.n8343 0.0214155
R62663 VSS.n8677 VSS.n8676 0.0214155
R62664 VSS.n8140 VSS.n8139 0.0214155
R62665 VSS.n18488 VSS.n18476 0.0212042
R62666 VSS.n14575 VSS.n14574 0.0212042
R62667 VSS.n14820 VSS.n14819 0.0212042
R62668 VSS.n16699 VSS.n16698 0.0212042
R62669 VSS.n16448 VSS.n16447 0.0212042
R62670 VSS.n15861 VSS.n15860 0.0212042
R62671 VSS.n15347 VSS.n15346 0.0212042
R62672 VSS.n8467 VSS.n8466 0.0212042
R62673 VSS.n8549 VSS.n8548 0.0212042
R62674 VSS.n8315 VSS.n8314 0.0212042
R62675 VSS.n8404 VSS.n8403 0.0212042
R62676 VSS.n8373 VSS.n8372 0.0212042
R62677 VSS.n19562 VSS.n19561 0.0212042
R62678 VSS.n19753 VSS.n19752 0.0212042
R62679 VSS.n19843 VSS.n19842 0.0212042
R62680 VSS.n2101 VSS.n2100 0.0212042
R62681 VSS.n841 VSS.n840 0.0212042
R62682 VSS.n1939 VSS.n1938 0.0212042
R62683 VSS.n1663 VSS.n1662 0.0212042
R62684 VSS.n8618 VSS.n8617 0.0212042
R62685 VSS.n8700 VSS.n8699 0.0212042
R62686 VSS.n8111 VSS.n8110 0.0212042
R62687 VSS.n8212 VSS.n8211 0.0212042
R62688 VSS.n8181 VSS.n8180 0.0212042
R62689 VSS.n17198 VSS.n17197 0.0212
R62690 VSS.n5903 VSS.n5902 0.0211145
R62691 VSS.n18667 VSS.n18666 0.020993
R62692 VSS.n14470 VSS.n14460 0.020993
R62693 VSS.n14675 VSS.n14674 0.020993
R62694 VSS.n17161 VSS.n17160 0.020993
R62695 VSS.n16869 VSS.n16868 0.020993
R62696 VSS.n16680 VSS.n16679 0.020993
R62697 VSS.n15718 VSS.n15705 0.020993
R62698 VSS.n15346 VSS.n15345 0.020993
R62699 VSS.n8466 VSS.n8465 0.020993
R62700 VSS.n8548 VSS.n8547 0.020993
R62701 VSS.n8314 VSS.n8313 0.020993
R62702 VSS.n8403 VSS.n8402 0.020993
R62703 VSS.n8374 VSS.n8373 0.020993
R62704 VSS.n19536 VSS.n19535 0.020993
R62705 VSS.n19727 VSS.n19726 0.020993
R62706 VSS.n19781 VSS.n19771 0.020993
R62707 VSS.n19862 VSS.n19861 0.020993
R62708 VSS.n2127 VSS.n2126 0.020993
R62709 VSS.n752 VSS.n751 0.020993
R62710 VSS.n1965 VSS.n1964 0.020993
R62711 VSS.n1662 VSS.n1661 0.020993
R62712 VSS.n8617 VSS.n8616 0.020993
R62713 VSS.n8699 VSS.n8698 0.020993
R62714 VSS.n8110 VSS.n8109 0.020993
R62715 VSS.n8211 VSS.n8210 0.020993
R62716 VSS.n8182 VSS.n8181 0.020993
R62717 VSS.n16666 VSS.n16643 0.0207817
R62718 VSS.n754 VSS.n753 0.0207817
R62719 VSS.n5656 VSS.n5654 0.0207703
R62720 VSS.n5536 VSS.n5535 0.0207703
R62721 VSS.n16041 VSS.n16040 0.0207703
R62722 VSS.n1020 VSS.n1019 0.0207703
R62723 VSS.n20908 VSS.n20907 0.0207703
R62724 VSS.n20923 VSS.n20921 0.0207703
R62725 VSS.n17160 VSS.n17131 0.0205704
R62726 VSS.n19863 VSS.n19862 0.0205704
R62727 VSS.n16500 VSS.n14993 0.0203592
R62728 VSS.n830 VSS.n829 0.0203592
R62729 VSS.n331 VSS.n330 0.0203552
R62730 VSS.n20979 VSS.n20976 0.0201277
R62731 VSS.n15406 VSS.n15405 0.0199366
R62732 VSS.n1722 VSS.n1721 0.0199366
R62733 VSS.n15647 VSS.n15646 0.0198883
R62734 VSS.n15620 VSS.n15618 0.0198883
R62735 VSS.n15597 VSS.n15596 0.0198883
R62736 VSS.n5707 VSS.n5705 0.0198883
R62737 VSS.n15438 VSS.n15436 0.0198883
R62738 VSS.n4656 VSS.n4655 0.01985
R62739 VSS.n12222 VSS.n12221 0.0196339
R62740 VSS.n10170 VSS.n10169 0.0196339
R62741 VSS.n15464 VSS.n15463 0.0193028
R62742 VSS.n1766 VSS.n1765 0.0193028
R62743 VSS.n22230 VSS.n22229 0.0192235
R62744 VSS.n21986 VSS.n21985 0.0192235
R62745 VSS.n14253 VSS.n14251 0.0191871
R62746 VSS.n13631 VSS.n13629 0.0191871
R62747 VSS.n22175 VSS.n22161 0.0191871
R62748 VSS.n21978 VSS.n21967 0.0191871
R62749 VSS.n15374 VSS.n15373 0.0191189
R62750 VSS.n21229 VSS.n21227 0.0191034
R62751 VSS.n11258 VSS.n11257 0.0191034
R62752 VSS.n4014 VSS.n4013 0.0191024
R62753 VSS.n4018 VSS.n4017 0.0191024
R62754 VSS.n4029 VSS.n4028 0.0191024
R62755 VSS.n4036 VSS.n4035 0.0191024
R62756 VSS.n4040 VSS.n4039 0.0191024
R62757 VSS.n2348 VSS.n2347 0.0191024
R62758 VSS.n2352 VSS.n2351 0.0191024
R62759 VSS.n2359 VSS.n2358 0.0191024
R62760 VSS.n2370 VSS.n2369 0.0191024
R62761 VSS.n2374 VSS.n2373 0.0191024
R62762 VSS.n17321 VSS.n17320 0.0191024
R62763 VSS.n17317 VSS.n17316 0.0191024
R62764 VSS.n11526 VSS.n11525 0.0191024
R62765 VSS.n11530 VSS.n11529 0.0191024
R62766 VSS.n11534 VSS.n11533 0.0191024
R62767 VSS.n11541 VSS.n11540 0.0191024
R62768 VSS.n11545 VSS.n11544 0.0191024
R62769 VSS.n11554 VSS.n11553 0.0191024
R62770 VSS.n11558 VSS.n11557 0.0191024
R62771 VSS.n11562 VSS.n11561 0.0191024
R62772 VSS.n11568 VSS.n11567 0.0191024
R62773 VSS.n11572 VSS.n11571 0.0191024
R62774 VSS.n11581 VSS.n11580 0.0191024
R62775 VSS.n11585 VSS.n11584 0.0191024
R62776 VSS.n11339 VSS.n11338 0.0191024
R62777 VSS.n11343 VSS.n11342 0.0191024
R62778 VSS.n11354 VSS.n11353 0.0191024
R62779 VSS.n11358 VSS.n11357 0.0191024
R62780 VSS.n11365 VSS.n11364 0.0191024
R62781 VSS.n5858 VSS.n5857 0.0191024
R62782 VSS.n5854 VSS.n5853 0.0191024
R62783 VSS.n5735 VSS.n5734 0.0191024
R62784 VSS.n5728 VSS.n5727 0.0191024
R62785 VSS.n5597 VSS.n5596 0.0191024
R62786 VSS.n5593 VSS.n5592 0.0191024
R62787 VSS.n5589 VSS.n5588 0.0191024
R62788 VSS.n5582 VSS.n5581 0.0191024
R62789 VSS.n5578 VSS.n5577 0.0191024
R62790 VSS.n5542 VSS.n5541 0.0191024
R62791 VSS.n9478 VSS.n9477 0.0191024
R62792 VSS.n9487 VSS.n9486 0.0191024
R62793 VSS.n9491 VSS.n9490 0.0191024
R62794 VSS.n9546 VSS.n9545 0.0191024
R62795 VSS.n9593 VSS.n9592 0.0191024
R62796 VSS.n9589 VSS.n9588 0.0191024
R62797 VSS.n9585 VSS.n9584 0.0191024
R62798 VSS.n9578 VSS.n9577 0.0191024
R62799 VSS.n9574 VSS.n9573 0.0191024
R62800 VSS.n9565 VSS.n9564 0.0191024
R62801 VSS.n9561 VSS.n9560 0.0191024
R62802 VSS.n9019 VSS.n9018 0.0191024
R62803 VSS.n9028 VSS.n9027 0.0191024
R62804 VSS.n9032 VSS.n9031 0.0191024
R62805 VSS.n9043 VSS.n9042 0.0191024
R62806 VSS.n9047 VSS.n9046 0.0191024
R62807 VSS.n9156 VSS.n9155 0.0191024
R62808 VSS.n9152 VSS.n9151 0.0191024
R62809 VSS.n9148 VSS.n9147 0.0191024
R62810 VSS.n9141 VSS.n9140 0.0191024
R62811 VSS.n9137 VSS.n9136 0.0191024
R62812 VSS.n9128 VSS.n9127 0.0191024
R62813 VSS.n9124 VSS.n9123 0.0191024
R62814 VSS.n9114 VSS.n9113 0.0191024
R62815 VSS.n9110 VSS.n9109 0.0191024
R62816 VSS.n9101 VSS.n9100 0.0191024
R62817 VSS.n9097 VSS.n9096 0.0191024
R62818 VSS.n13039 VSS.n13038 0.0191024
R62819 VSS.n13043 VSS.n13042 0.0191024
R62820 VSS.n13056 VSS.n13055 0.0191024
R62821 VSS.n13065 VSS.n13064 0.0191024
R62822 VSS.n13069 VSS.n13068 0.0191024
R62823 VSS.n13156 VSS.n13155 0.0191024
R62824 VSS.n13160 VSS.n13159 0.0191024
R62825 VSS.n13169 VSS.n13168 0.0191024
R62826 VSS.n13182 VSS.n13181 0.0191024
R62827 VSS.n13186 VSS.n13185 0.0191024
R62828 VSS.n12989 VSS.n12988 0.0191024
R62829 VSS.n12985 VSS.n12984 0.0191024
R62830 VSS.n12978 VSS.n12977 0.0191024
R62831 VSS.n12974 VSS.n12973 0.0191024
R62832 VSS.n12970 VSS.n12969 0.0191024
R62833 VSS.n12961 VSS.n12960 0.0191024
R62834 VSS.n12957 VSS.n12956 0.0191024
R62835 VSS.n12948 VSS.n12947 0.0191024
R62836 VSS.n12944 VSS.n12943 0.0191024
R62837 VSS.n12931 VSS.n12930 0.0191024
R62838 VSS.n12927 VSS.n12926 0.0191024
R62839 VSS.n12918 VSS.n12917 0.0191024
R62840 VSS.n12914 VSS.n12913 0.0191024
R62841 VSS.n12870 VSS.n12869 0.0191024
R62842 VSS.n12866 VSS.n12865 0.0191024
R62843 VSS.n12855 VSS.n12854 0.0191024
R62844 VSS.n12851 VSS.n12850 0.0191024
R62845 VSS.n12842 VSS.n12841 0.0191024
R62846 VSS.n12807 VSS.n12806 0.0191024
R62847 VSS.n12803 VSS.n12802 0.0191024
R62848 VSS.n12792 VSS.n12791 0.0191024
R62849 VSS.n12788 VSS.n12787 0.0191024
R62850 VSS.n12779 VSS.n12778 0.0191024
R62851 VSS.n12771 VSS.n12770 0.0191024
R62852 VSS.n12767 VSS.n12766 0.0191024
R62853 VSS.n12760 VSS.n12759 0.0191024
R62854 VSS.n12756 VSS.n12755 0.0191024
R62855 VSS.n12752 VSS.n12751 0.0191024
R62856 VSS.n12743 VSS.n12742 0.0191024
R62857 VSS.n12739 VSS.n12738 0.0191024
R62858 VSS.n12730 VSS.n12729 0.0191024
R62859 VSS.n12726 VSS.n12725 0.0191024
R62860 VSS.n12714 VSS.n12713 0.0191024
R62861 VSS.n12710 VSS.n12709 0.0191024
R62862 VSS.n12701 VSS.n12700 0.0191024
R62863 VSS.n12697 VSS.n12696 0.0191024
R62864 VSS.n18885 VSS.n18884 0.0191024
R62865 VSS.n18889 VSS.n18888 0.0191024
R62866 VSS.n18900 VSS.n18899 0.0191024
R62867 VSS.n18907 VSS.n18906 0.0191024
R62868 VSS.n18911 VSS.n18910 0.0191024
R62869 VSS.n2247 VSS.n2246 0.0191024
R62870 VSS.n2251 VSS.n2250 0.0191024
R62871 VSS.n2258 VSS.n2257 0.0191024
R62872 VSS.n2269 VSS.n2268 0.0191024
R62873 VSS.n2273 VSS.n2272 0.0191024
R62874 VSS.n14413 VSS.n14412 0.0191024
R62875 VSS.n14409 VSS.n14408 0.0191024
R62876 VSS.n15000 VSS.n14999 0.0191024
R62877 VSS.n15004 VSS.n15003 0.0191024
R62878 VSS.n15008 VSS.n15007 0.0191024
R62879 VSS.n15015 VSS.n15014 0.0191024
R62880 VSS.n15019 VSS.n15018 0.0191024
R62881 VSS.n15028 VSS.n15027 0.0191024
R62882 VSS.n15032 VSS.n15031 0.0191024
R62883 VSS.n15043 VSS.n15042 0.0191024
R62884 VSS.n15047 VSS.n15046 0.0191024
R62885 VSS.n15056 VSS.n15055 0.0191024
R62886 VSS.n15060 VSS.n15059 0.0191024
R62887 VSS.n15140 VSS.n15139 0.0191024
R62888 VSS.n15144 VSS.n15143 0.0191024
R62889 VSS.n15155 VSS.n15154 0.0191024
R62890 VSS.n15159 VSS.n15158 0.0191024
R62891 VSS.n15166 VSS.n15165 0.0191024
R62892 VSS.n16219 VSS.n16218 0.0191024
R62893 VSS.n16215 VSS.n16214 0.0191024
R62894 VSS.n16183 VSS.n16182 0.0191024
R62895 VSS.n16176 VSS.n16175 0.0191024
R62896 VSS.n16113 VSS.n16112 0.0191024
R62897 VSS.n16109 VSS.n16108 0.0191024
R62898 VSS.n16105 VSS.n16104 0.0191024
R62899 VSS.n16098 VSS.n16097 0.0191024
R62900 VSS.n16094 VSS.n16093 0.0191024
R62901 VSS.n16052 VSS.n16051 0.0191024
R62902 VSS.n9604 VSS.n9603 0.0191024
R62903 VSS.n9608 VSS.n9607 0.0191024
R62904 VSS.n9663 VSS.n9662 0.0191024
R62905 VSS.n9710 VSS.n9709 0.0191024
R62906 VSS.n9706 VSS.n9705 0.0191024
R62907 VSS.n9702 VSS.n9701 0.0191024
R62908 VSS.n9695 VSS.n9694 0.0191024
R62909 VSS.n9691 VSS.n9690 0.0191024
R62910 VSS.n9682 VSS.n9681 0.0191024
R62911 VSS.n9678 VSS.n9677 0.0191024
R62912 VSS.n9162 VSS.n9161 0.0191024
R62913 VSS.n9171 VSS.n9170 0.0191024
R62914 VSS.n9175 VSS.n9174 0.0191024
R62915 VSS.n9186 VSS.n9185 0.0191024
R62916 VSS.n9190 VSS.n9189 0.0191024
R62917 VSS.n9319 VSS.n9318 0.0191024
R62918 VSS.n9315 VSS.n9314 0.0191024
R62919 VSS.n9311 VSS.n9310 0.0191024
R62920 VSS.n9304 VSS.n9303 0.0191024
R62921 VSS.n9300 VSS.n9299 0.0191024
R62922 VSS.n9291 VSS.n9290 0.0191024
R62923 VSS.n9287 VSS.n9286 0.0191024
R62924 VSS.n9277 VSS.n9276 0.0191024
R62925 VSS.n9273 VSS.n9272 0.0191024
R62926 VSS.n9264 VSS.n9263 0.0191024
R62927 VSS.n9260 VSS.n9259 0.0191024
R62928 VSS.n21812 VSS.n21811 0.0191024
R62929 VSS.n21816 VSS.n21815 0.0191024
R62930 VSS.n21829 VSS.n21828 0.0191024
R62931 VSS.n21838 VSS.n21837 0.0191024
R62932 VSS.n21842 VSS.n21841 0.0191024
R62933 VSS.n2296 VSS.n2295 0.0191024
R62934 VSS.n2300 VSS.n2299 0.0191024
R62935 VSS.n2309 VSS.n2308 0.0191024
R62936 VSS.n2322 VSS.n2321 0.0191024
R62937 VSS.n2326 VSS.n2325 0.0191024
R62938 VSS.n20595 VSS.n20594 0.0191024
R62939 VSS.n20599 VSS.n20598 0.0191024
R62940 VSS.n20606 VSS.n20605 0.0191024
R62941 VSS.n20610 VSS.n20609 0.0191024
R62942 VSS.n20614 VSS.n20613 0.0191024
R62943 VSS.n20623 VSS.n20622 0.0191024
R62944 VSS.n20627 VSS.n20626 0.0191024
R62945 VSS.n20636 VSS.n20635 0.0191024
R62946 VSS.n20640 VSS.n20639 0.0191024
R62947 VSS.n20653 VSS.n20652 0.0191024
R62948 VSS.n20657 VSS.n20656 0.0191024
R62949 VSS.n20666 VSS.n20665 0.0191024
R62950 VSS.n20670 VSS.n20669 0.0191024
R62951 VSS.n20790 VSS.n20789 0.0191024
R62952 VSS.n20794 VSS.n20793 0.0191024
R62953 VSS.n20805 VSS.n20804 0.0191024
R62954 VSS.n20809 VSS.n20808 0.0191024
R62955 VSS.n20818 VSS.n20817 0.0191024
R62956 VSS.n21161 VSS.n21160 0.0191024
R62957 VSS.n21157 VSS.n21156 0.0191024
R62958 VSS.n21125 VSS.n21124 0.0191024
R62959 VSS.n21116 VSS.n21115 0.0191024
R62960 VSS.n21047 VSS.n21046 0.0191024
R62961 VSS.n21043 VSS.n21042 0.0191024
R62962 VSS.n21039 VSS.n21038 0.0191024
R62963 VSS.n21030 VSS.n21029 0.0191024
R62964 VSS.n21026 VSS.n21025 0.0191024
R62965 VSS.n6909 VSS.n6908 0.0191024
R62966 VSS.n6918 VSS.n6917 0.0191024
R62967 VSS.n6922 VSS.n6921 0.0191024
R62968 VSS.n6953 VSS.n6952 0.0191024
R62969 VSS.n7005 VSS.n7004 0.0191024
R62970 VSS.n7001 VSS.n7000 0.0191024
R62971 VSS.n6997 VSS.n6996 0.0191024
R62972 VSS.n6988 VSS.n6987 0.0191024
R62973 VSS.n6984 VSS.n6983 0.0191024
R62974 VSS.n6975 VSS.n6974 0.0191024
R62975 VSS.n6971 VSS.n6970 0.0191024
R62976 VSS.n6650 VSS.n6649 0.0191024
R62977 VSS.n6659 VSS.n6658 0.0191024
R62978 VSS.n6663 VSS.n6662 0.0191024
R62979 VSS.n6676 VSS.n6675 0.0191024
R62980 VSS.n6680 VSS.n6679 0.0191024
R62981 VSS.n6645 VSS.n6644 0.0191024
R62982 VSS.n6641 VSS.n6640 0.0191024
R62983 VSS.n6637 VSS.n6636 0.0191024
R62984 VSS.n6628 VSS.n6627 0.0191024
R62985 VSS.n6624 VSS.n6623 0.0191024
R62986 VSS.n6615 VSS.n6614 0.0191024
R62987 VSS.n6611 VSS.n6610 0.0191024
R62988 VSS.n6598 VSS.n6597 0.0191024
R62989 VSS.n6594 VSS.n6593 0.0191024
R62990 VSS.n6585 VSS.n6584 0.0191024
R62991 VSS.n6581 VSS.n6580 0.0191024
R62992 VSS.n19097 VSS.n19096 0.0191024
R62993 VSS.n19101 VSS.n19100 0.0191024
R62994 VSS.n19114 VSS.n19113 0.0191024
R62995 VSS.n19123 VSS.n19122 0.0191024
R62996 VSS.n19127 VSS.n19126 0.0191024
R62997 VSS.n17904 VSS.n17903 0.0191024
R62998 VSS.n17908 VSS.n17907 0.0191024
R62999 VSS.n17917 VSS.n17916 0.0191024
R63000 VSS.n17930 VSS.n17929 0.0191024
R63001 VSS.n17934 VSS.n17933 0.0191024
R63002 VSS.n20157 VSS.n20156 0.0191024
R63003 VSS.n20161 VSS.n20160 0.0191024
R63004 VSS.n20143 VSS.n20142 0.0191024
R63005 VSS.n20139 VSS.n20138 0.0191024
R63006 VSS.n20135 VSS.n20134 0.0191024
R63007 VSS.n20126 VSS.n20125 0.0191024
R63008 VSS.n20122 VSS.n20121 0.0191024
R63009 VSS.n20113 VSS.n20112 0.0191024
R63010 VSS.n20109 VSS.n20108 0.0191024
R63011 VSS.n20096 VSS.n20095 0.0191024
R63012 VSS.n20092 VSS.n20091 0.0191024
R63013 VSS.n20083 VSS.n20082 0.0191024
R63014 VSS.n20079 VSS.n20078 0.0191024
R63015 VSS.n2029 VSS.n2028 0.0191024
R63016 VSS.n2025 VSS.n2024 0.0191024
R63017 VSS.n2014 VSS.n2013 0.0191024
R63018 VSS.n2010 VSS.n2009 0.0191024
R63019 VSS.n2001 VSS.n2000 0.0191024
R63020 VSS.n1290 VSS.n1289 0.0191024
R63021 VSS.n1286 VSS.n1285 0.0191024
R63022 VSS.n1175 VSS.n1174 0.0191024
R63023 VSS.n1166 VSS.n1165 0.0191024
R63024 VSS.n1093 VSS.n1092 0.0191024
R63025 VSS.n1089 VSS.n1088 0.0191024
R63026 VSS.n1085 VSS.n1084 0.0191024
R63027 VSS.n1076 VSS.n1075 0.0191024
R63028 VSS.n1072 VSS.n1071 0.0191024
R63029 VSS.n1026 VSS.n1025 0.0191024
R63030 VSS.n6786 VSS.n6785 0.0191024
R63031 VSS.n6795 VSS.n6794 0.0191024
R63032 VSS.n6799 VSS.n6798 0.0191024
R63033 VSS.n6851 VSS.n6850 0.0191024
R63034 VSS.n6903 VSS.n6902 0.0191024
R63035 VSS.n6899 VSS.n6898 0.0191024
R63036 VSS.n6895 VSS.n6894 0.0191024
R63037 VSS.n6886 VSS.n6885 0.0191024
R63038 VSS.n6882 VSS.n6881 0.0191024
R63039 VSS.n6873 VSS.n6872 0.0191024
R63040 VSS.n6869 VSS.n6868 0.0191024
R63041 VSS.n6500 VSS.n6499 0.0191024
R63042 VSS.n6509 VSS.n6508 0.0191024
R63043 VSS.n6513 VSS.n6512 0.0191024
R63044 VSS.n6526 VSS.n6525 0.0191024
R63045 VSS.n6530 VSS.n6529 0.0191024
R63046 VSS.n6495 VSS.n6494 0.0191024
R63047 VSS.n6491 VSS.n6490 0.0191024
R63048 VSS.n6487 VSS.n6486 0.0191024
R63049 VSS.n6478 VSS.n6477 0.0191024
R63050 VSS.n6474 VSS.n6473 0.0191024
R63051 VSS.n6465 VSS.n6464 0.0191024
R63052 VSS.n6461 VSS.n6460 0.0191024
R63053 VSS.n6448 VSS.n6447 0.0191024
R63054 VSS.n6444 VSS.n6443 0.0191024
R63055 VSS.n6435 VSS.n6434 0.0191024
R63056 VSS.n6431 VSS.n6430 0.0191024
R63057 VSS.n21583 VSS.n21582 0.0191024
R63058 VSS.n21587 VSS.n21586 0.0191024
R63059 VSS.n21600 VSS.n21599 0.0191024
R63060 VSS.n21609 VSS.n21608 0.0191024
R63061 VSS.n21613 VSS.n21612 0.0191024
R63062 VSS.n21517 VSS.n21516 0.0191024
R63063 VSS.n21513 VSS.n21512 0.0191024
R63064 VSS.n21504 VSS.n21503 0.0191024
R63065 VSS.n21491 VSS.n21490 0.0191024
R63066 VSS.n21487 VSS.n21486 0.0191024
R63067 VSS.n21406 VSS.n21405 0.0191024
R63068 VSS.n21402 VSS.n21401 0.0191024
R63069 VSS.n21395 VSS.n21394 0.0191024
R63070 VSS.n21391 VSS.n21390 0.0191024
R63071 VSS.n21387 VSS.n21386 0.0191024
R63072 VSS.n21378 VSS.n21377 0.0191024
R63073 VSS.n21374 VSS.n21373 0.0191024
R63074 VSS.n21365 VSS.n21364 0.0191024
R63075 VSS.n21361 VSS.n21360 0.0191024
R63076 VSS.n21348 VSS.n21347 0.0191024
R63077 VSS.n21344 VSS.n21343 0.0191024
R63078 VSS.n21335 VSS.n21334 0.0191024
R63079 VSS.n21331 VSS.n21330 0.0191024
R63080 VSS.n21291 VSS.n21290 0.0191024
R63081 VSS.n21287 VSS.n21286 0.0191024
R63082 VSS.n21276 VSS.n21275 0.0191024
R63083 VSS.n21272 VSS.n21271 0.0191024
R63084 VSS.n21263 VSS.n21262 0.0191024
R63085 VSS.n7555 VSS.n7554 0.0191024
R63086 VSS.n7559 VSS.n7558 0.0191024
R63087 VSS.n7570 VSS.n7569 0.0191024
R63088 VSS.n7574 VSS.n7573 0.0191024
R63089 VSS.n7583 VSS.n7582 0.0191024
R63090 VSS.n7591 VSS.n7590 0.0191024
R63091 VSS.n7595 VSS.n7594 0.0191024
R63092 VSS.n7602 VSS.n7601 0.0191024
R63093 VSS.n7606 VSS.n7605 0.0191024
R63094 VSS.n7610 VSS.n7609 0.0191024
R63095 VSS.n7619 VSS.n7618 0.0191024
R63096 VSS.n7623 VSS.n7622 0.0191024
R63097 VSS.n7632 VSS.n7631 0.0191024
R63098 VSS.n7636 VSS.n7635 0.0191024
R63099 VSS.n7649 VSS.n7648 0.0191024
R63100 VSS.n7653 VSS.n7652 0.0191024
R63101 VSS.n7662 VSS.n7661 0.0191024
R63102 VSS.n7666 VSS.n7665 0.0191024
R63103 VSS.n7679 VSS.n7678 0.0191024
R63104 VSS.n7683 VSS.n7682 0.0191024
R63105 VSS.n7690 VSS.n7689 0.0191024
R63106 VSS.n7694 VSS.n7693 0.0191024
R63107 VSS.n7698 VSS.n7697 0.0191024
R63108 VSS.n7707 VSS.n7706 0.0191024
R63109 VSS.n7711 VSS.n7710 0.0191024
R63110 VSS.n7720 VSS.n7719 0.0191024
R63111 VSS.n7724 VSS.n7723 0.0191024
R63112 VSS.n7737 VSS.n7736 0.0191024
R63113 VSS.n7741 VSS.n7740 0.0191024
R63114 VSS.n7750 VSS.n7749 0.0191024
R63115 VSS.n7754 VSS.n7753 0.0191024
R63116 VSS.n7767 VSS.n7766 0.0191024
R63117 VSS.n7771 VSS.n7770 0.0191024
R63118 VSS.n7849 VSS.n7848 0.0191024
R63119 VSS.n7845 VSS.n7844 0.0191024
R63120 VSS.n7841 VSS.n7840 0.0191024
R63121 VSS.n7832 VSS.n7831 0.0191024
R63122 VSS.n7828 VSS.n7827 0.0191024
R63123 VSS.n7819 VSS.n7818 0.0191024
R63124 VSS.n7815 VSS.n7814 0.0191024
R63125 VSS.n7802 VSS.n7801 0.0191024
R63126 VSS.n7798 VSS.n7797 0.0191024
R63127 VSS.n7789 VSS.n7788 0.0191024
R63128 VSS.n7785 VSS.n7784 0.0191024
R63129 VSS.n3816 VSS.n3815 0.0191024
R63130 VSS.n3820 VSS.n3819 0.0191024
R63131 VSS.n3831 VSS.n3830 0.0191024
R63132 VSS.n3838 VSS.n3837 0.0191024
R63133 VSS.n3842 VSS.n3841 0.0191024
R63134 VSS.n4701 VSS.n4700 0.0191024
R63135 VSS.n4705 VSS.n4704 0.0191024
R63136 VSS.n4712 VSS.n4711 0.0191024
R63137 VSS.n4723 VSS.n4722 0.0191024
R63138 VSS.n4727 VSS.n4726 0.0191024
R63139 VSS.n11731 VSS.n11730 0.0191024
R63140 VSS.n11727 VSS.n11726 0.0191024
R63141 VSS.n11709 VSS.n11708 0.0191024
R63142 VSS.n11705 VSS.n11704 0.0191024
R63143 VSS.n11701 VSS.n11700 0.0191024
R63144 VSS.n11694 VSS.n11693 0.0191024
R63145 VSS.n11690 VSS.n11689 0.0191024
R63146 VSS.n11681 VSS.n11680 0.0191024
R63147 VSS.n11677 VSS.n11676 0.0191024
R63148 VSS.n11666 VSS.n11665 0.0191024
R63149 VSS.n11662 VSS.n11661 0.0191024
R63150 VSS.n11653 VSS.n11652 0.0191024
R63151 VSS.n11649 VSS.n11648 0.0191024
R63152 VSS.n11449 VSS.n11448 0.0191024
R63153 VSS.n11445 VSS.n11444 0.0191024
R63154 VSS.n11434 VSS.n11433 0.0191024
R63155 VSS.n11430 VSS.n11429 0.0191024
R63156 VSS.n11423 VSS.n11422 0.0191024
R63157 VSS.n11228 VSS.n11227 0.0191024
R63158 VSS.n11224 VSS.n11223 0.0191024
R63159 VSS.n11213 VSS.n11212 0.0191024
R63160 VSS.n11209 VSS.n11208 0.0191024
R63161 VSS.n11202 VSS.n11201 0.0191024
R63162 VSS.n11194 VSS.n11193 0.0191024
R63163 VSS.n11190 VSS.n11189 0.0191024
R63164 VSS.n6152 VSS.n6151 0.0191024
R63165 VSS.n6148 VSS.n6147 0.0191024
R63166 VSS.n6144 VSS.n6143 0.0191024
R63167 VSS.n6137 VSS.n6136 0.0191024
R63168 VSS.n6133 VSS.n6132 0.0191024
R63169 VSS.n6124 VSS.n6123 0.0191024
R63170 VSS.n6120 VSS.n6119 0.0191024
R63171 VSS.n6110 VSS.n6109 0.0191024
R63172 VSS.n6106 VSS.n6105 0.0191024
R63173 VSS.n6097 VSS.n6096 0.0191024
R63174 VSS.n6093 VSS.n6092 0.0191024
R63175 VSS.n6082 VSS.n6081 0.0191024
R63176 VSS.n6078 VSS.n6077 0.0191024
R63177 VSS.n6071 VSS.n6070 0.0191024
R63178 VSS.n6067 VSS.n6066 0.0191024
R63179 VSS.n6063 VSS.n6062 0.0191024
R63180 VSS.n6056 VSS.n6055 0.0191024
R63181 VSS.n6052 VSS.n6051 0.0191024
R63182 VSS.n6043 VSS.n6042 0.0191024
R63183 VSS.n6039 VSS.n6038 0.0191024
R63184 VSS.n6029 VSS.n6028 0.0191024
R63185 VSS.n6025 VSS.n6024 0.0191024
R63186 VSS.n6016 VSS.n6015 0.0191024
R63187 VSS.n6012 VSS.n6011 0.0191024
R63188 VSS.n6001 VSS.n6000 0.0191024
R63189 VSS.n5997 VSS.n5996 0.0191024
R63190 VSS.n5990 VSS.n5989 0.0191024
R63191 VSS.n5986 VSS.n5985 0.0191024
R63192 VSS.n5982 VSS.n5981 0.0191024
R63193 VSS.n5975 VSS.n5974 0.0191024
R63194 VSS.n5971 VSS.n5970 0.0191024
R63195 VSS.n5962 VSS.n5961 0.0191024
R63196 VSS.n5958 VSS.n5957 0.0191024
R63197 VSS.n5948 VSS.n5947 0.0191024
R63198 VSS.n5944 VSS.n5943 0.0191024
R63199 VSS.n5935 VSS.n5934 0.0191024
R63200 VSS.n5931 VSS.n5930 0.0191024
R63201 VSS.n3255 VSS.n3254 0.0191024
R63202 VSS.n3251 VSS.n3250 0.0191024
R63203 VSS.n2646 VSS.n2645 0.0191024
R63204 VSS.n2653 VSS.n2652 0.0191024
R63205 VSS.n2657 VSS.n2656 0.0191024
R63206 VSS.n671 VSS.n670 0.0191024
R63207 VSS.n675 VSS.n674 0.0191024
R63208 VSS.n666 VSS.n665 0.0191024
R63209 VSS.n662 VSS.n661 0.0191024
R63210 VSS.n658 VSS.n657 0.0191024
R63211 VSS.n651 VSS.n650 0.0191024
R63212 VSS.n647 VSS.n646 0.0191024
R63213 VSS.n638 VSS.n637 0.0191024
R63214 VSS.n634 VSS.n633 0.0191024
R63215 VSS.n624 VSS.n623 0.0191024
R63216 VSS.n620 VSS.n619 0.0191024
R63217 VSS.n611 VSS.n610 0.0191024
R63218 VSS.n607 VSS.n606 0.0191024
R63219 VSS.n567 VSS.n566 0.0191024
R63220 VSS.n563 VSS.n562 0.0191024
R63221 VSS.n552 VSS.n551 0.0191024
R63222 VSS.n548 VSS.n547 0.0191024
R63223 VSS.n541 VSS.n540 0.0191024
R63224 VSS.n508 VSS.n507 0.0191024
R63225 VSS.n504 VSS.n503 0.0191024
R63226 VSS.n493 VSS.n492 0.0191024
R63227 VSS.n489 VSS.n488 0.0191024
R63228 VSS.n482 VSS.n481 0.0191024
R63229 VSS.n474 VSS.n473 0.0191024
R63230 VSS.n470 VSS.n469 0.0191024
R63231 VSS.n10624 VSS.n10623 0.0191024
R63232 VSS.n10620 VSS.n10619 0.0191024
R63233 VSS.n10616 VSS.n10615 0.0191024
R63234 VSS.n10609 VSS.n10608 0.0191024
R63235 VSS.n10605 VSS.n10604 0.0191024
R63236 VSS.n10596 VSS.n10595 0.0191024
R63237 VSS.n10592 VSS.n10591 0.0191024
R63238 VSS.n10582 VSS.n10581 0.0191024
R63239 VSS.n10578 VSS.n10577 0.0191024
R63240 VSS.n10569 VSS.n10568 0.0191024
R63241 VSS.n10565 VSS.n10564 0.0191024
R63242 VSS.n18773 VSS.n18772 0.0190915
R63243 VSS.n16885 VSS.n16884 0.0190915
R63244 VSS.n19445 VSS.n19444 0.0190915
R63245 VSS.n20031 VSS.n20030 0.0190915
R63246 VSS.n16443 VSS.n16442 0.0190636
R63247 VSS.n19758 VSS.n19757 0.0190636
R63248 VSS.n19848 VSS.n19847 0.0190636
R63249 VSS.n20033 VSS.n20032 0.0190636
R63250 VSS.n2096 VSS.n2095 0.0190636
R63251 VSS.n2378 VSS.n2377 0.0189252
R63252 VSS.n11347 VSS.n11346 0.0189252
R63253 VSS.n13190 VSS.n13189 0.0189252
R63254 VSS.n12862 VSS.n12861 0.0189252
R63255 VSS.n12799 VSS.n12798 0.0189252
R63256 VSS.n2277 VSS.n2276 0.0189252
R63257 VSS.n15148 VSS.n15147 0.0189252
R63258 VSS.n2330 VSS.n2329 0.0189252
R63259 VSS.n20798 VSS.n20797 0.0189252
R63260 VSS.n17938 VSS.n17937 0.0189252
R63261 VSS.n2021 VSS.n2020 0.0189252
R63262 VSS.n21483 VSS.n21482 0.0189252
R63263 VSS.n21283 VSS.n21282 0.0189252
R63264 VSS.n7563 VSS.n7562 0.0189252
R63265 VSS.n4731 VSS.n4730 0.0189252
R63266 VSS.n11441 VSS.n11440 0.0189252
R63267 VSS.n11220 VSS.n11219 0.0189252
R63268 VSS.n559 VSS.n558 0.0189252
R63269 VSS.n500 VSS.n499 0.0189252
R63270 VSS.n203 VSS.n202 0.018852
R63271 VSS.n8351 VSS.n8350 0.0187841
R63272 VSS.n8159 VSS.n8158 0.0187841
R63273 VSS.n18208 VSS.n18207 0.018669
R63274 VSS.n15534 VSS.n15533 0.018669
R63275 VSS.n19648 VSS.n19647 0.018669
R63276 VSS.n1822 VSS.n1821 0.018669
R63277 VSS.n15325 VSS.n15324 0.0184577
R63278 VSS.n1641 VSS.n1640 0.0184577
R63279 VSS.n1690 VSS.n1689 0.0184525
R63280 VSS.n14570 VSS.n14569 0.0183973
R63281 VSS.n14825 VSS.n14824 0.0183973
R63282 VSS.n16883 VSS.n16882 0.0183973
R63283 VSS.n16694 VSS.n16693 0.0183973
R63284 VSS.n8347 VSS.n8346 0.0183973
R63285 VSS.n8149 VSS.n8148 0.0183973
R63286 VSS.n846 VSS.n845 0.0183973
R63287 VSS.n8156 VSS.n8149 0.0183973
R63288 VSS.n8348 VSS.n8347 0.0183973
R63289 VSS.n4010 VSS.n4009 0.0183937
R63290 VSS.n13035 VSS.n13034 0.0183937
R63291 VSS.n18881 VSS.n18880 0.0183937
R63292 VSS.n21808 VSS.n21807 0.0183937
R63293 VSS.n19093 VSS.n19092 0.0183937
R63294 VSS.n21579 VSS.n21578 0.0183937
R63295 VSS.n3812 VSS.n3811 0.0183937
R63296 VSS.n3259 VSS.n3258 0.0183937
R63297 VSS.n18815 VSS.n18814 0.0182575
R63298 VSS.n19487 VSS.n19486 0.0182575
R63299 VSS.n18391 VSS.n18390 0.0182465
R63300 VSS.n19631 VSS.n19630 0.0182465
R63301 VSS.n2344 VSS.n2343 0.0182165
R63302 VSS.n11350 VSS.n11349 0.0182165
R63303 VSS.n13152 VSS.n13151 0.0182165
R63304 VSS.n12859 VSS.n12858 0.0182165
R63305 VSS.n12796 VSS.n12795 0.0182165
R63306 VSS.n2243 VSS.n2242 0.0182165
R63307 VSS.n15151 VSS.n15150 0.0182165
R63308 VSS.n2292 VSS.n2291 0.0182165
R63309 VSS.n20801 VSS.n20800 0.0182165
R63310 VSS.n17900 VSS.n17899 0.0182165
R63311 VSS.n2018 VSS.n2017 0.0182165
R63312 VSS.n21521 VSS.n21520 0.0182165
R63313 VSS.n21280 VSS.n21279 0.0182165
R63314 VSS.n7566 VSS.n7565 0.0182165
R63315 VSS.n4697 VSS.n4696 0.0182165
R63316 VSS.n11438 VSS.n11437 0.0182165
R63317 VSS.n11217 VSS.n11216 0.0182165
R63318 VSS.n556 VSS.n555 0.0182165
R63319 VSS.n497 VSS.n496 0.0182165
R63320 VSS.n4044 VSS.n4043 0.0180394
R63321 VSS.n17313 VSS.n17312 0.0180394
R63322 VSS.n9550 VSS.n9549 0.0180394
R63323 VSS.n9051 VSS.n9050 0.0180394
R63324 VSS.n13073 VSS.n13072 0.0180394
R63325 VSS.n12981 VSS.n12980 0.0180394
R63326 VSS.n12763 VSS.n12762 0.0180394
R63327 VSS.n18915 VSS.n18914 0.0180394
R63328 VSS.n14405 VSS.n14404 0.0180394
R63329 VSS.n9667 VSS.n9666 0.0180394
R63330 VSS.n9194 VSS.n9193 0.0180394
R63331 VSS.n21846 VSS.n21845 0.0180394
R63332 VSS.n20603 VSS.n20602 0.0180394
R63333 VSS.n6957 VSS.n6956 0.0180394
R63334 VSS.n6684 VSS.n6683 0.0180394
R63335 VSS.n19131 VSS.n19130 0.0180394
R63336 VSS.n20165 VSS.n20164 0.0180394
R63337 VSS.n6855 VSS.n6854 0.0180394
R63338 VSS.n6534 VSS.n6533 0.0180394
R63339 VSS.n21617 VSS.n21616 0.0180394
R63340 VSS.n21398 VSS.n21397 0.0180394
R63341 VSS.n7599 VSS.n7598 0.0180394
R63342 VSS.n7687 VSS.n7686 0.0180394
R63343 VSS.n7775 VSS.n7774 0.0180394
R63344 VSS.n3846 VSS.n3845 0.0180394
R63345 VSS.n11723 VSS.n11722 0.0180394
R63346 VSS.n11186 VSS.n11185 0.0180394
R63347 VSS.n6074 VSS.n6073 0.0180394
R63348 VSS.n5993 VSS.n5992 0.0180394
R63349 VSS.n2661 VSS.n2660 0.0180394
R63350 VSS.n679 VSS.n678 0.0180394
R63351 VSS.n466 VSS.n465 0.0180394
R63352 VSS.n18756 VSS.n18755 0.0180352
R63353 VSS.n19279 VSS.n19237 0.0180352
R63354 VSS.n15295 VSS.n15294 0.0179734
R63355 VSS.n15510 VSS.n15509 0.0179734
R63356 VSS.n11549 VSS.n11548 0.0178622
R63357 VSS.n11577 VSS.n11576 0.0178622
R63358 VSS.n5574 VSS.n5573 0.0178622
R63359 VSS.n9483 VSS.n9482 0.0178622
R63360 VSS.n9570 VSS.n9569 0.0178622
R63361 VSS.n9024 VSS.n9023 0.0178622
R63362 VSS.n9133 VSS.n9132 0.0178622
R63363 VSS.n9105 VSS.n9104 0.0178622
R63364 VSS.n12953 VSS.n12952 0.0178622
R63365 VSS.n12922 VSS.n12921 0.0178622
R63366 VSS.n12735 VSS.n12734 0.0178622
R63367 VSS.n12705 VSS.n12704 0.0178622
R63368 VSS.n15023 VSS.n15022 0.0178622
R63369 VSS.n15052 VSS.n15051 0.0178622
R63370 VSS.n16090 VSS.n16089 0.0178622
R63371 VSS.n9600 VSS.n9599 0.0178622
R63372 VSS.n9687 VSS.n9686 0.0178622
R63373 VSS.n9167 VSS.n9166 0.0178622
R63374 VSS.n9296 VSS.n9295 0.0178622
R63375 VSS.n9268 VSS.n9267 0.0178622
R63376 VSS.n20631 VSS.n20630 0.0178622
R63377 VSS.n20662 VSS.n20661 0.0178622
R63378 VSS.n21022 VSS.n21021 0.0178622
R63379 VSS.n6914 VSS.n6913 0.0178622
R63380 VSS.n6980 VSS.n6979 0.0178622
R63381 VSS.n6655 VSS.n6654 0.0178622
R63382 VSS.n6620 VSS.n6619 0.0178622
R63383 VSS.n6589 VSS.n6588 0.0178622
R63384 VSS.n20118 VSS.n20117 0.0178622
R63385 VSS.n20087 VSS.n20086 0.0178622
R63386 VSS.n1068 VSS.n1067 0.0178622
R63387 VSS.n6791 VSS.n6790 0.0178622
R63388 VSS.n6878 VSS.n6877 0.0178622
R63389 VSS.n6505 VSS.n6504 0.0178622
R63390 VSS.n6470 VSS.n6469 0.0178622
R63391 VSS.n6439 VSS.n6438 0.0178622
R63392 VSS.n21370 VSS.n21369 0.0178622
R63393 VSS.n21339 VSS.n21338 0.0178622
R63394 VSS.n7627 VSS.n7626 0.0178622
R63395 VSS.n7658 VSS.n7657 0.0178622
R63396 VSS.n7715 VSS.n7714 0.0178622
R63397 VSS.n7746 VSS.n7745 0.0178622
R63398 VSS.n7824 VSS.n7823 0.0178622
R63399 VSS.n7793 VSS.n7792 0.0178622
R63400 VSS.n11686 VSS.n11685 0.0178622
R63401 VSS.n11657 VSS.n11656 0.0178622
R63402 VSS.n6129 VSS.n6128 0.0178622
R63403 VSS.n6101 VSS.n6100 0.0178622
R63404 VSS.n6048 VSS.n6047 0.0178622
R63405 VSS.n6020 VSS.n6019 0.0178622
R63406 VSS.n5967 VSS.n5966 0.0178622
R63407 VSS.n5939 VSS.n5938 0.0178622
R63408 VSS.n643 VSS.n642 0.0178622
R63409 VSS.n615 VSS.n614 0.0178622
R63410 VSS.n10601 VSS.n10600 0.0178622
R63411 VSS.n10573 VSS.n10572 0.0178622
R63412 VSS.n11550 VSS.n11549 0.017685
R63413 VSS.n11576 VSS.n11575 0.017685
R63414 VSS.n5573 VSS.n5572 0.017685
R63415 VSS.n9482 VSS.n9481 0.017685
R63416 VSS.n9569 VSS.n9568 0.017685
R63417 VSS.n9023 VSS.n9022 0.017685
R63418 VSS.n9132 VSS.n9131 0.017685
R63419 VSS.n9106 VSS.n9105 0.017685
R63420 VSS.n12952 VSS.n12951 0.017685
R63421 VSS.n12923 VSS.n12922 0.017685
R63422 VSS.n12734 VSS.n12733 0.017685
R63423 VSS.n12706 VSS.n12705 0.017685
R63424 VSS.n15024 VSS.n15023 0.017685
R63425 VSS.n15051 VSS.n15050 0.017685
R63426 VSS.n16089 VSS.n16088 0.017685
R63427 VSS.n9599 VSS.n9598 0.017685
R63428 VSS.n9686 VSS.n9685 0.017685
R63429 VSS.n9166 VSS.n9165 0.017685
R63430 VSS.n9295 VSS.n9294 0.017685
R63431 VSS.n9269 VSS.n9268 0.017685
R63432 VSS.n20632 VSS.n20631 0.017685
R63433 VSS.n20661 VSS.n20660 0.017685
R63434 VSS.n21021 VSS.n21020 0.017685
R63435 VSS.n6913 VSS.n6912 0.017685
R63436 VSS.n6979 VSS.n6978 0.017685
R63437 VSS.n6654 VSS.n6653 0.017685
R63438 VSS.n6619 VSS.n6618 0.017685
R63439 VSS.n6590 VSS.n6589 0.017685
R63440 VSS.n20117 VSS.n20116 0.017685
R63441 VSS.n20088 VSS.n20087 0.017685
R63442 VSS.n1067 VSS.n1066 0.017685
R63443 VSS.n6790 VSS.n6789 0.017685
R63444 VSS.n6877 VSS.n6876 0.017685
R63445 VSS.n6504 VSS.n6503 0.017685
R63446 VSS.n6469 VSS.n6468 0.017685
R63447 VSS.n6440 VSS.n6439 0.017685
R63448 VSS.n21369 VSS.n21368 0.017685
R63449 VSS.n21340 VSS.n21339 0.017685
R63450 VSS.n7628 VSS.n7627 0.017685
R63451 VSS.n7657 VSS.n7656 0.017685
R63452 VSS.n7716 VSS.n7715 0.017685
R63453 VSS.n7745 VSS.n7744 0.017685
R63454 VSS.n7823 VSS.n7822 0.017685
R63455 VSS.n7794 VSS.n7793 0.017685
R63456 VSS.n11685 VSS.n11684 0.017685
R63457 VSS.n11658 VSS.n11657 0.017685
R63458 VSS.n6128 VSS.n6127 0.017685
R63459 VSS.n6102 VSS.n6101 0.017685
R63460 VSS.n6047 VSS.n6046 0.017685
R63461 VSS.n6021 VSS.n6020 0.017685
R63462 VSS.n5966 VSS.n5965 0.017685
R63463 VSS.n5940 VSS.n5939 0.017685
R63464 VSS.n642 VSS.n641 0.017685
R63465 VSS.n616 VSS.n615 0.017685
R63466 VSS.n10600 VSS.n10599 0.017685
R63467 VSS.n10574 VSS.n10573 0.017685
R63468 VSS.n16343 VSS.n16338 0.0174947
R63469 VSS.n16302 VSS.n16299 0.0174947
R63470 VSS.n16267 VSS.n16264 0.0174947
R63471 VSS.n5705 VSS.n5702 0.0174947
R63472 VSS.n5697 VSS.n5696 0.0174947
R63473 VSS.n5765 VSS.n5759 0.0174947
R63474 VSS.n1431 VSS.n1426 0.0172553
R63475 VSS.n1385 VSS.n1382 0.0172553
R63476 VSS.n1351 VSS.n1348 0.0172553
R63477 VSS.n20976 VSS.n20971 0.0172553
R63478 VSS.n20965 VSS.n20961 0.0172553
R63479 VSS.n20966 VSS.n20965 0.0172553
R63480 VSS.n1219 VSS.n1218 0.0172553
R63481 VSS.n1218 VSS.n1214 0.0172553
R63482 VSS.n8660 VSS.n8659 0.0171062
R63483 VSS.n8509 VSS.n8508 0.0171062
R63484 VSS.n19008 VSS.n19006 0.0170278
R63485 VSS.n19010 VSS.n19008 0.0170278
R63486 VSS.n16428 VSS.n16426 0.0170278
R63487 VSS.n14968 VSS.n14966 0.0170278
R63488 VSS.n14939 VSS.n14937 0.0170278
R63489 VSS.n17171 VSS.n17168 0.0170278
R63490 VSS.n17171 VSS.n17170 0.0170278
R63491 VSS.n14665 VSS.n14663 0.0170278
R63492 VSS.n18245 VSS.n2146 0.0170278
R63493 VSS.n19378 VSS.n19374 0.0170278
R63494 VSS.n5696 VSS.n5692 0.017016
R63495 VSS.n5766 VSS.n5765 0.017016
R63496 VSS.n12223 VSS.n12222 0.0169764
R63497 VSS.n10171 VSS.n10170 0.0169764
R63498 VSS.n16545 VSS.n16544 0.0169489
R63499 VSS.n793 VSS.n792 0.0169489
R63500 VSS.n166 VSS.n165 0.0168408
R63501 VSS.n5629 VSS.n5628 0.0167992
R63502 VSS.n16151 VSS.n16150 0.0167992
R63503 VSS.n21079 VSS.n21078 0.0167992
R63504 VSS.n1131 VSS.n1130 0.0167992
R63505 VSS.n18813 VSS.n18812 0.0167676
R63506 VSS.n19485 VSS.n19484 0.0167676
R63507 VSS.n14883 VSS.n14882 0.0167379
R63508 VSS.n19954 VSS.n19953 0.0167379
R63509 VSS.n5657 VSS.n5656 0.0167162
R63510 VSS.n5535 VSS.n5533 0.0167162
R63511 VSS.n16077 VSS.n16076 0.0167162
R63512 VSS.n16040 VSS.n16038 0.0167162
R63513 VSS.n1046 VSS.n1045 0.0167162
R63514 VSS.n1019 VSS.n1017 0.0167162
R63515 VSS.n20924 VSS.n20923 0.0167162
R63516 VSS.n16912 VSS.n16911 0.0166324
R63517 VSS.n20004 VSS.n20003 0.0166324
R63518 VSS.n16925 VSS.n16924 0.0163158
R63519 VSS.n19991 VSS.n19990 0.0163158
R63520 VSS.n5739 VSS.n5738 0.0162677
R63521 VSS.n16187 VSS.n16186 0.0162677
R63522 VSS.n21129 VSS.n21128 0.0162677
R63523 VSS.n1179 VSS.n1178 0.0162677
R63524 VSS.n14870 VSS.n14869 0.0162103
R63525 VSS.n19941 VSS.n19940 0.0162103
R63526 VSS.n18917 VSS.n18916 0.0161472
R63527 VSS.n21848 VSS.n21847 0.0161472
R63528 VSS.n17033 VSS.n17032 0.0161047
R63529 VSS.n16584 VSS.n16583 0.0161047
R63530 VSS.n19902 VSS.n19901 0.0161047
R63531 VSS.n784 VSS.n783 0.0161047
R63532 VSS.n11592 VSS.n11591 0.0160906
R63533 VSS.n12905 VSS.n12904 0.0160906
R63534 VSS.n15067 VSS.n15066 0.0160906
R63535 VSS.n20679 VSS.n20678 0.0160906
R63536 VSS.n20070 VSS.n20069 0.0160906
R63537 VSS.n600 VSS.n599 0.0160906
R63538 VSS.n12652 VSS.n12651 0.0160769
R63539 VSS.n9082 VSS.n9081 0.0160299
R63540 VSS.n6566 VSS.n6565 0.0160299
R63541 VSS.n9246 VSS.n9245 0.0160299
R63542 VSS.n17074 VSS.n17073 0.0159992
R63543 VSS.n19891 VSS.n19890 0.0159992
R63544 VSS.n1932 VSS.n1931 0.0159869
R63545 VSS.n15674 VSS.n15673 0.0159869
R63546 VSS.n21480 VSS.n21479 0.0159134
R63547 VSS.n4757 VSS.n4756 0.0159134
R63548 VSS.n9828 VSS.n9827 0.0158846
R63549 VSS.n5850 VSS.n5849 0.0157362
R63550 VSS.n16211 VSS.n16210 0.0157362
R63551 VSS.n21153 VSS.n21152 0.0157362
R63552 VSS.n1282 VSS.n1281 0.0157362
R63553 VSS.n18446 VSS.n18445 0.0157113
R63554 VSS.n8487 VSS.n8486 0.0157113
R63555 VSS.n19593 VSS.n19592 0.0157113
R63556 VSS.n8638 VSS.n8637 0.0157113
R63557 VSS.n16537 VSS.n16536 0.0156825
R63558 VSS.n801 VSS.n800 0.0156825
R63559 VSS.n14395 VSS.n14394 0.0155982
R63560 VSS.n14428 VSS.n14427 0.0155982
R63561 VSS.n15069 VSS.n15068 0.0155982
R63562 VSS.n15102 VSS.n15101 0.0155982
R63563 VSS.n15172 VSS.n15171 0.0155982
R63564 VSS.n13359 VSS.n13358 0.0155982
R63565 VSS.n13410 VSS.n13409 0.0155982
R63566 VSS.n20681 VSS.n20680 0.0155982
R63567 VSS.n20732 VSS.n20731 0.0155982
R63568 VSS.n20824 VSS.n20823 0.0155982
R63569 VSS.n6937 VSS.n6936 0.0155982
R63570 VSS.n9066 VSS.n9065 0.0155982
R63571 VSS.n535 VSS.n534 0.0155982
R63572 VSS.n9079 VSS.n9066 0.0155982
R63573 VSS.n16904 VSS.n16903 0.015577
R63574 VSS.n20012 VSS.n20011 0.015577
R63575 VSS.n14563 VSS.n14562 0.015567
R63576 VSS.n14832 VSS.n14831 0.015567
R63577 VSS.n16876 VSS.n16875 0.015567
R63578 VSS.n16687 VSS.n16686 0.015567
R63579 VSS.n16436 VSS.n16435 0.015567
R63580 VSS.n19765 VSS.n19764 0.015567
R63581 VSS.n19855 VSS.n19854 0.015567
R63582 VSS.n20040 VSS.n20039 0.015567
R63583 VSS.n2089 VSS.n2088 0.015567
R63584 VSS.n853 VSS.n852 0.015567
R63585 VSS.n17245 VSS.n17244 0.0155658
R63586 VSS.n11739 VSS.n11738 0.0155658
R63587 VSS.n4927 VSS.n4926 0.0155658
R63588 VSS.n11460 VSS.n11459 0.0155658
R63589 VSS.n11245 VSS.n11244 0.0155658
R63590 VSS.n5552 VSS.n5551 0.0155591
R63591 VSS.n16062 VSS.n16061 0.0155591
R63592 VSS.n20997 VSS.n20996 0.0155591
R63593 VSS.n1039 VSS.n1038 0.0155591
R63594 VSS.n18173 VSS.n18172 0.0155
R63595 VSS.n19683 VSS.n19682 0.0155
R63596 VSS.n13075 VSS.n13074 0.0154808
R63597 VSS.n19133 VSS.n19132 0.0154808
R63598 VSS.n2662 VSS.n2641 0.0154808
R63599 VSS.n4046 VSS.n4045 0.0154808
R63600 VSS.n6416 VSS.n6415 0.0153635
R63601 VSS.n18720 VSS.n18719 0.0152887
R63602 VSS.n19202 VSS.n19201 0.0152887
R63603 VSS.n17079 VSS.n17078 0.0151547
R63604 VSS.n14862 VSS.n14861 0.0151547
R63605 VSS.n19886 VSS.n19885 0.0151547
R63606 VSS.n19933 VSS.n19932 0.0151547
R63607 VSS.n15309 VSS.n15308 0.0150946
R63608 VSS.n1628 VSS.n1627 0.0150946
R63609 VSS.n1621 VSS.n1619 0.0150946
R63610 VSS.n18804 VSS.n18803 0.0149435
R63611 VSS.n14891 VSS.n14890 0.0149435
R63612 VSS.n19476 VSS.n19475 0.0149435
R63613 VSS.n19962 VSS.n19961 0.0149435
R63614 VSS.n4660 VSS.n4659 0.0149
R63615 VSS.n18140 VSS.n18139 0.0148662
R63616 VSS.n19716 VSS.n19715 0.0148662
R63617 VSS.n12221 VSS.n12220 0.0148504
R63618 VSS.n10169 VSS.n10168 0.0148504
R63619 VSS.n18399 VSS.n18398 0.0148379
R63620 VSS.n19623 VSS.n19622 0.0148379
R63621 VSS.n5599 VSS.n5598 0.0147386
R63622 VSS.n16115 VSS.n16114 0.0147386
R63623 VSS.n21049 VSS.n21048 0.0147386
R63624 VSS.n1095 VSS.n1094 0.0147386
R63625 VSS.n7543 VSS.n7542 0.014713
R63626 VSS.n11239 VSS.n11238 0.014713
R63627 VSS.n18166 VSS.n18165 0.0146549
R63628 VSS.n19690 VSS.n19689 0.0146549
R63629 VSS.n14670 VSS.n14388 0.0146478
R63630 VSS.n17165 VSS.n14833 0.0146478
R63631 VSS.n16874 VSS.n16873 0.0146478
R63632 VSS.n16685 VSS.n16684 0.0146478
R63633 VSS.n16433 VSS.n14994 0.0146478
R63634 VSS.n18448 VSS.n18447 0.0146478
R63635 VSS.n18175 VSS.n18174 0.0146478
R63636 VSS.n18722 VSS.n18721 0.0146478
R63637 VSS.n8430 VSS.n8344 0.0146478
R63638 VSS.n8575 VSS.n8526 0.0146478
R63639 VSS.n8726 VSS.n8677 0.0146478
R63640 VSS.n8238 VSS.n8140 0.0146478
R63641 VSS.n19768 VSS.n19767 0.0146478
R63642 VSS.n19858 VSS.n19857 0.0146478
R63643 VSS.n20042 VSS.n2130 0.0146478
R63644 VSS.n2086 VSS.n739 0.0146478
R63645 VSS.n1969 VSS.n854 0.0146478
R63646 VSS.n19591 VSS.n19590 0.0146478
R63647 VSS.n19681 VSS.n19680 0.0146478
R63648 VSS.n19203 VSS.n19202 0.0146478
R63649 VSS.n8506 VSS.n8487 0.0146478
R63650 VSS.n8657 VSS.n8638 0.0146478
R63651 VSS.n18437 VSS.n18436 0.0146267
R63652 VSS.n19602 VSS.n19601 0.0146267
R63653 VSS.n6837 VSS.n6836 0.0146212
R63654 VSS.n9533 VSS.n9532 0.0146212
R63655 VSS.n9650 VSS.n9649 0.0146212
R63656 VSS.n18781 VSS.n18780 0.0145211
R63657 VSS.n16933 VSS.n16932 0.0145211
R63658 VSS.n19453 VSS.n19452 0.0145211
R63659 VSS.n19983 VSS.n19982 0.0145211
R63660 VSS.n21524 VSS.n21523 0.0144961
R63661 VSS.n4141 VSS.n2430 0.0144961
R63662 VSS.n16592 VSS.n16591 0.0144155
R63663 VSS.n776 VSS.n775 0.0144155
R63664 VSS.n16434 VSS.n16433 0.0143948
R63665 VSS.n14671 VSS.n14670 0.0143948
R63666 VSS.n17165 VSS.n17164 0.0143948
R63667 VSS.n16873 VSS.n16872 0.0143948
R63668 VSS.n16684 VSS.n16683 0.0143948
R63669 VSS.n18721 VSS.n18720 0.0143948
R63670 VSS.n18447 VSS.n18446 0.0143948
R63671 VSS.n18174 VSS.n18173 0.0143948
R63672 VSS.n8430 VSS.n8429 0.0143948
R63673 VSS.n8575 VSS.n8574 0.0143948
R63674 VSS.n8238 VSS.n8237 0.0143948
R63675 VSS.n8726 VSS.n8725 0.0143948
R63676 VSS.n19857 VSS.n19856 0.0143948
R63677 VSS.n19767 VSS.n19766 0.0143948
R63678 VSS.n1969 VSS.n1968 0.0143948
R63679 VSS.n2087 VSS.n2086 0.0143948
R63680 VSS.n20042 VSS.n20041 0.0143948
R63681 VSS.n19204 VSS.n19203 0.0143948
R63682 VSS.n19592 VSS.n19591 0.0143948
R63683 VSS.n19682 VSS.n19681 0.0143948
R63684 VSS.n8507 VSS.n8506 0.0143948
R63685 VSS.n8658 VSS.n8657 0.0143948
R63686 VSS.n18200 VSS.n18199 0.0143098
R63687 VSS.n17025 VSS.n17024 0.0143098
R63688 VSS.n19656 VSS.n19655 0.0143098
R63689 VSS.n19910 VSS.n19909 0.0143098
R63690 VSS.n18749 VSS.n18748 0.0142042
R63691 VSS.n19231 VSS.n19230 0.0142042
R63692 VSS.n21255 VSS.n21254 0.0141909
R63693 VSS.n21307 VSS.n21306 0.0141909
R63694 VSS.n21318 VSS.n21317 0.0141909
R63695 VSS.n21417 VSS.n21416 0.0141909
R63696 VSS.n21428 VSS.n21427 0.0141909
R63697 VSS.n17248 VSS.n17247 0.0141909
R63698 VSS.n11742 VSS.n11741 0.0141909
R63699 VSS.n4924 VSS.n4923 0.0141909
R63700 VSS.n11463 VSS.n11462 0.0141909
R63701 VSS.n11242 VSS.n11241 0.0141909
R63702 VSS.n21252 VSS.n21251 0.0141618
R63703 VSS.n21304 VSS.n21303 0.0141618
R63704 VSS.n21315 VSS.n21314 0.0141618
R63705 VSS.n21414 VSS.n21413 0.0141618
R63706 VSS.n21425 VSS.n21424 0.0141618
R63707 VSS.n9093 VSS.n9092 0.0141417
R63708 VSS.n15039 VSS.n15038 0.0141417
R63709 VSS.n21620 VSS.n21619 0.0141417
R63710 VSS.n3849 VSS.n3848 0.0141417
R63711 VSS.n11670 VSS.n11669 0.0141417
R63712 VSS.n141 VSS.n139 0.0140754
R63713 VSS.n139 VSS.n136 0.0140754
R63714 VSS.n110 VSS.n108 0.0140754
R63715 VSS.n108 VSS.n105 0.0140754
R63716 VSS.n78 VSS.n76 0.0140754
R63717 VSS.n76 VSS.n73 0.0140754
R63718 VSS.n53 VSS.n51 0.0140754
R63719 VSS.n51 VSS.n48 0.0140754
R63720 VSS.n48 VSS.n46 0.0140754
R63721 VSS.n46 VSS.n43 0.0140754
R63722 VSS.n211 VSS.n208 0.0140754
R63723 VSS.n213 VSS.n211 0.0140754
R63724 VSS.n216 VSS.n213 0.0140754
R63725 VSS.n218 VSS.n216 0.0140754
R63726 VSS.n241 VSS.n238 0.0140754
R63727 VSS.n243 VSS.n241 0.0140754
R63728 VSS.n273 VSS.n270 0.0140754
R63729 VSS.n275 VSS.n273 0.0140754
R63730 VSS.n305 VSS.n302 0.0140754
R63731 VSS.n307 VSS.n305 0.0140754
R63732 VSS.n329 VSS.n327 0.0140754
R63733 VSS.n1479 VSS.n856 0.0140754
R63734 VSS.n1479 VSS.n1476 0.0140754
R63735 VSS.n1476 VSS.n1474 0.0140754
R63736 VSS.n1469 VSS.n878 0.0140754
R63737 VSS.n878 VSS.n876 0.0140754
R63738 VSS.n876 VSS.n873 0.0140754
R63739 VSS.n873 VSS.n871 0.0140754
R63740 VSS.n871 VSS.n868 0.0140754
R63741 VSS.n868 VSS.n866 0.0140754
R63742 VSS.n866 VSS.n863 0.0140754
R63743 VSS.n863 VSS.n861 0.0140754
R63744 VSS.n449 VSS.n447 0.0140754
R63745 VSS.n452 VSS.n449 0.0140754
R63746 VSS.n454 VSS.n452 0.0140754
R63747 VSS.n457 VSS.n454 0.0140754
R63748 VSS.n459 VSS.n457 0.0140754
R63749 VSS.n21195 VSS.n459 0.0140754
R63750 VSS.n21197 VSS.n21195 0.0140754
R63751 VSS.n21200 VSS.n21197 0.0140754
R63752 VSS.n21206 VSS.n21204 0.0140754
R63753 VSS.n21209 VSS.n21206 0.0140754
R63754 VSS.n21211 VSS.n21209 0.0140754
R63755 VSS.n21214 VSS.n21211 0.0140754
R63756 VSS.n21216 VSS.n21214 0.0140754
R63757 VSS.n21219 VSS.n21216 0.0140754
R63758 VSS.n21221 VSS.n21219 0.0140754
R63759 VSS.n21224 VSS.n21221 0.0140754
R63760 VSS.n21231 VSS.n21229 0.0140754
R63761 VSS.n21233 VSS.n21231 0.0140754
R63762 VSS.n15185 VSS.n15183 0.0140754
R63763 VSS.n15188 VSS.n15185 0.0140754
R63764 VSS.n15190 VSS.n15188 0.0140754
R63765 VSS.n15193 VSS.n15190 0.0140754
R63766 VSS.n15195 VSS.n15193 0.0140754
R63767 VSS.n15914 VSS.n15195 0.0140754
R63768 VSS.n15914 VSS.n15911 0.0140754
R63769 VSS.n15911 VSS.n15909 0.0140754
R63770 VSS.n15905 VSS.n15200 0.0140754
R63771 VSS.n15200 VSS.n15198 0.0140754
R63772 VSS.n11257 VSS.n11255 0.0140754
R63773 VSS.n11265 VSS.n11263 0.0140754
R63774 VSS.n11268 VSS.n11265 0.0140754
R63775 VSS.n11270 VSS.n11268 0.0140754
R63776 VSS.n11273 VSS.n11270 0.0140754
R63777 VSS.n11275 VSS.n11273 0.0140754
R63778 VSS.n11278 VSS.n11275 0.0140754
R63779 VSS.n11280 VSS.n11278 0.0140754
R63780 VSS.n11282 VSS.n11280 0.0140754
R63781 VSS.n11289 VSS.n11287 0.0140754
R63782 VSS.n11292 VSS.n11289 0.0140754
R63783 VSS.n11294 VSS.n11292 0.0140754
R63784 VSS.n11297 VSS.n11294 0.0140754
R63785 VSS.n11299 VSS.n11297 0.0140754
R63786 VSS.n11308 VSS.n11299 0.0140754
R63787 VSS.n11308 VSS.n11305 0.0140754
R63788 VSS.n11305 VSS.n11303 0.0140754
R63789 VSS.n163 VSS.n161 0.013824
R63790 VSS.n11255 VSS.n11253 0.013824
R63791 VSS.n10552 VSS.n10551 0.0137198
R63792 VSS.n12684 VSS.n12683 0.0137198
R63793 VSS.n1465 VSS.n1464 0.0136815
R63794 VSS.n12821 VSS.n12820 0.0136815
R63795 VSS.n21190 VSS.n21189 0.0136815
R63796 VSS.n16382 VSS.n16381 0.0136815
R63797 VSS.n5881 VSS.n5880 0.0136815
R63798 VSS.n18700 VSS.n18699 0.0135986
R63799 VSS.n18742 VSS.n18741 0.0135986
R63800 VSS.n18420 VSS.n18412 0.0135986
R63801 VSS.n18193 VSS.n18192 0.0135986
R63802 VSS.n17125 VSS.n17124 0.0135986
R63803 VSS.n17069 VSS.n17068 0.0135986
R63804 VSS.n14875 VSS.n14874 0.0135986
R63805 VSS.n16917 VSS.n16916 0.0135986
R63806 VSS.n16579 VSS.n16578 0.0135986
R63807 VSS.n15525 VSS.n15524 0.0135986
R63808 VSS.n15335 VSS.n15334 0.0135986
R63809 VSS.n19182 VSS.n19181 0.0135986
R63810 VSS.n19224 VSS.n19223 0.0135986
R63811 VSS.n19609 VSS.n19608 0.0135986
R63812 VSS.n19663 VSS.n19662 0.0135986
R63813 VSS.n19870 VSS.n19869 0.0135986
R63814 VSS.n19896 VSS.n19895 0.0135986
R63815 VSS.n19946 VSS.n19945 0.0135986
R63816 VSS.n19999 VSS.n19998 0.0135986
R63817 VSS.n789 VSS.n788 0.0135986
R63818 VSS.n1813 VSS.n1812 0.0135986
R63819 VSS.n1651 VSS.n1650 0.0135986
R63820 VSS.n5651 VSS.n5650 0.013473
R63821 VSS.n5647 VSS.n5645 0.013473
R63822 VSS.n16031 VSS.n16029 0.013473
R63823 VSS.n16045 VSS.n16043 0.013473
R63824 VSS.n1006 VSS.n1004 0.013473
R63825 VSS.n20913 VSS.n20911 0.013473
R63826 VSS.n20918 VSS.n20917 0.013473
R63827 VSS.n13244 VSS.n13243 0.0134466
R63828 VSS.n13002 VSS.n13001 0.0134466
R63829 VSS.n12901 VSS.n12900 0.0134466
R63830 VSS.n12888 VSS.n12887 0.0134466
R63831 VSS.n12834 VSS.n12833 0.0134466
R63832 VSS.n13504 VSS.n13503 0.0134466
R63833 VSS.n2050 VSS.n2049 0.0134466
R63834 VSS.n2047 VSS.n2046 0.0134466
R63835 VSS.n880 VSS.n879 0.0134466
R63836 VSS.n596 VSS.n595 0.0134466
R63837 VSS.n583 VSS.n582 0.0134466
R63838 VSS.n12686 VSS.n12685 0.0134331
R63839 VSS.n10554 VSS.n10553 0.0134331
R63840 VSS.n16349 VSS.n16346 0.0134255
R63841 VSS.n16355 VSS.n16349 0.0134255
R63842 VSS.n16355 VSS.n16354 0.0134255
R63843 VSS.n15940 VSS.n15937 0.0134255
R63844 VSS.n15949 VSS.n15940 0.0134255
R63845 VSS.n15949 VSS.n15948 0.0134255
R63846 VSS.n15948 VSS.n15945 0.0134255
R63847 VSS.n15227 VSS.n15224 0.0134255
R63848 VSS.n15236 VSS.n15227 0.0134255
R63849 VSS.n15236 VSS.n15235 0.0134255
R63850 VSS.n15235 VSS.n15232 0.0134255
R63851 VSS.n15647 VSS.n15640 0.0134255
R63852 VSS.n1501 VSS.n1498 0.0134255
R63853 VSS.n1510 VSS.n1501 0.0134255
R63854 VSS.n1510 VSS.n1509 0.0134255
R63855 VSS.n1509 VSS.n1506 0.0134255
R63856 VSS.n1519 VSS.n1513 0.0134255
R63857 VSS.n913 VSS.n910 0.0134255
R63858 VSS.n922 VSS.n913 0.0134255
R63859 VSS.n922 VSS.n921 0.0134255
R63860 VSS.n921 VSS.n918 0.0134255
R63861 VSS.n1436 VSS.n1411 0.0134255
R63862 VSS.n1436 VSS.n1435 0.0134255
R63863 VSS.n1435 VSS.n1432 0.0134255
R63864 VSS.n16306 VSS.n16304 0.0134255
R63865 VSS.n16310 VSS.n16306 0.0134255
R63866 VSS.n16310 VSS.n16308 0.0134255
R63867 VSS.n15953 VSS.n15951 0.0134255
R63868 VSS.n15959 VSS.n15953 0.0134255
R63869 VSS.n15959 VSS.n15957 0.0134255
R63870 VSS.n15957 VSS.n15955 0.0134255
R63871 VSS.n15242 VSS.n15240 0.0134255
R63872 VSS.n15248 VSS.n15242 0.0134255
R63873 VSS.n15248 VSS.n15246 0.0134255
R63874 VSS.n15246 VSS.n15244 0.0134255
R63875 VSS.n15620 VSS.n15616 0.0134255
R63876 VSS.n1523 VSS.n1521 0.0134255
R63877 VSS.n1529 VSS.n1523 0.0134255
R63878 VSS.n1529 VSS.n1527 0.0134255
R63879 VSS.n1527 VSS.n1525 0.0134255
R63880 VSS.n1535 VSS.n1531 0.0134255
R63881 VSS.n926 VSS.n924 0.0134255
R63882 VSS.n932 VSS.n926 0.0134255
R63883 VSS.n932 VSS.n930 0.0134255
R63884 VSS.n930 VSS.n928 0.0134255
R63885 VSS.n1391 VSS.n1375 0.0134255
R63886 VSS.n1391 VSS.n1389 0.0134255
R63887 VSS.n1389 VSS.n1387 0.0134255
R63888 VSS.n16271 VSS.n16269 0.0134255
R63889 VSS.n16275 VSS.n16271 0.0134255
R63890 VSS.n16275 VSS.n16274 0.0134255
R63891 VSS.n15963 VSS.n15961 0.0134255
R63892 VSS.n15969 VSS.n15963 0.0134255
R63893 VSS.n15969 VSS.n15968 0.0134255
R63894 VSS.n15968 VSS.n15966 0.0134255
R63895 VSS.n15254 VSS.n15252 0.0134255
R63896 VSS.n15260 VSS.n15254 0.0134255
R63897 VSS.n15260 VSS.n15259 0.0134255
R63898 VSS.n15259 VSS.n15257 0.0134255
R63899 VSS.n15597 VSS.n15593 0.0134255
R63900 VSS.n1539 VSS.n1537 0.0134255
R63901 VSS.n1545 VSS.n1539 0.0134255
R63902 VSS.n1545 VSS.n1544 0.0134255
R63903 VSS.n1544 VSS.n1542 0.0134255
R63904 VSS.n1551 VSS.n1547 0.0134255
R63905 VSS.n936 VSS.n934 0.0134255
R63906 VSS.n942 VSS.n936 0.0134255
R63907 VSS.n942 VSS.n941 0.0134255
R63908 VSS.n941 VSS.n939 0.0134255
R63909 VSS.n1356 VSS.n1339 0.0134255
R63910 VSS.n1356 VSS.n1355 0.0134255
R63911 VSS.n1355 VSS.n1353 0.0134255
R63912 VSS.n5709 VSS.n5707 0.0134255
R63913 VSS.n5713 VSS.n5709 0.0134255
R63914 VSS.n5713 VSS.n5711 0.0134255
R63915 VSS.n5503 VSS.n5501 0.0134255
R63916 VSS.n5527 VSS.n5503 0.0134255
R63917 VSS.n5527 VSS.n5525 0.0134255
R63918 VSS.n5525 VSS.n5523 0.0134255
R63919 VSS.n5519 VSS.n5517 0.0134255
R63920 VSS.n5517 VSS.n5515 0.0134255
R63921 VSS.n5515 VSS.n5513 0.0134255
R63922 VSS.n5513 VSS.n5511 0.0134255
R63923 VSS.n5511 VSS.n5509 0.0134255
R63924 VSS.n5509 VSS.n5507 0.0134255
R63925 VSS.n5507 VSS.n5505 0.0134255
R63926 VSS.n15426 VSS.n15424 0.0134255
R63927 VSS.n15424 VSS.n15422 0.0134255
R63928 VSS.n15432 VSS.n15430 0.0134255
R63929 VSS.n15434 VSS.n15432 0.0134255
R63930 VSS.n15438 VSS.n15434 0.0134255
R63931 VSS.n1738 VSS.n1737 0.0134255
R63932 VSS.n1737 VSS.n1735 0.0134255
R63933 VSS.n1586 VSS.n1584 0.0134255
R63934 VSS.n1588 VSS.n1586 0.0134255
R63935 VSS.n1592 VSS.n1588 0.0134255
R63936 VSS.n974 VSS.n972 0.0134255
R63937 VSS.n980 VSS.n974 0.0134255
R63938 VSS.n980 VSS.n979 0.0134255
R63939 VSS.n979 VSS.n977 0.0134255
R63940 VSS.n1151 VSS.n1143 0.0134255
R63941 VSS.n1151 VSS.n1150 0.0134255
R63942 VSS.n1150 VSS.n1148 0.0134255
R63943 VSS.n21095 VSS.n21092 0.0134255
R63944 VSS.n21101 VSS.n21095 0.0134255
R63945 VSS.n21101 VSS.n21100 0.0134255
R63946 VSS.n20898 VSS.n20895 0.0134255
R63947 VSS.n20983 VSS.n20898 0.0134255
R63948 VSS.n20983 VSS.n20982 0.0134255
R63949 VSS.n20982 VSS.n20979 0.0134255
R63950 VSS.n5682 VSS.n5680 0.0134255
R63951 VSS.n5680 VSS.n5678 0.0134255
R63952 VSS.n16144 VSS.n16140 0.0134255
R63953 VSS.n16144 VSS.n16142 0.0134255
R63954 VSS.n15286 VSS.n15282 0.0134255
R63955 VSS.n15286 VSS.n15284 0.0134255
R63956 VSS.n1599 VSS.n1595 0.0134255
R63957 VSS.n1599 VSS.n1598 0.0134255
R63958 VSS.n1124 VSS.n1120 0.0134255
R63959 VSS.n1124 VSS.n1122 0.0134255
R63960 VSS.n20949 VSS.n20947 0.0134255
R63961 VSS.n20951 VSS.n20949 0.0134255
R63962 VSS.n5836 VSS.n5783 0.0134255
R63963 VSS.n5836 VSS.n5833 0.0134255
R63964 VSS.n5803 VSS.n5800 0.0134255
R63965 VSS.n5800 VSS.n5799 0.0134255
R63966 VSS.n15499 VSS.n15496 0.0134255
R63967 VSS.n15502 VSS.n15499 0.0134255
R63968 VSS.n15519 VSS.n15502 0.0134255
R63969 VSS.n15519 VSS.n15516 0.0134255
R63970 VSS.n1807 VSS.n1786 0.0134255
R63971 VSS.n1807 VSS.n1804 0.0134255
R63972 VSS.n1804 VSS.n1801 0.0134255
R63973 VSS.n1801 VSS.n1798 0.0134255
R63974 VSS.n1268 VSS.n1207 0.0134255
R63975 VSS.n1268 VSS.n1265 0.0134255
R63976 VSS.n1235 VSS.n1233 0.0134255
R63977 VSS.n1233 VSS.n1232 0.0134255
R63978 VSS.n18834 VSS.n18833 0.0133873
R63979 VSS.n19506 VSS.n19505 0.0133873
R63980 VSS.n17348 VSS.n17347 0.0133291
R63981 VSS.n17329 VSS.n17328 0.0133291
R63982 VSS.n11518 VSS.n11517 0.0133291
R63983 VSS.n11328 VSS.n11327 0.0133291
R63984 VSS.n11315 VSS.n11314 0.0133291
R63985 VSS.n13249 VSS.n13248 0.0133291
R63986 VSS.n12997 VSS.n12996 0.0133291
R63987 VSS.n12896 VSS.n12895 0.0133291
R63988 VSS.n12883 VSS.n12882 0.0133291
R63989 VSS.n12829 VSS.n12828 0.0133291
R63990 VSS.n14402 VSS.n14401 0.0133291
R63991 VSS.n14421 VSS.n14420 0.0133291
R63992 VSS.n15076 VSS.n15075 0.0133291
R63993 VSS.n15109 VSS.n15108 0.0133291
R63994 VSS.n15179 VSS.n15178 0.0133291
R63995 VSS.n13366 VSS.n13365 0.0133291
R63996 VSS.n13417 VSS.n13416 0.0133291
R63997 VSS.n20688 VSS.n20687 0.0133291
R63998 VSS.n20739 VSS.n20738 0.0133291
R63999 VSS.n20831 VSS.n20830 0.0133291
R64000 VSS.n13509 VSS.n13508 0.0133291
R64001 VSS.n20149 VSS.n20148 0.0133291
R64002 VSS.n2055 VSS.n2054 0.0133291
R64003 VSS.n2042 VSS.n2041 0.0133291
R64004 VSS.n885 VSS.n884 0.0133291
R64005 VSS.n591 VSS.n590 0.0133291
R64006 VSS.n578 VSS.n577 0.0133291
R64007 VSS.n528 VSS.n527 0.0133291
R64008 VSS.n9505 VSS.n9504 0.0132559
R64009 VSS.n9622 VSS.n9621 0.0132559
R64010 VSS.n6935 VSS.n6934 0.0132559
R64011 VSS.n6812 VSS.n6811 0.0132559
R64012 VSS.n16530 VSS.n16529 0.0131761
R64013 VSS.n808 VSS.n807 0.0131761
R64014 VSS.n17481 VSS.n17480 0.0130787
R64015 VSS.n13193 VSS.n13192 0.0130787
R64016 VSS.n18108 VSS.n18107 0.0130787
R64017 VSS.n2336 VSS.n2335 0.0130787
R64018 VSS.n17965 VSS.n17964 0.0130787
R64019 VSS.n148 VSS.n146 0.0130698
R64020 VSS.n130 VSS.n129 0.0130698
R64021 VSS.n117 VSS.n115 0.0130698
R64022 VSS.n99 VSS.n98 0.0130698
R64023 VSS.n85 VSS.n83 0.0130698
R64024 VSS.n67 VSS.n66 0.0130698
R64025 VSS.n232 VSS.n231 0.0130698
R64026 VSS.n250 VSS.n248 0.0130698
R64027 VSS.n264 VSS.n263 0.0130698
R64028 VSS.n282 VSS.n280 0.0130698
R64029 VSS.n296 VSS.n295 0.0130698
R64030 VSS.n314 VSS.n312 0.0130698
R64031 VSS.n520 VSS.n519 0.0130151
R64032 VSS.n1935 VSS.n1934 0.0129759
R64033 VSS.n15902 VSS.n15702 0.0129759
R64034 VSS.n14987 VSS.n14986 0.0129648
R64035 VSS.n823 VSS.n822 0.0129648
R64036 VSS.n4007 VSS.n4006 0.0129016
R64037 VSS.n13032 VSS.n13031 0.0129016
R64038 VSS.n12693 VSS.n12692 0.0129016
R64039 VSS.n18878 VSS.n18877 0.0129016
R64040 VSS.n21805 VSS.n21804 0.0129016
R64041 VSS.n19090 VSS.n19089 0.0129016
R64042 VSS.n21576 VSS.n21575 0.0129016
R64043 VSS.n3809 VSS.n3808 0.0129016
R64044 VSS.n3287 VSS.n3286 0.0129016
R64045 VSS.n10561 VSS.n10560 0.0129016
R64046 VSS.n17343 VSS.n17342 0.0127801
R64047 VSS.n17334 VSS.n17333 0.0127801
R64048 VSS.n11523 VSS.n11522 0.0127801
R64049 VSS.n11323 VSS.n11322 0.0127801
R64050 VSS.n11320 VSS.n11319 0.0127801
R64051 VSS.n16630 VSS.n16629 0.0127535
R64052 VSS.n15383 VSS.n15382 0.0127535
R64053 VSS.n768 VSS.n767 0.0127535
R64054 VSS.n1699 VSS.n1698 0.0127535
R64055 VSS.n1934 VSS.n1933 0.0127233
R64056 VSS.n15902 VSS.n15901 0.0127233
R64057 VSS.n19278 VSS.n19275 0.01265
R64058 VSS.n19285 VSS.n19282 0.01265
R64059 VSS.n19292 VSS.n19289 0.01265
R64060 VSS.n19299 VSS.n19296 0.01265
R64061 VSS.n19306 VSS.n19303 0.01265
R64062 VSS.n19313 VSS.n19310 0.01265
R64063 VSS.n19320 VSS.n19317 0.01265
R64064 VSS.n19327 VSS.n19324 0.01265
R64065 VSS.n19334 VSS.n19331 0.01265
R64066 VSS.n19341 VSS.n19338 0.01265
R64067 VSS.n19437 VSS.n19345 0.01265
R64068 VSS.n19435 VSS.n19433 0.01265
R64069 VSS.n19433 VSS.n19431 0.01265
R64070 VSS.n19431 VSS.n19429 0.01265
R64071 VSS.n19429 VSS.n19427 0.01265
R64072 VSS.n19427 VSS.n19425 0.01265
R64073 VSS.n19425 VSS.n19423 0.01265
R64074 VSS.n19423 VSS.n19421 0.01265
R64075 VSS.n19421 VSS.n19419 0.01265
R64076 VSS.n19419 VSS.n19417 0.01265
R64077 VSS.n19417 VSS.n19414 0.01265
R64078 VSS.n19414 VSS.n19412 0.01265
R64079 VSS.n19412 VSS.n19411 0.01265
R64080 VSS.n19393 VSS.n19391 0.01265
R64081 VSS.n19391 VSS.n19390 0.01265
R64082 VSS.n18665 VSS.n18662 0.01265
R64083 VSS.n18655 VSS.n18652 0.01265
R64084 VSS.n18648 VSS.n18645 0.01265
R64085 VSS.n18641 VSS.n18638 0.01265
R64086 VSS.n18634 VSS.n18631 0.01265
R64087 VSS.n18627 VSS.n18624 0.01265
R64088 VSS.n18620 VSS.n18617 0.01265
R64089 VSS.n18613 VSS.n18610 0.01265
R64090 VSS.n18606 VSS.n18603 0.01265
R64091 VSS.n18599 VSS.n18596 0.01265
R64092 VSS.n18592 VSS.n18589 0.01265
R64093 VSS.n18585 VSS.n18582 0.01265
R64094 VSS.n18578 VSS.n18575 0.01265
R64095 VSS.n18571 VSS.n18568 0.01265
R64096 VSS.n18564 VSS.n18555 0.01265
R64097 VSS.n18562 VSS.n18560 0.01265
R64098 VSS.n18550 VSS.n18547 0.01265
R64099 VSS.n18543 VSS.n18540 0.01265
R64100 VSS.n18536 VSS.n18533 0.01265
R64101 VSS.n18529 VSS.n18526 0.01265
R64102 VSS.n18522 VSS.n18519 0.01265
R64103 VSS.n18515 VSS.n18512 0.01265
R64104 VSS.n18508 VSS.n18505 0.01265
R64105 VSS.n18501 VSS.n18498 0.01265
R64106 VSS.n18494 VSS.n18491 0.01265
R64107 VSS.n18487 VSS.n18479 0.01265
R64108 VSS.n18487 VSS.n18486 0.01265
R64109 VSS.n18435 VSS.n18432 0.01265
R64110 VSS.n18419 VSS.n18416 0.01265
R64111 VSS.n18389 VSS.n18386 0.01265
R64112 VSS.n18358 VSS.n18355 0.01265
R64113 VSS.n18351 VSS.n18348 0.01265
R64114 VSS.n18344 VSS.n18341 0.01265
R64115 VSS.n18337 VSS.n18334 0.01265
R64116 VSS.n18330 VSS.n18327 0.01265
R64117 VSS.n18323 VSS.n18320 0.01265
R64118 VSS.n18316 VSS.n18313 0.01265
R64119 VSS.n18309 VSS.n18306 0.01265
R64120 VSS.n18302 VSS.n18217 0.01265
R64121 VSS.n18300 VSS.n18298 0.01265
R64122 VSS.n18298 VSS.n18296 0.01265
R64123 VSS.n18296 VSS.n18294 0.01265
R64124 VSS.n18294 VSS.n18292 0.01265
R64125 VSS.n18292 VSS.n18290 0.01265
R64126 VSS.n18290 VSS.n18288 0.01265
R64127 VSS.n18288 VSS.n18286 0.01265
R64128 VSS.n18286 VSS.n18284 0.01265
R64129 VSS.n18284 VSS.n18282 0.01265
R64130 VSS.n18282 VSS.n18280 0.01265
R64131 VSS.n18280 VSS.n18278 0.01265
R64132 VSS.n18278 VSS.n18276 0.01265
R64133 VSS.n18276 VSS.n18274 0.01265
R64134 VSS.n18274 VSS.n18272 0.01265
R64135 VSS.n18254 VSS.n18252 0.01265
R64136 VSS.n18252 VSS.n18251 0.01265
R64137 VSS.n16867 VSS.n16861 0.01265
R64138 VSS.n16867 VSS.n16864 0.01265
R64139 VSS.n16854 VSS.n16853 0.01265
R64140 VSS.n16847 VSS.n16844 0.01265
R64141 VSS.n16840 VSS.n16839 0.01265
R64142 VSS.n16833 VSS.n16830 0.01265
R64143 VSS.n16826 VSS.n16825 0.01265
R64144 VSS.n16819 VSS.n16816 0.01265
R64145 VSS.n16812 VSS.n16811 0.01265
R64146 VSS.n16805 VSS.n16802 0.01265
R64147 VSS.n16798 VSS.n16797 0.01265
R64148 VSS.n16791 VSS.n16788 0.01265
R64149 VSS.n16784 VSS.n16783 0.01265
R64150 VSS.n16777 VSS.n16774 0.01265
R64151 VSS.n16770 VSS.n16769 0.01265
R64152 VSS.n16760 VSS.n16758 0.01265
R64153 VSS.n16758 VSS.n16757 0.01265
R64154 VSS.n16749 VSS.n16746 0.01265
R64155 VSS.n16742 VSS.n16741 0.01265
R64156 VSS.n16735 VSS.n16732 0.01265
R64157 VSS.n16728 VSS.n16727 0.01265
R64158 VSS.n16721 VSS.n16718 0.01265
R64159 VSS.n16714 VSS.n16713 0.01265
R64160 VSS.n16707 VSS.n16704 0.01265
R64161 VSS.n14949 VSS.n14946 0.01265
R64162 VSS.n14952 VSS.n14949 0.01265
R64163 VSS.n14955 VSS.n14952 0.01265
R64164 VSS.n14958 VSS.n14955 0.01265
R64165 VSS.n14959 VSS.n14958 0.01265
R64166 VSS.n19780 VSS.n19777 0.01265
R64167 VSS.n14681 VSS.n14678 0.01265
R64168 VSS.n14688 VSS.n14685 0.01265
R64169 VSS.n19789 VSS.n19786 0.01265
R64170 VSS.n14696 VSS.n14693 0.01265
R64171 VSS.n19797 VSS.n19794 0.01265
R64172 VSS.n14704 VSS.n14701 0.01265
R64173 VSS.n14711 VSS.n14708 0.01265
R64174 VSS.n14718 VSS.n14715 0.01265
R64175 VSS.n19807 VSS.n19804 0.01265
R64176 VSS.n14726 VSS.n14723 0.01265
R64177 VSS.n19815 VSS.n19812 0.01265
R64178 VSS.n19822 VSS.n19819 0.01265
R64179 VSS.n19829 VSS.n19826 0.01265
R64180 VSS.n14807 VSS.n14733 0.01265
R64181 VSS.n14806 VSS.n14804 0.01265
R64182 VSS.n14804 VSS.n14802 0.01265
R64183 VSS.n14802 VSS.n14800 0.01265
R64184 VSS.n14800 VSS.n14799 0.01265
R64185 VSS.n14799 VSS.n14797 0.01265
R64186 VSS.n14797 VSS.n14795 0.01265
R64187 VSS.n14795 VSS.n14793 0.01265
R64188 VSS.n14793 VSS.n14792 0.01265
R64189 VSS.n14792 VSS.n14790 0.01265
R64190 VSS.n14790 VSS.n14788 0.01265
R64191 VSS.n14788 VSS.n14786 0.01265
R64192 VSS.n14786 VSS.n14785 0.01265
R64193 VSS.n14785 VSS.n14783 0.01265
R64194 VSS.n14783 VSS.n14781 0.01265
R64195 VSS.n14781 VSS.n14779 0.01265
R64196 VSS.n14779 VSS.n14778 0.01265
R64197 VSS.n14778 VSS.n14776 0.01265
R64198 VSS.n14776 VSS.n14774 0.01265
R64199 VSS.n14774 VSS.n14772 0.01265
R64200 VSS.n14772 VSS.n14771 0.01265
R64201 VSS.n14771 VSS.n14769 0.01265
R64202 VSS.n14769 VSS.n14767 0.01265
R64203 VSS.n14469 VSS.n14466 0.01265
R64204 VSS.n14476 VSS.n14473 0.01265
R64205 VSS.n14483 VSS.n14480 0.01265
R64206 VSS.n14490 VSS.n14487 0.01265
R64207 VSS.n14497 VSS.n14494 0.01265
R64208 VSS.n14504 VSS.n14501 0.01265
R64209 VSS.n14511 VSS.n14508 0.01265
R64210 VSS.n14518 VSS.n14515 0.01265
R64211 VSS.n14525 VSS.n14522 0.01265
R64212 VSS.n14532 VSS.n14529 0.01265
R64213 VSS.n14539 VSS.n14536 0.01265
R64214 VSS.n14546 VSS.n14543 0.01265
R64215 VSS.n14553 VSS.n14550 0.01265
R64216 VSS.n14560 VSS.n14557 0.01265
R64217 VSS.n14587 VSS.n14450 0.01265
R64218 VSS.n14593 VSS.n14590 0.01265
R64219 VSS.n14596 VSS.n14593 0.01265
R64220 VSS.n14599 VSS.n14596 0.01265
R64221 VSS.n14602 VSS.n14599 0.01265
R64222 VSS.n14605 VSS.n14602 0.01265
R64223 VSS.n14608 VSS.n14605 0.01265
R64224 VSS.n14611 VSS.n14608 0.01265
R64225 VSS.n14614 VSS.n14611 0.01265
R64226 VSS.n14617 VSS.n14614 0.01265
R64227 VSS.n14620 VSS.n14617 0.01265
R64228 VSS.n14623 VSS.n14620 0.01265
R64229 VSS.n14626 VSS.n14623 0.01265
R64230 VSS.n14629 VSS.n14626 0.01265
R64231 VSS.n14632 VSS.n14629 0.01265
R64232 VSS.n14635 VSS.n14632 0.01265
R64233 VSS.n14638 VSS.n14635 0.01265
R64234 VSS.n14641 VSS.n14638 0.01265
R64235 VSS.n14644 VSS.n14641 0.01265
R64236 VSS.n14647 VSS.n14644 0.01265
R64237 VSS.n14650 VSS.n14647 0.01265
R64238 VSS.n14653 VSS.n14650 0.01265
R64239 VSS.n14654 VSS.n14653 0.01265
R64240 VSS.n17159 VSS.n17137 0.01265
R64241 VSS.n17159 VSS.n17157 0.01265
R64242 VSS.n17115 VSS.n17113 0.01265
R64243 VSS.n17064 VSS.n17063 0.01265
R64244 VSS.n17008 VSS.n17006 0.01265
R64245 VSS.n16968 VSS.n16966 0.01265
R64246 VSS.n16966 VSS.n16964 0.01265
R64247 VSS.n16678 VSS.n16672 0.01265
R64248 VSS.n16678 VSS.n16676 0.01265
R64249 VSS.n16665 VSS.n16663 0.01265
R64250 VSS.n16628 VSS.n16625 0.01265
R64251 VSS.n16576 VSS.n16574 0.01265
R64252 VSS.n16521 VSS.n16518 0.01265
R64253 VSS.n16507 VSS.n16505 0.01265
R64254 VSS.n16505 VSS.n16503 0.01265
R64255 VSS.n16498 VSS.n16496 0.01265
R64256 VSS.n16491 VSS.n16489 0.01265
R64257 VSS.n16484 VSS.n16482 0.01265
R64258 VSS.n16477 VSS.n16475 0.01265
R64259 VSS.n16470 VSS.n16468 0.01265
R64260 VSS.n16463 VSS.n16461 0.01265
R64261 VSS.n16456 VSS.n16454 0.01265
R64262 VSS.n16409 VSS.n16406 0.01265
R64263 VSS.n16412 VSS.n16409 0.01265
R64264 VSS.n16415 VSS.n16412 0.01265
R64265 VSS.n16418 VSS.n16415 0.01265
R64266 VSS.n16419 VSS.n16418 0.01265
R64267 VSS.n15717 VSS.n15711 0.01265
R64268 VSS.n15717 VSS.n15716 0.01265
R64269 VSS.n15724 VSS.n15722 0.01265
R64270 VSS.n15731 VSS.n15730 0.01265
R64271 VSS.n15738 VSS.n15736 0.01265
R64272 VSS.n15745 VSS.n15744 0.01265
R64273 VSS.n15752 VSS.n15750 0.01265
R64274 VSS.n15759 VSS.n15758 0.01265
R64275 VSS.n15766 VSS.n15764 0.01265
R64276 VSS.n15773 VSS.n15772 0.01265
R64277 VSS.n15780 VSS.n15778 0.01265
R64278 VSS.n15787 VSS.n15786 0.01265
R64279 VSS.n15794 VSS.n15792 0.01265
R64280 VSS.n15801 VSS.n15800 0.01265
R64281 VSS.n15808 VSS.n15806 0.01265
R64282 VSS.n15822 VSS.n15816 0.01265
R64283 VSS.n15822 VSS.n15820 0.01265
R64284 VSS.n15829 VSS.n15828 0.01265
R64285 VSS.n15836 VSS.n15834 0.01265
R64286 VSS.n15843 VSS.n15842 0.01265
R64287 VSS.n15850 VSS.n15848 0.01265
R64288 VSS.n15869 VSS.n15866 0.01265
R64289 VSS.n15872 VSS.n15869 0.01265
R64290 VSS.n15875 VSS.n15872 0.01265
R64291 VSS.n15878 VSS.n15875 0.01265
R64292 VSS.n15881 VSS.n15878 0.01265
R64293 VSS.n15884 VSS.n15881 0.01265
R64294 VSS.n15887 VSS.n15884 0.01265
R64295 VSS.n15890 VSS.n15887 0.01265
R64296 VSS.n15893 VSS.n15890 0.01265
R64297 VSS.n15894 VSS.n15893 0.01265
R64298 VSS.n9530 VSS.n9505 0.0125559
R64299 VSS.n17341 VSS.n17340 0.0125559
R64300 VSS.n17336 VSS.n17335 0.0125559
R64301 VSS.n11593 VSS.n11524 0.0125559
R64302 VSS.n11512 VSS.n4859 0.0125559
R64303 VSS.n11370 VSS.n11321 0.0125559
R64304 VSS.n13242 VSS.n13241 0.0125559
R64305 VSS.n13252 VSS.n13251 0.0125559
R64306 VSS.n13254 VSS.n13003 0.0125559
R64307 VSS.n12999 VSS.n12993 0.0125559
R64308 VSS.n12903 VSS.n12902 0.0125559
R64309 VSS.n12893 VSS.n12892 0.0125559
R64310 VSS.n12890 VSS.n12889 0.0125559
R64311 VSS.n12880 VSS.n12879 0.0125559
R64312 VSS.n12836 VSS.n12835 0.0125559
R64313 VSS.n12826 VSS.n12825 0.0125559
R64314 VSS.n12797 VSS.n12796 0.0125559
R64315 VSS.n12861 VSS.n12860 0.0125559
R64316 VSS.n12979 VSS.n12978 0.0125559
R64317 VSS.n13033 VSS.n13032 0.0125559
R64318 VSS.n13150 VSS.n13149 0.0125559
R64319 VSS.n13191 VSS.n13190 0.0125559
R64320 VSS.n17482 VSS.n2378 0.0125559
R64321 VSS.n9647 VSS.n9622 0.0125559
R64322 VSS.n9244 VSS.n9243 0.0125559
R64323 VSS.n14431 VSS.n14403 0.0125559
R64324 VSS.n14419 VSS.n14418 0.0125559
R64325 VSS.n15098 VSS.n15077 0.0125559
R64326 VSS.n15131 VSS.n15110 0.0125559
R64327 VSS.n16387 VSS.n15180 0.0125559
R64328 VSS.n2242 VSS.n2241 0.0125559
R64329 VSS.n14999 VSS.n682 0.0125559
R64330 VSS.n15149 VSS.n15148 0.0125559
R64331 VSS.n18106 VSS.n2277 0.0125559
R64332 VSS.n18880 VSS.n18879 0.0125559
R64333 VSS.n13406 VSS.n13367 0.0125559
R64334 VSS.n13420 VSS.n13418 0.0125559
R64335 VSS.n20728 VSS.n20689 0.0125559
R64336 VSS.n20779 VSS.n20740 0.0125559
R64337 VSS.n20871 VSS.n20832 0.0125559
R64338 VSS.n20605 VSS.n20604 0.0125559
R64339 VSS.n20799 VSS.n20798 0.0125559
R64340 VSS.n2337 VSS.n2330 0.0125559
R64341 VSS.n21806 VSS.n21805 0.0125559
R64342 VSS.n2290 VSS.n2289 0.0125559
R64343 VSS.n9226 VSS.n9195 0.0125559
R64344 VSS.n6564 VSS.n6563 0.0125559
R64345 VSS.n6561 VSS.n6548 0.0125559
R64346 VSS.n6834 VSS.n6812 0.0125559
R64347 VSS.n6414 VSS.n6413 0.0125559
R64348 VSS.n13502 VSS.n13501 0.0125559
R64349 VSS.n13512 VSS.n13511 0.0125559
R64350 VSS.n13514 VSS.n13436 0.0125559
R64351 VSS.n20152 VSS.n20151 0.0125559
R64352 VSS.n20068 VSS.n734 0.0125559
R64353 VSS.n2058 VSS.n2057 0.0125559
R64354 VSS.n2060 VSS.n2048 0.0125559
R64355 VSS.n2039 VSS.n2038 0.0125559
R64356 VSS.n1995 VSS.n744 0.0125559
R64357 VSS.n888 VSS.n887 0.0125559
R64358 VSS.n20166 VSS.n20143 0.0125559
R64359 VSS.n2019 VSS.n2018 0.0125559
R64360 VSS.n17966 VSS.n17938 0.0125559
R64361 VSS.n19091 VSS.n19090 0.0125559
R64362 VSS.n17898 VSS.n17897 0.0125559
R64363 VSS.n7565 VSS.n7564 0.0125559
R64364 VSS.n21282 VSS.n21281 0.0125559
R64365 VSS.n21396 VSS.n21395 0.0125559
R64366 VSS.n21481 VSS.n21480 0.0125559
R64367 VSS.n21523 VSS.n21522 0.0125559
R64368 VSS.n21577 VSS.n21576 0.0125559
R64369 VSS.n21618 VSS.n21617 0.0125559
R64370 VSS.n9320 VSS.n9194 0.0125559
R64371 VSS.n7850 VSS.n7775 0.0125559
R64372 VSS.n9157 VSS.n9051 0.0125559
R64373 VSS.n6685 VSS.n6645 0.0125559
R64374 VSS.n6535 VSS.n6495 0.0125559
R64375 VSS.n9711 VSS.n9667 0.0125559
R64376 VSS.n6904 VSS.n6855 0.0125559
R64377 VSS.n7006 VSS.n6957 0.0125559
R64378 VSS.n7688 VSS.n7687 0.0125559
R64379 VSS.n9594 VSS.n9550 0.0125559
R64380 VSS.n7600 VSS.n7599 0.0125559
R64381 VSS.n12762 VSS.n12761 0.0125559
R64382 VSS.n3811 VSS.n3810 0.0125559
R64383 VSS.n3848 VSS.n3847 0.0125559
R64384 VSS.n4755 VSS.n4731 0.0125559
R64385 VSS.n11721 VSS.n11709 0.0125559
R64386 VSS.n11440 VSS.n11439 0.0125559
R64387 VSS.n11219 VSS.n11218 0.0125559
R64388 VSS.n11184 VSS.n6152 0.0125559
R64389 VSS.n6073 VSS.n6072 0.0125559
R64390 VSS.n5992 VSS.n5991 0.0125559
R64391 VSS.n4695 VSS.n2430 0.0125559
R64392 VSS.n3288 VSS.n3259 0.0125559
R64393 VSS.n598 VSS.n597 0.0125559
R64394 VSS.n588 VSS.n587 0.0125559
R64395 VSS.n585 VSS.n584 0.0125559
R64396 VSS.n575 VSS.n574 0.0125559
R64397 VSS.n526 VSS.n525 0.0125559
R64398 VSS.n499 VSS.n498 0.0125559
R64399 VSS.n10625 VSS.n10624 0.0125559
R64400 VSS.n558 VSS.n557 0.0125559
R64401 VSS.n680 VSS.n666 0.0125559
R64402 VSS.n17441 VSS.n17440 0.0125472
R64403 VSS.n13232 VSS.n13231 0.0125472
R64404 VSS.n2192 VSS.n2191 0.0125472
R64405 VSS.n13349 VSS.n13348 0.0125472
R64406 VSS.n13492 VSS.n13491 0.0125472
R64407 VSS.n18711 VSS.n18710 0.0125423
R64408 VSS.n18734 VSS.n18733 0.0125423
R64409 VSS.n18449 VSS.n18448 0.0125423
R64410 VSS.n18176 VSS.n18175 0.0125423
R64411 VSS.n19193 VSS.n19192 0.0125423
R64412 VSS.n19216 VSS.n19215 0.0125423
R64413 VSS.n19590 VSS.n19589 0.0125423
R64414 VSS.n19680 VSS.n19679 0.0125423
R64415 VSS.n5688 VSS.n5686 0.0124681
R64416 VSS.n5673 VSS.n5672 0.0124681
R64417 VSS.n16016 VSS.n16015 0.0124681
R64418 VSS.n16007 VSS.n16006 0.0124681
R64419 VSS.n997 VSS.n996 0.0124681
R64420 VSS.n988 VSS.n987 0.0124681
R64421 VSS.n20942 VSS.n20941 0.0124681
R64422 VSS.n20957 VSS.n20955 0.0124681
R64423 VSS.n5775 VSS.n5774 0.0124681
R64424 VSS.n5827 VSS.n5826 0.0124681
R64425 VSS.n5810 VSS.n5807 0.0124681
R64426 VSS.n1199 VSS.n1198 0.0124681
R64427 VSS.n1257 VSS.n1256 0.0124681
R64428 VSS.n1241 VSS.n1239 0.0124681
R64429 VSS.n1226 VSS.n1225 0.0124681
R64430 VSS.n5549 VSS.n5548 0.0124644
R64431 VSS.n9558 VSS.n9557 0.0124644
R64432 VSS.n9121 VSS.n9120 0.0124644
R64433 VSS.n15035 VSS.n15034 0.0124644
R64434 VSS.n16059 VSS.n16058 0.0124644
R64435 VSS.n9675 VSS.n9674 0.0124644
R64436 VSS.n9284 VSS.n9283 0.0124644
R64437 VSS.n11674 VSS.n11673 0.0124644
R64438 VSS.n6117 VSS.n6116 0.0124644
R64439 VSS.n6036 VSS.n6035 0.0124644
R64440 VSS.n5955 VSS.n5954 0.0124644
R64441 VSS.n631 VSS.n630 0.0124644
R64442 VSS.n10589 VSS.n10588 0.0124644
R64443 VSS.n19251 VSS.n19248 0.012425
R64444 VSS.n19268 VSS.n19267 0.012425
R64445 VSS.n16986 VSS.n16985 0.012425
R64446 VSS.n16974 VSS.n16972 0.012425
R64447 VSS.n9063 VSS.n9060 0.0124231
R64448 VSS.n9060 VSS.n9057 0.0124231
R64449 VSS.n9078 VSS.n9069 0.0124231
R64450 VSS.n9078 VSS.n9075 0.0124231
R64451 VSS.n9075 VSS.n9072 0.0124231
R64452 VSS.n9236 VSS.n9233 0.0124231
R64453 VSS.n9242 VSS.n9236 0.0124231
R64454 VSS.n9242 VSS.n9239 0.0124231
R64455 VSS.n9225 VSS.n9222 0.0124231
R64456 VSS.n9222 VSS.n9219 0.0124231
R64457 VSS.n9213 VSS.n9210 0.0124231
R64458 VSS.n9210 VSS.n9207 0.0124231
R64459 VSS.n9207 VSS.n9204 0.0124231
R64460 VSS.n9204 VSS.n9201 0.0124231
R64461 VSS.n8146 VSS.n8143 0.0124231
R64462 VSS.n8155 VSS.n8152 0.0124231
R64463 VSS.n6392 VSS.n6389 0.0124231
R64464 VSS.n6398 VSS.n6392 0.0124231
R64465 VSS.n6398 VSS.n6397 0.0124231
R64466 VSS.n6406 VSS.n6403 0.0124231
R64467 VSS.n6412 VSS.n6406 0.0124231
R64468 VSS.n6541 VSS.n6538 0.0124231
R64469 VSS.n6547 VSS.n6541 0.0124231
R64470 VSS.n6547 VSS.n6544 0.0124231
R64471 VSS.n6560 VSS.n6557 0.0124231
R64472 VSS.n6557 VSS.n6554 0.0124231
R64473 VSS.n9511 VSS.n9508 0.0124231
R64474 VSS.n9514 VSS.n9511 0.0124231
R64475 VSS.n9517 VSS.n9514 0.0124231
R64476 VSS.n9529 VSS.n9517 0.0124231
R64477 VSS.n9529 VSS.n9526 0.0124231
R64478 VSS.n9526 VSS.n9523 0.0124231
R64479 VSS.n9628 VSS.n9625 0.0124231
R64480 VSS.n9631 VSS.n9628 0.0124231
R64481 VSS.n9634 VSS.n9631 0.0124231
R64482 VSS.n9646 VSS.n9634 0.0124231
R64483 VSS.n9646 VSS.n9643 0.0124231
R64484 VSS.n9643 VSS.n9640 0.0124231
R64485 VSS.n8493 VSS.n8490 0.0124231
R64486 VSS.n8505 VSS.n8493 0.0124231
R64487 VSS.n8505 VSS.n8502 0.0124231
R64488 VSS.n8502 VSS.n8499 0.0124231
R64489 VSS.n8644 VSS.n8641 0.0124231
R64490 VSS.n8656 VSS.n8644 0.0124231
R64491 VSS.n8656 VSS.n8653 0.0124231
R64492 VSS.n8653 VSS.n8650 0.0124231
R64493 VSS.n6818 VSS.n6815 0.0124231
R64494 VSS.n6833 VSS.n6818 0.0124231
R64495 VSS.n6833 VSS.n6830 0.0124231
R64496 VSS.n6830 VSS.n6827 0.0124231
R64497 VSS.n6827 VSS.n6824 0.0124231
R64498 VSS.n6824 VSS.n6821 0.0124231
R64499 VSS.n12615 VSS.n12612 0.0124231
R64500 VSS.n12618 VSS.n12615 0.0124231
R64501 VSS.n12621 VSS.n12618 0.0124231
R64502 VSS.n12624 VSS.n12621 0.0124231
R64503 VSS.n12627 VSS.n12624 0.0124231
R64504 VSS.n12630 VSS.n12627 0.0124231
R64505 VSS.n17472 VSS.n17471 0.0123701
R64506 VSS.n13202 VSS.n13201 0.0123701
R64507 VSS.n2223 VSS.n2222 0.0123701
R64508 VSS.n13319 VSS.n13318 0.0123701
R64509 VSS.n17949 VSS.n17948 0.0123701
R64510 VSS.n18796 VSS.n18795 0.012331
R64511 VSS.n18455 VSS.n18454 0.012331
R64512 VSS.n18185 VSS.n18184 0.012331
R64513 VSS.n17116 VSS.n17085 0.012331
R64514 VSS.n19468 VSS.n19467 0.012331
R64515 VSS.n19584 VSS.n19583 0.012331
R64516 VSS.n19671 VSS.n19670 0.012331
R64517 VSS.n19879 VSS.n19878 0.012331
R64518 VSS.n9594 VSS.n9593 0.0123034
R64519 VSS.n11370 VSS.n11369 0.0123034
R64520 VSS.n11513 VSS.n11512 0.0123034
R64521 VSS.n11593 VSS.n11592 0.0123034
R64522 VSS.n17337 VSS.n17336 0.0123034
R64523 VSS.n17340 VSS.n17339 0.0123034
R64524 VSS.n13151 VSS.n13150 0.0123034
R64525 VSS.n12761 VSS.n12760 0.0123034
R64526 VSS.n12798 VSS.n12797 0.0123034
R64527 VSS.n12827 VSS.n12826 0.0123034
R64528 VSS.n12837 VSS.n12836 0.0123034
R64529 VSS.n12881 VSS.n12880 0.0123034
R64530 VSS.n12891 VSS.n12890 0.0123034
R64531 VSS.n12894 VSS.n12893 0.0123034
R64532 VSS.n12904 VSS.n12903 0.0123034
R64533 VSS.n12999 VSS.n12998 0.0123034
R64534 VSS.n13254 VSS.n13253 0.0123034
R64535 VSS.n13251 VSS.n13250 0.0123034
R64536 VSS.n13241 VSS.n13240 0.0123034
R64537 VSS.n12980 VSS.n12979 0.0123034
R64538 VSS.n12860 VSS.n12859 0.0123034
R64539 VSS.n13034 VSS.n13033 0.0123034
R64540 VSS.n17482 VSS.n17481 0.0123034
R64541 VSS.n13192 VSS.n13191 0.0123034
R64542 VSS.n15150 VSS.n15149 0.0123034
R64543 VSS.n9711 VSS.n9710 0.0123034
R64544 VSS.n14431 VSS.n14430 0.0123034
R64545 VSS.n14418 VSS.n14417 0.0123034
R64546 VSS.n14404 VSS.n682 0.0123034
R64547 VSS.n15099 VSS.n15098 0.0123034
R64548 VSS.n15132 VSS.n15131 0.0123034
R64549 VSS.n16387 VSS.n16386 0.0123034
R64550 VSS.n2241 VSS.n2240 0.0123034
R64551 VSS.n18879 VSS.n18878 0.0123034
R64552 VSS.n18107 VSS.n18106 0.0123034
R64553 VSS.n2291 VSS.n2290 0.0123034
R64554 VSS.n20800 VSS.n20799 0.0123034
R64555 VSS.n13407 VSS.n13406 0.0123034
R64556 VSS.n13420 VSS.n13419 0.0123034
R64557 VSS.n20729 VSS.n20728 0.0123034
R64558 VSS.n20780 VSS.n20779 0.0123034
R64559 VSS.n20872 VSS.n20871 0.0123034
R64560 VSS.n20604 VSS.n20603 0.0123034
R64561 VSS.n21807 VSS.n21806 0.0123034
R64562 VSS.n2337 VSS.n2336 0.0123034
R64563 VSS.n17899 VSS.n17898 0.0123034
R64564 VSS.n20166 VSS.n20165 0.0123034
R64565 VSS.n20151 VSS.n20150 0.0123034
R64566 VSS.n13514 VSS.n13513 0.0123034
R64567 VSS.n13511 VSS.n13510 0.0123034
R64568 VSS.n13501 VSS.n13500 0.0123034
R64569 VSS.n887 VSS.n886 0.0123034
R64570 VSS.n1996 VSS.n1995 0.0123034
R64571 VSS.n2020 VSS.n2019 0.0123034
R64572 VSS.n2040 VSS.n2039 0.0123034
R64573 VSS.n2060 VSS.n2059 0.0123034
R64574 VSS.n2057 VSS.n2056 0.0123034
R64575 VSS.n20069 VSS.n20068 0.0123034
R64576 VSS.n19092 VSS.n19091 0.0123034
R64577 VSS.n17966 VSS.n17965 0.0123034
R64578 VSS.n21522 VSS.n21521 0.0123034
R64579 VSS.n7601 VSS.n7600 0.0123034
R64580 VSS.n7689 VSS.n7688 0.0123034
R64581 VSS.n7564 VSS.n7563 0.0123034
R64582 VSS.n21397 VSS.n21396 0.0123034
R64583 VSS.n21281 VSS.n21280 0.0123034
R64584 VSS.n21482 VSS.n21481 0.0123034
R64585 VSS.n21619 VSS.n21618 0.0123034
R64586 VSS.n21578 VSS.n21577 0.0123034
R64587 VSS.n7850 VSS.n7849 0.0123034
R64588 VSS.n9320 VSS.n9319 0.0123034
R64589 VSS.n9157 VSS.n9156 0.0123034
R64590 VSS.n6685 VSS.n6684 0.0123034
R64591 VSS.n6535 VSS.n6534 0.0123034
R64592 VSS.n7006 VSS.n7005 0.0123034
R64593 VSS.n6904 VSS.n6903 0.0123034
R64594 VSS.n4696 VSS.n4695 0.0123034
R64595 VSS.n11439 VSS.n11438 0.0123034
R64596 VSS.n5991 VSS.n5990 0.0123034
R64597 VSS.n3810 VSS.n3809 0.0123034
R64598 VSS.n11722 VSS.n11721 0.0123034
R64599 VSS.n11185 VSS.n11184 0.0123034
R64600 VSS.n6072 VSS.n6071 0.0123034
R64601 VSS.n3847 VSS.n3846 0.0123034
R64602 VSS.n11218 VSS.n11217 0.0123034
R64603 VSS.n4756 VSS.n4755 0.0123034
R64604 VSS.n3288 VSS.n3287 0.0123034
R64605 VSS.n576 VSS.n575 0.0123034
R64606 VSS.n586 VSS.n585 0.0123034
R64607 VSS.n589 VSS.n588 0.0123034
R64608 VSS.n599 VSS.n598 0.0123034
R64609 VSS.n680 VSS.n679 0.0123034
R64610 VSS.n557 VSS.n556 0.0123034
R64611 VSS.n525 VSS.n524 0.0123034
R64612 VSS.n498 VSS.n497 0.0123034
R64613 VSS.n9531 VSS.n9530 0.0123034
R64614 VSS.n9648 VSS.n9647 0.0123034
R64615 VSS.n6835 VSS.n6834 0.0123034
R64616 VSS.n6563 VSS.n6562 0.0123034
R64617 VSS.n6562 VSS.n6561 0.0123034
R64618 VSS.n6413 VSS.n6400 0.0123034
R64619 VSS.n9243 VSS.n9227 0.0123034
R64620 VSS.n9227 VSS.n9226 0.0123034
R64621 VSS.n14238 VSS.n14237 0.0122524
R64622 VSS.n18379 VSS.n18378 0.0122
R64623 VSS.n16563 VSS.n16561 0.0122
R64624 VSS.n15320 VSS.n15319 0.0120643
R64625 VSS.n8536 VSS.n8535 0.0120643
R64626 VSS.n8391 VSS.n8390 0.0120643
R64627 VSS.n8390 VSS.n8389 0.0120643
R64628 VSS.n8535 VSS.n8534 0.0120643
R64629 VSS.n15321 VSS.n15320 0.0120643
R64630 VSS.n1636 VSS.n1635 0.0120643
R64631 VSS.n8687 VSS.n8686 0.0120643
R64632 VSS.n8199 VSS.n8198 0.0120643
R64633 VSS.n8686 VSS.n8685 0.0120643
R64634 VSS.n8198 VSS.n8197 0.0120643
R64635 VSS.n1637 VSS.n1636 0.0120643
R64636 VSS.n17109 VSS.n17108 0.011975
R64637 VSS.n17052 VSS.n17050 0.011975
R64638 VSS.n16954 VSS.n16952 0.011975
R64639 VSS.n14914 VSS.n14911 0.011975
R64640 VSS.n4008 VSS.n4007 0.0119309
R64641 VSS.n17350 VSS.n17338 0.0119309
R64642 VSS.n17326 VSS.n17325 0.0119309
R64643 VSS.n17312 VSS.n681 0.0119309
R64644 VSS.n11515 VSS.n11514 0.0119309
R64645 VSS.n11331 VSS.n11330 0.0119309
R64646 VSS.n11348 VSS.n11347 0.0119309
R64647 VSS.n11312 VSS.n11311 0.0119309
R64648 VSS.n17350 VSS.n17349 0.0119309
R64649 VSS.n17327 VSS.n17326 0.0119309
R64650 VSS.n11516 VSS.n11515 0.0119309
R64651 VSS.n11330 VSS.n11329 0.0119309
R64652 VSS.n11313 VSS.n11312 0.0119309
R64653 VSS.n4211 VSS.n4210 0.0119309
R64654 VSS.n11349 VSS.n11348 0.0119309
R64655 VSS.n11525 VSS.n681 0.0119309
R64656 VSS.n4009 VSS.n4008 0.0119309
R64657 VSS.n6399 VSS.n6380 0.0119309
R64658 VSS.n6400 VSS.n6399 0.0119309
R64659 VSS.n16637 VSS.n16636 0.0119085
R64660 VSS.n761 VSS.n760 0.0119085
R64661 VSS.n2429 VSS.n2428 0.0117632
R64662 VSS.n19399 VSS.n19397 0.01175
R64663 VSS.n19385 VSS.n19384 0.01175
R64664 VSS.n18267 VSS.n18266 0.01175
R64665 VSS.n16657 VSS.n16655 0.01175
R64666 VSS.n16621 VSS.n16620 0.01175
R64667 VSS.n18723 VSS.n18722 0.0116972
R64668 VSS.n17010 VSS.n17009 0.0116972
R64669 VSS.n14898 VSS.n14897 0.0116972
R64670 VSS.n8479 VSS.n8478 0.0116972
R64671 VSS.n19205 VSS.n19204 0.0116972
R64672 VSS.n19925 VSS.n19924 0.0116972
R64673 VSS.n19969 VSS.n19968 0.0116972
R64674 VSS.n8630 VSS.n8629 0.0116972
R64675 VSS.n21700 VSS.n21699 0.0116937
R64676 VSS.n367 VSS.n366 0.0116937
R64677 VSS.n21916 VSS.n21915 0.0116937
R64678 VSS.n14568 VSS.n14567 0.0115386
R64679 VSS.n14827 VSS.n14826 0.0115386
R64680 VSS.n16881 VSS.n16880 0.0115386
R64681 VSS.n16692 VSS.n16691 0.0115386
R64682 VSS.n16441 VSS.n16440 0.0115386
R64683 VSS.n16442 VSS.n16441 0.0115386
R64684 VSS.n14569 VSS.n14568 0.0115386
R64685 VSS.n14826 VSS.n14825 0.0115386
R64686 VSS.n16882 VSS.n16881 0.0115386
R64687 VSS.n16693 VSS.n16692 0.0115386
R64688 VSS.n19760 VSS.n19759 0.0115386
R64689 VSS.n19850 VSS.n19849 0.0115386
R64690 VSS.n20035 VSS.n20034 0.0115386
R64691 VSS.n2094 VSS.n2093 0.0115386
R64692 VSS.n848 VSS.n847 0.0115386
R64693 VSS.n19849 VSS.n19848 0.0115386
R64694 VSS.n19759 VSS.n19758 0.0115386
R64695 VSS.n847 VSS.n846 0.0115386
R64696 VSS.n2095 VSS.n2094 0.0115386
R64697 VSS.n20034 VSS.n20033 0.0115386
R64698 VSS.n17151 VSS.n17149 0.011525
R64699 VSS.n17002 VSS.n17001 0.011525
R64700 VSS.n16995 VSS.n16993 0.011525
R64701 VSS.n18824 VSS.n18823 0.0114859
R64702 VSS.n18406 VSS.n18405 0.0114859
R64703 VSS.n17009 VSS.n14834 0.0114859
R64704 VSS.n19496 VSS.n19495 0.0114859
R64705 VSS.n19616 VSS.n19615 0.0114859
R64706 VSS.n19926 VSS.n19925 0.0114859
R64707 VSS.n3987 VSS.n3986 0.0114843
R64708 VSS.n5842 VSS.n5841 0.0114843
R64709 VSS.n5562 VSS.n5561 0.0114843
R64710 VSS.n13013 VSS.n13012 0.0114843
R64711 VSS.n12592 VSS.n12591 0.0114843
R64712 VSS.n12583 VSS.n12582 0.0114843
R64713 VSS.n12577 VSS.n12576 0.0114843
R64714 VSS.n12562 VSS.n12561 0.0114843
R64715 VSS.n12553 VSS.n12552 0.0114843
R64716 VSS.n12516 VSS.n12515 0.0114843
R64717 VSS.n12507 VSS.n12506 0.0114843
R64718 VSS.n12326 VSS.n12325 0.0114843
R64719 VSS.n12317 VSS.n12316 0.0114843
R64720 VSS.n12308 VSS.n12307 0.0114843
R64721 VSS.n12282 VSS.n12281 0.0114843
R64722 VSS.n12273 VSS.n12272 0.0114843
R64723 VSS.n12259 VSS.n12258 0.0114843
R64724 VSS.n12250 VSS.n12249 0.0114843
R64725 VSS.n11971 VSS.n11970 0.0114843
R64726 VSS.n11964 VSS.n11963 0.0114843
R64727 VSS.n11935 VSS.n11934 0.0114843
R64728 VSS.n11928 VSS.n11927 0.0114843
R64729 VSS.n11912 VSS.n11911 0.0114843
R64730 VSS.n11881 VSS.n11880 0.0114843
R64731 VSS.n11874 VSS.n11873 0.0114843
R64732 VSS.n11865 VSS.n11864 0.0114843
R64733 VSS.n11841 VSS.n11840 0.0114843
R64734 VSS.n11832 VSS.n11831 0.0114843
R64735 VSS.n11818 VSS.n11817 0.0114843
R64736 VSS.n11809 VSS.n11808 0.0114843
R64737 VSS.n18858 VSS.n18857 0.0114843
R64738 VSS.n16203 VSS.n16202 0.0114843
R64739 VSS.n16072 VSS.n16071 0.0114843
R64740 VSS.n21786 VSS.n21785 0.0114843
R64741 VSS.n21145 VSS.n21144 0.0114843
R64742 VSS.n21011 VSS.n21010 0.0114843
R64743 VSS.n19071 VSS.n19070 0.0114843
R64744 VSS.n1274 VSS.n1273 0.0114843
R64745 VSS.n1057 VSS.n1056 0.0114843
R64746 VSS.n21554 VSS.n21553 0.0114843
R64747 VSS.n21534 VSS.n21533 0.0114843
R64748 VSS.n21470 VSS.n21469 0.0114843
R64749 VSS.n3787 VSS.n3786 0.0114843
R64750 VSS.n4150 VSS.n4149 0.0114843
R64751 VSS.n4766 VSS.n4765 0.0114843
R64752 VSS.n3267 VSS.n3266 0.0114843
R64753 VSS.n10526 VSS.n10525 0.0114843
R64754 VSS.n10518 VSS.n10517 0.0114843
R64755 VSS.n10512 VSS.n10511 0.0114843
R64756 VSS.n10506 VSS.n10505 0.0114843
R64757 VSS.n10498 VSS.n10497 0.0114843
R64758 VSS.n10461 VSS.n10460 0.0114843
R64759 VSS.n10453 VSS.n10452 0.0114843
R64760 VSS.n10272 VSS.n10271 0.0114843
R64761 VSS.n10264 VSS.n10263 0.0114843
R64762 VSS.n10256 VSS.n10255 0.0114843
R64763 VSS.n10230 VSS.n10229 0.0114843
R64764 VSS.n10222 VSS.n10221 0.0114843
R64765 VSS.n10207 VSS.n10206 0.0114843
R64766 VSS.n10199 VSS.n10198 0.0114843
R64767 VSS.n9974 VSS.n9973 0.0114843
R64768 VSS.n9967 VSS.n9966 0.0114843
R64769 VSS.n9936 VSS.n9935 0.0114843
R64770 VSS.n9929 VSS.n9928 0.0114843
R64771 VSS.n9913 VSS.n9912 0.0114843
R64772 VSS.n8943 VSS.n8942 0.0114843
R64773 VSS.n8787 VSS.n8786 0.0114843
R64774 VSS.n15701 VSS.n15700 0.0113101
R64775 VSS.n4066 VSS.n4065 0.0113071
R64776 VSS.n13094 VSS.n13093 0.0113071
R64777 VSS.n12674 VSS.n12673 0.0113071
R64778 VSS.n12525 VSS.n12524 0.0113071
R64779 VSS.n12265 VSS.n12264 0.0113071
R64780 VSS.n11919 VSS.n11918 0.0113071
R64781 VSS.n11895 VSS.n11894 0.0113071
R64782 VSS.n18937 VSS.n18936 0.0113071
R64783 VSS.n21867 VSS.n21866 0.0113071
R64784 VSS.n19152 VSS.n19151 0.0113071
R64785 VSS.n21436 VSS.n21435 0.0113071
R64786 VSS.n17392 VSS.n17391 0.0113071
R64787 VSS.n2622 VSS.n2621 0.0113071
R64788 VSS.n10542 VSS.n10541 0.0113071
R64789 VSS.n10470 VSS.n10469 0.0113071
R64790 VSS.n10213 VSS.n10212 0.0113071
R64791 VSS.n9920 VSS.n9919 0.0113071
R64792 VSS.n14205 VSS.n14204 0.0113
R64793 VSS.n19406 VSS.n19405 0.0113
R64794 VSS.n18260 VSS.n18258 0.0113
R64795 VSS.n16615 VSS.n16613 0.0113
R64796 VSS.n16514 VSS.n16513 0.0113
R64797 VSS.n18679 VSS.n18678 0.0112746
R64798 VSS.n19524 VSS.n19523 0.0112746
R64799 VSS.n8517 VSS.n8516 0.0112232
R64800 VSS.n8518 VSS.n8517 0.0112232
R64801 VSS.n8669 VSS.n8668 0.0112232
R64802 VSS.n8668 VSS.n8667 0.0112232
R64803 VSS.n11790 VSS.n11789 0.0111514
R64804 VSS.n1467 VSS.n889 0.0111514
R64805 VSS.n21192 VSS.n20873 0.0111514
R64806 VSS.n12823 VSS.n12822 0.0111514
R64807 VSS.n16385 VSS.n16384 0.0111514
R64808 VSS.n11309 VSS.n5882 0.0111514
R64809 VSS.n523 VSS.n522 0.0111514
R64810 VSS.n8895 VSS.n8894 0.0111514
R64811 VSS.n8893 VSS.n8892 0.0111514
R64812 VSS.n8890 VSS.n8889 0.0111514
R64813 VSS.n11787 VSS.n11786 0.0111514
R64814 VSS.n11791 VSS.n11790 0.0111514
R64815 VSS.n9543 VSS.n9542 0.0111389
R64816 VSS.n9660 VSS.n9659 0.0111389
R64817 VSS.n11849 VSS.n11848 0.0111299
R64818 VSS.n11826 VSS.n11825 0.0111299
R64819 VSS.n17103 VSS.n17101 0.011075
R64820 VSS.n17059 VSS.n17058 0.011075
R64821 VSS.n16960 VSS.n16959 0.011075
R64822 VSS.n14923 VSS.n14922 0.011075
R64823 VSS.n18473 VSS.n18472 0.0110634
R64824 VSS.n19566 VSS.n19565 0.0110634
R64825 VSS.n12298 VSS.n12297 0.0109528
R64826 VSS.n12240 VSS.n12239 0.0109528
R64827 VSS.n11949 VSS.n11948 0.0109528
R64828 VSS.n11793 VSS.n11792 0.0109528
R64829 VSS.n21651 VSS.n21650 0.0109528
R64830 VSS.n3880 VSS.n3879 0.0109528
R64831 VSS.n10246 VSS.n10245 0.0109528
R64832 VSS.n10189 VSS.n10188 0.0109528
R64833 VSS.n9951 VSS.n9950 0.0109528
R64834 VSS.n8896 VSS.n8895 0.0109528
R64835 VSS.n11792 VSS.n11791 0.0108992
R64836 VSS.n11788 VSS.n11787 0.0108992
R64837 VSS.n1467 VSS.n1466 0.0108992
R64838 VSS.n12824 VSS.n12823 0.0108992
R64839 VSS.n21192 VSS.n21191 0.0108992
R64840 VSS.n16384 VSS.n16383 0.0108992
R64841 VSS.n11310 VSS.n11309 0.0108992
R64842 VSS.n522 VSS.n521 0.0108992
R64843 VSS.n11789 VSS.n11788 0.0108992
R64844 VSS.n8894 VSS.n8893 0.0108992
R64845 VSS.n8892 VSS.n8891 0.0108992
R64846 VSS.n8891 VSS.n8890 0.0108992
R64847 VSS.n9868 VSS.n9867 0.0108846
R64848 VSS.n10298 VSS.n10293 0.0108846
R64849 VSS.n10299 VSS.n10298 0.0108846
R64850 VSS.n10448 VSS.n10323 0.0108846
R64851 VSS.n10448 VSS.n10441 0.0108846
R64852 VSS.n10417 VSS.n10416 0.0108846
R64853 VSS.n10416 VSS.n10411 0.0108846
R64854 VSS.n10355 VSS.n10354 0.0108846
R64855 VSS.n10354 VSS.n10349 0.0108846
R64856 VSS.n10333 VSS.n10332 0.0108846
R64857 VSS.n10332 VSS.n10327 0.0108846
R64858 VSS.n10327 VSS.n10326 0.0108846
R64859 VSS.n10163 VSS.n9976 0.0108846
R64860 VSS.n10163 VSS.n10156 0.0108846
R64861 VSS.n10132 VSS.n10131 0.0108846
R64862 VSS.n10131 VSS.n10126 0.0108846
R64863 VSS.n10070 VSS.n10069 0.0108846
R64864 VSS.n10069 VSS.n10064 0.0108846
R64865 VSS.n10016 VSS.n10015 0.0108846
R64866 VSS.n10015 VSS.n10010 0.0108846
R64867 VSS.n12672 VSS.n12657 0.0108846
R64868 VSS.n12352 VSS.n12347 0.0108846
R64869 VSS.n12353 VSS.n12352 0.0108846
R64870 VSS.n12502 VSS.n12377 0.0108846
R64871 VSS.n12502 VSS.n12495 0.0108846
R64872 VSS.n12471 VSS.n12470 0.0108846
R64873 VSS.n12470 VSS.n12465 0.0108846
R64874 VSS.n12409 VSS.n12408 0.0108846
R64875 VSS.n12408 VSS.n12403 0.0108846
R64876 VSS.n12387 VSS.n12386 0.0108846
R64877 VSS.n12386 VSS.n12381 0.0108846
R64878 VSS.n12381 VSS.n12380 0.0108846
R64879 VSS.n12214 VSS.n11973 0.0108846
R64880 VSS.n12214 VSS.n12207 0.0108846
R64881 VSS.n12183 VSS.n12182 0.0108846
R64882 VSS.n12182 VSS.n12177 0.0108846
R64883 VSS.n12121 VSS.n12120 0.0108846
R64884 VSS.n12120 VSS.n12115 0.0108846
R64885 VSS.n12067 VSS.n12066 0.0108846
R64886 VSS.n12066 VSS.n12061 0.0108846
R64887 VSS.n18788 VSS.n18787 0.0108521
R64888 VSS.n18797 VSS.n18796 0.0108521
R64889 VSS.n18454 VSS.n18453 0.0108521
R64890 VSS.n18184 VSS.n18183 0.0108521
R64891 VSS.n18148 VSS.n18147 0.0108521
R64892 VSS.n17117 VSS.n17116 0.0108521
R64893 VSS.n19460 VSS.n19459 0.0108521
R64894 VSS.n19469 VSS.n19468 0.0108521
R64895 VSS.n19585 VSS.n19584 0.0108521
R64896 VSS.n19672 VSS.n19671 0.0108521
R64897 VSS.n19708 VSS.n19707 0.0108521
R64898 VSS.n19878 VSS.n19877 0.0108521
R64899 VSS.n18370 VSS.n18367 0.01085
R64900 VSS.n16569 VSS.n16568 0.01085
R64901 VSS.n11564 VSS.n11563 0.0107895
R64902 VSS.n5546 VSS.n5545 0.0107895
R64903 VSS.n9555 VSS.n9554 0.0107895
R64904 VSS.n9118 VSS.n9117 0.0107895
R64905 VSS.n16056 VSS.n16055 0.0107895
R64906 VSS.n9672 VSS.n9671 0.0107895
R64907 VSS.n9281 VSS.n9280 0.0107895
R64908 VSS.n6114 VSS.n6113 0.0107895
R64909 VSS.n6033 VSS.n6032 0.0107895
R64910 VSS.n5952 VSS.n5951 0.0107895
R64911 VSS.n628 VSS.n627 0.0107895
R64912 VSS.n10586 VSS.n10585 0.0107895
R64913 VSS.n11411 VSS.n11409 0.0107778
R64914 VSS.n20842 VSS.n20841 0.0107778
R64915 VSS.n11473 VSS.n11472 0.0107778
R64916 VSS.n20750 VSS.n20749 0.0107778
R64917 VSS.n11634 VSS.n11632 0.0107778
R64918 VSS.n20699 VSS.n20698 0.0107778
R64919 VSS.n17235 VSS.n17234 0.0107778
R64920 VSS.n13258 VSS.n13257 0.0107778
R64921 VSS.n17380 VSS.n17378 0.0107778
R64922 VSS.n13377 VSS.n13376 0.0107778
R64923 VSS.n5608 VSS.n5607 0.0107756
R64924 VSS.n12544 VSS.n12543 0.0107756
R64925 VSS.n16124 VSS.n16123 0.0107756
R64926 VSS.n21058 VSS.n21057 0.0107756
R64927 VSS.n1104 VSS.n1103 0.0107756
R64928 VSS.n21631 VSS.n21630 0.0107756
R64929 VSS.n3859 VSS.n3858 0.0107756
R64930 VSS.n10489 VSS.n10488 0.0107756
R64931 VSS.n6939 VSS.n6938 0.010723
R64932 VSS.n6938 VSS.n6937 0.010723
R64933 VSS.n11537 VSS.n11536 0.010701
R64934 VSS.n11589 VSS.n11588 0.010701
R64935 VSS.n5586 VSS.n5585 0.010701
R64936 VSS.n9582 VSS.n9581 0.010701
R64937 VSS.n9145 VSS.n9144 0.010701
R64938 VSS.n15011 VSS.n15010 0.010701
R64939 VSS.n16102 VSS.n16101 0.010701
R64940 VSS.n9699 VSS.n9698 0.010701
R64941 VSS.n9308 VSS.n9307 0.010701
R64942 VSS.n15064 VSS.n15063 0.010701
R64943 VSS.n9179 VSS.n9178 0.010701
R64944 VSS.n9036 VSS.n9035 0.010701
R64945 VSS.n11698 VSS.n11697 0.010701
R64946 VSS.n6141 VSS.n6140 0.010701
R64947 VSS.n6060 VSS.n6059 0.010701
R64948 VSS.n5979 VSS.n5978 0.010701
R64949 VSS.n5927 VSS.n5926 0.010701
R64950 VSS.n6008 VSS.n6007 0.010701
R64951 VSS.n11645 VSS.n11644 0.010701
R64952 VSS.n6089 VSS.n6088 0.010701
R64953 VSS.n655 VSS.n654 0.010701
R64954 VSS.n603 VSS.n602 0.010701
R64955 VSS.n10613 VSS.n10612 0.010701
R64956 VSS.n10529 VSS.n10528 0.0106923
R64957 VSS.n10380 VSS.n10379 0.0106923
R64958 VSS.n10363 VSS.n10362 0.0106923
R64959 VSS.n10095 VSS.n10094 0.0106923
R64960 VSS.n10078 VSS.n10077 0.0106923
R64961 VSS.n10003 VSS.n10002 0.0106923
R64962 VSS.n9986 VSS.n9985 0.0106923
R64963 VSS.n12595 VSS.n12594 0.0106923
R64964 VSS.n12434 VSS.n12433 0.0106923
R64965 VSS.n12417 VSS.n12416 0.0106923
R64966 VSS.n12146 VSS.n12145 0.0106923
R64967 VSS.n12129 VSS.n12128 0.0106923
R64968 VSS.n12054 VSS.n12053 0.0106923
R64969 VSS.n12037 VSS.n12036 0.0106923
R64970 VSS.n11984 VSS.n11983 0.0106727
R64971 VSS.n18712 VSS.n18711 0.0106408
R64972 VSS.n16940 VSS.n16939 0.0106408
R64973 VSS.n16897 VSS.n16896 0.0106408
R64974 VSS.n19194 VSS.n19193 0.0106408
R64975 VSS.n19976 VSS.n19975 0.0106408
R64976 VSS.n20019 VSS.n20018 0.0106408
R64977 VSS.n19259 VSS.n19256 0.010625
R64978 VSS.n19260 VSS.n19259 0.010625
R64979 VSS.n16981 VSS.n16980 0.010625
R64980 VSS.n16980 VSS.n16978 0.010625
R64981 VSS.n4032 VSS.n4031 0.0106125
R64982 VSS.n2367 VSS.n2366 0.0106125
R64983 VSS.n5861 VSS.n5860 0.0106125
R64984 VSS.n11336 VSS.n11335 0.0106125
R64985 VSS.n18903 VSS.n18902 0.0106125
R64986 VSS.n2266 VSS.n2265 0.0106125
R64987 VSS.n15137 VSS.n15136 0.0106125
R64988 VSS.n16222 VSS.n16221 0.0106125
R64989 VSS.n9256 VSS.n9255 0.0106125
R64990 VSS.n3834 VSS.n3833 0.0106125
R64991 VSS.n4720 VSS.n4719 0.0106125
R64992 VSS.n11452 VSS.n11451 0.0106125
R64993 VSS.n11231 VSS.n11230 0.0106125
R64994 VSS.n2649 VSS.n2648 0.0106125
R64995 VSS.n570 VSS.n569 0.0106125
R64996 VSS.n511 VSS.n510 0.0106125
R64997 VSS.n3998 VSS.n3997 0.0105984
R64998 VSS.n4210 VSS.n4209 0.0105984
R64999 VSS.n13023 VSS.n13022 0.0105984
R65000 VSS.n13149 VSS.n13148 0.0105984
R65001 VSS.n11950 VSS.n11949 0.0105984
R65002 VSS.n18869 VSS.n18868 0.0105984
R65003 VSS.n2240 VSS.n2239 0.0105984
R65004 VSS.n21796 VSS.n21795 0.0105984
R65005 VSS.n2289 VSS.n2288 0.0105984
R65006 VSS.n19081 VSS.n19080 0.0105984
R65007 VSS.n17897 VSS.n17896 0.0105984
R65008 VSS.n21567 VSS.n21566 0.0105984
R65009 VSS.n3800 VSS.n3799 0.0105984
R65010 VSS.n3278 VSS.n3277 0.0105984
R65011 VSS.n9952 VSS.n9951 0.0105984
R65012 VSS.n8869 VSS.n8868 0.01057
R65013 VSS.n149 VSS.n148 0.0105559
R65014 VSS.n129 VSS.n127 0.0105559
R65015 VSS.n118 VSS.n117 0.0105559
R65016 VSS.n98 VSS.n96 0.0105559
R65017 VSS.n86 VSS.n85 0.0105559
R65018 VSS.n66 VSS.n64 0.0105559
R65019 VSS.n231 VSS.n229 0.0105559
R65020 VSS.n251 VSS.n250 0.0105559
R65021 VSS.n263 VSS.n261 0.0105559
R65022 VSS.n283 VSS.n282 0.0105559
R65023 VSS.n295 VSS.n293 0.0105559
R65024 VSS.n315 VSS.n314 0.0105559
R65025 VSS.n17243 VSS.n17242 0.0105466
R65026 VSS.n11737 VSS.n11736 0.0105466
R65027 VSS.n4929 VSS.n4928 0.0105466
R65028 VSS.n11458 VSS.n11457 0.0105466
R65029 VSS.n11247 VSS.n11246 0.0105466
R65030 VSS.n11248 VSS.n11247 0.0105466
R65031 VSS.n11457 VSS.n11456 0.0105466
R65032 VSS.n4930 VSS.n4929 0.0105466
R65033 VSS.n11736 VSS.n11735 0.0105466
R65034 VSS.n17242 VSS.n17241 0.0105466
R65035 VSS.n21430 VSS.n21429 0.0105264
R65036 VSS.n21422 VSS.n21421 0.0105264
R65037 VSS.n21419 VSS.n21418 0.0105264
R65038 VSS.n21411 VSS.n21410 0.0105264
R65039 VSS.n21320 VSS.n21319 0.0105264
R65040 VSS.n21312 VSS.n21311 0.0105264
R65041 VSS.n21309 VSS.n21308 0.0105264
R65042 VSS.n21301 VSS.n21300 0.0105264
R65043 VSS.n21257 VSS.n21256 0.0105264
R65044 VSS.n21249 VSS.n21248 0.0105264
R65045 VSS.n21247 VSS.n21246 0.0105264
R65046 VSS.n21431 VSS.n21430 0.0105264
R65047 VSS.n21423 VSS.n21422 0.0105264
R65048 VSS.n21420 VSS.n21419 0.0105264
R65049 VSS.n21412 VSS.n21411 0.0105264
R65050 VSS.n21321 VSS.n21320 0.0105264
R65051 VSS.n21313 VSS.n21312 0.0105264
R65052 VSS.n21310 VSS.n21309 0.0105264
R65053 VSS.n21302 VSS.n21301 0.0105264
R65054 VSS.n21258 VSS.n21257 0.0105264
R65055 VSS.n21250 VSS.n21249 0.0105264
R65056 VSS.n21246 VSS.n445 0.0105264
R65057 VSS.n17387 VSS.n17386 0.0105264
R65058 VSS.n17240 VSS.n17239 0.0105264
R65059 VSS.n11641 VSS.n11640 0.0105264
R65060 VSS.n11465 VSS.n4931 0.0105264
R65061 VSS.n11418 VSS.n11417 0.0105264
R65062 VSS.n11250 VSS.n11240 0.0105264
R65063 VSS.n17386 VSS.n17249 0.0105264
R65064 VSS.n17239 VSS.n11743 0.0105264
R65065 VSS.n11640 VSS.n4797 0.0105264
R65066 VSS.n11465 VSS.n11464 0.0105264
R65067 VSS.n11417 VSS.n5414 0.0105264
R65068 VSS.n11250 VSS.n11249 0.0105264
R65069 VSS.n3984 VSS.n3983 0.010524
R65070 VSS.n11362 VSS.n11361 0.010524
R65071 VSS.n5731 VSS.n5730 0.010524
R65072 VSS.n2356 VSS.n2355 0.010524
R65073 VSS.n18855 VSS.n18854 0.010524
R65074 VSS.n2255 VSS.n2254 0.010524
R65075 VSS.n16179 VSS.n16178 0.010524
R65076 VSS.n15163 VSS.n15162 0.010524
R65077 VSS.n3784 VSS.n3783 0.010524
R65078 VSS.n4709 VSS.n4708 0.010524
R65079 VSS.n11205 VSS.n11204 0.010524
R65080 VSS.n11426 VSS.n11425 0.010524
R65081 VSS.n3264 VSS.n3263 0.010524
R65082 VSS.n485 VSS.n484 0.010524
R65083 VSS.n544 VSS.n543 0.010524
R65084 VSS.n3366 VSS.n3365 0.0105
R65085 VSS.n3405 VSS.n3404 0.0105
R65086 VSS.n3404 VSS.n3403 0.0105
R65087 VSS.n3403 VSS.n3402 0.0105
R65088 VSS.n3413 VSS.n3412 0.0105
R65089 VSS.n3417 VSS.n3416 0.0105
R65090 VSS.n3489 VSS.n3488 0.0105
R65091 VSS.n3501 VSS.n3500 0.0105
R65092 VSS.n3500 VSS.n3499 0.0105
R65093 VSS.n3499 VSS.n3498 0.0105
R65094 VSS.n3508 VSS.n3507 0.0105
R65095 VSS.n3546 VSS.n3545 0.0105
R65096 VSS.n3603 VSS.n3602 0.0105
R65097 VSS.n3224 VSS.n3222 0.0105
R65098 VSS.n3226 VSS.n3224 0.0105
R65099 VSS.n3228 VSS.n3226 0.0105
R65100 VSS.n3231 VSS.n3228 0.0105
R65101 VSS.n3307 VSS.n3305 0.0105
R65102 VSS.n3309 VSS.n3307 0.0105
R65103 VSS.n3311 VSS.n3309 0.0105
R65104 VSS.n3314 VSS.n3311 0.0105
R65105 VSS.n3345 VSS.n3343 0.0105
R65106 VSS.n3347 VSS.n3345 0.0105
R65107 VSS.n3349 VSS.n3347 0.0105
R65108 VSS.n3351 VSS.n3349 0.0105
R65109 VSS.n3353 VSS.n3351 0.0105
R65110 VSS.n3355 VSS.n3353 0.0105
R65111 VSS.n3357 VSS.n3355 0.0105
R65112 VSS.n3359 VSS.n3357 0.0105
R65113 VSS.n3361 VSS.n3359 0.0105
R65114 VSS.n3363 VSS.n3361 0.0105
R65115 VSS.n3367 VSS.n3363 0.0105
R65116 VSS.n3368 VSS.n3367 0.0105
R65117 VSS.n3399 VSS.n3397 0.0105
R65118 VSS.n3401 VSS.n3399 0.0105
R65119 VSS.n3406 VSS.n3401 0.0105
R65120 VSS.n3407 VSS.n3406 0.0105
R65121 VSS.n3408 VSS.n3407 0.0105
R65122 VSS.n3409 VSS.n3408 0.0105
R65123 VSS.n3411 VSS.n3409 0.0105
R65124 VSS.n3414 VSS.n3411 0.0105
R65125 VSS.n3415 VSS.n3414 0.0105
R65126 VSS.n3418 VSS.n3415 0.0105
R65127 VSS.n3419 VSS.n3418 0.0105
R65128 VSS.n3421 VSS.n3419 0.0105
R65129 VSS.n3487 VSS.n3485 0.0105
R65130 VSS.n3490 VSS.n3487 0.0105
R65131 VSS.n3491 VSS.n3490 0.0105
R65132 VSS.n3493 VSS.n3491 0.0105
R65133 VSS.n3495 VSS.n3493 0.0105
R65134 VSS.n3497 VSS.n3495 0.0105
R65135 VSS.n3502 VSS.n3497 0.0105
R65136 VSS.n3503 VSS.n3502 0.0105
R65137 VSS.n3504 VSS.n3503 0.0105
R65138 VSS.n3505 VSS.n3504 0.0105
R65139 VSS.n3509 VSS.n3505 0.0105
R65140 VSS.n3510 VSS.n3509 0.0105
R65141 VSS.n3547 VSS.n3544 0.0105
R65142 VSS.n3548 VSS.n3547 0.0105
R65143 VSS.n3550 VSS.n3548 0.0105
R65144 VSS.n3552 VSS.n3550 0.0105
R65145 VSS.n3554 VSS.n3552 0.0105
R65146 VSS.n3556 VSS.n3554 0.0105
R65147 VSS.n3558 VSS.n3556 0.0105
R65148 VSS.n3560 VSS.n3558 0.0105
R65149 VSS.n3562 VSS.n3560 0.0105
R65150 VSS.n3564 VSS.n3562 0.0105
R65151 VSS.n3566 VSS.n3564 0.0105
R65152 VSS.n3569 VSS.n3566 0.0105
R65153 VSS.n3605 VSS.n3604 0.0105
R65154 VSS.n3607 VSS.n3605 0.0105
R65155 VSS.n3609 VSS.n3607 0.0105
R65156 VSS.n3612 VSS.n3609 0.0105
R65157 VSS.n3648 VSS.n3646 0.0105
R65158 VSS.n3650 VSS.n3648 0.0105
R65159 VSS.n3652 VSS.n3650 0.0105
R65160 VSS.n4022 VSS.n4021 0.0104355
R65161 VSS.n18893 VSS.n18892 0.0104355
R65162 VSS.n3824 VSS.n3823 0.0104355
R65163 VSS.n3247 VSS.n3246 0.0104355
R65164 VSS.n18686 VSS.n18685 0.0104296
R65165 VSS.n18450 VSS.n18449 0.0104296
R65166 VSS.n17018 VSS.n17017 0.0104296
R65167 VSS.n19518 VSS.n19517 0.0104296
R65168 VSS.n19589 VSS.n19588 0.0104296
R65169 VSS.n19917 VSS.n19916 0.0104296
R65170 VSS.n4204 VSS.n4203 0.0104213
R65171 VSS.n13143 VSS.n13142 0.0104213
R65172 VSS.n11800 VSS.n11799 0.0104213
R65173 VSS.n2234 VSS.n2233 0.0104213
R65174 VSS.n2283 VSS.n2282 0.0104213
R65175 VSS.n17891 VSS.n17890 0.0104213
R65176 VSS.n21671 VSS.n21670 0.0104213
R65177 VSS.n4132 VSS.n4131 0.0104213
R65178 VSS.n8903 VSS.n8902 0.0104213
R65179 VSS.n18371 VSS.n18370 0.0104
R65180 VSS.n16568 VSS.n16566 0.0104
R65181 VSS.n4021 VSS.n4020 0.010347
R65182 VSS.n18892 VSS.n18891 0.010347
R65183 VSS.n3823 VSS.n3822 0.010347
R65184 VSS.n3248 VSS.n3247 0.010347
R65185 VSS.n444 VSS.n443 0.0103395
R65186 VSS.n427 VSS.n426 0.0103395
R65187 VSS.n410 VSS.n409 0.0103395
R65188 VSS.n14281 VSS.n393 0.0103395
R65189 VSS.n392 VSS.n391 0.0103395
R65190 VSS.n10307 VSS.n10306 0.0103077
R65191 VSS.n10425 VSS.n10424 0.0103077
R65192 VSS.n10140 VSS.n10139 0.0103077
R65193 VSS.n10048 VSS.n10047 0.0103077
R65194 VSS.n10033 VSS.n10032 0.0103077
R65195 VSS.n12361 VSS.n12360 0.0103077
R65196 VSS.n12479 VSS.n12478 0.0103077
R65197 VSS.n12191 VSS.n12190 0.0103077
R65198 VSS.n12099 VSS.n12098 0.0103077
R65199 VSS.n12084 VSS.n12083 0.0103077
R65200 VSS.n3207 VSS.n3206 0.0102887
R65201 VSS.n5548 VSS.n5547 0.010282
R65202 VSS.n12940 VSS.n12939 0.010282
R65203 VSS.n12721 VSS.n12720 0.010282
R65204 VSS.n12939 VSS.n12938 0.010282
R65205 VSS.n16058 VSS.n16057 0.010282
R65206 VSS.n15036 VSS.n15035 0.010282
R65207 VSS.n20644 VSS.n20643 0.010282
R65208 VSS.n20992 VSS.n20991 0.010282
R65209 VSS.n6967 VSS.n6966 0.010282
R65210 VSS.n6607 VSS.n6606 0.010282
R65211 VSS.n20645 VSS.n20644 0.010282
R65212 VSS.n20105 VSS.n20104 0.010282
R65213 VSS.n1034 VSS.n1033 0.010282
R65214 VSS.n6865 VSS.n6864 0.010282
R65215 VSS.n6457 VSS.n6456 0.010282
R65216 VSS.n20104 VSS.n20103 0.010282
R65217 VSS.n21357 VSS.n21356 0.010282
R65218 VSS.n7641 VSS.n7640 0.010282
R65219 VSS.n7729 VSS.n7728 0.010282
R65220 VSS.n7810 VSS.n7809 0.010282
R65221 VSS.n21356 VSS.n21355 0.010282
R65222 VSS.n9283 VSS.n9282 0.010282
R65223 VSS.n9120 VSS.n9119 0.010282
R65224 VSS.n7811 VSS.n7810 0.010282
R65225 VSS.n6606 VSS.n6605 0.010282
R65226 VSS.n6456 VSS.n6455 0.010282
R65227 VSS.n9674 VSS.n9673 0.010282
R65228 VSS.n9557 VSS.n9556 0.010282
R65229 VSS.n7728 VSS.n7727 0.010282
R65230 VSS.n6966 VSS.n6965 0.010282
R65231 VSS.n6864 VSS.n6863 0.010282
R65232 VSS.n12722 VSS.n12721 0.010282
R65233 VSS.n7640 VSS.n7639 0.010282
R65234 VSS.n1035 VSS.n1034 0.010282
R65235 VSS.n20993 VSS.n20992 0.010282
R65236 VSS.n6116 VSS.n6115 0.010282
R65237 VSS.n11673 VSS.n11672 0.010282
R65238 VSS.n6035 VSS.n6034 0.010282
R65239 VSS.n5954 VSS.n5953 0.010282
R65240 VSS.n10588 VSS.n10587 0.010282
R65241 VSS.n630 VSS.n629 0.010282
R65242 VSS.n11361 VSS.n11360 0.0102585
R65243 VSS.n5732 VSS.n5731 0.0102585
R65244 VSS.n2355 VSS.n2354 0.0102585
R65245 VSS.n3983 VSS.n3982 0.0102585
R65246 VSS.n18854 VSS.n18853 0.0102585
R65247 VSS.n2254 VSS.n2253 0.0102585
R65248 VSS.n15162 VSS.n15161 0.0102585
R65249 VSS.n16180 VSS.n16179 0.0102585
R65250 VSS.n3783 VSS.n3782 0.0102585
R65251 VSS.n4708 VSS.n4707 0.0102585
R65252 VSS.n11427 VSS.n11426 0.0102585
R65253 VSS.n11206 VSS.n11205 0.0102585
R65254 VSS.n3263 VSS.n3262 0.0102585
R65255 VSS.n545 VSS.n544 0.0102585
R65256 VSS.n486 VSS.n485 0.0102585
R65257 VSS.n12291 VSS.n12290 0.0102441
R65258 VSS.n11943 VSS.n11942 0.0102441
R65259 VSS.n11904 VSS.n11903 0.0102441
R65260 VSS.n10239 VSS.n10238 0.0102441
R65261 VSS.n9945 VSS.n9944 0.0102441
R65262 VSS.n9904 VSS.n9903 0.0102441
R65263 VSS.n18469 VSS.n18468 0.0102183
R65264 VSS.n19570 VSS.n19569 0.0102183
R65265 VSS.n17104 VSS.n17103 0.010175
R65266 VSS.n17058 VSS.n17056 0.010175
R65267 VSS.n16959 VSS.n16957 0.010175
R65268 VSS.n14922 VSS.n14919 0.010175
R65269 VSS.n4033 VSS.n4032 0.01017
R65270 VSS.n2366 VSS.n2365 0.01017
R65271 VSS.n11335 VSS.n11334 0.01017
R65272 VSS.n5862 VSS.n5861 0.01017
R65273 VSS.n18904 VSS.n18903 0.01017
R65274 VSS.n2265 VSS.n2264 0.01017
R65275 VSS.n16223 VSS.n16222 0.01017
R65276 VSS.n15136 VSS.n15135 0.01017
R65277 VSS.n3835 VSS.n3834 0.01017
R65278 VSS.n4719 VSS.n4718 0.01017
R65279 VSS.n11453 VSS.n11452 0.01017
R65280 VSS.n11232 VSS.n11231 0.01017
R65281 VSS.n2650 VSS.n2649 0.01017
R65282 VSS.n571 VSS.n570 0.01017
R65283 VSS.n512 VSS.n511 0.01017
R65284 VSS.n11416 VSS.n5477 0.0101595
R65285 VSS.n11466 VSS.n4922 0.0101595
R65286 VSS.n11639 VSS.n4858 0.0101595
R65287 VSS.n17238 VSS.n11744 0.0101595
R65288 VSS.n17385 VSS.n17310 0.0101595
R65289 VSS.n11538 VSS.n11537 0.0100815
R65290 VSS.n9581 VSS.n9580 0.0100815
R65291 VSS.n9035 VSS.n9034 0.0100815
R65292 VSS.n11588 VSS.n11587 0.0100815
R65293 VSS.n15063 VSS.n15062 0.0100815
R65294 VSS.n9178 VSS.n9177 0.0100815
R65295 VSS.n15012 VSS.n15011 0.0100815
R65296 VSS.n9307 VSS.n9306 0.0100815
R65297 VSS.n9144 VSS.n9143 0.0100815
R65298 VSS.n9257 VSS.n9256 0.0100815
R65299 VSS.n9698 VSS.n9697 0.0100815
R65300 VSS.n16101 VSS.n16100 0.0100815
R65301 VSS.n5585 VSS.n5584 0.0100815
R65302 VSS.n11646 VSS.n11645 0.0100815
R65303 VSS.n6090 VSS.n6089 0.0100815
R65304 VSS.n6059 VSS.n6058 0.0100815
R65305 VSS.n6009 VSS.n6008 0.0100815
R65306 VSS.n5928 VSS.n5927 0.0100815
R65307 VSS.n5978 VSS.n5977 0.0100815
R65308 VSS.n6140 VSS.n6139 0.0100815
R65309 VSS.n11697 VSS.n11696 0.0100815
R65310 VSS.n604 VSS.n603 0.0100815
R65311 VSS.n10612 VSS.n10611 0.0100815
R65312 VSS.n654 VSS.n653 0.0100815
R65313 VSS.n5689 VSS.n5688 0.0100745
R65314 VSS.n5672 VSS.n5670 0.0100745
R65315 VSS.n16015 VSS.n16013 0.0100745
R65316 VSS.n996 VSS.n994 0.0100745
R65317 VSS.n987 VSS.n985 0.0100745
R65318 VSS.n20941 VSS.n20939 0.0100745
R65319 VSS.n20958 VSS.n20957 0.0100745
R65320 VSS.n5774 VSS.n5771 0.0100745
R65321 VSS.n5826 VSS.n5823 0.0100745
R65322 VSS.n5811 VSS.n5810 0.0100745
R65323 VSS.n15479 VSS.n15478 0.0100745
R65324 VSS.n1198 VSS.n1195 0.0100745
R65325 VSS.n1256 VSS.n1253 0.0100745
R65326 VSS.n1242 VSS.n1241 0.0100745
R65327 VSS.n1225 VSS.n1223 0.0100745
R65328 VSS.n16444 VSS.n16443 0.0100303
R65329 VSS.n19847 VSS.n19846 0.0100303
R65330 VSS.n19757 VSS.n19756 0.0100303
R65331 VSS.n2097 VSS.n2096 0.0100303
R65332 VSS.n20032 VSS.n20031 0.0100303
R65333 VSS.n11565 VSS.n11564 0.00999298
R65334 VSS.n5545 VSS.n5544 0.00999298
R65335 VSS.n16055 VSS.n16054 0.00999298
R65336 VSS.n9280 VSS.n9279 0.00999298
R65337 VSS.n9117 VSS.n9116 0.00999298
R65338 VSS.n9671 VSS.n9670 0.00999298
R65339 VSS.n9554 VSS.n9553 0.00999298
R65340 VSS.n6113 VSS.n6112 0.00999298
R65341 VSS.n6032 VSS.n6031 0.00999298
R65342 VSS.n5951 VSS.n5950 0.00999298
R65343 VSS.n10585 VSS.n10584 0.00999298
R65344 VSS.n627 VSS.n626 0.00999298
R65345 VSS.n19405 VSS.n19403 0.00995
R65346 VSS.n18261 VSS.n18260 0.00995
R65347 VSS.n16663 VSS.n16661 0.00995
R65348 VSS.n16616 VSS.n16615 0.00995
R65349 VSS.n16513 VSS.n16511 0.00995
R65350 VSS.n4167 VSS.n4166 0.00994444
R65351 VSS.n21709 VSS.n21708 0.00994444
R65352 VSS.n17403 VSS.n17402 0.00994444
R65353 VSS.n13285 VSS.n13284 0.00994444
R65354 VSS.n4109 VSS.n4108 0.00994444
R65355 VSS.n21905 VSS.n21904 0.00994444
R65356 VSS.n3450 VSS.n3449 0.00993662
R65357 VSS.n3454 VSS.n3453 0.00993662
R65358 VSS.n12682 VSS.n12681 0.0099291
R65359 VSS.n10550 VSS.n10549 0.0099291
R65360 VSS.n10551 VSS.n10550 0.0099291
R65361 VSS.n12683 VSS.n12682 0.0099291
R65362 VSS.n10277 VSS.n10276 0.00992308
R65363 VSS.n10286 VSS.n10285 0.00992308
R65364 VSS.n10404 VSS.n10403 0.00992308
R65365 VSS.n10395 VSS.n10394 0.00992308
R65366 VSS.n10119 VSS.n10118 0.00992308
R65367 VSS.n10110 VSS.n10109 0.00992308
R65368 VSS.n12331 VSS.n12330 0.00992308
R65369 VSS.n12340 VSS.n12339 0.00992308
R65370 VSS.n12458 VSS.n12457 0.00992308
R65371 VSS.n12449 VSS.n12448 0.00992308
R65372 VSS.n12170 VSS.n12169 0.00992308
R65373 VSS.n12161 VSS.n12160 0.00992308
R65374 VSS.n12022 VSS.n12021 0.00992308
R65375 VSS.n12013 VSS.n12012 0.00992308
R65376 VSS.n8350 VSS.n8349 0.00989057
R65377 VSS.n8158 VSS.n8157 0.00989057
R65378 VSS.n9495 VSS.n9494 0.00988976
R65379 VSS.n9612 VSS.n9611 0.00988976
R65380 VSS.n6926 VSS.n6925 0.00988976
R65381 VSS.n6803 VSS.n6802 0.00988976
R65382 VSS.n17201 VSS.n17200 0.00987905
R65383 VSS.n14397 VSS.n14396 0.00984086
R65384 VSS.n14426 VSS.n14425 0.00984086
R65385 VSS.n15071 VSS.n15070 0.00984086
R65386 VSS.n15104 VSS.n15103 0.00984086
R65387 VSS.n15174 VSS.n15173 0.00984086
R65388 VSS.n14396 VSS.n14395 0.00984086
R65389 VSS.n14427 VSS.n14426 0.00984086
R65390 VSS.n15070 VSS.n15069 0.00984086
R65391 VSS.n15103 VSS.n15102 0.00984086
R65392 VSS.n15173 VSS.n15172 0.00984086
R65393 VSS.n13361 VSS.n13360 0.00984086
R65394 VSS.n13412 VSS.n13411 0.00984086
R65395 VSS.n20683 VSS.n20682 0.00984086
R65396 VSS.n20734 VSS.n20733 0.00984086
R65397 VSS.n20826 VSS.n20825 0.00984086
R65398 VSS.n13360 VSS.n13359 0.00984086
R65399 VSS.n13411 VSS.n13410 0.00984086
R65400 VSS.n20682 VSS.n20681 0.00984086
R65401 VSS.n20733 VSS.n20732 0.00984086
R65402 VSS.n20825 VSS.n20824 0.00984086
R65403 VSS.n533 VSS.n532 0.00984086
R65404 VSS.n534 VSS.n533 0.00984086
R65405 VSS.n16629 VSS.n16598 0.00979577
R65406 VSS.n769 VSS.n768 0.00979577
R65407 DVSS VSS.n19435 0.009725
R65408 DVSS VSS.n18562 0.009725
R65409 DVSS VSS.n18300 0.009725
R65410 DVSS VSS.n16760 0.009725
R65411 DVSS VSS.n14806 0.009725
R65412 VSS.n14590 DVSS 0.009725
R65413 VSS.n17157 VSS.n17155 0.009725
R65414 VSS.n17152 VSS.n17151 0.009725
R65415 VSS.n17001 VSS.n16999 0.009725
R65416 VSS.n16996 VSS.n16995 0.009725
R65417 VSS.n15816 DVSS 0.009725
R65418 VSS.n4055 VSS.n4054 0.0097126
R65419 VSS.n13084 VSS.n13083 0.0097126
R65420 VSS.n18926 VSS.n18925 0.0097126
R65421 VSS.n21857 VSS.n21856 0.0097126
R65422 VSS.n19142 VSS.n19141 0.0097126
R65423 VSS.n2633 VSS.n2632 0.0097126
R65424 VSS.n14571 VSS.n14570 0.00969863
R65425 VSS.n14824 VSS.n14823 0.00969863
R65426 VSS.n16884 VSS.n16883 0.00969863
R65427 VSS.n16695 VSS.n16694 0.00969863
R65428 VSS.n8349 VSS.n8348 0.00969863
R65429 VSS.n8346 VSS.n8345 0.00969863
R65430 VSS.n845 VSS.n844 0.00969863
R65431 VSS.n8157 VSS.n8156 0.00969863
R65432 VSS.n8148 VSS.n8147 0.00969863
R65433 VSS.n15663 VSS.n15662 0.00964533
R65434 VSS.n15652 VSS.n15651 0.00964533
R65435 VSS.n15636 VSS.n15635 0.00964533
R65436 VSS.n15625 VSS.n15624 0.00964533
R65437 VSS.n15613 VSS.n15612 0.00964533
R65438 VSS.n15602 VSS.n15601 0.00964533
R65439 VSS.n15590 VSS.n15589 0.00964533
R65440 VSS.n15571 VSS.n15570 0.00964533
R65441 VSS.n15556 VSS.n15555 0.00964533
R65442 VSS.n15441 VSS.n15440 0.00964533
R65443 VSS.n15415 VSS.n15414 0.00964533
R65444 VSS.n15572 VSS.n15571 0.00964533
R65445 VSS.n15637 VSS.n15636 0.00964533
R65446 VSS.n15626 VSS.n15625 0.00964533
R65447 VSS.n15614 VSS.n15613 0.00964533
R65448 VSS.n15603 VSS.n15602 0.00964533
R65449 VSS.n15591 VSS.n15590 0.00964533
R65450 VSS.n15653 VSS.n15652 0.00964533
R65451 VSS.n15664 VSS.n15663 0.00964533
R65452 VSS.n15416 VSS.n15415 0.00964533
R65453 VSS.n15442 VSS.n15441 0.00964533
R65454 VSS.n15557 VSS.n15556 0.00964533
R65455 VSS.n1921 VSS.n1920 0.00964533
R65456 VSS.n1910 VSS.n1909 0.00964533
R65457 VSS.n1904 VSS.n1903 0.00964533
R65458 VSS.n1893 VSS.n1892 0.00964533
R65459 VSS.n1887 VSS.n1886 0.00964533
R65460 VSS.n1876 VSS.n1875 0.00964533
R65461 VSS.n1870 VSS.n1869 0.00964533
R65462 VSS.n1859 VSS.n1858 0.00964533
R65463 VSS.n1844 VSS.n1843 0.00964533
R65464 VSS.n1743 VSS.n1742 0.00964533
R65465 VSS.n1731 VSS.n1730 0.00964533
R65466 VSS.n1860 VSS.n1859 0.00964533
R65467 VSS.n1905 VSS.n1904 0.00964533
R65468 VSS.n1894 VSS.n1893 0.00964533
R65469 VSS.n1888 VSS.n1887 0.00964533
R65470 VSS.n1877 VSS.n1876 0.00964533
R65471 VSS.n1871 VSS.n1870 0.00964533
R65472 VSS.n1911 VSS.n1910 0.00964533
R65473 VSS.n1922 VSS.n1921 0.00964533
R65474 VSS.n1845 VSS.n1844 0.00964533
R65475 VSS.n1732 VSS.n1731 0.00964533
R65476 VSS.n1744 VSS.n1743 0.00964533
R65477 VSS.n18814 VSS.n18813 0.00962875
R65478 VSS.n19486 VSS.n19485 0.00962875
R65479 VSS.n13745 VSS.n13744 0.00962857
R65480 VSS.n13751 VSS.n13750 0.00962857
R65481 VSS.n13769 VSS.n13768 0.00962857
R65482 VSS.n13793 VSS.n13792 0.00962857
R65483 VSS.n13835 VSS.n13834 0.00962857
R65484 VSS.n13839 VSS.n13838 0.00962857
R65485 VSS.n13844 VSS.n13843 0.00962857
R65486 VSS.n13843 VSS.n13842 0.00962857
R65487 VSS.n13851 VSS.n13670 0.00962857
R65488 VSS.n13670 VSS.n13668 0.00962857
R65489 VSS.n13668 VSS.n13666 0.00962857
R65490 VSS.n14240 VSS.n14239 0.00962857
R65491 VSS.n14239 VSS.n14230 0.00962857
R65492 VSS.n14230 VSS.n14228 0.00962857
R65493 VSS.n14228 VSS.n14226 0.00962857
R65494 VSS.n14226 VSS.n14224 0.00962857
R65495 VSS.n14224 VSS.n14222 0.00962857
R65496 VSS.n14222 VSS.n14220 0.00962857
R65497 VSS.n14220 VSS.n14218 0.00962857
R65498 VSS.n14218 VSS.n14216 0.00962857
R65499 VSS.n14216 VSS.n14214 0.00962857
R65500 VSS.n13681 VSS.n13679 0.00962857
R65501 VSS.n13683 VSS.n13681 0.00962857
R65502 VSS.n13685 VSS.n13683 0.00962857
R65503 VSS.n13687 VSS.n13685 0.00962857
R65504 VSS.n13689 VSS.n13687 0.00962857
R65505 VSS.n13691 VSS.n13689 0.00962857
R65506 VSS.n13693 VSS.n13691 0.00962857
R65507 VSS.n13695 VSS.n13693 0.00962857
R65508 VSS.n13697 VSS.n13695 0.00962857
R65509 VSS.n13699 VSS.n13697 0.00962857
R65510 VSS.n13701 VSS.n13699 0.00962857
R65511 VSS.n13703 VSS.n13701 0.00962857
R65512 VSS.n13705 VSS.n13703 0.00962857
R65513 VSS.n13707 VSS.n13705 0.00962857
R65514 VSS.n13709 VSS.n13707 0.00962857
R65515 VSS.n13711 VSS.n13709 0.00962857
R65516 VSS.n13713 VSS.n13711 0.00962857
R65517 VSS.n13715 VSS.n13713 0.00962857
R65518 VSS.n13717 VSS.n13715 0.00962857
R65519 VSS.n13719 VSS.n13717 0.00962857
R65520 VSS.n13721 VSS.n13719 0.00962857
R65521 VSS.n13723 VSS.n13721 0.00962857
R65522 VSS.n13725 VSS.n13723 0.00962857
R65523 VSS.n13727 VSS.n13725 0.00962857
R65524 VSS.n13729 VSS.n13727 0.00962857
R65525 VSS.n13731 VSS.n13729 0.00962857
R65526 VSS.n13733 VSS.n13731 0.00962857
R65527 VSS.n13735 VSS.n13733 0.00962857
R65528 VSS.n13737 VSS.n13735 0.00962857
R65529 VSS.n13739 VSS.n13737 0.00962857
R65530 VSS.n13741 VSS.n13739 0.00962857
R65531 VSS.n13743 VSS.n13741 0.00962857
R65532 VSS.n13746 VSS.n13743 0.00962857
R65533 VSS.n13747 VSS.n13746 0.00962857
R65534 VSS.n13749 VSS.n13747 0.00962857
R65535 VSS.n13752 VSS.n13749 0.00962857
R65536 VSS.n13753 VSS.n13752 0.00962857
R65537 VSS.n13755 VSS.n13753 0.00962857
R65538 VSS.n13757 VSS.n13755 0.00962857
R65539 VSS.n13759 VSS.n13757 0.00962857
R65540 VSS.n13761 VSS.n13759 0.00962857
R65541 VSS.n13763 VSS.n13761 0.00962857
R65542 VSS.n13765 VSS.n13763 0.00962857
R65543 VSS.n13767 VSS.n13765 0.00962857
R65544 VSS.n13770 VSS.n13767 0.00962857
R65545 VSS.n13771 VSS.n13770 0.00962857
R65546 VSS.n13773 VSS.n13771 0.00962857
R65547 VSS.n13775 VSS.n13773 0.00962857
R65548 VSS.n13777 VSS.n13775 0.00962857
R65549 VSS.n13779 VSS.n13777 0.00962857
R65550 VSS.n13781 VSS.n13779 0.00962857
R65551 VSS.n13783 VSS.n13781 0.00962857
R65552 VSS.n13785 VSS.n13783 0.00962857
R65553 VSS.n13787 VSS.n13785 0.00962857
R65554 VSS.n13789 VSS.n13787 0.00962857
R65555 VSS.n13791 VSS.n13789 0.00962857
R65556 VSS.n13794 VSS.n13791 0.00962857
R65557 VSS.n13795 VSS.n13794 0.00962857
R65558 VSS.n13797 VSS.n13795 0.00962857
R65559 VSS.n13799 VSS.n13797 0.00962857
R65560 VSS.n13801 VSS.n13799 0.00962857
R65561 VSS.n13803 VSS.n13801 0.00962857
R65562 VSS.n13805 VSS.n13803 0.00962857
R65563 VSS.n13807 VSS.n13805 0.00962857
R65564 VSS.n13809 VSS.n13807 0.00962857
R65565 VSS.n13811 VSS.n13809 0.00962857
R65566 VSS.n13813 VSS.n13811 0.00962857
R65567 VSS.n13815 VSS.n13813 0.00962857
R65568 VSS.n13817 VSS.n13815 0.00962857
R65569 VSS.n13819 VSS.n13817 0.00962857
R65570 VSS.n13821 VSS.n13819 0.00962857
R65571 VSS.n13823 VSS.n13821 0.00962857
R65572 VSS.n13825 VSS.n13823 0.00962857
R65573 VSS.n13827 VSS.n13825 0.00962857
R65574 VSS.n13829 VSS.n13827 0.00962857
R65575 VSS.n13831 VSS.n13829 0.00962857
R65576 VSS.n13833 VSS.n13831 0.00962857
R65577 VSS.n13836 VSS.n13833 0.00962857
R65578 VSS.n13837 VSS.n13836 0.00962857
R65579 VSS.n13840 VSS.n13837 0.00962857
R65580 VSS.n13841 VSS.n13840 0.00962857
R65581 VSS.n13845 VSS.n13841 0.00962857
R65582 VSS.n13846 VSS.n13845 0.00962857
R65583 VSS.n13847 VSS.n13846 0.00962857
R65584 VSS.n13849 VSS.n13847 0.00962857
R65585 VSS.n2583 VSS.n2582 0.00962857
R65586 VSS.n2698 VSS.n2697 0.00962857
R65587 VSS.n2697 VSS.n2696 0.00962857
R65588 VSS.n2696 VSS.n2695 0.00962857
R65589 VSS.n2751 VSS.n2750 0.00962857
R65590 VSS.n2750 VSS.n2749 0.00962857
R65591 VSS.n2749 VSS.n2748 0.00962857
R65592 VSS.n2748 VSS.n2747 0.00962857
R65593 VSS.n2747 VSS.n2746 0.00962857
R65594 VSS.n2746 VSS.n2745 0.00962857
R65595 VSS.n2745 VSS.n2744 0.00962857
R65596 VSS.n2744 VSS.n2743 0.00962857
R65597 VSS.n2743 VSS.n2742 0.00962857
R65598 VSS.n2742 VSS.n2741 0.00962857
R65599 VSS.n2741 VSS.n2740 0.00962857
R65600 VSS.n2740 VSS.n2739 0.00962857
R65601 VSS.n2801 VSS.n2800 0.00962857
R65602 VSS.n2800 VSS.n2799 0.00962857
R65603 VSS.n2897 VSS.n2896 0.00962857
R65604 VSS.n2896 VSS.n2895 0.00962857
R65605 VSS.n2895 VSS.n2894 0.00962857
R65606 VSS.n2905 VSS.n2904 0.00962857
R65607 VSS.n2975 VSS.n2974 0.00962857
R65608 VSS.n3071 VSS.n3070 0.00962857
R65609 VSS.n2581 VSS.n2579 0.00962857
R65610 VSS.n2584 VSS.n2581 0.00962857
R65611 VSS.n2585 VSS.n2584 0.00962857
R65612 VSS.n2587 VSS.n2585 0.00962857
R65613 VSS.n2700 VSS.n2699 0.00962857
R65614 VSS.n2701 VSS.n2700 0.00962857
R65615 VSS.n2702 VSS.n2701 0.00962857
R65616 VSS.n2704 VSS.n2702 0.00962857
R65617 VSS.n2753 VSS.n2752 0.00962857
R65618 VSS.n2754 VSS.n2753 0.00962857
R65619 VSS.n2755 VSS.n2754 0.00962857
R65620 VSS.n2756 VSS.n2755 0.00962857
R65621 VSS.n2757 VSS.n2756 0.00962857
R65622 VSS.n2758 VSS.n2757 0.00962857
R65623 VSS.n2759 VSS.n2758 0.00962857
R65624 VSS.n2760 VSS.n2759 0.00962857
R65625 VSS.n2761 VSS.n2760 0.00962857
R65626 VSS.n2762 VSS.n2761 0.00962857
R65627 VSS.n2763 VSS.n2762 0.00962857
R65628 VSS.n2764 VSS.n2763 0.00962857
R65629 VSS.n2803 VSS.n2802 0.00962857
R65630 VSS.n2804 VSS.n2803 0.00962857
R65631 VSS.n2806 VSS.n2804 0.00962857
R65632 VSS.n2808 VSS.n2806 0.00962857
R65633 VSS.n2810 VSS.n2808 0.00962857
R65634 VSS.n2812 VSS.n2810 0.00962857
R65635 VSS.n2814 VSS.n2812 0.00962857
R65636 VSS.n2816 VSS.n2814 0.00962857
R65637 VSS.n2818 VSS.n2816 0.00962857
R65638 VSS.n2820 VSS.n2818 0.00962857
R65639 VSS.n2822 VSS.n2820 0.00962857
R65640 VSS.n2824 VSS.n2822 0.00962857
R65641 VSS.n2899 VSS.n2898 0.00962857
R65642 VSS.n2900 VSS.n2899 0.00962857
R65643 VSS.n2901 VSS.n2900 0.00962857
R65644 VSS.n2903 VSS.n2901 0.00962857
R65645 VSS.n2906 VSS.n2903 0.00962857
R65646 VSS.n2907 VSS.n2906 0.00962857
R65647 VSS.n2909 VSS.n2907 0.00962857
R65648 VSS.n2911 VSS.n2909 0.00962857
R65649 VSS.n2913 VSS.n2911 0.00962857
R65650 VSS.n2915 VSS.n2913 0.00962857
R65651 VSS.n2917 VSS.n2915 0.00962857
R65652 VSS.n2920 VSS.n2917 0.00962857
R65653 VSS.n2961 VSS.n2959 0.00962857
R65654 VSS.n2963 VSS.n2961 0.00962857
R65655 VSS.n2965 VSS.n2963 0.00962857
R65656 VSS.n2967 VSS.n2965 0.00962857
R65657 VSS.n2969 VSS.n2967 0.00962857
R65658 VSS.n2971 VSS.n2969 0.00962857
R65659 VSS.n2973 VSS.n2971 0.00962857
R65660 VSS.n2976 VSS.n2973 0.00962857
R65661 VSS.n2977 VSS.n2976 0.00962857
R65662 VSS.n2979 VSS.n2977 0.00962857
R65663 VSS.n2981 VSS.n2979 0.00962857
R65664 VSS.n2984 VSS.n2981 0.00962857
R65665 VSS.n3025 VSS.n3023 0.00962857
R65666 VSS.n3027 VSS.n3025 0.00962857
R65667 VSS.n3029 VSS.n3027 0.00962857
R65668 VSS.n3032 VSS.n3029 0.00962857
R65669 VSS.n3073 VSS.n3072 0.00962857
R65670 VSS.n3075 VSS.n3073 0.00962857
R65671 VSS.n3077 VSS.n3075 0.00962857
R65672 VSS.n4980 VSS.n4979 0.00962857
R65673 VSS.n4979 VSS.n4978 0.00962857
R65674 VSS.n4978 VSS.n4977 0.00962857
R65675 VSS.n5044 VSS.n5043 0.00962857
R65676 VSS.n5052 VSS.n5051 0.00962857
R65677 VSS.n5059 VSS.n5058 0.00962857
R65678 VSS.n5058 VSS.n5057 0.00962857
R65679 VSS.n5092 VSS.n5091 0.00962857
R65680 VSS.n4982 VSS.n4981 0.00962857
R65681 VSS.n4983 VSS.n4982 0.00962857
R65682 VSS.n4984 VSS.n4983 0.00962857
R65683 VSS.n4986 VSS.n4984 0.00962857
R65684 VSS.n5010 VSS.n5008 0.00962857
R65685 VSS.n5012 VSS.n5010 0.00962857
R65686 VSS.n5014 VSS.n5012 0.00962857
R65687 VSS.n5016 VSS.n5014 0.00962857
R65688 VSS.n5040 VSS.n5038 0.00962857
R65689 VSS.n5042 VSS.n5040 0.00962857
R65690 VSS.n5045 VSS.n5042 0.00962857
R65691 VSS.n5046 VSS.n5045 0.00962857
R65692 VSS.n5048 VSS.n5046 0.00962857
R65693 VSS.n5050 VSS.n5048 0.00962857
R65694 VSS.n5053 VSS.n5050 0.00962857
R65695 VSS.n5054 VSS.n5053 0.00962857
R65696 VSS.n5056 VSS.n5054 0.00962857
R65697 VSS.n5060 VSS.n5056 0.00962857
R65698 VSS.n5061 VSS.n5060 0.00962857
R65699 VSS.n5062 VSS.n5061 0.00962857
R65700 VSS.n5086 VSS.n5084 0.00962857
R65701 VSS.n5088 VSS.n5086 0.00962857
R65702 VSS.n5090 VSS.n5088 0.00962857
R65703 VSS.n5093 VSS.n5090 0.00962857
R65704 VSS.n5094 VSS.n5093 0.00962857
R65705 VSS.n5096 VSS.n5094 0.00962857
R65706 VSS.n5098 VSS.n5096 0.00962857
R65707 VSS.n5100 VSS.n5098 0.00962857
R65708 VSS.n5102 VSS.n5100 0.00962857
R65709 VSS.n5104 VSS.n5102 0.00962857
R65710 VSS.n5106 VSS.n5104 0.00962857
R65711 VSS.n5109 VSS.n5106 0.00962857
R65712 VSS.n5166 VSS.n5164 0.00962857
R65713 VSS.n5168 VSS.n5166 0.00962857
R65714 VSS.n5170 VSS.n5168 0.00962857
R65715 VSS.n5172 VSS.n5170 0.00962857
R65716 VSS.n5174 VSS.n5172 0.00962857
R65717 VSS.n5176 VSS.n5174 0.00962857
R65718 VSS.n5178 VSS.n5176 0.00962857
R65719 VSS.n5180 VSS.n5178 0.00962857
R65720 VSS.n5182 VSS.n5180 0.00962857
R65721 VSS.n5184 VSS.n5182 0.00962857
R65722 VSS.n5186 VSS.n5184 0.00962857
R65723 VSS.n5189 VSS.n5186 0.00962857
R65724 VSS.n5217 VSS.n5215 0.00962857
R65725 VSS.n5219 VSS.n5217 0.00962857
R65726 VSS.n5221 VSS.n5219 0.00962857
R65727 VSS.n5223 VSS.n5221 0.00962857
R65728 VSS.n5225 VSS.n5223 0.00962857
R65729 VSS.n5227 VSS.n5225 0.00962857
R65730 VSS.n5229 VSS.n5227 0.00962857
R65731 VSS.n5231 VSS.n5229 0.00962857
R65732 VSS.n5233 VSS.n5231 0.00962857
R65733 VSS.n5235 VSS.n5233 0.00962857
R65734 VSS.n5237 VSS.n5235 0.00962857
R65735 VSS.n5240 VSS.n5237 0.00962857
R65736 VSS.n5268 VSS.n5266 0.00962857
R65737 VSS.n5270 VSS.n5268 0.00962857
R65738 VSS.n5272 VSS.n5270 0.00962857
R65739 VSS.n5275 VSS.n5272 0.00962857
R65740 VSS.n5303 VSS.n5301 0.00962857
R65741 VSS.n5305 VSS.n5303 0.00962857
R65742 VSS.n5307 VSS.n5305 0.00962857
R65743 VSS.n7410 VSS.n7409 0.00962857
R65744 VSS.n7348 VSS.n7347 0.00962857
R65745 VSS.n7336 VSS.n7335 0.00962857
R65746 VSS.n7330 VSS.n7329 0.00962857
R65747 VSS.n7329 VSS.n7328 0.00962857
R65748 VSS.n7328 VSS.n7327 0.00962857
R65749 VSS.n7294 VSS.n7293 0.00962857
R65750 VSS.n7196 VSS.n7195 0.00962857
R65751 VSS.n7195 VSS.n7194 0.00962857
R65752 VSS.n7151 VSS.n7150 0.00962857
R65753 VSS.n7150 VSS.n7149 0.00962857
R65754 VSS.n7149 VSS.n7148 0.00962857
R65755 VSS.n7148 VSS.n7147 0.00962857
R65756 VSS.n7147 VSS.n7146 0.00962857
R65757 VSS.n7146 VSS.n7145 0.00962857
R65758 VSS.n7137 VSS.n7136 0.00962857
R65759 VSS.n7136 VSS.n7135 0.00962857
R65760 VSS.n7135 VSS.n7134 0.00962857
R65761 VSS.n7134 VSS.n7133 0.00962857
R65762 VSS.n7094 VSS.n7093 0.00962857
R65763 VSS.n7093 VSS.n7092 0.00962857
R65764 VSS.n7088 VSS.n7087 0.00962857
R65765 VSS.n7057 VSS.n7056 0.00962857
R65766 VSS.n7056 VSS.n7055 0.00962857
R65767 VSS.n7417 VSS.n7415 0.00962857
R65768 VSS.n7415 VSS.n7413 0.00962857
R65769 VSS.n7413 VSS.n7411 0.00962857
R65770 VSS.n7411 VSS.n7408 0.00962857
R65771 VSS.n7387 VSS.n7385 0.00962857
R65772 VSS.n7385 VSS.n7383 0.00962857
R65773 VSS.n7383 VSS.n7381 0.00962857
R65774 VSS.n7381 VSS.n7379 0.00962857
R65775 VSS.n7349 VSS.n7346 0.00962857
R65776 VSS.n7346 VSS.n7345 0.00962857
R65777 VSS.n7345 VSS.n7343 0.00962857
R65778 VSS.n7343 VSS.n7341 0.00962857
R65779 VSS.n7341 VSS.n7339 0.00962857
R65780 VSS.n7339 VSS.n7337 0.00962857
R65781 VSS.n7337 VSS.n7334 0.00962857
R65782 VSS.n7334 VSS.n7333 0.00962857
R65783 VSS.n7333 VSS.n7331 0.00962857
R65784 VSS.n7331 VSS.n7326 0.00962857
R65785 VSS.n7326 VSS.n7325 0.00962857
R65786 VSS.n7325 VSS.n7324 0.00962857
R65787 VSS.n7295 VSS.n7292 0.00962857
R65788 VSS.n7292 VSS.n7291 0.00962857
R65789 VSS.n7291 VSS.n7289 0.00962857
R65790 VSS.n7289 VSS.n7287 0.00962857
R65791 VSS.n7287 VSS.n7285 0.00962857
R65792 VSS.n7285 VSS.n7283 0.00962857
R65793 VSS.n7283 VSS.n7281 0.00962857
R65794 VSS.n7281 VSS.n7279 0.00962857
R65795 VSS.n7279 VSS.n7277 0.00962857
R65796 VSS.n7277 VSS.n7275 0.00962857
R65797 VSS.n7275 VSS.n7273 0.00962857
R65798 VSS.n7273 VSS.n7271 0.00962857
R65799 VSS.n7213 VSS.n7211 0.00962857
R65800 VSS.n7211 VSS.n7209 0.00962857
R65801 VSS.n7209 VSS.n7207 0.00962857
R65802 VSS.n7207 VSS.n7205 0.00962857
R65803 VSS.n7205 VSS.n7203 0.00962857
R65804 VSS.n7203 VSS.n7201 0.00962857
R65805 VSS.n7201 VSS.n7199 0.00962857
R65806 VSS.n7199 VSS.n7197 0.00962857
R65807 VSS.n7197 VSS.n7193 0.00962857
R65808 VSS.n7193 VSS.n7192 0.00962857
R65809 VSS.n7192 VSS.n7191 0.00962857
R65810 VSS.n7191 VSS.n7189 0.00962857
R65811 VSS.n7154 VSS.n7152 0.00962857
R65812 VSS.n7152 VSS.n7144 0.00962857
R65813 VSS.n7144 VSS.n7143 0.00962857
R65814 VSS.n7143 VSS.n7142 0.00962857
R65815 VSS.n7142 VSS.n7141 0.00962857
R65816 VSS.n7141 VSS.n7140 0.00962857
R65817 VSS.n7140 VSS.n7139 0.00962857
R65818 VSS.n7139 VSS.n7138 0.00962857
R65819 VSS.n7138 VSS.n7132 0.00962857
R65820 VSS.n7132 VSS.n7131 0.00962857
R65821 VSS.n7131 VSS.n7130 0.00962857
R65822 VSS.n7130 VSS.n7129 0.00962857
R65823 VSS.n7095 VSS.n7091 0.00962857
R65824 VSS.n7091 VSS.n7090 0.00962857
R65825 VSS.n7090 VSS.n7089 0.00962857
R65826 VSS.n7089 VSS.n7085 0.00962857
R65827 VSS.n7059 VSS.n7058 0.00962857
R65828 VSS.n7058 VSS.n7049 0.00962857
R65829 VSS.n7050 VSS.n7049 0.00962857
R65830 VSS.n4668 VSS.n4667 0.00962857
R65831 VSS.n4470 VSS.n4469 0.00962857
R65832 VSS.n4681 VSS.n4679 0.00962857
R65833 VSS.n4679 VSS.n4677 0.00962857
R65834 VSS.n4677 VSS.n4675 0.00962857
R65835 VSS.n4675 VSS.n4673 0.00962857
R65836 VSS.n4650 VSS.n4649 0.00962857
R65837 VSS.n4649 VSS.n4647 0.00962857
R65838 VSS.n4647 VSS.n4645 0.00962857
R65839 VSS.n4645 VSS.n4643 0.00962857
R65840 VSS.n4643 VSS.n4641 0.00962857
R65841 VSS.n4641 VSS.n4639 0.00962857
R65842 VSS.n4617 VSS.n4615 0.00962857
R65843 VSS.n4615 VSS.n4613 0.00962857
R65844 VSS.n4613 VSS.n4611 0.00962857
R65845 VSS.n4611 VSS.n4609 0.00962857
R65846 VSS.n4609 VSS.n4607 0.00962857
R65847 VSS.n4607 VSS.n4605 0.00962857
R65848 VSS.n4605 VSS.n4603 0.00962857
R65849 VSS.n4603 VSS.n4601 0.00962857
R65850 VSS.n4601 VSS.n4599 0.00962857
R65851 VSS.n4599 VSS.n4597 0.00962857
R65852 VSS.n4597 VSS.n4595 0.00962857
R65853 VSS.n4595 VSS.n4593 0.00962857
R65854 VSS.n4571 VSS.n4569 0.00962857
R65855 VSS.n4569 VSS.n4567 0.00962857
R65856 VSS.n4567 VSS.n4565 0.00962857
R65857 VSS.n4565 VSS.n4563 0.00962857
R65858 VSS.n4563 VSS.n4561 0.00962857
R65859 VSS.n4561 VSS.n4559 0.00962857
R65860 VSS.n4559 VSS.n4557 0.00962857
R65861 VSS.n4557 VSS.n4555 0.00962857
R65862 VSS.n4555 VSS.n4553 0.00962857
R65863 VSS.n4553 VSS.n4551 0.00962857
R65864 VSS.n4551 VSS.n4549 0.00962857
R65865 VSS.n4549 VSS.n4547 0.00962857
R65866 VSS.n4491 VSS.n4489 0.00962857
R65867 VSS.n4489 VSS.n4487 0.00962857
R65868 VSS.n4487 VSS.n4485 0.00962857
R65869 VSS.n4485 VSS.n4483 0.00962857
R65870 VSS.n4483 VSS.n4481 0.00962857
R65871 VSS.n4481 VSS.n4479 0.00962857
R65872 VSS.n4479 VSS.n4477 0.00962857
R65873 VSS.n4477 VSS.n4475 0.00962857
R65874 VSS.n4475 VSS.n4473 0.00962857
R65875 VSS.n4473 VSS.n4471 0.00962857
R65876 VSS.n4471 VSS.n4468 0.00962857
R65877 VSS.n4468 VSS.n4467 0.00962857
R65878 VSS.n4440 VSS.n4438 0.00962857
R65879 VSS.n4438 VSS.n4436 0.00962857
R65880 VSS.n4436 VSS.n4434 0.00962857
R65881 VSS.n4434 VSS.n4432 0.00962857
R65882 VSS.n4432 VSS.n4430 0.00962857
R65883 VSS.n4430 VSS.n4428 0.00962857
R65884 VSS.n4428 VSS.n4426 0.00962857
R65885 VSS.n4426 VSS.n4424 0.00962857
R65886 VSS.n4424 VSS.n4422 0.00962857
R65887 VSS.n4422 VSS.n4420 0.00962857
R65888 VSS.n4420 VSS.n4418 0.00962857
R65889 VSS.n4418 VSS.n4416 0.00962857
R65890 VSS.n4389 VSS.n4387 0.00962857
R65891 VSS.n4387 VSS.n4385 0.00962857
R65892 VSS.n4385 VSS.n4383 0.00962857
R65893 VSS.n4383 VSS.n4381 0.00962857
R65894 VSS.n4354 VSS.n4352 0.00962857
R65895 VSS.n4352 VSS.n4350 0.00962857
R65896 VSS.n4350 VSS.n4348 0.00962857
R65897 VSS.n17599 VSS.n17597 0.00962857
R65898 VSS.n17597 VSS.n17595 0.00962857
R65899 VSS.n17595 VSS.n17593 0.00962857
R65900 VSS.n17593 VSS.n17591 0.00962857
R65901 VSS.n17576 VSS.n17574 0.00962857
R65902 VSS.n17574 VSS.n17567 0.00962857
R65903 VSS.n17567 VSS.n17566 0.00962857
R65904 VSS.n17566 VSS.n17565 0.00962857
R65905 VSS.n17565 VSS.n17564 0.00962857
R65906 VSS.n17564 VSS.n17563 0.00962857
R65907 VSS.n17530 VSS.n17516 0.00962857
R65908 VSS.n17516 VSS.n17515 0.00962857
R65909 VSS.n17515 VSS.n17514 0.00962857
R65910 VSS.n17514 VSS.n17513 0.00962857
R65911 VSS.n17513 VSS.n17512 0.00962857
R65912 VSS.n17512 VSS.n17511 0.00962857
R65913 VSS.n17511 VSS.n17510 0.00962857
R65914 VSS.n17510 VSS.n17509 0.00962857
R65915 VSS.n17509 VSS.n17508 0.00962857
R65916 VSS.n17508 VSS.n17507 0.00962857
R65917 VSS.n17507 VSS.n17506 0.00962857
R65918 VSS.n17506 VSS.n17505 0.00962857
R65919 VSS.n18096 VSS.n18092 0.00962857
R65920 VSS.n18092 VSS.n18091 0.00962857
R65921 VSS.n18091 VSS.n18090 0.00962857
R65922 VSS.n18090 VSS.n18088 0.00962857
R65923 VSS.n18088 VSS.n18086 0.00962857
R65924 VSS.n18086 VSS.n18084 0.00962857
R65925 VSS.n18084 VSS.n18082 0.00962857
R65926 VSS.n18082 VSS.n18080 0.00962857
R65927 VSS.n18080 VSS.n18078 0.00962857
R65928 VSS.n18078 VSS.n18076 0.00962857
R65929 VSS.n18076 VSS.n18074 0.00962857
R65930 VSS.n18074 VSS.n18072 0.00962857
R65931 VSS.n18006 VSS.n18004 0.00962857
R65932 VSS.n18004 VSS.n18001 0.00962857
R65933 VSS.n18001 VSS.n18000 0.00962857
R65934 VSS.n18000 VSS.n17998 0.00962857
R65935 VSS.n17998 VSS.n17995 0.00962857
R65936 VSS.n17995 VSS.n17994 0.00962857
R65937 VSS.n17994 VSS.n17992 0.00962857
R65938 VSS.n17992 VSS.n17990 0.00962857
R65939 VSS.n17990 VSS.n17988 0.00962857
R65940 VSS.n17988 VSS.n17986 0.00962857
R65941 VSS.n17986 VSS.n17984 0.00962857
R65942 VSS.n17984 VSS.n17982 0.00962857
R65943 VSS.n17852 VSS.n17850 0.00962857
R65944 VSS.n17850 VSS.n17848 0.00962857
R65945 VSS.n17848 VSS.n17846 0.00962857
R65946 VSS.n17846 VSS.n17844 0.00962857
R65947 VSS.n17844 VSS.n17842 0.00962857
R65948 VSS.n17842 VSS.n17839 0.00962857
R65949 VSS.n17839 VSS.n17838 0.00962857
R65950 VSS.n17838 VSS.n17836 0.00962857
R65951 VSS.n17836 VSS.n17834 0.00962857
R65952 VSS.n17834 VSS.n17832 0.00962857
R65953 VSS.n17832 VSS.n17830 0.00962857
R65954 VSS.n17830 VSS.n17828 0.00962857
R65955 VSS.n17791 VSS.n17789 0.00962857
R65956 VSS.n17789 VSS.n17787 0.00962857
R65957 VSS.n17787 VSS.n17784 0.00962857
R65958 VSS.n17784 VSS.n17783 0.00962857
R65959 VSS.n17746 VSS.n17744 0.00962857
R65960 VSS.n17744 VSS.n17742 0.00962857
R65961 VSS.n17742 VSS.n17740 0.00962857
R65962 VSS.n17573 VSS.n17572 0.00962857
R65963 VSS.n17572 VSS.n17571 0.00962857
R65964 VSS.n17571 VSS.n17570 0.00962857
R65965 VSS.n17570 VSS.n17569 0.00962857
R65966 VSS.n17569 VSS.n17568 0.00962857
R65967 VSS.n17529 VSS.n17528 0.00962857
R65968 VSS.n17528 VSS.n17527 0.00962857
R65969 VSS.n17527 VSS.n17526 0.00962857
R65970 VSS.n17526 VSS.n17525 0.00962857
R65971 VSS.n17525 VSS.n17524 0.00962857
R65972 VSS.n17524 VSS.n17523 0.00962857
R65973 VSS.n17523 VSS.n17522 0.00962857
R65974 VSS.n17522 VSS.n17521 0.00962857
R65975 VSS.n17521 VSS.n17520 0.00962857
R65976 VSS.n17520 VSS.n17519 0.00962857
R65977 VSS.n17519 VSS.n17518 0.00962857
R65978 VSS.n17518 VSS.n17517 0.00962857
R65979 VSS.n18095 VSS.n18094 0.00962857
R65980 VSS.n18094 VSS.n18093 0.00962857
R65981 VSS.n18003 VSS.n18002 0.00962857
R65982 VSS.n17997 VSS.n17996 0.00962857
R65983 VSS.n17841 VSS.n17840 0.00962857
R65984 VSS.n17786 VSS.n17785 0.00962857
R65985 VSS.n22003 VSS.n22002 0.00962857
R65986 VSS.n21992 VSS.n21991 0.00962857
R65987 VSS.n21994 VSS.n21993 0.00962857
R65988 VSS.n13950 VSS.n13949 0.00962857
R65989 VSS.n13954 VSS.n13953 0.00962857
R65990 VSS.n13955 VSS.n13954 0.00962857
R65991 VSS.n13956 VSS.n13955 0.00962857
R65992 VSS.n14102 VSS.n14101 0.00962857
R65993 VSS.n14098 VSS.n14097 0.00962857
R65994 VSS.n14094 VSS.n14093 0.00962857
R65995 VSS.n13958 VSS.n13957 0.00962857
R65996 VSS.n13959 VSS.n13958 0.00962857
R65997 VSS.n13967 VSS.n13966 0.00962857
R65998 VSS.n14038 VSS.n14037 0.00962857
R65999 VSS.n13978 VSS.n13977 0.00962857
R66000 VSS.n13979 VSS.n13978 0.00962857
R66001 VSS.n14029 VSS.n14028 0.00962857
R66002 VSS.n14018 VSS.n14017 0.00962857
R66003 VSS.n14019 VSS.n14018 0.00962857
R66004 VSS.n14020 VSS.n14019 0.00962857
R66005 VSS.n14014 VSS.n14013 0.00962857
R66006 VSS.n13985 VSS.n13984 0.00962857
R66007 VSS.n13999 VSS.n13998 0.00962857
R66008 VSS.n14000 VSS.n13999 0.00962857
R66009 VSS.n22257 VSS.n22256 0.00962857
R66010 VSS.n22007 VSS.n22005 0.00962857
R66011 VSS.n22005 VSS.n22004 0.00962857
R66012 VSS.n22004 VSS.n22001 0.00962857
R66013 VSS.n22001 VSS.n22000 0.00962857
R66014 VSS.n22000 VSS.n21998 0.00962857
R66015 VSS.n21998 VSS.n21997 0.00962857
R66016 VSS.n21997 VSS.n21996 0.00962857
R66017 VSS.n21996 VSS.n21995 0.00962857
R66018 VSS.n14118 VSS.n14117 0.00962857
R66019 VSS.n14117 VSS.n14116 0.00962857
R66020 VSS.n14116 VSS.n14114 0.00962857
R66021 VSS.n14114 VSS.n14113 0.00962857
R66022 VSS.n14113 VSS.n14111 0.00962857
R66023 VSS.n14111 VSS.n14110 0.00962857
R66024 VSS.n14110 VSS.n14109 0.00962857
R66025 VSS.n14109 VSS.n14108 0.00962857
R66026 VSS.n14108 VSS.n14107 0.00962857
R66027 VSS.n14107 VSS.n14106 0.00962857
R66028 VSS.n14106 VSS.n14104 0.00962857
R66029 VSS.n14104 VSS.n14103 0.00962857
R66030 VSS.n14103 VSS.n14100 0.00962857
R66031 VSS.n14100 VSS.n14099 0.00962857
R66032 VSS.n14099 VSS.n14096 0.00962857
R66033 VSS.n14096 VSS.n14095 0.00962857
R66034 VSS.n14095 VSS.n14092 0.00962857
R66035 VSS.n14092 VSS.n14091 0.00962857
R66036 VSS.n14091 VSS.n14090 0.00962857
R66037 VSS.n14090 VSS.n14089 0.00962857
R66038 VSS.n14089 VSS.n14087 0.00962857
R66039 VSS.n14087 VSS.n14086 0.00962857
R66040 VSS.n14086 VSS.n14084 0.00962857
R66041 VSS.n14084 VSS.n14083 0.00962857
R66042 VSS.n14083 VSS.n14081 0.00962857
R66043 VSS.n14081 VSS.n14080 0.00962857
R66044 VSS.n14080 VSS.n14078 0.00962857
R66045 VSS.n14078 VSS.n14077 0.00962857
R66046 VSS.n14077 VSS.n14075 0.00962857
R66047 VSS.n14075 VSS.n14074 0.00962857
R66048 VSS.n14074 VSS.n14072 0.00962857
R66049 VSS.n14072 VSS.n14071 0.00962857
R66050 VSS.n14071 VSS.n14070 0.00962857
R66051 VSS.n14070 VSS.n14069 0.00962857
R66052 VSS.n14069 VSS.n14067 0.00962857
R66053 VSS.n14067 VSS.n14066 0.00962857
R66054 VSS.n14066 VSS.n14064 0.00962857
R66055 VSS.n14064 VSS.n14063 0.00962857
R66056 VSS.n14063 VSS.n14061 0.00962857
R66057 VSS.n14061 VSS.n14060 0.00962857
R66058 VSS.n14060 VSS.n14058 0.00962857
R66059 VSS.n14058 VSS.n14057 0.00962857
R66060 VSS.n14057 VSS.n14055 0.00962857
R66061 VSS.n14055 VSS.n14054 0.00962857
R66062 VSS.n14054 VSS.n14052 0.00962857
R66063 VSS.n14052 VSS.n14051 0.00962857
R66064 VSS.n14051 VSS.n14049 0.00962857
R66065 VSS.n14049 VSS.n14048 0.00962857
R66066 VSS.n14048 VSS.n14046 0.00962857
R66067 VSS.n14046 VSS.n14045 0.00962857
R66068 VSS.n14045 VSS.n14043 0.00962857
R66069 VSS.n14043 VSS.n14042 0.00962857
R66070 VSS.n14042 VSS.n14040 0.00962857
R66071 VSS.n14040 VSS.n14039 0.00962857
R66072 VSS.n14039 VSS.n14036 0.00962857
R66073 VSS.n14036 VSS.n14035 0.00962857
R66074 VSS.n14035 VSS.n14034 0.00962857
R66075 VSS.n14034 VSS.n14033 0.00962857
R66076 VSS.n14033 VSS.n14031 0.00962857
R66077 VSS.n14031 VSS.n14030 0.00962857
R66078 VSS.n14030 VSS.n14027 0.00962857
R66079 VSS.n14027 VSS.n14026 0.00962857
R66080 VSS.n14026 VSS.n14024 0.00962857
R66081 VSS.n14024 VSS.n14023 0.00962857
R66082 VSS.n14023 VSS.n14022 0.00962857
R66083 VSS.n14022 VSS.n14021 0.00962857
R66084 VSS.n14021 VSS.n14016 0.00962857
R66085 VSS.n14016 VSS.n14015 0.00962857
R66086 VSS.n14015 VSS.n14012 0.00962857
R66087 VSS.n14012 VSS.n14011 0.00962857
R66088 VSS.n14011 VSS.n14009 0.00962857
R66089 VSS.n14009 VSS.n14008 0.00962857
R66090 VSS.n14008 VSS.n14006 0.00962857
R66091 VSS.n14006 VSS.n14005 0.00962857
R66092 VSS.n14005 VSS.n14004 0.00962857
R66093 VSS.n14004 VSS.n14003 0.00962857
R66094 VSS.n14003 VSS.n14002 0.00962857
R66095 VSS.n14002 VSS.n14001 0.00962857
R66096 VSS.n14001 VSS.n13997 0.00962857
R66097 VSS.n13997 VSS.n13996 0.00962857
R66098 VSS.n13996 VSS.n13994 0.00962857
R66099 VSS.n13994 VSS.n13993 0.00962857
R66100 VSS.n13993 VSS.n13991 0.00962857
R66101 VSS.n13991 VSS.n13990 0.00962857
R66102 VSS.n13990 VSS.n0 0.00962857
R66103 VSS.n22265 VSS.n2 0.00962857
R66104 VSS.n22107 VSS.n2 0.00962857
R66105 VSS.n22258 VSS.n22107 0.00962857
R66106 VSS.n20837 VSS.n444 0.00959676
R66107 VSS.n20745 VSS.n427 0.00959676
R66108 VSS.n20694 VSS.n410 0.00959676
R66109 VSS.n13255 VSS.n393 0.00959676
R66110 VSS.n13372 VSS.n392 0.00959676
R66111 VSS.n6949 VSS.n6948 0.00957614
R66112 VSS.n6847 VSS.n6846 0.00957614
R66113 VSS.n9659 VSS.n9658 0.00957614
R66114 VSS.n9542 VSS.n9541 0.00957614
R66115 VSS.n6948 VSS.n6947 0.00957614
R66116 VSS.n6846 VSS.n6845 0.00957614
R66117 VSS.n13679 VSS.n13677 0.00956429
R66118 VSS.n13949 VSS.n13948 0.00956429
R66119 VSS.n14119 VSS.n14118 0.00956429
R66120 VSS.n54 VSS.n53 0.00955028
R66121 VSS.n43 VSS.n41 0.00955028
R66122 VSS.n208 VSS.n206 0.00955028
R66123 VSS.n219 VSS.n218 0.00955028
R66124 VSS.n10316 VSS.n10315 0.00953846
R66125 VSS.n10434 VSS.n10433 0.00953846
R66126 VSS.n10342 VSS.n10341 0.00953846
R66127 VSS.n10149 VSS.n10148 0.00953846
R66128 VSS.n10057 VSS.n10056 0.00953846
R66129 VSS.n10024 VSS.n10023 0.00953846
R66130 VSS.n12370 VSS.n12369 0.00953846
R66131 VSS.n12488 VSS.n12487 0.00953846
R66132 VSS.n12396 VSS.n12395 0.00953846
R66133 VSS.n12200 VSS.n12199 0.00953846
R66134 VSS.n12108 VSS.n12107 0.00953846
R66135 VSS.n12075 VSS.n12074 0.00953846
R66136 VSS.n9843 VSS.n9842 0.00953846
R66137 VSS.n3967 VSS.n3966 0.00953543
R66138 VSS.n13113 VSS.n13112 0.00953543
R66139 VSS.n18958 VSS.n18957 0.00953543
R66140 VSS.n21765 VSS.n21764 0.00953543
R66141 VSS.n19050 VSS.n19049 0.00953543
R66142 VSS.n2601 VSS.n2600 0.00953543
R66143 VSS.n2515 VSS.n2514 0.00952778
R66144 VSS.n3941 VSS.n3940 0.00952778
R66145 VSS.n17200 VSS.n17199 0.00950322
R66146 VSS.n4658 VSS.n4657 0.00950322
R66147 VSS.n14146 VSS.n14145 0.0095
R66148 VSS.n14184 VSS.n14183 0.0095
R66149 VSS.n19400 VSS.n19399 0.0095
R66150 VSS.n19384 VSS.n19383 0.0095
R66151 VSS.n18266 VSS.n18264 0.0095
R66152 VSS.n16658 VSS.n16657 0.0095
R66153 VSS.n16620 VSS.n16618 0.0095
R66154 VSS.n16508 VSS.n16507 0.0095
R66155 VSS.n17214 VSS.n17213 0.00945304
R66156 VSS.n3230 VSS.n3229 0.00944366
R66157 VSS.n3313 VSS.n3312 0.00944366
R66158 VSS.n3365 VSS.n3364 0.00944366
R66159 VSS.n2928 VSS.n2927 0.00943572
R66160 VSS.n2992 VSS.n2991 0.00943572
R66161 VSS.n3040 VSS.n3039 0.00943572
R66162 VSS.n2555 VSS.n2554 0.00943572
R66163 VSS.n5194 VSS.n5193 0.00943572
R66164 VSS.n5245 VSS.n5244 0.00943572
R66165 VSS.n4966 VSS.n4965 0.00943572
R66166 VSS.n7079 VSS.n7078 0.00943572
R66167 VSS.n4459 VSS.n4458 0.00943572
R66168 VSS.n4408 VSS.n4407 0.00943572
R66169 VSS.n4373 VSS.n4372 0.00943572
R66170 VSS.n4319 VSS.n4318 0.00943572
R66171 VSS.n17972 VSS.n17971 0.00943572
R66172 VSS.n17818 VSS.n17817 0.00943572
R66173 VSS.n17773 VSS.n17772 0.00943572
R66174 VSS.n17709 VSS.n17708 0.00943572
R66175 VSS.n5653 VSS.n5651 0.00941892
R66176 VSS.n16029 VSS.n16028 0.00941892
R66177 VSS.n16043 VSS.n16042 0.00941892
R66178 VSS.n1004 VSS.n1003 0.00941892
R66179 VSS.n1022 VSS.n1011 0.00941892
R66180 VSS.n20911 VSS.n20910 0.00941892
R66181 VSS.n20920 VSS.n20918 0.00941892
R66182 VSS.n18421 VSS.n18420 0.00937324
R66183 VSS.n19608 VSS.n19607 0.00937324
R66184 VSS.n2724 VSS.n2723 0.00937143
R66185 VSS.n2784 VSS.n2783 0.00937143
R66186 VSS.n4946 VSS.n4945 0.00937143
R66187 VSS.n17544 VSS.n17543 0.00937143
R66188 VSS.n17486 VSS.n17485 0.00937143
R66189 VSS.n11985 VSS.n11984 0.0093706
R66190 VSS.n3955 VSS.n3954 0.00935827
R66191 VSS.n13125 VSS.n13124 0.00935827
R66192 VSS.n11857 VSS.n11856 0.00935827
R66193 VSS.n18970 VSS.n18969 0.00935827
R66194 VSS.n21753 VSS.n21752 0.00935827
R66195 VSS.n19038 VSS.n19037 0.00935827
R66196 VSS.n9868 VSS.n9852 0.00934615
R66197 VSS.n12672 VSS.n12656 0.00934615
R66198 VSS.n8887 VSS.n8886 0.00934615
R66199 VSS.n11994 VSS.n11980 0.00934615
R66200 VSS.n12635 VSS.n12634 0.00934615
R66201 VSS.n5108 VSS.n5107 0.00930714
R66202 VSS.n7270 VSS.n7269 0.00930714
R66203 VSS.n4546 VSS.n4545 0.00930714
R66204 VSS.n8870 VSS.n8869 0.00928172
R66205 VSS.n17108 VSS.n17106 0.009275
R66206 VSS.n17053 VSS.n17052 0.009275
R66207 VSS.n16955 VSS.n16954 0.009275
R66208 VSS.n14915 VSS.n14914 0.009275
R66209 VSS.n3201 VSS.n3200 0.00923239
R66210 VSS.n4205 VSS.n4204 0.0091811
R66211 VSS.n17450 VSS.n17449 0.0091811
R66212 VSS.n13144 VSS.n13143 0.0091811
R66213 VSS.n13224 VSS.n13223 0.0091811
R66214 VSS.n12232 VSS.n12231 0.0091811
R66215 VSS.n11956 VSS.n11955 0.0091811
R66216 VSS.n11889 VSS.n11888 0.0091811
R66217 VSS.n2235 VSS.n2234 0.0091811
R66218 VSS.n2201 VSS.n2200 0.0091811
R66219 VSS.n2284 VSS.n2283 0.0091811
R66220 VSS.n13341 VSS.n13340 0.0091811
R66221 VSS.n17892 VSS.n17891 0.0091811
R66222 VSS.n13484 VSS.n13483 0.0091811
R66223 VSS.n10180 VSS.n10179 0.0091811
R66224 VSS.n9958 VSS.n9957 0.0091811
R66225 VSS.n18464 VSS.n18463 0.00916197
R66226 VSS.n19575 VSS.n19574 0.00916197
R66227 VSS.n4659 VSS.n4658 0.00915406
R66228 VSS.n9870 VSS.n9869 0.00915385
R66229 VSS.n10372 VSS.n10371 0.00915385
R66230 VSS.n10371 VSS.n10370 0.00915385
R66231 VSS.n10087 VSS.n10086 0.00915385
R66232 VSS.n10086 VSS.n10085 0.00915385
R66233 VSS.n9995 VSS.n9994 0.00915385
R66234 VSS.n9994 VSS.n9993 0.00915385
R66235 VSS.n11771 VSS.n11770 0.00915385
R66236 VSS.n12426 VSS.n12425 0.00915385
R66237 VSS.n12425 VSS.n12424 0.00915385
R66238 VSS.n12138 VSS.n12137 0.00915385
R66239 VSS.n12137 VSS.n12136 0.00915385
R66240 VSS.n12046 VSS.n12045 0.00915385
R66241 VSS.n12045 VSS.n12044 0.00915385
R66242 VSS.n15373 VSS.n15372 0.00912168
R66243 VSS.n18696 VSS.n18695 0.00911913
R66244 VSS.n16890 VSS.n16889 0.00911913
R66245 VSS.n15546 VSS.n15545 0.00911913
R66246 VSS.n15456 VSS.n15455 0.00911913
R66247 VSS.n15360 VSS.n15359 0.00911913
R66248 VSS.n15317 VSS.n15316 0.00911913
R66249 VSS.n8562 VSS.n8561 0.00911913
R66250 VSS.n8532 VSS.n8531 0.00911913
R66251 VSS.n8327 VSS.n8326 0.00911913
R66252 VSS.n8417 VSS.n8416 0.00911913
R66253 VSS.n8387 VSS.n8386 0.00911913
R66254 VSS.n8360 VSS.n8359 0.00911913
R66255 VSS.n15455 VSS.n15454 0.00911913
R66256 VSS.n16889 VSS.n16888 0.00911913
R66257 VSS.n18695 VSS.n18694 0.00911913
R66258 VSS.n15547 VSS.n15546 0.00911913
R66259 VSS.n8416 VSS.n8415 0.00911913
R66260 VSS.n8386 VSS.n8385 0.00911913
R66261 VSS.n8361 VSS.n8360 0.00911913
R66262 VSS.n8561 VSS.n8560 0.00911913
R66263 VSS.n8531 VSS.n8530 0.00911913
R66264 VSS.n8328 VSS.n8327 0.00911913
R66265 VSS.n15318 VSS.n15317 0.00911913
R66266 VSS.n15359 VSS.n15358 0.00911913
R66267 VSS.n19178 VSS.n19177 0.00911913
R66268 VSS.n20026 VSS.n20025 0.00911913
R66269 VSS.n1834 VSS.n1833 0.00911913
R66270 VSS.n1758 VSS.n1757 0.00911913
R66271 VSS.n1675 VSS.n1674 0.00911913
R66272 VSS.n1632 VSS.n1631 0.00911913
R66273 VSS.n8713 VSS.n8712 0.00911913
R66274 VSS.n8683 VSS.n8682 0.00911913
R66275 VSS.n8123 VSS.n8122 0.00911913
R66276 VSS.n8225 VSS.n8224 0.00911913
R66277 VSS.n8195 VSS.n8194 0.00911913
R66278 VSS.n8169 VSS.n8168 0.00911913
R66279 VSS.n8168 VSS.n8167 0.00911913
R66280 VSS.n8712 VSS.n8711 0.00911913
R66281 VSS.n8682 VSS.n8681 0.00911913
R66282 VSS.n8124 VSS.n8123 0.00911913
R66283 VSS.n8224 VSS.n8223 0.00911913
R66284 VSS.n8194 VSS.n8193 0.00911913
R66285 VSS.n1633 VSS.n1632 0.00911913
R66286 VSS.n1676 VSS.n1675 0.00911913
R66287 VSS.n1757 VSS.n1756 0.00911913
R66288 VSS.n20027 VSS.n20026 0.00911913
R66289 VSS.n19177 VSS.n19176 0.00911913
R66290 VSS.n1835 VSS.n1834 0.00911913
R66291 VSS.n15293 VSS.n15292 0.00911702
R66292 VSS.n1595 VSS.n1593 0.00911702
R66293 VSS.n1602 VSS.n1601 0.00911702
R66294 VSS.n15496 VSS.n15493 0.00911702
R66295 VSS.n15516 VSS.n15513 0.00911702
R66296 VSS.n1786 VSS.n1783 0.00911702
R66297 VSS.n1798 VSS.n1795 0.00911702
R66298 VSS.n2857 VSS.n2856 0.00911429
R66299 VSS.n2861 VSS.n2860 0.00911429
R66300 VSS.n5133 VSS.n5132 0.00911429
R66301 VSS.n5137 VSS.n5136 0.00911429
R66302 VSS.n7243 VSS.n7242 0.00911429
R66303 VSS.n7241 VSS.n7240 0.00911429
R66304 VSS.n4520 VSS.n4519 0.00911429
R66305 VSS.n4518 VSS.n4517 0.00911429
R66306 VSS.n18037 VSS.n18036 0.00911429
R66307 VSS.n18039 VSS.n18038 0.00911429
R66308 VSS.n4173 VSS.n4171 0.00911111
R66309 VSS.n4176 VSS.n4173 0.00911111
R66310 VSS.n4182 VSS.n4180 0.00911111
R66311 VSS.n4186 VSS.n4182 0.00911111
R66312 VSS.n4186 VSS.n4184 0.00911111
R66313 VSS.n4192 VSS.n4190 0.00911111
R66314 VSS.n4197 VSS.n4192 0.00911111
R66315 VSS.n18983 VSS.n18981 0.00911111
R66316 VSS.n18985 VSS.n18983 0.00911111
R66317 VSS.n18990 VSS.n2164 0.00911111
R66318 VSS.n18992 VSS.n18990 0.00911111
R66319 VSS.n18994 VSS.n18992 0.00911111
R66320 VSS.n19000 VSS.n18998 0.00911111
R66321 VSS.n19002 VSS.n19000 0.00911111
R66322 VSS.n19004 VSS.n19002 0.00911111
R66323 VSS.n19006 VSS.n19004 0.00911111
R66324 VSS.n19012 VSS.n19010 0.00911111
R66325 VSS.n19014 VSS.n19012 0.00911111
R66326 VSS.n19016 VSS.n19014 0.00911111
R66327 VSS.n19018 VSS.n19016 0.00911111
R66328 VSS.n19024 VSS.n19022 0.00911111
R66329 VSS.n19026 VSS.n19024 0.00911111
R66330 VSS.n17884 VSS.n17875 0.00911111
R66331 VSS.n17884 VSS.n17882 0.00911111
R66332 VSS.n17882 VSS.n17880 0.00911111
R66333 VSS.n21739 VSS.n21737 0.00911111
R66334 VSS.n21741 VSS.n21739 0.00911111
R66335 VSS.n21733 VSS.n349 0.00911111
R66336 VSS.n21733 VSS.n21731 0.00911111
R66337 VSS.n21731 VSS.n21729 0.00911111
R66338 VSS.n21725 VSS.n21723 0.00911111
R66339 VSS.n21723 VSS.n21721 0.00911111
R66340 VSS.n21721 VSS.n21719 0.00911111
R66341 VSS.n21719 VSS.n21717 0.00911111
R66342 VSS.n21717 VSS.n21715 0.00911111
R66343 VSS.n21715 VSS.n21713 0.00911111
R66344 VSS.n11406 VSS.n11403 0.00911111
R66345 VSS.n11403 VSS.n11401 0.00911111
R66346 VSS.n11401 VSS.n11398 0.00911111
R66347 VSS.n11398 VSS.n11396 0.00911111
R66348 VSS.n11396 VSS.n11393 0.00911111
R66349 VSS.n11393 VSS.n11391 0.00911111
R66350 VSS.n11387 VSS.n11385 0.00911111
R66351 VSS.n11385 VSS.n11383 0.00911111
R66352 VSS.n11383 VSS.n11381 0.00911111
R66353 VSS.n11381 VSS.n11379 0.00911111
R66354 VSS.n11379 VSS.n11377 0.00911111
R66355 VSS.n11377 VSS.n11375 0.00911111
R66356 VSS.n14998 VSS.n14996 0.00911111
R66357 VSS.n16389 VSS.n14998 0.00911111
R66358 VSS.n16391 VSS.n16389 0.00911111
R66359 VSS.n16393 VSS.n16391 0.00911111
R66360 VSS.n16395 VSS.n16393 0.00911111
R66361 VSS.n16397 VSS.n16395 0.00911111
R66362 VSS.n16403 VSS.n16401 0.00911111
R66363 VSS.n16432 VSS.n16403 0.00911111
R66364 VSS.n16432 VSS.n16430 0.00911111
R66365 VSS.n16430 VSS.n16428 0.00911111
R66366 VSS.n748 VSS.n746 0.00911111
R66367 VSS.n1971 VSS.n748 0.00911111
R66368 VSS.n1973 VSS.n1971 0.00911111
R66369 VSS.n1975 VSS.n1973 0.00911111
R66370 VSS.n1981 VSS.n1979 0.00911111
R66371 VSS.n1983 VSS.n1981 0.00911111
R66372 VSS.n1985 VSS.n1983 0.00911111
R66373 VSS.n1994 VSS.n1985 0.00911111
R66374 VSS.n1994 VSS.n1992 0.00911111
R66375 VSS.n1992 VSS.n1990 0.00911111
R66376 VSS.n20836 VSS.n20834 0.00911111
R66377 VSS.n20870 VSS.n20836 0.00911111
R66378 VSS.n20870 VSS.n20868 0.00911111
R66379 VSS.n20868 VSS.n20866 0.00911111
R66380 VSS.n20866 VSS.n20864 0.00911111
R66381 VSS.n20864 VSS.n20862 0.00911111
R66382 VSS.n20858 VSS.n20856 0.00911111
R66383 VSS.n20856 VSS.n20854 0.00911111
R66384 VSS.n20854 VSS.n20852 0.00911111
R66385 VSS.n20852 VSS.n20850 0.00911111
R66386 VSS.n20850 VSS.n20848 0.00911111
R66387 VSS.n20848 VSS.n20846 0.00911111
R66388 VSS.n11480 VSS.n11478 0.00911111
R66389 VSS.n11483 VSS.n11480 0.00911111
R66390 VSS.n11485 VSS.n11483 0.00911111
R66391 VSS.n11488 VSS.n11485 0.00911111
R66392 VSS.n11490 VSS.n11488 0.00911111
R66393 VSS.n11492 VSS.n11490 0.00911111
R66394 VSS.n11498 VSS.n11496 0.00911111
R66395 VSS.n11500 VSS.n11498 0.00911111
R66396 VSS.n11502 VSS.n11500 0.00911111
R66397 VSS.n11511 VSS.n11502 0.00911111
R66398 VSS.n11511 VSS.n11509 0.00911111
R66399 VSS.n11509 VSS.n11507 0.00911111
R66400 VSS.n15114 VSS.n15112 0.00911111
R66401 VSS.n15130 VSS.n15114 0.00911111
R66402 VSS.n15130 VSS.n15128 0.00911111
R66403 VSS.n15128 VSS.n15126 0.00911111
R66404 VSS.n15126 VSS.n15124 0.00911111
R66405 VSS.n15124 VSS.n15122 0.00911111
R66406 VSS.n15118 VSS.n15116 0.00911111
R66407 VSS.n15116 VSS.n14972 0.00911111
R66408 VSS.n14972 VSS.n14970 0.00911111
R66409 VSS.n14970 VSS.n14968 0.00911111
R66410 VSS.n743 VSS.n741 0.00911111
R66411 VSS.n2085 VSS.n743 0.00911111
R66412 VSS.n2085 VSS.n2083 0.00911111
R66413 VSS.n2083 VSS.n2081 0.00911111
R66414 VSS.n2077 VSS.n2075 0.00911111
R66415 VSS.n2075 VSS.n2073 0.00911111
R66416 VSS.n2073 VSS.n2071 0.00911111
R66417 VSS.n2071 VSS.n2069 0.00911111
R66418 VSS.n2069 VSS.n2067 0.00911111
R66419 VSS.n2067 VSS.n2065 0.00911111
R66420 VSS.n20744 VSS.n20742 0.00911111
R66421 VSS.n20778 VSS.n20744 0.00911111
R66422 VSS.n20778 VSS.n20776 0.00911111
R66423 VSS.n20776 VSS.n20774 0.00911111
R66424 VSS.n20774 VSS.n20772 0.00911111
R66425 VSS.n20772 VSS.n20770 0.00911111
R66426 VSS.n20766 VSS.n20764 0.00911111
R66427 VSS.n20764 VSS.n20762 0.00911111
R66428 VSS.n20762 VSS.n20760 0.00911111
R66429 VSS.n20760 VSS.n20758 0.00911111
R66430 VSS.n20758 VSS.n20756 0.00911111
R66431 VSS.n20756 VSS.n20754 0.00911111
R66432 VSS.n11629 VSS.n11626 0.00911111
R66433 VSS.n11626 VSS.n11624 0.00911111
R66434 VSS.n11624 VSS.n11621 0.00911111
R66435 VSS.n11621 VSS.n11619 0.00911111
R66436 VSS.n11619 VSS.n11616 0.00911111
R66437 VSS.n11616 VSS.n11614 0.00911111
R66438 VSS.n11610 VSS.n11608 0.00911111
R66439 VSS.n11608 VSS.n11606 0.00911111
R66440 VSS.n11606 VSS.n11604 0.00911111
R66441 VSS.n11604 VSS.n11602 0.00911111
R66442 VSS.n11602 VSS.n11600 0.00911111
R66443 VSS.n11600 VSS.n11598 0.00911111
R66444 VSS.n15081 VSS.n15079 0.00911111
R66445 VSS.n15097 VSS.n15081 0.00911111
R66446 VSS.n15097 VSS.n15095 0.00911111
R66447 VSS.n15095 VSS.n15093 0.00911111
R66448 VSS.n15093 VSS.n15091 0.00911111
R66449 VSS.n15091 VSS.n15089 0.00911111
R66450 VSS.n15085 VSS.n15083 0.00911111
R66451 VSS.n15083 VSS.n14943 0.00911111
R66452 VSS.n14943 VSS.n14941 0.00911111
R66453 VSS.n14941 VSS.n14939 0.00911111
R66454 VSS.n738 VSS.n736 0.00911111
R66455 VSS.n20044 VSS.n738 0.00911111
R66456 VSS.n20046 VSS.n20044 0.00911111
R66457 VSS.n20048 VSS.n20046 0.00911111
R66458 VSS.n20054 VSS.n20052 0.00911111
R66459 VSS.n20056 VSS.n20054 0.00911111
R66460 VSS.n20058 VSS.n20056 0.00911111
R66461 VSS.n20067 VSS.n20058 0.00911111
R66462 VSS.n20067 VSS.n20065 0.00911111
R66463 VSS.n20065 VSS.n20063 0.00911111
R66464 VSS.n20693 VSS.n20691 0.00911111
R66465 VSS.n20727 VSS.n20693 0.00911111
R66466 VSS.n20727 VSS.n20725 0.00911111
R66467 VSS.n20725 VSS.n20723 0.00911111
R66468 VSS.n20723 VSS.n20721 0.00911111
R66469 VSS.n20721 VSS.n20719 0.00911111
R66470 VSS.n20715 VSS.n20713 0.00911111
R66471 VSS.n20713 VSS.n20711 0.00911111
R66472 VSS.n20711 VSS.n20709 0.00911111
R66473 VSS.n20709 VSS.n20707 0.00911111
R66474 VSS.n20707 VSS.n20705 0.00911111
R66475 VSS.n20705 VSS.n20703 0.00911111
R66476 VSS.n17232 VSS.n17184 0.00911111
R66477 VSS.n17184 VSS.n17183 0.00911111
R66478 VSS.n14343 VSS.n14341 0.00911111
R66479 VSS.n14343 VSS.n14342 0.00911111
R66480 VSS.n14349 VSS.n14348 0.00911111
R66481 VSS.n14348 VSS.n14347 0.00911111
R66482 VSS.n14359 VSS.n14358 0.00911111
R66483 VSS.n14382 VSS.n14380 0.00911111
R66484 VSS.n14383 VSS.n14382 0.00911111
R66485 VSS.n14384 VSS.n14383 0.00911111
R66486 VSS.n14387 VSS.n14386 0.00911111
R66487 VSS.n17166 VSS.n14387 0.00911111
R66488 VSS.n17167 VSS.n17166 0.00911111
R66489 VSS.n17168 VSS.n17167 0.00911111
R66490 VSS.n17170 VSS.n17169 0.00911111
R66491 VSS.n17169 VSS.n2131 0.00911111
R66492 VSS.n13519 VSS.n2131 0.00911111
R66493 VSS.n13520 VSS.n13519 0.00911111
R66494 VSS.n13523 VSS.n13522 0.00911111
R66495 VSS.n13525 VSS.n13523 0.00911111
R66496 VSS.n13525 VSS.n13524 0.00911111
R66497 VSS.n13431 VSS.n13428 0.00911111
R66498 VSS.n13278 VSS.n13277 0.00911111
R66499 VSS.n13421 VSS.n13278 0.00911111
R66500 VSS.n13273 VSS.n13272 0.00911111
R66501 VSS.n13268 VSS.n11769 0.00911111
R66502 VSS.n13266 VSS.n13265 0.00911111
R66503 VSS.n13265 VSS.n13264 0.00911111
R66504 VSS.n13264 VSS.n13263 0.00911111
R66505 VSS.n13263 VSS.n13262 0.00911111
R66506 VSS.n13262 VSS.n13261 0.00911111
R66507 VSS.n13261 VSS.n13260 0.00911111
R66508 VSS.n17375 VSS.n17372 0.00911111
R66509 VSS.n17372 VSS.n17370 0.00911111
R66510 VSS.n17366 VSS.n17364 0.00911111
R66511 VSS.n17364 VSS.n17362 0.00911111
R66512 VSS.n17362 VSS.n17360 0.00911111
R66513 VSS.n17360 VSS.n17358 0.00911111
R66514 VSS.n17358 VSS.n17356 0.00911111
R66515 VSS.n17356 VSS.n17354 0.00911111
R66516 VSS.n14392 VSS.n14390 0.00911111
R66517 VSS.n14433 VSS.n14392 0.00911111
R66518 VSS.n14435 VSS.n14433 0.00911111
R66519 VSS.n14437 VSS.n14435 0.00911111
R66520 VSS.n14439 VSS.n14437 0.00911111
R66521 VSS.n14441 VSS.n14439 0.00911111
R66522 VSS.n14447 VSS.n14445 0.00911111
R66523 VSS.n14669 VSS.n14447 0.00911111
R66524 VSS.n14669 VSS.n14667 0.00911111
R66525 VSS.n14667 VSS.n14665 0.00911111
R66526 VSS.n2135 VSS.n2133 0.00911111
R66527 VSS.n2137 VSS.n2135 0.00911111
R66528 VSS.n13438 VSS.n2137 0.00911111
R66529 VSS.n13440 VSS.n13438 0.00911111
R66530 VSS.n13446 VSS.n13444 0.00911111
R66531 VSS.n13448 VSS.n13446 0.00911111
R66532 VSS.n13450 VSS.n13448 0.00911111
R66533 VSS.n13459 VSS.n13450 0.00911111
R66534 VSS.n13459 VSS.n13457 0.00911111
R66535 VSS.n13457 VSS.n13455 0.00911111
R66536 VSS.n13371 VSS.n13369 0.00911111
R66537 VSS.n13405 VSS.n13371 0.00911111
R66538 VSS.n13405 VSS.n13403 0.00911111
R66539 VSS.n13403 VSS.n13401 0.00911111
R66540 VSS.n13401 VSS.n13399 0.00911111
R66541 VSS.n13399 VSS.n13397 0.00911111
R66542 VSS.n13393 VSS.n13391 0.00911111
R66543 VSS.n13391 VSS.n13389 0.00911111
R66544 VSS.n13389 VSS.n13387 0.00911111
R66545 VSS.n13387 VSS.n13385 0.00911111
R66546 VSS.n13385 VSS.n13383 0.00911111
R66547 VSS.n13383 VSS.n13381 0.00911111
R66548 VSS.n17409 VSS.n17407 0.00911111
R66549 VSS.n17412 VSS.n17409 0.00911111
R66550 VSS.n17418 VSS.n17416 0.00911111
R66551 VSS.n17420 VSS.n17418 0.00911111
R66552 VSS.n17422 VSS.n17420 0.00911111
R66553 VSS.n17424 VSS.n17422 0.00911111
R66554 VSS.n17426 VSS.n17424 0.00911111
R66555 VSS.n17431 VSS.n17426 0.00911111
R66556 VSS.n18113 VSS.n18111 0.00911111
R66557 VSS.n18115 VSS.n18113 0.00911111
R66558 VSS.n18117 VSS.n18115 0.00911111
R66559 VSS.n18119 VSS.n18117 0.00911111
R66560 VSS.n18121 VSS.n18119 0.00911111
R66561 VSS.n18123 VSS.n18121 0.00911111
R66562 VSS.n18129 VSS.n18127 0.00911111
R66563 VSS.n18137 VSS.n18129 0.00911111
R66564 VSS.n18137 VSS.n18134 0.00911111
R66565 VSS.n18134 VSS.n18132 0.00911111
R66566 VSS.n2146 VSS.n2144 0.00911111
R66567 VSS.n2144 VSS.n2142 0.00911111
R66568 VSS.n2142 VSS.n2139 0.00911111
R66569 VSS.n13465 VSS.n13463 0.00911111
R66570 VSS.n13471 VSS.n13465 0.00911111
R66571 VSS.n13471 VSS.n13469 0.00911111
R66572 VSS.n13469 VSS.n13467 0.00911111
R66573 VSS.n17962 VSS.n17957 0.00911111
R66574 VSS.n13282 VSS.n13280 0.00911111
R66575 VSS.n13314 VSS.n13282 0.00911111
R66576 VSS.n13314 VSS.n13312 0.00911111
R66577 VSS.n13312 VSS.n13310 0.00911111
R66578 VSS.n13310 VSS.n13308 0.00911111
R66579 VSS.n13308 VSS.n13306 0.00911111
R66580 VSS.n13302 VSS.n13301 0.00911111
R66581 VSS.n13301 VSS.n13299 0.00911111
R66582 VSS.n13299 VSS.n13296 0.00911111
R66583 VSS.n13296 VSS.n13294 0.00911111
R66584 VSS.n13294 VSS.n13291 0.00911111
R66585 VSS.n13291 VSS.n13289 0.00911111
R66586 VSS.n4105 VSS.n4104 0.00911111
R66587 VSS.n4104 VSS.n4102 0.00911111
R66588 VSS.n4102 VSS.n4099 0.00911111
R66589 VSS.n4099 VSS.n4097 0.00911111
R66590 VSS.n4097 VSS.n4094 0.00911111
R66591 VSS.n4094 VSS.n4092 0.00911111
R66592 VSS.n4087 VSS.n4085 0.00911111
R66593 VSS.n4085 VSS.n4083 0.00911111
R66594 VSS.n4083 VSS.n4081 0.00911111
R66595 VSS.n4081 VSS.n4079 0.00911111
R66596 VSS.n4079 VSS.n4077 0.00911111
R66597 VSS.n4077 VSS.n4075 0.00911111
R66598 VSS.n2169 VSS.n2167 0.00911111
R66599 VSS.n2171 VSS.n2169 0.00911111
R66600 VSS.n2173 VSS.n2171 0.00911111
R66601 VSS.n2175 VSS.n2173 0.00911111
R66602 VSS.n2177 VSS.n2175 0.00911111
R66603 VSS.n18850 VSS.n2177 0.00911111
R66604 VSS.n18846 VSS.n18844 0.00911111
R66605 VSS.n18844 VSS.n18842 0.00911111
R66606 VSS.n18842 VSS.n2181 0.00911111
R66607 VSS.n2181 VSS.n2179 0.00911111
R66608 VSS.n19374 VSS.n19372 0.00911111
R66609 VSS.n19372 VSS.n19172 0.00911111
R66610 VSS.n19172 VSS.n19170 0.00911111
R66611 VSS.n19170 VSS.n19168 0.00911111
R66612 VSS.n19164 VSS.n19162 0.00911111
R66613 VSS.n19162 VSS.n19160 0.00911111
R66614 VSS.n19160 VSS.n2160 0.00911111
R66615 VSS.n2160 VSS.n2158 0.00911111
R66616 VSS.n2158 VSS.n2156 0.00911111
R66617 VSS.n2156 VSS.n2154 0.00911111
R66618 VSS.n346 VSS.n344 0.00911111
R66619 VSS.n21875 VSS.n346 0.00911111
R66620 VSS.n21877 VSS.n21875 0.00911111
R66621 VSS.n21879 VSS.n21877 0.00911111
R66622 VSS.n21881 VSS.n21879 0.00911111
R66623 VSS.n21883 VSS.n21881 0.00911111
R66624 VSS.n21889 VSS.n21887 0.00911111
R66625 VSS.n21892 VSS.n21889 0.00911111
R66626 VSS.n21894 VSS.n21892 0.00911111
R66627 VSS.n21897 VSS.n21894 0.00911111
R66628 VSS.n21899 VSS.n21897 0.00911111
R66629 VSS.n21901 VSS.n21899 0.00911111
R66630 VSS.n8508 VSS.n8507 0.00905176
R66631 VSS.n8659 VSS.n8658 0.00905176
R66632 VSS.n18378 VSS.n18375 0.00905
R66633 VSS.n16564 VSS.n16563 0.00905
R66634 VSS.n161 VSS.n159 0.00904749
R66635 VSS.n327 VSS.n325 0.00904749
R66636 VSS.n3999 VSS.n3998 0.00900394
R66637 VSS.n13024 VSS.n13023 0.00900394
R66638 VSS.n18870 VSS.n18869 0.00900394
R66639 VSS.n21797 VSS.n21796 0.00900394
R66640 VSS.n19082 VSS.n19081 0.00900394
R66641 VSS.n21568 VSS.n21567 0.00900394
R66642 VSS.n3801 VSS.n3800 0.00900394
R66643 VSS.n3279 VSS.n3278 0.00900394
R66644 VSS.n16522 VSS.n14973 0.0089507
R66645 VSS.n816 VSS.n815 0.0089507
R66646 VSS.n4657 VSS.n4656 0.00885505
R66647 VSS.n17199 VSS.n17198 0.00885505
R66648 VSS.n3975 VSS.n3974 0.00882677
R66649 VSS.n4209 VSS.n4208 0.00882677
R66650 VSS.n13106 VSS.n13105 0.00882677
R66651 VSS.n13148 VSS.n13147 0.00882677
R66652 VSS.n18950 VSS.n18949 0.00882677
R66653 VSS.n2239 VSS.n2238 0.00882677
R66654 VSS.n21772 VSS.n21771 0.00882677
R66655 VSS.n2288 VSS.n2287 0.00882677
R66656 VSS.n19057 VSS.n19056 0.00882677
R66657 VSS.n17896 VSS.n17895 0.00882677
R66658 VSS.n21632 VSS.n21631 0.00882677
R66659 VSS.n3860 VSS.n3859 0.00882677
R66660 VSS.n2609 VSS.n2608 0.00882677
R66661 VSS.n19252 VSS.n19251 0.008825
R66662 VSS.n19267 VSS.n19264 0.008825
R66663 VSS.n16985 VSS.n16983 0.008825
R66664 VSS.n16975 VSS.n16974 0.008825
R66665 VSS.n1689 VSS.n1688 0.00878984
R66666 VSS.n17188 VSS.n17187 0.0087865
R66667 VSS.n17194 VSS.n17193 0.0087865
R66668 VSS.n17208 VSS.n17207 0.0087865
R66669 VSS.n10315 VSS.n10314 0.00876923
R66670 VSS.n10433 VSS.n10432 0.00876923
R66671 VSS.n10341 VSS.n10340 0.00876923
R66672 VSS.n10148 VSS.n10147 0.00876923
R66673 VSS.n10056 VSS.n10055 0.00876923
R66674 VSS.n10025 VSS.n10024 0.00876923
R66675 VSS.n12369 VSS.n12368 0.00876923
R66676 VSS.n12487 VSS.n12486 0.00876923
R66677 VSS.n12395 VSS.n12394 0.00876923
R66678 VSS.n12199 VSS.n12198 0.00876923
R66679 VSS.n12107 VSS.n12106 0.00876923
R66680 VSS.n12076 VSS.n12075 0.00876923
R66681 VSS.n3507 VSS.n3506 0.00866901
R66682 VSS.n3568 VSS.n3567 0.00866901
R66683 VSS.n3611 VSS.n3610 0.00866901
R66684 VSS.n3676 VSS.n3212 0.00866901
R66685 VSS.n3951 VSS.n3950 0.00864961
R66686 VSS.n13129 VSS.n13128 0.00864961
R66687 VSS.n12241 VSS.n12240 0.00864961
R66688 VSS.n18974 VSS.n18973 0.00864961
R66689 VSS.n21749 VSS.n21748 0.00864961
R66690 VSS.n19034 VSS.n19033 0.00864961
R66691 VSS.n10190 VSS.n10189 0.00864961
R66692 VSS.n18432 VSS.n18431 0.0086
R66693 VSS.n18363 VSS.n18362 0.0086
R66694 VSS.n16574 VSS.n16572 0.0086
R66695 VSS.n18916 VSS.n18915 0.00857235
R66696 VSS.n21847 VSS.n21846 0.00857235
R66697 VSS.n142 VSS.n141 0.00854469
R66698 VSS.n136 VSS.n134 0.00854469
R66699 VSS.n111 VSS.n110 0.00854469
R66700 VSS.n105 VSS.n103 0.00854469
R66701 VSS.n79 VSS.n78 0.00854469
R66702 VSS.n73 VSS.n71 0.00854469
R66703 VSS.n238 VSS.n236 0.00854469
R66704 VSS.n244 VSS.n243 0.00854469
R66705 VSS.n270 VSS.n268 0.00854469
R66706 VSS.n276 VSS.n275 0.00854469
R66707 VSS.n302 VSS.n300 0.00854469
R66708 VSS.n308 VSS.n307 0.00854469
R66709 VSS.n3651 DVSS 0.00852817
R66710 DVSS VSS.n3652 0.00852817
R66711 VSS.n9081 VSS.n9080 0.00851368
R66712 VSS.n9245 VSS.n9244 0.00851368
R66713 VSS.n6565 VSS.n6564 0.00851368
R66714 VSS.n1933 VSS.n1932 0.0084922
R66715 VSS.n15702 VSS.n15674 0.0084922
R66716 VSS.n11848 VSS.n11847 0.00847244
R66717 VSS.n8998 VSS.n8997 0.00847244
R66718 VSS.n2547 VSS.n2546 0.00847143
R66719 VSS.n4949 VSS.n4948 0.00847143
R66720 VSS.n7065 VSS.n7064 0.00847143
R66721 VSS.n7527 VSS.n7526 0.00847143
R66722 VSS.n4313 VSS.n4312 0.00847143
R66723 VSS.n17703 VSS.n17702 0.00847143
R66724 VSS.n13947 VSS.n13946 0.00847143
R66725 VSS.n10278 VSS.n10277 0.00838462
R66726 VSS.n10285 VSS.n10284 0.00838462
R66727 VSS.n10403 VSS.n10402 0.00838462
R66728 VSS.n10396 VSS.n10395 0.00838462
R66729 VSS.n10118 VSS.n10117 0.00838462
R66730 VSS.n10111 VSS.n10110 0.00838462
R66731 VSS.n8955 VSS.n8954 0.00838462
R66732 VSS.n8964 VSS.n8963 0.00838462
R66733 VSS.n12332 VSS.n12331 0.00838462
R66734 VSS.n12339 VSS.n12338 0.00838462
R66735 VSS.n12457 VSS.n12456 0.00838462
R66736 VSS.n12450 VSS.n12449 0.00838462
R66737 VSS.n12169 VSS.n12168 0.00838462
R66738 VSS.n12162 VSS.n12161 0.00838462
R66739 VSS.n12021 VSS.n12020 0.00838462
R66740 VSS.n12014 VSS.n12013 0.00838462
R66741 VSS.n9831 VSS.n9830 0.00838462
R66742 VSS.n9852 VSS.n9851 0.00838462
R66743 VSS.n12656 VSS.n12648 0.00838462
R66744 VSS.n12655 VSS.n12654 0.00838462
R66745 VSS.n17099 VSS.n17098 0.008375
R66746 VSS.n17063 VSS.n17061 0.008375
R66747 VSS.n16964 VSS.n16962 0.008375
R66748 VSS.n14928 VSS.n14927 0.008375
R66749 VSS.n16523 VSS.n16522 0.0083169
R66750 VSS.n815 VSS.n814 0.0083169
R66751 VSS.n9080 VSS.n9079 0.00829908
R66752 VSS.n9065 VSS.n9064 0.00829908
R66753 VSS.n14394 VSS.n14393 0.00829908
R66754 VSS.n14429 VSS.n14428 0.00829908
R66755 VSS.n15068 VSS.n15067 0.00829908
R66756 VSS.n15101 VSS.n15100 0.00829908
R66757 VSS.n15171 VSS.n15170 0.00829908
R66758 VSS.n13358 VSS.n13357 0.00829908
R66759 VSS.n13409 VSS.n13408 0.00829908
R66760 VSS.n20680 VSS.n20679 0.00829908
R66761 VSS.n20731 VSS.n20730 0.00829908
R66762 VSS.n20823 VSS.n20822 0.00829908
R66763 VSS.n536 VSS.n535 0.00829908
R66764 VSS.n6936 VSS.n6935 0.00829908
R66765 VSS.n21446 VSS.n21445 0.00829528
R66766 VSS.n4789 VSS.n4788 0.00829528
R66767 VSS.n14562 VSS.n14388 0.00828229
R66768 VSS.n14833 VSS.n14832 0.00828229
R66769 VSS.n16875 VSS.n16874 0.00828229
R66770 VSS.n16686 VSS.n16685 0.00828229
R66771 VSS.n16435 VSS.n16434 0.00828229
R66772 VSS.n19766 VSS.n19765 0.00828229
R66773 VSS.n19856 VSS.n19855 0.00828229
R66774 VSS.n20041 VSS.n20040 0.00828229
R66775 VSS.n2088 VSS.n2087 0.00828229
R66776 VSS.n854 VSS.n853 0.00828229
R66777 VSS.n5870 VSS.n5869 0.00825207
R66778 VSS.n5718 VSS.n5717 0.00825207
R66779 VSS.n5638 VSS.n5637 0.00825207
R66780 VSS.n16371 VSS.n16370 0.00825207
R66781 VSS.n16360 VSS.n16359 0.00825207
R66782 VSS.n16326 VSS.n16325 0.00825207
R66783 VSS.n16315 VSS.n16314 0.00825207
R66784 VSS.n16291 VSS.n16290 0.00825207
R66785 VSS.n16280 VSS.n16279 0.00825207
R66786 VSS.n16255 VSS.n16254 0.00825207
R66787 VSS.n16245 VSS.n16244 0.00825207
R66788 VSS.n16231 VSS.n16230 0.00825207
R66789 VSS.n16166 VSS.n16165 0.00825207
R66790 VSS.n16160 VSS.n16159 0.00825207
R66791 VSS.n16244 VSS.n16241 0.00825207
R66792 VSS.n16327 VSS.n16326 0.00825207
R66793 VSS.n16316 VSS.n16315 0.00825207
R66794 VSS.n16292 VSS.n16291 0.00825207
R66795 VSS.n16281 VSS.n16280 0.00825207
R66796 VSS.n16256 VSS.n16255 0.00825207
R66797 VSS.n16361 VSS.n16360 0.00825207
R66798 VSS.n16372 VSS.n16371 0.00825207
R66799 VSS.n5639 VSS.n5638 0.00825207
R66800 VSS.n16161 VSS.n16160 0.00825207
R66801 VSS.n5719 VSS.n5718 0.00825207
R66802 VSS.n16167 VSS.n16166 0.00825207
R66803 VSS.n5871 VSS.n5870 0.00825207
R66804 VSS.n16232 VSS.n16231 0.00825207
R66805 VSS.n21175 VSS.n21174 0.00825207
R66806 VSS.n21106 VSS.n21105 0.00825207
R66807 VSS.n21088 VSS.n21087 0.00825207
R66808 VSS.n21176 VSS.n21175 0.00825207
R66809 VSS.n21089 VSS.n21088 0.00825207
R66810 VSS.n21107 VSS.n21106 0.00825207
R66811 VSS.n1452 VSS.n1451 0.00825207
R66812 VSS.n1441 VSS.n1440 0.00825207
R66813 VSS.n1407 VSS.n1406 0.00825207
R66814 VSS.n1396 VSS.n1395 0.00825207
R66815 VSS.n1372 VSS.n1371 0.00825207
R66816 VSS.n1361 VSS.n1360 0.00825207
R66817 VSS.n1336 VSS.n1335 0.00825207
R66818 VSS.n1325 VSS.n1324 0.00825207
R66819 VSS.n1310 VSS.n1309 0.00825207
R66820 VSS.n1156 VSS.n1155 0.00825207
R66821 VSS.n1140 VSS.n1139 0.00825207
R66822 VSS.n1326 VSS.n1325 0.00825207
R66823 VSS.n1408 VSS.n1407 0.00825207
R66824 VSS.n1397 VSS.n1396 0.00825207
R66825 VSS.n1373 VSS.n1372 0.00825207
R66826 VSS.n1362 VSS.n1361 0.00825207
R66827 VSS.n1337 VSS.n1336 0.00825207
R66828 VSS.n1442 VSS.n1441 0.00825207
R66829 VSS.n1453 VSS.n1452 0.00825207
R66830 VSS.n1311 VSS.n1310 0.00825207
R66831 VSS.n1141 VSS.n1140 0.00825207
R66832 VSS.n1157 VSS.n1156 0.00825207
R66833 VSS.n13074 VSS.n13073 0.00824041
R66834 VSS.n19132 VSS.n19131 0.00824041
R66835 VSS.n2662 VSS.n2661 0.00824041
R66836 VSS.n4045 VSS.n4044 0.0082404
R66837 VSS.n6415 VSS.n6414 0.00818173
R66838 VSS.n3422 VSS.n3421 0.00817606
R66839 VSS.n5683 VSS.n5682 0.00815957
R66840 VSS.n5678 VSS.n5676 0.00815957
R66841 VSS.n20947 VSS.n20945 0.00815957
R66842 VSS.n20952 VSS.n20951 0.00815957
R66843 VSS.n5783 VSS.n5780 0.00815957
R66844 VSS.n5833 VSS.n5830 0.00815957
R66845 VSS.n5804 VSS.n5803 0.00815957
R66846 VSS.n5799 VSS.n5796 0.00815957
R66847 VSS.n1207 VSS.n1204 0.00815957
R66848 VSS.n1265 VSS.n1262 0.00815957
R66849 VSS.n1236 VSS.n1235 0.00815957
R66850 VSS.n1232 VSS.n1230 0.00815957
R66851 VSS.n19411 VSS.n19409 0.00815
R66852 VSS.n18255 VSS.n18254 0.00815
R66853 VSS.n16610 VSS.n16609 0.00815
R66854 VSS.n16518 VSS.n16517 0.00815
R66855 VSS.n12673 VSS.n12606 0.00811811
R66856 VSS.n10541 VSS.n10540 0.00811811
R66857 VSS.n3485 VSS.n3483 0.00803521
R66858 VSS.n10308 VSS.n10307 0.008
R66859 VSS.n10426 VSS.n10425 0.008
R66860 VSS.n10334 VSS.n10333 0.008
R66861 VSS.n10141 VSS.n10140 0.008
R66862 VSS.n10049 VSS.n10048 0.008
R66863 VSS.n10032 VSS.n10031 0.008
R66864 VSS.n21704 VSS.n21702 0.008
R66865 VSS.n11413 VSS.n11411 0.008
R66866 VSS.n20841 VSS.n20839 0.008
R66867 VSS.n20839 VSS.n20837 0.008
R66868 VSS.n11472 VSS.n11470 0.008
R66869 VSS.n20749 VSS.n20747 0.008
R66870 VSS.n20747 VSS.n20745 0.008
R66871 VSS.n11636 VSS.n11634 0.008
R66872 VSS.n20698 VSS.n20696 0.008
R66873 VSS.n20696 VSS.n20694 0.008
R66874 VSS.n17236 VSS.n17235 0.008
R66875 VSS.n13257 VSS.n13256 0.008
R66876 VSS.n13256 VSS.n13255 0.008
R66877 VSS.n17382 VSS.n17380 0.008
R66878 VSS.n13376 VSS.n13374 0.008
R66879 VSS.n13374 VSS.n13372 0.008
R66880 VSS.n371 VSS.n369 0.008
R66881 VSS.n12362 VSS.n12361 0.008
R66882 VSS.n12480 VSS.n12479 0.008
R66883 VSS.n12388 VSS.n12387 0.008
R66884 VSS.n12192 VSS.n12191 0.008
R66885 VSS.n12100 VSS.n12099 0.008
R66886 VSS.n12083 VSS.n12082 0.008
R66887 VSS.n21914 VSS.n21912 0.008
R66888 VSS.n2919 VSS.n2918 0.00795714
R66889 VSS.n2983 VSS.n2982 0.00795714
R66890 VSS.n3031 VSS.n3030 0.00795714
R66891 VSS.n5188 VSS.n5187 0.00795714
R66892 VSS.n5239 VSS.n5238 0.00795714
R66893 VSS.n5274 VSS.n5273 0.00795714
R66894 VSS.n7087 VSS.n7086 0.00795714
R66895 VSS.n4466 VSS.n4465 0.00795714
R66896 VSS.n4415 VSS.n4414 0.00795714
R66897 VSS.n4380 VSS.n4379 0.00795714
R66898 VSS.n4346 VSS.n4212 0.00795714
R66899 VSS.n17981 VSS.n17980 0.00795714
R66900 VSS.n17827 VSS.n17826 0.00795714
R66901 VSS.n17782 VSS.n17781 0.00795714
R66902 VSS.n17738 VSS.n17714 0.00795714
R66903 VSS.n12299 VSS.n12298 0.00794094
R66904 VSS.n10247 VSS.n10246 0.00794094
R66905 VSS.n17146 VSS.n17145 0.007925
R66906 VSS.n17006 VSS.n17004 0.007925
R66907 VSS.n16991 VSS.n16990 0.007925
R66908 VSS.n3238 VSS.n3237 0.00789437
R66909 VSS.n3321 VSS.n3320 0.00789437
R66910 VSS.n3375 VSS.n3374 0.00789437
R66911 VSS.n3437 VSS.n3436 0.00789437
R66912 VSS.n3469 VSS.n3468 0.00789437
R66913 VSS.n3204 VSS.n3203 0.00789437
R66914 VSS.n5598 VSS.n5597 0.00786815
R66915 VSS.n16114 VSS.n16113 0.00786815
R66916 VSS.n21048 VSS.n21047 0.00786815
R66917 VSS.n1094 VSS.n1093 0.00786815
R66918 VSS.n2520 VSS.n2518 0.00786111
R66919 VSS.n11415 VSS.n11413 0.00786111
R66920 VSS.n11470 VSS.n11468 0.00786111
R66921 VSS.n11638 VSS.n11636 0.00786111
R66922 VSS.n17237 VSS.n17236 0.00786111
R66923 VSS.n17384 VSS.n17382 0.00786111
R66924 VSS.n17398 VSS.n17396 0.00786111
R66925 VSS.n4118 VSS.n4116 0.00786111
R66926 VSS.n13848 VSS 0.00782857
R66927 VSS VSS.n13849 0.00782857
R66928 VSS.n3076 DVSS 0.00782857
R66929 DVSS VSS.n3077 0.00782857
R66930 VSS.n5306 DVSS 0.00782857
R66931 DVSS VSS.n5307 0.00782857
R66932 VSS.n7055 DVSS 0.00782857
R66933 DVSS VSS.n7050 0.00782857
R66934 VSS.n4347 DVSS 0.00782857
R66935 VSS.n4348 DVSS 0.00782857
R66936 VSS.n17740 DVSS 0.00782857
R66937 VSS.n17739 DVSS 0.00782857
R66938 VSS VSS.n22263 0.00782857
R66939 VSS VSS.n0 0.00782857
R66940 VSS.n13009 VSS.n13008 0.00781054
R66941 VSS.n13047 VSS.n13046 0.00781054
R66942 VSS.n13060 VSS.n13059 0.00781054
R66943 VSS.n13164 VSS.n13163 0.00781054
R66944 VSS.n13178 VSS.n13177 0.00781054
R66945 VSS.n12965 VSS.n12964 0.00781054
R66946 VSS.n12936 VSS.n12935 0.00781054
R66947 VSS.n12909 VSS.n12908 0.00781054
R66948 VSS.n12874 VSS.n12873 0.00781054
R66949 VSS.n12846 VSS.n12845 0.00781054
R66950 VSS.n12811 VSS.n12810 0.00781054
R66951 VSS.n12783 VSS.n12782 0.00781054
R66952 VSS.n12747 VSS.n12746 0.00781054
R66953 VSS.n12718 VSS.n12717 0.00781054
R66954 VSS.n13165 VSS.n13164 0.00781054
R66955 VSS.n12784 VSS.n12783 0.00781054
R66956 VSS.n12935 VSS.n12934 0.00781054
R66957 VSS.n12966 VSS.n12965 0.00781054
R66958 VSS.n12910 VSS.n12909 0.00781054
R66959 VSS.n12875 VSS.n12874 0.00781054
R66960 VSS.n12847 VSS.n12846 0.00781054
R66961 VSS.n13048 VSS.n13047 0.00781054
R66962 VSS.n13061 VSS.n13060 0.00781054
R66963 VSS.n13008 VSS.n13007 0.00781054
R66964 VSS.n12812 VSS.n12811 0.00781054
R66965 VSS.n13177 VSS.n13176 0.00781054
R66966 VSS.n21782 VSS.n21781 0.00781054
R66967 VSS.n21820 VSS.n21819 0.00781054
R66968 VSS.n21833 VSS.n21832 0.00781054
R66969 VSS.n2304 VSS.n2303 0.00781054
R66970 VSS.n2318 VSS.n2317 0.00781054
R66971 VSS.n20619 VSS.n20618 0.00781054
R66972 VSS.n20648 VSS.n20647 0.00781054
R66973 VSS.n20675 VSS.n20674 0.00781054
R66974 VSS.n20786 VSS.n20785 0.00781054
R66975 VSS.n20814 VSS.n20813 0.00781054
R66976 VSS.n21165 VSS.n21164 0.00781054
R66977 VSS.n21120 VSS.n21119 0.00781054
R66978 VSS.n21035 VSS.n21034 0.00781054
R66979 VSS.n20988 VSS.n20987 0.00781054
R66980 VSS.n6993 VSS.n6992 0.00781054
R66981 VSS.n6963 VSS.n6962 0.00781054
R66982 VSS.n6667 VSS.n6666 0.00781054
R66983 VSS.n6633 VSS.n6632 0.00781054
R66984 VSS.n6603 VSS.n6602 0.00781054
R66985 VSS.n6577 VSS.n6576 0.00781054
R66986 VSS.n2305 VSS.n2304 0.00781054
R66987 VSS.n21121 VSS.n21120 0.00781054
R66988 VSS.n20649 VSS.n20648 0.00781054
R66989 VSS.n20618 VSS.n20617 0.00781054
R66990 VSS.n20674 VSS.n20673 0.00781054
R66991 VSS.n20785 VSS.n20784 0.00781054
R66992 VSS.n20813 VSS.n20812 0.00781054
R66993 VSS.n21821 VSS.n21820 0.00781054
R66994 VSS.n21834 VSS.n21833 0.00781054
R66995 VSS.n21781 VSS.n21780 0.00781054
R66996 VSS.n2317 VSS.n2316 0.00781054
R66997 VSS.n21166 VSS.n21165 0.00781054
R66998 VSS.n19067 VSS.n19066 0.00781054
R66999 VSS.n19105 VSS.n19104 0.00781054
R67000 VSS.n19118 VSS.n19117 0.00781054
R67001 VSS.n17912 VSS.n17911 0.00781054
R67002 VSS.n17926 VSS.n17925 0.00781054
R67003 VSS.n20130 VSS.n20129 0.00781054
R67004 VSS.n20101 VSS.n20100 0.00781054
R67005 VSS.n20074 VSS.n20073 0.00781054
R67006 VSS.n2034 VSS.n2033 0.00781054
R67007 VSS.n2006 VSS.n2005 0.00781054
R67008 VSS.n1294 VSS.n1293 0.00781054
R67009 VSS.n1170 VSS.n1169 0.00781054
R67010 VSS.n1081 VSS.n1080 0.00781054
R67011 VSS.n1030 VSS.n1029 0.00781054
R67012 VSS.n6891 VSS.n6890 0.00781054
R67013 VSS.n6861 VSS.n6860 0.00781054
R67014 VSS.n6517 VSS.n6516 0.00781054
R67015 VSS.n6483 VSS.n6482 0.00781054
R67016 VSS.n6453 VSS.n6452 0.00781054
R67017 VSS.n6427 VSS.n6426 0.00781054
R67018 VSS.n17913 VSS.n17912 0.00781054
R67019 VSS.n1171 VSS.n1170 0.00781054
R67020 VSS.n20100 VSS.n20099 0.00781054
R67021 VSS.n20131 VSS.n20130 0.00781054
R67022 VSS.n20075 VSS.n20074 0.00781054
R67023 VSS.n2033 VSS.n2032 0.00781054
R67024 VSS.n2005 VSS.n2004 0.00781054
R67025 VSS.n19106 VSS.n19105 0.00781054
R67026 VSS.n19119 VSS.n19118 0.00781054
R67027 VSS.n19066 VSS.n19065 0.00781054
R67028 VSS.n17925 VSS.n17924 0.00781054
R67029 VSS.n1295 VSS.n1294 0.00781054
R67030 VSS.n21550 VSS.n21549 0.00781054
R67031 VSS.n21591 VSS.n21590 0.00781054
R67032 VSS.n21604 VSS.n21603 0.00781054
R67033 VSS.n21509 VSS.n21508 0.00781054
R67034 VSS.n21495 VSS.n21494 0.00781054
R67035 VSS.n21382 VSS.n21381 0.00781054
R67036 VSS.n21353 VSS.n21352 0.00781054
R67037 VSS.n21326 VSS.n21325 0.00781054
R67038 VSS.n21295 VSS.n21294 0.00781054
R67039 VSS.n21267 VSS.n21266 0.00781054
R67040 VSS.n7551 VSS.n7550 0.00781054
R67041 VSS.n7579 VSS.n7578 0.00781054
R67042 VSS.n7615 VSS.n7614 0.00781054
R67043 VSS.n7645 VSS.n7644 0.00781054
R67044 VSS.n7670 VSS.n7669 0.00781054
R67045 VSS.n7703 VSS.n7702 0.00781054
R67046 VSS.n7733 VSS.n7732 0.00781054
R67047 VSS.n7759 VSS.n7758 0.00781054
R67048 VSS.n7836 VSS.n7835 0.00781054
R67049 VSS.n7806 VSS.n7805 0.00781054
R67050 VSS.n7781 VSS.n7780 0.00781054
R67051 VSS.n21508 VSS.n21507 0.00781054
R67052 VSS.n7578 VSS.n7577 0.00781054
R67053 VSS.n7550 VSS.n7549 0.00781054
R67054 VSS.n21352 VSS.n21351 0.00781054
R67055 VSS.n21383 VSS.n21382 0.00781054
R67056 VSS.n21327 VSS.n21326 0.00781054
R67057 VSS.n21296 VSS.n21295 0.00781054
R67058 VSS.n21268 VSS.n21267 0.00781054
R67059 VSS.n21592 VSS.n21591 0.00781054
R67060 VSS.n21605 VSS.n21604 0.00781054
R67061 VSS.n21549 VSS.n21548 0.00781054
R67062 VSS.n21496 VSS.n21495 0.00781054
R67063 VSS.n6426 VSS.n6425 0.00781054
R67064 VSS.n7837 VSS.n7836 0.00781054
R67065 VSS.n6632 VSS.n6631 0.00781054
R67066 VSS.n6482 VSS.n6481 0.00781054
R67067 VSS.n7807 VSS.n7806 0.00781054
R67068 VSS.n6602 VSS.n6601 0.00781054
R67069 VSS.n6452 VSS.n6451 0.00781054
R67070 VSS.n6576 VSS.n6575 0.00781054
R67071 VSS.n7780 VSS.n7779 0.00781054
R67072 VSS.n7702 VSS.n7701 0.00781054
R67073 VSS.n6992 VSS.n6991 0.00781054
R67074 VSS.n6890 VSS.n6889 0.00781054
R67075 VSS.n7732 VSS.n7731 0.00781054
R67076 VSS.n6962 VSS.n6961 0.00781054
R67077 VSS.n6860 VSS.n6859 0.00781054
R67078 VSS.n7758 VSS.n7757 0.00781054
R67079 VSS.n6668 VSS.n6667 0.00781054
R67080 VSS.n6518 VSS.n6517 0.00781054
R67081 VSS.n7671 VSS.n7670 0.00781054
R67082 VSS.n1031 VSS.n1030 0.00781054
R67083 VSS.n20989 VSS.n20988 0.00781054
R67084 VSS.n12719 VSS.n12718 0.00781054
R67085 VSS.n7644 VSS.n7643 0.00781054
R67086 VSS.n12748 VSS.n12747 0.00781054
R67087 VSS.n7614 VSS.n7613 0.00781054
R67088 VSS.n21034 VSS.n21033 0.00781054
R67089 VSS.n1080 VSS.n1079 0.00781054
R67090 VSS.n6836 VSS.n6835 0.00780945
R67091 VSS.n9532 VSS.n9531 0.00780945
R67092 VSS.n9649 VSS.n9648 0.00780945
R67093 VSS.n15311 VSS.n15309 0.0077973
R67094 VSS.n15315 VSS.n15312 0.0077973
R67095 VSS.n1629 VSS.n1628 0.0077973
R67096 VSS.n1619 VSS.n1618 0.0077973
R67097 VSS.n14156 VSS.n14155 0.00779557
R67098 VSS.n14200 VSS.n14199 0.00779557
R67099 VSS.n14188 VSS.n14187 0.0077955
R67100 VSS.n14141 VSS.n14140 0.00779539
R67101 VSS.n14134 VSS.n14133 0.00779449
R67102 VSS.n14171 VSS.n14170 0.00779449
R67103 VSS.n14160 VSS.n14159 0.00779416
R67104 VSS.n14196 VSS.n14195 0.00779416
R67105 VSS.n14152 VSS.n14151 0.00779335
R67106 VSS.n14137 VSS.n14136 0.00779236
R67107 VSS.n17190 VSS.n17189 0.0077918
R67108 VSS.n17196 VSS.n17195 0.0077918
R67109 VSS.n17204 VSS.n17203 0.0077918
R67110 VSS.n17210 VSS.n17209 0.0077918
R67111 VSS.n17216 VSS.n17215 0.0077918
R67112 VSS.n3946 VSS.n2450 0.00776378
R67113 VSS.n13134 VSS.n13133 0.00776378
R67114 VSS.n18979 VSS.n18978 0.00776378
R67115 VSS.n21744 VSS.n21743 0.00776378
R67116 VSS.n19029 VSS.n19028 0.00776378
R67117 VSS.n19394 VSS.n19393 0.0077
R67118 VSS.n19390 VSS.n19388 0.0077
R67119 VSS.n18272 VSS.n18270 0.0077
R67120 VSS.n16652 VSS.n16651 0.0077
R67121 VSS.n16625 VSS.n16623 0.0077
R67122 VSS.n18159 VSS.n18158 0.0076831
R67123 VSS.n19697 VSS.n19696 0.0076831
R67124 VSS.n15475 VSS.n15474 0.0076451
R67125 VSS.n15474 VSS.n15473 0.0076451
R67126 VSS.n1776 VSS.n1775 0.0076451
R67127 VSS.n1777 VSS.n1776 0.0076451
R67128 VSS.n9878 VSS.n9877 0.00761538
R67129 VSS.n10379 VSS.n10378 0.00761538
R67130 VSS.n10364 VSS.n10363 0.00761538
R67131 VSS.n10094 VSS.n10093 0.00761538
R67132 VSS.n10079 VSS.n10078 0.00761538
R67133 VSS.n10002 VSS.n10001 0.00761538
R67134 VSS.n9987 VSS.n9986 0.00761538
R67135 VSS.n11779 VSS.n11778 0.00761538
R67136 VSS.n12433 VSS.n12432 0.00761538
R67137 VSS.n12418 VSS.n12417 0.00761538
R67138 VSS.n12145 VSS.n12144 0.00761538
R67139 VSS.n12130 VSS.n12129 0.00761538
R67140 VSS.n12053 VSS.n12052 0.00761538
R67141 VSS.n12038 VSS.n12037 0.00761538
R67142 VSS.n13661 VSS.n13660 0.00757143
R67143 VSS.n22256 VSS.n22255 0.00757143
R67144 VSS.n5110 VSS.n5109 0.00750714
R67145 VSS.n7271 VSS.n7268 0.00750714
R67146 VSS.n4547 VSS.n4544 0.00750714
R67147 VSS.n17113 VSS.n17111 0.007475
R67148 VSS.n17047 VSS.n17046 0.007475
R67149 VSS.n14907 VSS.n14906 0.007475
R67150 VSS.n12534 VSS.n12533 0.00740945
R67151 VSS.n21643 VSS.n21642 0.00740945
R67152 VSS.n3872 VSS.n3871 0.00740945
R67153 VSS.n10479 VSS.n10478 0.00740945
R67154 VSS.n5164 VSS.n5162 0.00737857
R67155 VSS.n7214 VSS.n7213 0.00737857
R67156 VSS.n4492 VSS.n4491 0.00737857
R67157 VSS.n12685 VSS.n12684 0.00735992
R67158 VSS.n10553 VSS.n10552 0.00735992
R67159 VSS.n1466 VSS.n1465 0.00733971
R67160 VSS.n12822 VSS.n12821 0.00733971
R67161 VSS.n21191 VSS.n21190 0.00733971
R67162 VSS.n7542 VSS.n445 0.00733971
R67163 VSS.n16383 VSS.n16382 0.00733971
R67164 VSS.n5882 VSS.n5881 0.00733971
R67165 VSS.n11240 VSS.n11239 0.00733971
R67166 VSS.n14241 VSS.n14240 0.00731429
R67167 VSS.n21989 VSS.n21988 0.00731429
R67168 VSS.n13615 VSS.n13614 0.00725
R67169 VSS.n18386 VSS.n18383 0.00725
R67170 VSS.n18251 VSS.n18250 0.00725
R67171 VSS.n16558 VSS.n16557 0.00725
R67172 VSS.n2669 VSS.n2668 0.00725
R67173 VSS.n2713 VSS.n2712 0.00725
R67174 VSS.n2773 VSS.n2772 0.00725
R67175 VSS.n2843 VSS.n2842 0.00725
R67176 VSS.n3003 VSS.n3002 0.00725
R67177 VSS.n3051 VSS.n3050 0.00725
R67178 VSS.n2550 VSS.n2549 0.00725
R67179 VSS.n2825 VSS.n2824 0.00725
R67180 VSS.n4992 VSS.n4991 0.00725
R67181 VSS.n5022 VSS.n5021 0.00725
R67182 VSS.n5068 VSS.n5067 0.00725
R67183 VSS.n5122 VSS.n5121 0.00725
R67184 VSS.n5150 VSS.n5149 0.00725
R67185 VSS.n4952 VSS.n4951 0.00725
R67186 VSS.n7402 VSS.n7401 0.00725
R67187 VSS.n7370 VSS.n7369 0.00725
R67188 VSS.n7316 VSS.n7315 0.00725
R67189 VSS.n7254 VSS.n7253 0.00725
R67190 VSS.n7228 VSS.n7227 0.00725
R67191 VSS.n4632 VSS.n4631 0.00725
R67192 VSS.n4586 VSS.n4585 0.00725
R67193 VSS.n4532 VSS.n4531 0.00725
R67194 VSS.n4504 VSS.n4503 0.00725
R67195 VSS.n4316 VSS.n4315 0.00725
R67196 VSS.n18072 VSS.n18070 0.00725
R67197 VSS.n17555 VSS.n17554 0.00725
R67198 VSS.n17497 VSS.n17496 0.00725
R67199 VSS.n18053 VSS.n18052 0.00725
R67200 VSS.n17706 VSS.n17705 0.00725
R67201 VSS.n14127 VSS.n14126 0.00725
R67202 VSS.n12535 VSS.n12534 0.00723228
R67203 VSS.n10480 VSS.n10479 0.00723228
R67204 VSS.n10323 VSS.n10322 0.00723077
R67205 VSS.n10441 VSS.n10440 0.00723077
R67206 VSS.n10349 VSS.n10348 0.00723077
R67207 VSS.n10156 VSS.n10155 0.00723077
R67208 VSS.n10064 VSS.n10063 0.00723077
R67209 VSS.n10017 VSS.n10016 0.00723077
R67210 VSS.n12377 VSS.n12376 0.00723077
R67211 VSS.n12495 VSS.n12494 0.00723077
R67212 VSS.n12403 VSS.n12402 0.00723077
R67213 VSS.n12207 VSS.n12206 0.00723077
R67214 VSS.n12115 VSS.n12114 0.00723077
R67215 VSS.n12068 VSS.n12067 0.00723077
R67216 VSS.n15395 VSS.n15394 0.00722377
R67217 VSS.n15396 VSS.n15395 0.00722377
R67218 VSS.n1711 VSS.n1710 0.00722377
R67219 VSS.n1712 VSS.n1711 0.00722377
R67220 VSS.n13243 VSS.n13242 0.00722225
R67221 VSS.n13003 VSS.n13002 0.00722225
R67222 VSS.n12902 VSS.n12901 0.00722225
R67223 VSS.n12889 VSS.n12888 0.00722225
R67224 VSS.n12835 VSS.n12834 0.00722225
R67225 VSS.n13503 VSS.n13502 0.00722225
R67226 VSS.n13436 VSS.n13435 0.00722225
R67227 VSS.n2049 VSS.n734 0.00722225
R67228 VSS.n2048 VSS.n2047 0.00722225
R67229 VSS.n879 VSS.n744 0.00722225
R67230 VSS.n597 VSS.n596 0.00722225
R67231 VSS.n584 VSS.n583 0.00722225
R67232 VSS.n3232 VSS.n3231 0.00719014
R67233 VSS.n3315 VSS.n3314 0.00719014
R67234 VSS.n3369 VSS.n3368 0.00719014
R67235 VSS.n17349 VSS.n17348 0.00716351
R67236 VSS.n17328 VSS.n17327 0.00716351
R67237 VSS.n11517 VSS.n11516 0.00716351
R67238 VSS.n11329 VSS.n11328 0.00716351
R67239 VSS.n11314 VSS.n11313 0.00716351
R67240 VSS.n13250 VSS.n13249 0.00716351
R67241 VSS.n12998 VSS.n12997 0.00716351
R67242 VSS.n12895 VSS.n12894 0.00716351
R67243 VSS.n12882 VSS.n12881 0.00716351
R67244 VSS.n12828 VSS.n12827 0.00716351
R67245 VSS.n14403 VSS.n14402 0.00716351
R67246 VSS.n14420 VSS.n14419 0.00716351
R67247 VSS.n15077 VSS.n15076 0.00716351
R67248 VSS.n15110 VSS.n15109 0.00716351
R67249 VSS.n15180 VSS.n15179 0.00716351
R67250 VSS.n13367 VSS.n13366 0.00716351
R67251 VSS.n13418 VSS.n13417 0.00716351
R67252 VSS.n20689 VSS.n20688 0.00716351
R67253 VSS.n20740 VSS.n20739 0.00716351
R67254 VSS.n20832 VSS.n20831 0.00716351
R67255 VSS.n13510 VSS.n13509 0.00716351
R67256 VSS.n20150 VSS.n20149 0.00716351
R67257 VSS.n2056 VSS.n2055 0.00716351
R67258 VSS.n2041 VSS.n2040 0.00716351
R67259 VSS.n886 VSS.n885 0.00716351
R67260 VSS.n590 VSS.n589 0.00716351
R67261 VSS.n577 VSS.n576 0.00716351
R67262 VSS.n527 VSS.n526 0.00716351
R67263 VSS.n17215 VSS.n17214 0.00706681
R67264 VSS.n17203 VSS.n17202 0.00706681
R67265 VSS.n17195 VSS.n17194 0.00706681
R67266 VSS.n17189 VSS.n17188 0.00706681
R67267 VSS.n17209 VSS.n17208 0.00706681
R67268 VSS.n18468 VSS.n18467 0.0070493
R67269 VSS.n16894 VSS.n16893 0.0070493
R67270 VSS.n19571 VSS.n19570 0.0070493
R67271 VSS.n20022 VSS.n20021 0.0070493
R67272 VSS.n19244 VSS.n19243 0.007025
R67273 VSS.n19275 VSS.n19272 0.007025
R67274 VSS.n16990 VSS.n16989 0.007025
R67275 VSS.n16969 VSS.n16968 0.007025
R67276 VSS.n521 VSS.n520 0.00700754
R67277 VSS.n2898 VSS.n2893 0.00699286
R67278 VSS.n18007 VSS.n18006 0.00699286
R67279 VSS.n3544 VSS.n3542 0.00690845
R67280 VSS.n3604 VSS.n3601 0.00690845
R67281 VSS.n3646 VSS.n3644 0.00690845
R67282 VSS.n17342 VSS.n17341 0.00689005
R67283 VSS.n17335 VSS.n17334 0.00689005
R67284 VSS.n11524 VSS.n11523 0.00689005
R67285 VSS.n11322 VSS.n4859 0.00689005
R67286 VSS.n11321 VSS.n11320 0.00689005
R67287 VSS.n21679 VSS.n21678 0.00687795
R67288 VSS.n4140 VSS.n4139 0.00687795
R67289 VSS.n4987 VSS.n4986 0.00686429
R67290 VSS.n5017 VSS.n5016 0.00686429
R67291 VSS.n5063 VSS.n5062 0.00686429
R67292 VSS.n7408 VSS.n7407 0.00686429
R67293 VSS.n4639 VSS.n4637 0.00686429
R67294 VSS.n4593 VSS.n4591 0.00686429
R67295 VSS.n9886 VSS.n9885 0.00684615
R67296 VSS.n10293 VSS.n10292 0.00684615
R67297 VSS.n10411 VSS.n10410 0.00684615
R67298 VSS.n10388 VSS.n10387 0.00684615
R67299 VSS.n10126 VSS.n10125 0.00684615
R67300 VSS.n10103 VSS.n10102 0.00684615
R67301 VSS.n9978 VSS.n9977 0.00684615
R67302 VSS.n12565 VSS.n12564 0.00684615
R67303 VSS.n12347 VSS.n12346 0.00684615
R67304 VSS.n12465 VSS.n12464 0.00684615
R67305 VSS.n12442 VSS.n12441 0.00684615
R67306 VSS.n12177 VSS.n12176 0.00684615
R67307 VSS.n12154 VSS.n12153 0.00684615
R67308 VSS.n12029 VSS.n12028 0.00684615
R67309 VSS.n9847 VSS.n9846 0.00684615
R67310 VSS.n12639 VSS.n12638 0.00684615
R67311 VSS.n14175 VSS.n14174 0.0068424
R67312 VSS.n14174 VSS.n14173 0.0068424
R67313 VSS.n18416 VSS.n18413 0.0068
R67314 VSS.n165 VSS.n164 0.00678492
R67315 VSS.n11251 VSS.n5903 0.00678492
R67316 VSS.n5477 VSS.n5476 0.00668725
R67317 VSS.n4922 VSS.n4921 0.00668725
R67318 VSS.n4858 VSS.n4857 0.00668725
R67319 VSS.n14291 VSS.n11744 0.00668725
R67320 VSS.n17310 VSS.n17309 0.00668725
R67321 VSS.n14214 VSS.n14209 0.00667143
R67322 VSS.n5215 VSS.n5213 0.00667143
R67323 VSS.n5266 VSS.n5264 0.00667143
R67324 VSS.n5301 VSS.n5299 0.00667143
R67325 VSS.n7060 VSS.n7059 0.00667143
R67326 VSS.n4441 VSS.n4440 0.00667143
R67327 VSS.n4390 VSS.n4389 0.00667143
R67328 VSS.n4355 VSS.n4354 0.00667143
R67329 VSS.n13945 VSS.n13944 0.00667143
R67330 VSS.n16940 VSS.n14903 0.00662676
R67331 VSS.n19975 VSS.n19974 0.00662676
R67332 VSS.n14163 VSS.n14162 0.00661798
R67333 VSS.n14192 VSS.n14191 0.00661798
R67334 VSS.n14193 VSS.n14192 0.00661798
R67335 VSS.n17223 VSS.n17222 0.00661798
R67336 VSS.n7379 VSS.n7377 0.00660714
R67337 VSS.n7324 VSS.n7323 0.00660714
R67338 VSS.n5748 VSS.n5747 0.0065738
R67339 VSS.n16196 VSS.n16195 0.0065738
R67340 VSS.n16197 VSS.n16196 0.0065738
R67341 VSS.n5749 VSS.n5748 0.0065738
R67342 VSS.n21138 VSS.n21137 0.0065738
R67343 VSS.n21139 VSS.n21138 0.0065738
R67344 VSS.n1188 VSS.n1187 0.0065738
R67345 VSS.n1189 VSS.n1188 0.0065738
R67346 VSS.n8878 VSS.n8877 0.00656106
R67347 VSS.n8885 VSS.n8884 0.00656106
R67348 VSS.n8884 VSS.n8883 0.00656106
R67349 VSS.n11978 VSS.n11977 0.00656106
R67350 VSS.n11979 VSS.n11978 0.00656106
R67351 VSS.n11993 VSS.n11992 0.00656106
R67352 VSS.n17463 VSS.n17462 0.00652362
R67353 VSS.n13211 VSS.n13210 0.00652362
R67354 VSS.n2214 VSS.n2213 0.00652362
R67355 VSS.n13328 VSS.n13327 0.00652362
R67356 VSS.n17940 VSS.n17939 0.00652362
R67357 VSS.n21459 VSS.n21458 0.00652362
R67358 VSS.n4776 VSS.n4775 0.00652362
R67359 VSS.n10790 VSS.n8785 0.0065
R67360 VSS.n10905 VSS.n8100 0.0065
R67361 VSS.n10650 VSS.n10649 0.0065
R67362 VSS.n10782 VSS.n10771 0.0065
R67363 VSS.n11025 VSS.n11024 0.0065
R67364 VSS.n10787 VSS.n10782 0.0065
R67365 VSS.n10651 VSS.n10650 0.0065
R67366 VSS.n10886 VSS.n10885 0.0065
R67367 VSS.n10885 VSS.n10880 0.0065
R67368 VSS.n11024 VSS.n11023 0.0065
R67369 VSS.n9802 VSS.n9410 0.0065
R67370 VSS.n8785 VSS.n8453 0.0065
R67371 VSS.n8100 VSS.n6784 0.0065
R67372 VSS.n7999 VSS.n7906 0.0065
R67373 VSS.n10654 VSS.n9802 0.0065
R67374 VSS.n10300 VSS.n10299 0.00646154
R67375 VSS.n10418 VSS.n10417 0.00646154
R67376 VSS.n10133 VSS.n10132 0.00646154
R67377 VSS.n10041 VSS.n10040 0.00646154
R67378 VSS.n10040 VSS.n10039 0.00646154
R67379 VSS.n12354 VSS.n12353 0.00646154
R67380 VSS.n12472 VSS.n12471 0.00646154
R67381 VSS.n12184 VSS.n12183 0.00646154
R67382 VSS.n12092 VSS.n12091 0.00646154
R67383 VSS.n12091 VSS.n12090 0.00646154
R67384 VSS.n15319 VSS.n15318 0.00641549
R67385 VSS.n19519 VSS.n19518 0.00641549
R67386 VSS.n17222 VSS.n17221 0.00639353
R67387 VSS.n17229 VSS.n17228 0.00639353
R67388 VSS.n14151 VSS.n14150 0.00639353
R67389 VSS.n7155 VSS.n7154 0.00635
R67390 VSS.n7096 VSS.n7095 0.00635
R67391 VSS.n21447 VSS.n21446 0.00634646
R67392 VSS.n4788 VSS.n4787 0.00634646
R67393 VSS.n21429 VSS.n21428 0.00628209
R67394 VSS.n21418 VSS.n21417 0.00628209
R67395 VSS.n21319 VSS.n21318 0.00628209
R67396 VSS.n21308 VSS.n21307 0.00628209
R67397 VSS.n21256 VSS.n21255 0.00628209
R67398 VSS.n17249 VSS.n17248 0.00628209
R67399 VSS.n11743 VSS.n11742 0.00628209
R67400 VSS.n4923 VSS.n4797 0.00628209
R67401 VSS.n11464 VSS.n11463 0.00628209
R67402 VSS.n11241 VSS.n5414 0.00628209
R67403 VSS.n21424 VSS.n21423 0.0062233
R67404 VSS.n21413 VSS.n21412 0.0062233
R67405 VSS.n21314 VSS.n21313 0.0062233
R67406 VSS.n21303 VSS.n21302 0.0062233
R67407 VSS.n21251 VSS.n21250 0.0062233
R67408 VSS.n17244 VSS.n17243 0.0062233
R67409 VSS.n11738 VSS.n11737 0.0062233
R67410 VSS.n4928 VSS.n4927 0.0062233
R67411 VSS.n11459 VSS.n11458 0.0062233
R67412 VSS.n11246 VSS.n11245 0.0062233
R67413 VSS.n5619 VSS.n5618 0.00622032
R67414 VSS.n16135 VSS.n16134 0.00622032
R67415 VSS.n16136 VSS.n16135 0.00622032
R67416 VSS.n5620 VSS.n5619 0.00622032
R67417 VSS.n21069 VSS.n21068 0.00622032
R67418 VSS.n21070 VSS.n21069 0.00622032
R67419 VSS.n1115 VSS.n1114 0.00622032
R67420 VSS.n1116 VSS.n1115 0.00622032
R67421 VSS.n8465 VSS.n8464 0.00620423
R67422 VSS.n8547 VSS.n8546 0.00620423
R67423 VSS.n8313 VSS.n8312 0.00620423
R67424 VSS.n8402 VSS.n8401 0.00620423
R67425 VSS.n8375 VSS.n8374 0.00620423
R67426 VSS.n8616 VSS.n8615 0.00620423
R67427 VSS.n8698 VSS.n8697 0.00620423
R67428 VSS.n8109 VSS.n8108 0.00620423
R67429 VSS.n8210 VSS.n8209 0.00620423
R67430 VSS.n8183 VSS.n8182 0.00620423
R67431 VSS.n5658 VSS.n5657 0.00617568
R67432 VSS.n5533 VSS.n5532 0.00617568
R67433 VSS.n16078 VSS.n16077 0.00617568
R67434 VSS.n16038 VSS.n16037 0.00617568
R67435 VSS.n1047 VSS.n1046 0.00617568
R67436 VSS.n1017 VSS.n1016 0.00617568
R67437 VSS.n21001 VSS.n20999 0.00617568
R67438 VSS.n20927 VSS.n20924 0.00617568
R67439 VSS.n18486 VSS.n18485 0.00616099
R67440 VSS.n14960 VSS.n14959 0.00616099
R67441 VSS.n14767 VSS.n14766 0.00616099
R67442 VSS.n14655 VSS.n14654 0.00616099
R67443 VSS.n14929 VSS.n14928 0.00616099
R67444 VSS.n16420 VSS.n16419 0.00616099
R67445 VSS.n15895 VSS.n15894 0.00616099
R67446 VSS.n5190 VSS.n5189 0.00615714
R67447 VSS.n5241 VSS.n5240 0.00615714
R67448 VSS.n5276 VSS.n5275 0.00615714
R67449 VSS.n5310 VSS.n5309 0.00615714
R67450 VSS.n7085 VSS.n7084 0.00615714
R67451 VSS.n7053 VSS.n7052 0.00615714
R67452 VSS.n4467 VSS.n4464 0.00615714
R67453 VSS.n4416 VSS.n4413 0.00615714
R67454 VSS.n4381 VSS.n4378 0.00615714
R67455 VSS.n19247 VSS.n19244 0.006125
R67456 VSS.n19272 VSS.n19271 0.006125
R67457 VSS.n16989 VSS.n16988 0.006125
R67458 VSS.n16971 VSS.n16969 0.006125
R67459 VSS.n9887 VSS.n9886 0.00607692
R67460 VSS.n10387 VSS.n10386 0.00607692
R67461 VSS.n10356 VSS.n10355 0.00607692
R67462 VSS.n10102 VSS.n10101 0.00607692
R67463 VSS.n10071 VSS.n10070 0.00607692
R67464 VSS.n10010 VSS.n10009 0.00607692
R67465 VSS.n9979 VSS.n9978 0.00607692
R67466 VSS.n12566 VSS.n12565 0.00607692
R67467 VSS.n12441 VSS.n12440 0.00607692
R67468 VSS.n12410 VSS.n12409 0.00607692
R67469 VSS.n12153 VSS.n12152 0.00607692
R67470 VSS.n12122 VSS.n12121 0.00607692
R67471 VSS.n12061 VSS.n12060 0.00607692
R67472 VSS.n12030 VSS.n12029 0.00607692
R67473 VSS.n9846 VSS.n9845 0.00607692
R67474 VSS.n12638 VSS.n12637 0.00607692
R67475 VSS.n19243 VSS.n19242 0.00607384
R67476 VSS.n18662 VSS.n18661 0.00607384
R67477 VSS.n16861 VSS.n16860 0.00607384
R67478 VSS.n19777 VSS.n19776 0.00607384
R67479 VSS.n14466 VSS.n14465 0.00607384
R67480 VSS.n17137 VSS.n17136 0.00607384
R67481 VSS.n16672 VSS.n16671 0.00607384
R67482 VSS.n15711 VSS.n15710 0.00607384
R67483 VSS.n145 VSS.n142 0.00603073
R67484 VSS.n134 VSS.n133 0.00603073
R67485 VSS.n114 VSS.n111 0.00603073
R67486 VSS.n103 VSS.n102 0.00603073
R67487 VSS.n82 VSS.n79 0.00603073
R67488 VSS.n71 VSS.n70 0.00603073
R67489 VSS.n236 VSS.n235 0.00603073
R67490 VSS.n247 VSS.n244 0.00603073
R67491 VSS.n268 VSS.n267 0.00603073
R67492 VSS.n279 VSS.n276 0.00603073
R67493 VSS.n300 VSS.n299 0.00603073
R67494 VSS.n311 VSS.n308 0.00603073
R67495 VSS.n342 VSS.n337 0.00603073
R67496 VSS.n21243 VSS.n21240 0.00603073
R67497 VSS.n18436 VSS.n18425 0.00599296
R67498 VSS.n14901 VSS.n14900 0.00599296
R67499 VSS.n16578 VSS.n16577 0.00599296
R67500 VSS.n15348 VSS.n15347 0.00599296
R67501 VSS.n8468 VSS.n8467 0.00599296
R67502 VSS.n8485 VSS.n8484 0.00599296
R67503 VSS.n8550 VSS.n8549 0.00599296
R67504 VSS.n8316 VSS.n8315 0.00599296
R67505 VSS.n8405 VSS.n8404 0.00599296
R67506 VSS.n8372 VSS.n8371 0.00599296
R67507 VSS.n8356 VSS.n8355 0.00599296
R67508 VSS.n19603 VSS.n19602 0.00599296
R67509 VSS.n19972 VSS.n19971 0.00599296
R67510 VSS.n790 VSS.n789 0.00599296
R67511 VSS.n1664 VSS.n1663 0.00599296
R67512 VSS.n8619 VSS.n8618 0.00599296
R67513 VSS.n8636 VSS.n8635 0.00599296
R67514 VSS.n8701 VSS.n8700 0.00599296
R67515 VSS.n8112 VSS.n8111 0.00599296
R67516 VSS.n8213 VSS.n8212 0.00599296
R67517 VSS.n8180 VSS.n8179 0.00599296
R67518 VSS.n8164 VSS.n8163 0.00599296
R67519 VSS.n3950 VSS.n3949 0.00599213
R67520 VSS.n13130 VSS.n13129 0.00599213
R67521 VSS.n11896 VSS.n11895 0.00599213
R67522 VSS.n18975 VSS.n18974 0.00599213
R67523 VSS.n21748 VSS.n21747 0.00599213
R67524 VSS.n19033 VSS.n19032 0.00599213
R67525 VSS.n9895 VSS.n9894 0.00599213
R67526 VSS.n4981 VSS.n4976 0.00596429
R67527 VSS.n5008 VSS.n5006 0.00596429
R67528 VSS.n5038 VSS.n5036 0.00596429
R67529 VSS.n5084 VSS.n5082 0.00596429
R67530 VSS.n7418 VSS.n7417 0.00596429
R67531 VSS.n7388 VSS.n7387 0.00596429
R67532 VSS.n4618 VSS.n4617 0.00596429
R67533 VSS.n4572 VSS.n4571 0.00596429
R67534 VSS.n14195 VSS.n14194 0.00594456
R67535 VSS.n8881 VSS.n8880 0.00594375
R67536 VSS.n3432 VSS.n3431 0.00592254
R67537 VSS.n3475 VSS.n3474 0.00592254
R67538 VSS.n14168 VSS.n14167 0.0059
R67539 VSS.n18383 VSS.n18382 0.0059
R67540 VSS.n16560 VSS.n16558 0.0059
R67541 VSS.n2588 VSS.n2587 0.0059
R67542 VSS.n2705 VSS.n2704 0.0059
R67543 VSS.n2765 VSS.n2764 0.0059
R67544 VSS.n17563 VSS.n17562 0.0059
R67545 VSS.n17505 VSS.n17504 0.0059
R67546 VSS.n13108 VSS.n13107 0.00587205
R67547 VSS.n11975 VSS.n11974 0.00584085
R67548 VSS.n11980 VSS.n11979 0.00581245
R67549 VSS.n11992 VSS.n11985 0.00581245
R67550 VSS.n8877 VSS.n8870 0.00581245
R67551 VSS.n8886 VSS.n8885 0.00581245
R67552 VSS.n11977 VSS.n11976 0.00581245
R67553 VSS.n8883 VSS.n8882 0.00581245
R67554 VSS.n18717 VSS.n18716 0.00578169
R67555 VSS.n18732 VSS.n18731 0.00578169
R67556 VSS.n18755 VSS.n18754 0.00578169
R67557 VSS.n18169 VSS.n18168 0.00578169
R67558 VSS.n17083 VSS.n17082 0.00578169
R67559 VSS.n14900 VSS.n14899 0.00578169
R67560 VSS.n8525 VSS.n8524 0.00578169
R67561 VSS.n8343 VSS.n8342 0.00578169
R67562 VSS.n19199 VSS.n19198 0.00578169
R67563 VSS.n19214 VSS.n19213 0.00578169
R67564 VSS.n19237 VSS.n19236 0.00578169
R67565 VSS.n19687 VSS.n19686 0.00578169
R67566 VSS.n19882 VSS.n19881 0.00578169
R67567 VSS.n19971 VSS.n19970 0.00578169
R67568 VSS.n8676 VSS.n8675 0.00578169
R67569 VSS.n8139 VSS.n8138 0.00578169
R67570 VSS.n5685 VSS.n5683 0.00576596
R67571 VSS.n5676 VSS.n5675 0.00576596
R67572 VSS.n16019 VSS.n16017 0.00576596
R67573 VSS.n16009 VSS.n16004 0.00576596
R67574 VSS.n1000 VSS.n998 0.00576596
R67575 VSS.n990 VSS.n981 0.00576596
R67576 VSS.n20945 VSS.n20944 0.00576596
R67577 VSS.n20954 VSS.n20952 0.00576596
R67578 VSS.n5780 VSS.n5779 0.00576596
R67579 VSS.n5830 VSS.n5829 0.00576596
R67580 VSS.n5805 VSS.n5804 0.00576596
R67581 VSS.n5796 VSS.n5795 0.00576596
R67582 VSS.n1204 VSS.n1203 0.00576596
R67583 VSS.n1262 VSS.n1261 0.00576596
R67584 VSS.n1238 VSS.n1236 0.00576596
R67585 VSS.n18485 VSS.n18484 0.0057309
R67586 VSS.n14962 VSS.n14960 0.0057309
R67587 VSS.n14766 VSS.n14765 0.0057309
R67588 VSS.n14657 VSS.n14655 0.0057309
R67589 VSS.n14931 VSS.n14929 0.0057309
R67590 VSS.n16422 VSS.n16420 0.0057309
R67591 VSS.n15897 VSS.n15895 0.0057309
R67592 VSS.n14172 VSS.n14171 0.00572004
R67593 VSS.n4673 VSS.n4671 0.00570714
R67594 VSS.n22008 VSS.n22007 0.00567998
R67595 VSS.n17111 VSS.n17110 0.005675
R67596 VSS.n17049 VSS.n17047 0.005675
R67597 VSS.n16951 VSS.n16950 0.005675
R67598 VSS.n14910 VSS.n14907 0.005675
R67599 VSS.n2959 VSS.n2957 0.00564286
R67600 VSS.n3023 VSS.n3021 0.00564286
R67601 VSS.n3072 VSS.n3069 0.00564286
R67602 VSS.n17853 VSS.n17852 0.00564286
R67603 VSS.n17792 VSS.n17791 0.00564286
R67604 VSS.n17747 VSS.n17746 0.00564286
R67605 VSS.n3511 VSS.n3510 0.00564085
R67606 VSS.n3570 VSS.n3569 0.00564085
R67607 VSS.n3613 VSS.n3612 0.00564085
R67608 VSS.n18685 VSS.n18684 0.00560681
R67609 VSS.n19242 VSS.n19241 0.00559337
R67610 VSS.n18661 VSS.n18660 0.00559337
R67611 VSS.n16860 VSS.n16859 0.00559337
R67612 VSS.n19776 VSS.n19775 0.00559337
R67613 VSS.n14465 VSS.n14464 0.00559337
R67614 VSS.n17136 VSS.n17135 0.00559337
R67615 VSS.n16671 VSS.n16670 0.00559337
R67616 VSS.n15710 VSS.n15709 0.00559337
R67617 VSS.n4666 VSS.n4650 0.00557857
R67618 VSS.n14877 VSS.n14876 0.00557042
R67619 VSS.n16528 VSS.n16527 0.00557042
R67620 VSS.n19948 VSS.n19947 0.00557042
R67621 VSS.n810 VSS.n809 0.00557042
R67622 VSS.n159 VSS.n158 0.00552793
R67623 VSS.n325 VSS.n324 0.00552793
R67624 VSS.n13229 VSS.n13228 0.00551772
R67625 VSS.n13346 VSS.n13345 0.00551772
R67626 VSS.n13489 VSS.n13488 0.00551772
R67627 VSS.n12720 VSS.n12719 0.00546063
R67628 VSS.n14180 VSS.n14179 0.00545
R67629 VSS.n13671 VSS.n13612 0.00545
R67630 VSS.n19396 VSS.n19394 0.00545
R67631 VSS.n19388 VSS.n19387 0.00545
R67632 VSS.n19382 VSS.n19380 0.00545
R67633 VSS.n18270 VSS.n18269 0.00545
R67634 VSS.n16654 VSS.n16652 0.00545
R67635 VSS.n16623 VSS.n16622 0.00545
R67636 VSS.n4942 VSS.n4941 0.00545
R67637 VSS.n4996 VSS.n4995 0.00545
R67638 VSS.n5026 VSS.n5025 0.00545
R67639 VSS.n5072 VSS.n5071 0.00545
R67640 VSS.n5117 VSS.n5116 0.00545
R67641 VSS.n5156 VSS.n5155 0.00545
R67642 VSS.n5206 VSS.n5205 0.00545
R67643 VSS.n5257 VSS.n5256 0.00545
R67644 VSS.n5292 VSS.n5291 0.00545
R67645 VSS.n4960 VSS.n4959 0.00545
R67646 VSS.n5913 VSS.n5912 0.00545
R67647 VSS.n7399 VSS.n7398 0.00545
R67648 VSS.n7260 VSS.n7259 0.00545
R67649 VSS.n7223 VSS.n7222 0.00545
R67650 VSS.n7069 VSS.n7068 0.00545
R67651 VSS.n7531 VSS.n7530 0.00545
R67652 VSS.n4629 VSS.n4628 0.00545
R67653 VSS.n4583 VSS.n4582 0.00545
R67654 VSS.n4538 VSS.n4537 0.00545
R67655 VSS.n4499 VSS.n4498 0.00545
R67656 VSS.n4449 VSS.n4448 0.00545
R67657 VSS.n4398 VSS.n4397 0.00545
R67658 VSS.n4363 VSS.n4362 0.00545
R67659 VSS.n14121 VSS.n14120 0.00545
R67660 VSS.n13666 VSS.n13664 0.00543435
R67661 VSS.n22259 VSS.n22258 0.00543435
R67662 VSS.n5659 VSS.n5658 0.00536486
R67663 VSS.n5532 VSS.n5530 0.00536486
R67664 VSS.n16078 VSS.n16073 0.00536486
R67665 VSS.n16037 VSS.n16035 0.00536486
R67666 VSS.n1047 VSS.n1042 0.00536486
R67667 VSS.n1016 VSS.n1014 0.00536486
R67668 VSS.n21001 VSS.n20998 0.00536486
R67669 VSS.n20928 VSS.n20927 0.00536486
R67670 VSS.n3305 VSS.n3303 0.00535915
R67671 VSS.n3343 VSS.n3341 0.00535915
R67672 VSS.n3397 VSS.n3395 0.00535915
R67673 VSS.n3675 VSS.n3674 0.00535915
R67674 VSS.n17081 VSS.n17080 0.00535915
R67675 VSS.n17016 VSS.n17015 0.00535915
R67676 VSS.n16916 VSS.n16915 0.00535915
R67677 VSS.n16633 VSS.n16632 0.00535915
R67678 VSS.n19884 VSS.n19883 0.00535915
R67679 VSS.n19919 VSS.n19918 0.00535915
R67680 VSS.n20000 VSS.n19999 0.00535915
R67681 VSS.n765 VSS.n764 0.00535915
R67682 VSS.n21244 VSS.n21243 0.00535333
R67683 VSS.n13198 VSS.n13197 0.00534055
R67684 VSS.n17953 VSS.n17952 0.00534055
R67685 VSS.n18138 VSS.n2182 0.00532561
R67686 VSS.n18164 VSS.n18163 0.00532561
R67687 VSS.n18171 VSS.n18170 0.00532561
R67688 VSS.n18146 VSS.n18145 0.00532561
R67689 VSS.n19685 VSS.n19684 0.00532561
R67690 VSS.n19710 VSS.n19709 0.00532561
R67691 VSS.n10535 VSS.n10534 0.00530769
R67692 VSS.n9892 VSS.n9887 0.00530769
R67693 VSS.n10386 VSS.n10385 0.00530769
R67694 VSS.n10361 VSS.n10356 0.00530769
R67695 VSS.n10101 VSS.n10100 0.00530769
R67696 VSS.n10076 VSS.n10071 0.00530769
R67697 VSS.n10009 VSS.n10008 0.00530769
R67698 VSS.n9984 VSS.n9979 0.00530769
R67699 VSS.n8888 VSS.n8887 0.00530769
R67700 VSS.n12601 VSS.n12600 0.00530769
R67701 VSS.n12571 VSS.n12566 0.00530769
R67702 VSS.n12440 VSS.n12439 0.00530769
R67703 VSS.n12415 VSS.n12410 0.00530769
R67704 VSS.n12152 VSS.n12151 0.00530769
R67705 VSS.n12127 VSS.n12122 0.00530769
R67706 VSS.n12060 VSS.n12059 0.00530769
R67707 VSS.n12035 VSS.n12030 0.00530769
R67708 VSS.n11995 VSS.n11994 0.00530769
R67709 VSS.n9845 VSS.n9844 0.00530769
R67710 VSS.n12637 VSS.n12636 0.00530769
R67711 VSS.n11551 VSS.n11550 0.00528346
R67712 VSS.n11575 VSS.n11574 0.00528346
R67713 VSS.n9481 VSS.n9480 0.00528346
R67714 VSS.n9568 VSS.n9567 0.00528346
R67715 VSS.n9022 VSS.n9021 0.00528346
R67716 VSS.n9131 VSS.n9130 0.00528346
R67717 VSS.n9107 VSS.n9106 0.00528346
R67718 VSS.n12951 VSS.n12950 0.00528346
R67719 VSS.n12924 VSS.n12923 0.00528346
R67720 VSS.n12733 VSS.n12732 0.00528346
R67721 VSS.n12707 VSS.n12706 0.00528346
R67722 VSS.n12503 VSS.n12326 0.00528346
R67723 VSS.n18953 VSS.n18952 0.00528346
R67724 VSS.n15025 VSS.n15024 0.00528346
R67725 VSS.n15050 VSS.n15049 0.00528346
R67726 VSS.n9598 VSS.n9597 0.00528346
R67727 VSS.n9685 VSS.n9684 0.00528346
R67728 VSS.n9165 VSS.n9164 0.00528346
R67729 VSS.n9294 VSS.n9293 0.00528346
R67730 VSS.n9270 VSS.n9269 0.00528346
R67731 VSS.n20633 VSS.n20632 0.00528346
R67732 VSS.n20660 VSS.n20659 0.00528346
R67733 VSS.n6912 VSS.n6911 0.00528346
R67734 VSS.n6978 VSS.n6977 0.00528346
R67735 VSS.n6653 VSS.n6652 0.00528346
R67736 VSS.n6618 VSS.n6617 0.00528346
R67737 VSS.n6591 VSS.n6590 0.00528346
R67738 VSS.n20116 VSS.n20115 0.00528346
R67739 VSS.n20089 VSS.n20088 0.00528346
R67740 VSS.n6789 VSS.n6788 0.00528346
R67741 VSS.n6876 VSS.n6875 0.00528346
R67742 VSS.n6503 VSS.n6502 0.00528346
R67743 VSS.n6468 VSS.n6467 0.00528346
R67744 VSS.n6441 VSS.n6440 0.00528346
R67745 VSS.n21368 VSS.n21367 0.00528346
R67746 VSS.n21341 VSS.n21340 0.00528346
R67747 VSS.n7629 VSS.n7628 0.00528346
R67748 VSS.n7656 VSS.n7655 0.00528346
R67749 VSS.n7717 VSS.n7716 0.00528346
R67750 VSS.n7744 VSS.n7743 0.00528346
R67751 VSS.n7822 VSS.n7821 0.00528346
R67752 VSS.n7795 VSS.n7794 0.00528346
R67753 VSS.n11684 VSS.n11683 0.00528346
R67754 VSS.n11659 VSS.n11658 0.00528346
R67755 VSS.n6127 VSS.n6126 0.00528346
R67756 VSS.n6103 VSS.n6102 0.00528346
R67757 VSS.n6046 VSS.n6045 0.00528346
R67758 VSS.n6022 VSS.n6021 0.00528346
R67759 VSS.n5965 VSS.n5964 0.00528346
R67760 VSS.n5941 VSS.n5940 0.00528346
R67761 VSS.n641 VSS.n640 0.00528346
R67762 VSS.n617 VSS.n616 0.00528346
R67763 VSS.n10599 VSS.n10598 0.00528346
R67764 VSS.n10575 VSS.n10574 0.00528346
R67765 VSS.n10449 VSS.n10272 0.00528346
R67766 VSS.n8882 VSS.n8881 0.00527824
R67767 VSS.n7251 VSS.n7250 0.00525714
R67768 VSS.n17213 VSS.n17212 0.00522582
R67769 VSS.n18404 VSS.n18403 0.0052251
R67770 VSS.n19618 VSS.n19617 0.0052251
R67771 VSS.n17148 VSS.n17146 0.005225
R67772 VSS.n17004 VSS.n17003 0.005225
R67773 VSS.n2521 VSS.n2520 0.00522222
R67774 VSS.n21705 VSS.n21704 0.00522222
R67775 VSS.n17399 VSS.n17398 0.00522222
R67776 VSS.n372 VSS.n371 0.00522222
R67777 VSS.n4116 VSS.n4114 0.00522222
R67778 VSS.n21912 VSS.n21910 0.00522222
R67779 VSS.n3296 VSS.n3295 0.00521831
R67780 VSS.n3334 VSS.n3333 0.00521831
R67781 VSS.n3388 VSS.n3387 0.00521831
R67782 VSS.n3668 VSS.n3667 0.00521831
R67783 VSS.n21455 VSS.n21454 0.00520602
R67784 VSS.n7189 VSS.n7187 0.00519286
R67785 VSS.n7129 VSS.n7128 0.00519286
R67786 VSS.n11976 VSS.n11975 0.0051892
R67787 VSS.n14564 VSS.n14563 0.00518499
R67788 VSS.n14831 VSS.n14830 0.00518499
R67789 VSS.n16877 VSS.n16876 0.00518499
R67790 VSS.n16688 VSS.n16687 0.00518499
R67791 VSS.n16437 VSS.n16436 0.00518499
R67792 VSS.n15427 VSS.n15416 0.00518499
R67793 VSS.n19764 VSS.n19763 0.00518499
R67794 VSS.n19854 VSS.n19853 0.00518499
R67795 VSS.n20039 VSS.n20038 0.00518499
R67796 VSS.n2090 VSS.n2089 0.00518499
R67797 VSS.n852 VSS.n851 0.00518499
R67798 VSS.n3523 VSS.n3522 0.00514789
R67799 VSS.n3582 VSS.n3581 0.00514789
R67800 VSS.n3625 VSS.n3624 0.00514789
R67801 VSS.n18726 VSS.n18725 0.00514789
R67802 VSS.n18727 VSS.n18726 0.00514789
R67803 VSS.n18731 VSS.n18730 0.00514789
R67804 VSS.n18790 VSS.n18789 0.00514789
R67805 VSS.n18802 VSS.n18801 0.00514789
R67806 VSS.n18207 VSS.n18206 0.00514789
R67807 VSS.n16594 VSS.n16593 0.00514789
R67808 VSS.n15523 VSS.n15522 0.00514789
R67809 VSS.n8482 VSS.n8481 0.00514789
R67810 VSS.n19208 VSS.n19207 0.00514789
R67811 VSS.n19209 VSS.n19208 0.00514789
R67812 VSS.n19213 VSS.n19212 0.00514789
R67813 VSS.n19462 VSS.n19461 0.00514789
R67814 VSS.n19474 VSS.n19473 0.00514789
R67815 VSS.n19649 VSS.n19648 0.00514789
R67816 VSS.n774 VSS.n773 0.00514789
R67817 VSS.n1811 VSS.n1810 0.00514789
R67818 VSS.n8633 VSS.n8632 0.00514789
R67819 VSS.n7232 VSS.n7231 0.00512857
R67820 VSS.n18786 VSS.n18785 0.0051193
R67821 VSS.n19458 VSS.n19457 0.0051193
R67822 VSS.n17020 VSS.n17019 0.00511916
R67823 VSS.n19915 VSS.n19914 0.00511916
R67824 VSS.n11548 VSS.n11547 0.0051063
R67825 VSS.n11578 VSS.n11577 0.0051063
R67826 VSS.n5575 VSS.n5574 0.0051063
R67827 VSS.n9484 VSS.n9483 0.0051063
R67828 VSS.n9571 VSS.n9570 0.0051063
R67829 VSS.n9025 VSS.n9024 0.0051063
R67830 VSS.n9134 VSS.n9133 0.0051063
R67831 VSS.n9104 VSS.n9103 0.0051063
R67832 VSS.n9087 VSS.n9086 0.0051063
R67833 VSS.n12954 VSS.n12953 0.0051063
R67834 VSS.n12921 VSS.n12920 0.0051063
R67835 VSS.n12736 VSS.n12735 0.0051063
R67836 VSS.n12704 VSS.n12703 0.0051063
R67837 VSS.n15022 VSS.n15021 0.0051063
R67838 VSS.n15053 VSS.n15052 0.0051063
R67839 VSS.n16091 VSS.n16090 0.0051063
R67840 VSS.n9601 VSS.n9600 0.0051063
R67841 VSS.n9688 VSS.n9687 0.0051063
R67842 VSS.n9168 VSS.n9167 0.0051063
R67843 VSS.n9297 VSS.n9296 0.0051063
R67844 VSS.n9267 VSS.n9266 0.0051063
R67845 VSS.n9251 VSS.n9250 0.0051063
R67846 VSS.n20630 VSS.n20629 0.0051063
R67847 VSS.n20663 VSS.n20662 0.0051063
R67848 VSS.n21023 VSS.n21022 0.0051063
R67849 VSS.n6915 VSS.n6914 0.0051063
R67850 VSS.n6981 VSS.n6980 0.0051063
R67851 VSS.n6656 VSS.n6655 0.0051063
R67852 VSS.n6621 VSS.n6620 0.0051063
R67853 VSS.n6588 VSS.n6587 0.0051063
R67854 VSS.n6571 VSS.n6570 0.0051063
R67855 VSS.n20119 VSS.n20118 0.0051063
R67856 VSS.n20086 VSS.n20085 0.0051063
R67857 VSS.n1069 VSS.n1068 0.0051063
R67858 VSS.n6792 VSS.n6791 0.0051063
R67859 VSS.n6879 VSS.n6878 0.0051063
R67860 VSS.n6506 VSS.n6505 0.0051063
R67861 VSS.n6471 VSS.n6470 0.0051063
R67862 VSS.n6438 VSS.n6437 0.0051063
R67863 VSS.n6421 VSS.n6420 0.0051063
R67864 VSS.n21371 VSS.n21370 0.0051063
R67865 VSS.n21338 VSS.n21337 0.0051063
R67866 VSS.n7626 VSS.n7625 0.0051063
R67867 VSS.n7659 VSS.n7658 0.0051063
R67868 VSS.n7714 VSS.n7713 0.0051063
R67869 VSS.n7747 VSS.n7746 0.0051063
R67870 VSS.n7825 VSS.n7824 0.0051063
R67871 VSS.n7792 VSS.n7791 0.0051063
R67872 VSS.n11687 VSS.n11686 0.0051063
R67873 VSS.n11656 VSS.n11655 0.0051063
R67874 VSS.n6130 VSS.n6129 0.0051063
R67875 VSS.n6100 VSS.n6099 0.0051063
R67876 VSS.n6049 VSS.n6048 0.0051063
R67877 VSS.n6019 VSS.n6018 0.0051063
R67878 VSS.n5968 VSS.n5967 0.0051063
R67879 VSS.n5938 VSS.n5937 0.0051063
R67880 VSS.n644 VSS.n643 0.0051063
R67881 VSS.n614 VSS.n613 0.0051063
R67882 VSS.n10602 VSS.n10601 0.0051063
R67883 VSS.n10572 VSS.n10571 0.0051063
R67884 VSS.n3217 VSS.n3215 0.00507746
R67885 VSS.n3222 VSS.n3220 0.00507746
R67886 VSS.n4974 VSS.n4943 0.00506429
R67887 VSS.n5003 VSS.n5002 0.00506429
R67888 VSS.n5033 VSS.n5032 0.00506429
R67889 VSS.n5079 VSS.n5078 0.00506429
R67890 VSS.n5923 VSS.n5922 0.00506429
R67891 VSS.n7392 VSS.n7391 0.00506429
R67892 VSS.n4622 VSS.n4621 0.00506429
R67893 VSS.n4576 VSS.n4575 0.00506429
R67894 VSS.n15440 VSS.n15439 0.00504436
R67895 VSS.n14567 VSS.n14566 0.00504436
R67896 VSS.n14828 VSS.n14827 0.00504436
R67897 VSS.n16880 VSS.n16879 0.00504436
R67898 VSS.n16691 VSS.n16690 0.00504436
R67899 VSS.n16440 VSS.n16439 0.00504436
R67900 VSS.n19761 VSS.n19760 0.00504436
R67901 VSS.n19851 VSS.n19850 0.00504436
R67902 VSS.n20036 VSS.n20035 0.00504436
R67903 VSS.n2093 VSS.n2092 0.00504436
R67904 VSS.n849 VSS.n848 0.00504436
R67905 VSS.n1742 VSS.n1741 0.00504436
R67906 VSS.n56 VSS.n54 0.00502514
R67907 VSS.n41 VSS.n40 0.00502514
R67908 VSS.n206 VSS.n205 0.00502514
R67909 VSS.n222 VSS.n219 0.00502514
R67910 VSS.n332 VSS.n331 0.00502514
R67911 VSS.n337 VSS.n333 0.00502514
R67912 VSS.n19409 VSS.n19408 0.005
R67913 VSS.n18257 VSS.n18255 0.005
R67914 VSS.n16612 VSS.n16610 0.005
R67915 VSS.n16517 VSS.n16516 0.005
R67916 VSS.n5199 VSS.n5198 0.005
R67917 VSS.n5250 VSS.n5249 0.005
R67918 VSS.n5284 VSS.n5283 0.005
R67919 VSS.n4969 VSS.n4968 0.005
R67920 VSS.n7076 VSS.n7075 0.005
R67921 VSS.n7541 VSS.n7540 0.005
R67922 VSS.n4456 VSS.n4455 0.005
R67923 VSS.n4405 VSS.n4404 0.005
R67924 VSS.n4370 VSS.n4369 0.005
R67925 VSS.n15697 VSS.n15696 0.005
R67926 VSS.n3774 VSS.n3773 0.00494444
R67927 VSS.n3773 VSS.n3772 0.00494444
R67928 VSS.n3772 VSS.n3771 0.00494444
R67929 VSS.n3771 VSS.n3770 0.00494444
R67930 VSS.n3770 VSS.n3769 0.00494444
R67931 VSS.n3769 VSS.n3768 0.00494444
R67932 VSS.n3768 VSS.n3767 0.00494444
R67933 VSS.n3767 VSS.n3766 0.00494444
R67934 VSS.n3766 VSS.n3765 0.00494444
R67935 VSS.n3765 VSS.n3764 0.00494444
R67936 VSS.n3764 VSS.n3763 0.00494444
R67937 VSS.n3763 VSS.n3762 0.00494444
R67938 VSS.n3762 VSS.n3761 0.00494444
R67939 VSS.n3761 VSS.n3760 0.00494444
R67940 VSS.n3760 VSS.n3759 0.00494444
R67941 VSS.n3759 VSS.n3758 0.00494444
R67942 VSS.n3758 VSS.n3757 0.00494444
R67943 VSS.n3757 VSS.n3756 0.00494444
R67944 VSS.n3756 VSS.n3755 0.00494444
R67945 VSS.n3755 VSS.n3754 0.00494444
R67946 VSS.n3754 VSS.n3753 0.00494444
R67947 VSS.n3753 VSS.n3752 0.00494444
R67948 VSS.n3752 VSS.n3751 0.00494444
R67949 VSS.n3751 VSS.n3750 0.00494444
R67950 VSS.n3750 VSS.n3749 0.00494444
R67951 VSS.n3749 VSS.n3748 0.00494444
R67952 VSS.n3748 VSS.n3747 0.00494444
R67953 VSS.n3747 VSS.n3746 0.00494444
R67954 VSS.n3746 VSS.n3745 0.00494444
R67955 VSS.n3745 VSS.n3744 0.00494444
R67956 VSS.n3744 VSS.n3743 0.00494444
R67957 VSS.n3743 VSS.n3742 0.00494444
R67958 VSS.n3742 VSS.n3741 0.00494444
R67959 VSS.n3741 VSS.n3740 0.00494444
R67960 VSS.n3740 VSS.n3739 0.00494444
R67961 VSS.n3739 VSS.n3738 0.00494444
R67962 VSS.n3738 VSS.n3737 0.00494444
R67963 VSS.n3737 VSS.n3736 0.00494444
R67964 VSS.n3736 VSS.n3735 0.00494444
R67965 VSS.n3735 VSS.n3734 0.00494444
R67966 VSS.n3734 VSS.n3733 0.00494444
R67967 VSS.n3733 VSS.n3732 0.00494444
R67968 VSS.n3732 VSS.n3731 0.00494444
R67969 VSS.n3731 VSS.n3730 0.00494444
R67970 VSS.n3730 VSS.n3729 0.00494444
R67971 VSS.n3729 VSS.n3728 0.00494444
R67972 VSS.n3728 VSS.n3727 0.00494444
R67973 VSS.n3727 VSS.n3726 0.00494444
R67974 VSS.n3726 VSS.n3725 0.00494444
R67975 VSS.n3725 VSS.n3724 0.00494444
R67976 VSS.n3724 VSS.n3723 0.00494444
R67977 VSS.n3723 VSS.n3722 0.00494444
R67978 VSS.n3722 VSS.n3721 0.00494444
R67979 VSS.n3721 VSS.n3720 0.00494444
R67980 VSS.n3720 VSS.n3719 0.00494444
R67981 VSS.n3719 VSS.n3718 0.00494444
R67982 VSS.n3718 VSS.n3717 0.00494444
R67983 VSS.n3717 VSS.n3716 0.00494444
R67984 VSS.n3716 VSS.n3715 0.00494444
R67985 VSS.n3715 VSS.n3714 0.00494444
R67986 VSS.n3714 VSS.n3713 0.00494444
R67987 VSS.n3713 VSS.n3712 0.00494444
R67988 VSS.n3712 VSS.n3711 0.00494444
R67989 VSS.n3711 VSS.n3710 0.00494444
R67990 VSS.n3710 VSS.n3709 0.00494444
R67991 VSS.n3709 VSS.n3708 0.00494444
R67992 VSS.n3708 VSS.n3707 0.00494444
R67993 VSS.n3707 VSS.n3706 0.00494444
R67994 VSS.n3706 VSS.n3705 0.00494444
R67995 VSS.n3705 VSS.n3704 0.00494444
R67996 VSS.n3704 VSS.n3703 0.00494444
R67997 VSS.n3703 VSS.n3702 0.00494444
R67998 VSS.n3702 VSS.n3701 0.00494444
R67999 VSS.n3701 VSS.n3700 0.00494444
R68000 VSS.n3700 VSS.n3699 0.00494444
R68001 VSS.n3699 VSS.n3698 0.00494444
R68002 VSS.n3698 VSS.n3697 0.00494444
R68003 VSS.n3697 VSS.n3696 0.00494444
R68004 VSS.n3696 VSS.n3695 0.00494444
R68005 VSS.n3695 VSS.n3694 0.00494444
R68006 VSS.n3694 VSS.n3693 0.00494444
R68007 VSS.n3693 VSS.n3692 0.00494444
R68008 VSS.n3692 VSS.n3691 0.00494444
R68009 VSS.n3691 VSS.n3690 0.00494444
R68010 VSS.n3690 VSS.n3689 0.00494444
R68011 VSS.n3689 VSS.n3688 0.00494444
R68012 VSS.n3688 VSS.n3687 0.00494444
R68013 VSS.n3687 VSS.n3686 0.00494444
R68014 VSS.n3686 VSS.n3685 0.00494444
R68015 VSS.n3685 VSS.n3684 0.00494444
R68016 VSS.n3684 VSS.n3683 0.00494444
R68017 VSS.n3683 VSS.n3682 0.00494444
R68018 VSS.n3682 VSS.n3681 0.00494444
R68019 VSS.n3681 VSS.n3680 0.00494444
R68020 VSS.n3680 VSS.n3679 0.00494444
R68021 VSS.n3679 VSS.n3678 0.00494444
R68022 VSS.n3678 VSS.n3677 0.00494444
R68023 VSS.n3210 VSS.n3209 0.00494444
R68024 VSS.n3209 VSS.n3208 0.00494444
R68025 VSS.n18715 VSS.n18714 0.00493662
R68026 VSS.n18410 VSS.n18409 0.00493662
R68027 VSS.n18152 VSS.n18151 0.00493662
R68028 VSS.n17123 VSS.n17122 0.00493662
R68029 VSS.n14860 VSS.n14859 0.00493662
R68030 VSS.n14874 VSS.n14873 0.00493662
R68031 VSS.n19197 VSS.n19196 0.00493662
R68032 VSS.n19612 VSS.n19611 0.00493662
R68033 VSS.n19704 VSS.n19703 0.00493662
R68034 VSS.n19872 VSS.n19871 0.00493662
R68035 VSS.n19931 VSS.n19930 0.00493662
R68036 VSS.n19945 VSS.n19944 0.00493662
R68037 VSS.n3082 VSS.n3081 0.00493571
R68038 VSS.n5198 VSS.n5197 0.00493571
R68039 VSS.n5249 VSS.n5248 0.00493571
R68040 VSS.n5283 VSS.n5282 0.00493571
R68041 VSS.n4970 VSS.n4969 0.00493571
R68042 VSS.n7350 VSS.n7349 0.00493571
R68043 VSS.n7296 VSS.n7295 0.00493571
R68044 VSS.n7077 VSS.n7076 0.00493571
R68045 VSS.n7541 VSS.n7521 0.00493571
R68046 VSS.n4457 VSS.n4456 0.00493571
R68047 VSS.n4406 VSS.n4405 0.00493571
R68048 VSS.n4371 VSS.n4370 0.00493571
R68049 VSS.n4345 VSS.n4344 0.00493571
R68050 VSS.n17737 VSS.n17736 0.00493571
R68051 VSS.n4004 VSS.n4003 0.00492913
R68052 VSS.n4043 VSS.n4042 0.00492913
R68053 VSS.n17445 VSS.n17444 0.00492913
R68054 VSS.n17314 VSS.n17313 0.00492913
R68055 VSS.n9549 VSS.n9548 0.00492913
R68056 VSS.n9050 VSS.n9049 0.00492913
R68057 VSS.n13029 VSS.n13028 0.00492913
R68058 VSS.n13072 VSS.n13071 0.00492913
R68059 VSS.n12982 VSS.n12981 0.00492913
R68060 VSS.n12764 VSS.n12763 0.00492913
R68061 VSS.n12602 VSS.n12593 0.00492913
R68062 VSS.n12563 VSS.n12562 0.00492913
R68063 VSS.n12272 VSS.n12271 0.00492913
R68064 VSS.n12248 VSS.n12247 0.00492913
R68065 VSS.n11927 VSS.n11926 0.00492913
R68066 VSS.n11902 VSS.n11901 0.00492913
R68067 VSS.n11843 VSS.n11842 0.00492913
R68068 VSS.n11819 VSS.n11818 0.00492913
R68069 VSS.n18875 VSS.n18874 0.00492913
R68070 VSS.n18914 VSS.n18913 0.00492913
R68071 VSS.n2196 VSS.n2195 0.00492913
R68072 VSS.n14406 VSS.n14405 0.00492913
R68073 VSS.n9666 VSS.n9665 0.00492913
R68074 VSS.n9193 VSS.n9192 0.00492913
R68075 VSS.n21802 VSS.n21801 0.00492913
R68076 VSS.n21845 VSS.n21844 0.00492913
R68077 VSS.n20602 VSS.n20601 0.00492913
R68078 VSS.n6956 VSS.n6955 0.00492913
R68079 VSS.n6683 VSS.n6682 0.00492913
R68080 VSS.n19087 VSS.n19086 0.00492913
R68081 VSS.n19130 VSS.n19129 0.00492913
R68082 VSS.n20164 VSS.n20163 0.00492913
R68083 VSS.n6854 VSS.n6853 0.00492913
R68084 VSS.n6533 VSS.n6532 0.00492913
R68085 VSS.n21573 VSS.n21572 0.00492913
R68086 VSS.n21616 VSS.n21615 0.00492913
R68087 VSS.n21399 VSS.n21398 0.00492913
R68088 VSS.n7598 VSS.n7597 0.00492913
R68089 VSS.n7686 VSS.n7685 0.00492913
R68090 VSS.n7774 VSS.n7773 0.00492913
R68091 VSS.n3806 VSS.n3805 0.00492913
R68092 VSS.n3845 VSS.n3844 0.00492913
R68093 VSS.n11724 VSS.n11723 0.00492913
R68094 VSS.n11187 VSS.n11186 0.00492913
R68095 VSS.n6075 VSS.n6074 0.00492913
R68096 VSS.n5994 VSS.n5993 0.00492913
R68097 VSS.n3284 VSS.n3283 0.00492913
R68098 VSS.n2660 VSS.n2659 0.00492913
R68099 VSS.n678 VSS.n677 0.00492913
R68100 VSS.n467 VSS.n466 0.00492913
R68101 VSS.n10536 VSS.n10527 0.00492913
R68102 VSS.n10507 VSS.n10506 0.00492913
R68103 VSS.n10221 VSS.n10220 0.00492913
R68104 VSS.n10197 VSS.n10196 0.00492913
R68105 VSS.n9928 VSS.n9927 0.00492913
R68106 VSS.n9902 VSS.n9901 0.00492913
R68107 VSS.n9002 VSS.n9001 0.00492913
R68108 VSS.n8929 VSS.n8928 0.00492913
R68109 VSS.n10305 VSS.n10300 0.00492308
R68110 VSS.n10423 VSS.n10418 0.00492308
R68111 VSS.n10138 VSS.n10133 0.00492308
R68112 VSS.n10046 VSS.n10041 0.00492308
R68113 VSS.n10039 VSS.n10038 0.00492308
R68114 VSS.n12359 VSS.n12354 0.00492308
R68115 VSS.n12477 VSS.n12472 0.00492308
R68116 VSS.n12189 VSS.n12184 0.00492308
R68117 VSS.n12097 VSS.n12092 0.00492308
R68118 VSS.n12090 VSS.n12089 0.00492308
R68119 VSS.n17207 VSS.n17206 0.00489325
R68120 VSS.n17193 VSS.n17192 0.00489325
R68121 VSS.n17187 VSS.n17186 0.00489325
R68122 VSS.n3195 VSS.n3194 0.0048662
R68123 VSS.n14179 VSS.n14178 0.00482175
R68124 VSS.n14178 VSS.n14177 0.00482175
R68125 VSS.n14140 VSS.n14139 0.00482175
R68126 VSS.n15290 VSS.n15288 0.00480851
R68127 VSS.n15297 VSS.n15293 0.00480851
R68128 VSS.n1607 VSS.n1602 0.00480851
R68129 VSS.n15493 VSS.n15492 0.00480851
R68130 VSS.n1795 VSS.n1794 0.00480851
R68131 VSS.n2572 VSS.n2571 0.00480714
R68132 VSS.n4975 VSS.n4974 0.00480714
R68133 VSS.n5005 VSS.n5003 0.00480714
R68134 VSS.n5035 VSS.n5033 0.00480714
R68135 VSS.n5081 VSS.n5079 0.00480714
R68136 VSS.n7419 VSS.n5923 0.00480714
R68137 VSS.n7391 VSS.n7390 0.00480714
R68138 VSS.n7358 VSS.n7357 0.00480714
R68139 VSS.n7304 VSS.n7303 0.00480714
R68140 VSS.n4621 VSS.n4620 0.00480714
R68141 VSS.n4575 VSS.n4574 0.00480714
R68142 VSS.n4338 VSS.n4337 0.00480714
R68143 VSS.n17730 VSS.n17729 0.00480714
R68144 VSS.n3658 VSS.n3657 0.00479577
R68145 VSS.n18430 VSS.n18427 0.004775
R68146 VSS.n17100 VSS.n17099 0.004775
R68147 VSS.n17061 VSS.n17060 0.004775
R68148 VSS.n16962 VSS.n16961 0.004775
R68149 VSS.n14927 VSS.n14926 0.004775
R68150 VSS.n171 VSS.n170 0.00477374
R68151 VSS.n167 VSS.n166 0.00477374
R68152 VSS.n20362 VSS.n20361 0.00476
R68153 VSS.n20361 VSS.n20360 0.00476
R68154 VSS.n20360 VSS.n20359 0.00476
R68155 VSS.n20359 VSS.n20358 0.00476
R68156 VSS.n20329 VSS.n20328 0.00476
R68157 VSS.n20281 VSS.n20280 0.00476
R68158 VSS.n20280 VSS.n20279 0.00476
R68159 VSS.n20279 VSS.n20278 0.00476
R68160 VSS.n20278 VSS.n20277 0.00476
R68161 VSS.n20277 VSS.n20276 0.00476
R68162 VSS.n20276 VSS.n20275 0.00476
R68163 VSS.n20275 VSS.n20274 0.00476
R68164 VSS.n20274 VSS.n20273 0.00476
R68165 VSS.n20273 VSS.n20272 0.00476
R68166 VSS.n20272 VSS.n20271 0.00476
R68167 VSS.n20201 VSS.n20200 0.00476
R68168 VSS.n20200 VSS.n20199 0.00476
R68169 VSS.n20199 VSS.n20198 0.00476
R68170 VSS.n20191 VSS.n20190 0.00476
R68171 VSS.n20185 VSS.n20184 0.00476
R68172 VSS.n696 VSS.n695 0.00476
R68173 VSS.n20393 VSS.n20391 0.00476
R68174 VSS.n20391 VSS.n20389 0.00476
R68175 VSS.n20389 VSS.n20387 0.00476
R68176 VSS.n20387 VSS.n20385 0.00476
R68177 VSS.n20363 VSS.n20357 0.00476
R68178 VSS.n20357 VSS.n20356 0.00476
R68179 VSS.n20356 VSS.n20355 0.00476
R68180 VSS.n20355 VSS.n20354 0.00476
R68181 VSS.n20332 VSS.n20330 0.00476
R68182 VSS.n20330 VSS.n20327 0.00476
R68183 VSS.n20327 VSS.n20326 0.00476
R68184 VSS.n20326 VSS.n20324 0.00476
R68185 VSS.n20324 VSS.n20322 0.00476
R68186 VSS.n20322 VSS.n20320 0.00476
R68187 VSS.n20320 VSS.n20318 0.00476
R68188 VSS.n20318 VSS.n20316 0.00476
R68189 VSS.n20316 VSS.n20314 0.00476
R68190 VSS.n20314 VSS.n20312 0.00476
R68191 VSS.n20312 VSS.n20310 0.00476
R68192 VSS.n20310 VSS.n20308 0.00476
R68193 VSS.n20286 VSS.n20284 0.00476
R68194 VSS.n20284 VSS.n20282 0.00476
R68195 VSS.n20282 VSS.n20270 0.00476
R68196 VSS.n20270 VSS.n20269 0.00476
R68197 VSS.n20269 VSS.n20268 0.00476
R68198 VSS.n20268 VSS.n20267 0.00476
R68199 VSS.n20267 VSS.n20266 0.00476
R68200 VSS.n20266 VSS.n20265 0.00476
R68201 VSS.n20265 VSS.n20264 0.00476
R68202 VSS.n20264 VSS.n20263 0.00476
R68203 VSS.n20263 VSS.n20262 0.00476
R68204 VSS.n20262 VSS.n20261 0.00476
R68205 VSS.n20202 VSS.n20197 0.00476
R68206 VSS.n20197 VSS.n20196 0.00476
R68207 VSS.n20196 VSS.n20195 0.00476
R68208 VSS.n20195 VSS.n20194 0.00476
R68209 VSS.n20194 VSS.n20192 0.00476
R68210 VSS.n20192 VSS.n20189 0.00476
R68211 VSS.n20189 VSS.n20188 0.00476
R68212 VSS.n20188 VSS.n20186 0.00476
R68213 VSS.n20186 VSS.n20183 0.00476
R68214 VSS.n20183 VSS.n20182 0.00476
R68215 VSS.n20182 VSS.n20180 0.00476
R68216 VSS.n20180 VSS.n20178 0.00476
R68217 VSS.n717 VSS.n715 0.00476
R68218 VSS.n715 VSS.n713 0.00476
R68219 VSS.n713 VSS.n711 0.00476
R68220 VSS.n711 VSS.n709 0.00476
R68221 VSS.n709 VSS.n707 0.00476
R68222 VSS.n707 VSS.n705 0.00476
R68223 VSS.n705 VSS.n703 0.00476
R68224 VSS.n703 VSS.n701 0.00476
R68225 VSS.n701 VSS.n699 0.00476
R68226 VSS.n699 VSS.n697 0.00476
R68227 VSS.n697 VSS.n694 0.00476
R68228 VSS.n694 VSS.n693 0.00476
R68229 VSS.n20577 VSS.n20576 0.00476
R68230 VSS.n20576 VSS.n20575 0.00476
R68231 VSS.n20575 VSS.n20574 0.00476
R68232 VSS.n20574 VSS.n20573 0.00476
R68233 VSS.n20555 VSS.n20554 0.00476
R68234 VSS.n20554 VSS.n20553 0.00476
R68235 VSS.n20553 VSS.n20552 0.00476
R68236 VSS.n10698 VSS.n10697 0.00476
R68237 VSS.n10756 VSS.n10755 0.00476
R68238 VSS.n10786 VSS.n10785 0.00476
R68239 VSS.n10785 VSS.n10784 0.00476
R68240 VSS.n10784 VSS.n10783 0.00476
R68241 VSS.n10799 VSS.n10798 0.00476
R68242 VSS.n10798 VSS.n10797 0.00476
R68243 VSS.n10797 VSS.n10796 0.00476
R68244 VSS.n10796 VSS.n10795 0.00476
R68245 VSS.n10895 VSS.n10894 0.00476
R68246 VSS.n10894 VSS.n10893 0.00476
R68247 VSS.n10893 VSS.n10892 0.00476
R68248 VSS.n10892 VSS.n10891 0.00476
R68249 VSS.n10891 VSS.n10890 0.00476
R68250 VSS.n10890 VSS.n10889 0.00476
R68251 VSS.n10889 VSS.n10888 0.00476
R68252 VSS.n10888 VSS.n10887 0.00476
R68253 VSS.n10909 VSS.n10908 0.00476
R68254 VSS.n10908 VSS.n10907 0.00476
R68255 VSS.n10907 VSS.n10906 0.00476
R68256 VSS.n10956 VSS.n10955 0.00476
R68257 VSS.n10962 VSS.n10961 0.00476
R68258 VSS.n10967 VSS.n10966 0.00476
R68259 VSS.n10966 VSS.n10965 0.00476
R68260 VSS.n10975 VSS.n10974 0.00476
R68261 VSS.n10974 VSS.n10973 0.00476
R68262 VSS.n10973 VSS.n10972 0.00476
R68263 VSS.n10972 VSS.n10971 0.00476
R68264 VSS.n11078 VSS.n6348 0.00476
R68265 VSS.n11078 VSS.n11077 0.00476
R68266 VSS.n9770 VSS.n9769 0.00476
R68267 VSS.n9714 VSS.n9713 0.00476
R68268 VSS.n10781 VSS.n10780 0.00476
R68269 VSS.n10780 VSS.n10779 0.00476
R68270 VSS.n10779 VSS.n10778 0.00476
R68271 VSS.n10778 VSS.n10777 0.00476
R68272 VSS.n10777 VSS.n10776 0.00476
R68273 VSS.n10776 VSS.n10775 0.00476
R68274 VSS.n10775 VSS.n10774 0.00476
R68275 VSS.n10774 VSS.n10773 0.00476
R68276 VSS.n8592 VSS.n8591 0.00476
R68277 VSS.n8591 VSS.n8590 0.00476
R68278 VSS.n8590 VSS.n8589 0.00476
R68279 VSS.n8589 VSS.n8588 0.00476
R68280 VSS.n8588 VSS.n8587 0.00476
R68281 VSS.n8587 VSS.n8586 0.00476
R68282 VSS.n8586 VSS.n8585 0.00476
R68283 VSS.n8585 VSS.n8584 0.00476
R68284 VSS.n10884 VSS.n10883 0.00476
R68285 VSS.n10883 VSS.n10882 0.00476
R68286 VSS.n10882 VSS.n10881 0.00476
R68287 VSS.n8058 VSS.n8057 0.00476
R68288 VSS.n8057 VSS.n8056 0.00476
R68289 VSS.n8056 VSS.n8055 0.00476
R68290 VSS.n8055 VSS.n8054 0.00476
R68291 VSS.n8054 VSS.n8053 0.00476
R68292 VSS.n8053 VSS.n8052 0.00476
R68293 VSS.n8052 VSS.n8051 0.00476
R68294 VSS.n8051 VSS.n8050 0.00476
R68295 VSS.n8040 VSS.n8039 0.00476
R68296 VSS.n7997 VSS.n7996 0.00476
R68297 VSS.n7957 VSS.n7956 0.00476
R68298 VSS.n7956 VSS.n7955 0.00476
R68299 VSS.n7955 VSS.n7954 0.00476
R68300 VSS.n7954 VSS.n7953 0.00476
R68301 VSS.n9011 VSS.n9010 0.00476
R68302 VSS.n9325 VSS.n9324 0.00476
R68303 VSS.n9324 VSS.n9323 0.00476
R68304 VSS.n10770 VSS.n10769 0.00476
R68305 VSS.n10769 VSS.n10768 0.00476
R68306 VSS.n10768 VSS.n10767 0.00476
R68307 VSS.n10767 VSS.n10766 0.00476
R68308 VSS.n10766 VSS.n10765 0.00476
R68309 VSS.n10765 VSS.n10764 0.00476
R68310 VSS.n10764 VSS.n10763 0.00476
R68311 VSS.n10763 VSS.n10762 0.00476
R68312 VSS.n8255 VSS.n8254 0.00476
R68313 VSS.n8254 VSS.n8253 0.00476
R68314 VSS.n8253 VSS.n8252 0.00476
R68315 VSS.n8252 VSS.n8251 0.00476
R68316 VSS.n8251 VSS.n8250 0.00476
R68317 VSS.n8250 VSS.n8249 0.00476
R68318 VSS.n8241 VSS.n8240 0.00476
R68319 VSS.n10879 VSS.n10878 0.00476
R68320 VSS.n10878 VSS.n10877 0.00476
R68321 VSS.n10877 VSS.n10876 0.00476
R68322 VSS.n6744 VSS.n6743 0.00476
R68323 VSS.n6743 VSS.n6742 0.00476
R68324 VSS.n6742 VSS.n6741 0.00476
R68325 VSS.n6734 VSS.n6733 0.00476
R68326 VSS.n6733 VSS.n6732 0.00476
R68327 VSS.n7904 VSS.n7903 0.00476
R68328 VSS.n8822 VSS.n8820 0.00476
R68329 VSS.n8824 VSS.n8822 0.00476
R68330 VSS.n8826 VSS.n8824 0.00476
R68331 VSS.n8828 VSS.n8826 0.00476
R68332 VSS.n9009 VSS.n9008 0.00476
R68333 VSS.n9012 VSS.n9009 0.00476
R68334 VSS.n9014 VSS.n9012 0.00476
R68335 VSS.n9380 VSS.n9378 0.00476
R68336 VSS.n9378 VSS.n9376 0.00476
R68337 VSS.n9376 VSS.n9374 0.00476
R68338 VSS.n9374 VSS.n9372 0.00476
R68339 VSS.n9372 VSS.n9370 0.00476
R68340 VSS.n9370 VSS.n9368 0.00476
R68341 VSS.n9368 VSS.n9366 0.00476
R68342 VSS.n9366 VSS.n9364 0.00476
R68343 VSS.n9364 VSS.n9362 0.00476
R68344 VSS.n9362 VSS.n9360 0.00476
R68345 VSS.n9360 VSS.n9358 0.00476
R68346 VSS.n9358 VSS.n9356 0.00476
R68347 VSS.n9326 VSS.n9322 0.00476
R68348 VSS.n9322 VSS.n9321 0.00476
R68349 VSS.n8452 VSS.n8451 0.00476
R68350 VSS.n8451 VSS.n8450 0.00476
R68351 VSS.n8450 VSS.n8449 0.00476
R68352 VSS.n8449 VSS.n8448 0.00476
R68353 VSS.n8448 VSS.n8447 0.00476
R68354 VSS.n8447 VSS.n8446 0.00476
R68355 VSS.n8446 VSS.n8445 0.00476
R68356 VSS.n8445 VSS.n8444 0.00476
R68357 VSS.n8256 VSS.n8248 0.00476
R68358 VSS.n8248 VSS.n8247 0.00476
R68359 VSS.n8247 VSS.n8246 0.00476
R68360 VSS.n8246 VSS.n8245 0.00476
R68361 VSS.n8245 VSS.n8244 0.00476
R68362 VSS.n8244 VSS.n8243 0.00476
R68363 VSS.n8243 VSS.n8242 0.00476
R68364 VSS.n8242 VSS.n8239 0.00476
R68365 VSS.n6783 VSS.n6782 0.00476
R68366 VSS.n6782 VSS.n6781 0.00476
R68367 VSS.n6781 VSS.n6780 0.00476
R68368 VSS.n6745 VSS.n6740 0.00476
R68369 VSS.n6740 VSS.n6739 0.00476
R68370 VSS.n6739 VSS.n6738 0.00476
R68371 VSS.n6738 VSS.n6737 0.00476
R68372 VSS.n6737 VSS.n6735 0.00476
R68373 VSS.n6735 VSS.n6731 0.00476
R68374 VSS.n6731 VSS.n6730 0.00476
R68375 VSS.n6730 VSS.n6729 0.00476
R68376 VSS.n6729 VSS.n6727 0.00476
R68377 VSS.n6727 VSS.n6725 0.00476
R68378 VSS.n6725 VSS.n6723 0.00476
R68379 VSS.n6723 VSS.n6721 0.00476
R68380 VSS.n7905 VSS.n7902 0.00476
R68381 VSS.n7902 VSS.n7901 0.00476
R68382 VSS.n7901 VSS.n7899 0.00476
R68383 VSS.n7865 VSS.n7863 0.00476
R68384 VSS.n7863 VSS.n7862 0.00476
R68385 VSS.n7862 VSS.n7861 0.00476
R68386 VSS.n9435 VSS.n9433 0.00476
R68387 VSS.n9437 VSS.n9435 0.00476
R68388 VSS.n9439 VSS.n9437 0.00476
R68389 VSS.n9441 VSS.n9439 0.00476
R68390 VSS.n9472 VSS.n9470 0.00476
R68391 VSS.n9474 VSS.n9472 0.00476
R68392 VSS.n9476 VSS.n9474 0.00476
R68393 VSS.n9771 VSS.n9768 0.00476
R68394 VSS.n9768 VSS.n9767 0.00476
R68395 VSS.n9767 VSS.n9765 0.00476
R68396 VSS.n9765 VSS.n9763 0.00476
R68397 VSS.n9763 VSS.n9761 0.00476
R68398 VSS.n9761 VSS.n9759 0.00476
R68399 VSS.n9759 VSS.n9757 0.00476
R68400 VSS.n9757 VSS.n9755 0.00476
R68401 VSS.n9755 VSS.n9753 0.00476
R68402 VSS.n9753 VSS.n9751 0.00476
R68403 VSS.n9751 VSS.n9749 0.00476
R68404 VSS.n9749 VSS.n9747 0.00476
R68405 VSS.n9717 VSS.n9715 0.00476
R68406 VSS.n9715 VSS.n9712 0.00476
R68407 VSS.n8784 VSS.n8783 0.00476
R68408 VSS.n8783 VSS.n8782 0.00476
R68409 VSS.n8782 VSS.n8781 0.00476
R68410 VSS.n8781 VSS.n8780 0.00476
R68411 VSS.n8780 VSS.n8779 0.00476
R68412 VSS.n8779 VSS.n8778 0.00476
R68413 VSS.n8778 VSS.n8777 0.00476
R68414 VSS.n8777 VSS.n8776 0.00476
R68415 VSS.n8593 VSS.n8583 0.00476
R68416 VSS.n8583 VSS.n8582 0.00476
R68417 VSS.n8582 VSS.n8581 0.00476
R68418 VSS.n8581 VSS.n8580 0.00476
R68419 VSS.n8580 VSS.n8579 0.00476
R68420 VSS.n8579 VSS.n8578 0.00476
R68421 VSS.n8578 VSS.n8577 0.00476
R68422 VSS.n8577 VSS.n8576 0.00476
R68423 VSS.n8099 VSS.n8098 0.00476
R68424 VSS.n8098 VSS.n8097 0.00476
R68425 VSS.n8097 VSS.n8096 0.00476
R68426 VSS.n8061 VSS.n8059 0.00476
R68427 VSS.n8059 VSS.n8049 0.00476
R68428 VSS.n8049 VSS.n8048 0.00476
R68429 VSS.n8048 VSS.n8047 0.00476
R68430 VSS.n8047 VSS.n8046 0.00476
R68431 VSS.n8046 VSS.n8045 0.00476
R68432 VSS.n8045 VSS.n8044 0.00476
R68433 VSS.n8044 VSS.n8043 0.00476
R68434 VSS.n8043 VSS.n8042 0.00476
R68435 VSS.n8042 VSS.n8041 0.00476
R68436 VSS.n8041 VSS.n8038 0.00476
R68437 VSS.n8038 VSS.n8037 0.00476
R68438 VSS.n7998 VSS.n7995 0.00476
R68439 VSS.n7995 VSS.n7994 0.00476
R68440 VSS.n7994 VSS.n7992 0.00476
R68441 VSS.n7958 VSS.n7907 0.00476
R68442 VSS.n7942 VSS.n7907 0.00476
R68443 VSS.n7943 VSS.n7942 0.00476
R68444 VSS.n7944 VSS.n7943 0.00476
R68445 VSS.n9810 VSS.n9808 0.00476
R68446 VSS.n9812 VSS.n9810 0.00476
R68447 VSS.n9814 VSS.n9812 0.00476
R68448 VSS.n9816 VSS.n9814 0.00476
R68449 VSS.n10645 VSS.n10643 0.00476
R68450 VSS.n10647 VSS.n10645 0.00476
R68451 VSS.n10653 VSS.n10647 0.00476
R68452 VSS.n10696 VSS.n10694 0.00476
R68453 VSS.n10699 VSS.n10696 0.00476
R68454 VSS.n10700 VSS.n10699 0.00476
R68455 VSS.n10702 VSS.n10700 0.00476
R68456 VSS.n10704 VSS.n10702 0.00476
R68457 VSS.n10706 VSS.n10704 0.00476
R68458 VSS.n10708 VSS.n10706 0.00476
R68459 VSS.n10710 VSS.n10708 0.00476
R68460 VSS.n10712 VSS.n10710 0.00476
R68461 VSS.n10714 VSS.n10712 0.00476
R68462 VSS.n10716 VSS.n10714 0.00476
R68463 VSS.n10718 VSS.n10716 0.00476
R68464 VSS.n10758 VSS.n10757 0.00476
R68465 VSS.n10760 VSS.n10758 0.00476
R68466 VSS.n10789 VSS.n10760 0.00476
R68467 VSS.n10792 VSS.n10791 0.00476
R68468 VSS.n10793 VSS.n10792 0.00476
R68469 VSS.n10794 VSS.n10793 0.00476
R68470 VSS.n10800 VSS.n10794 0.00476
R68471 VSS.n10801 VSS.n10800 0.00476
R68472 VSS.n10802 VSS.n10801 0.00476
R68473 VSS.n10803 VSS.n10802 0.00476
R68474 VSS.n10804 VSS.n10803 0.00476
R68475 VSS.n10897 VSS.n10896 0.00476
R68476 VSS.n10898 VSS.n10897 0.00476
R68477 VSS.n10899 VSS.n10898 0.00476
R68478 VSS.n10900 VSS.n10899 0.00476
R68479 VSS.n10901 VSS.n10900 0.00476
R68480 VSS.n10902 VSS.n10901 0.00476
R68481 VSS.n10903 VSS.n10902 0.00476
R68482 VSS.n10904 VSS.n10903 0.00476
R68483 VSS.n10911 VSS.n10910 0.00476
R68484 VSS.n10912 VSS.n10911 0.00476
R68485 VSS.n10913 VSS.n10912 0.00476
R68486 VSS.n10958 VSS.n10957 0.00476
R68487 VSS.n10960 VSS.n10958 0.00476
R68488 VSS.n10963 VSS.n10960 0.00476
R68489 VSS.n10964 VSS.n10963 0.00476
R68490 VSS.n10968 VSS.n10964 0.00476
R68491 VSS.n10969 VSS.n10968 0.00476
R68492 VSS.n10970 VSS.n10969 0.00476
R68493 VSS.n10976 VSS.n10970 0.00476
R68494 VSS.n10977 VSS.n10976 0.00476
R68495 VSS.n10978 VSS.n10977 0.00476
R68496 VSS.n10979 VSS.n10978 0.00476
R68497 VSS.n10980 VSS.n10979 0.00476
R68498 VSS.n11032 VSS.n11030 0.00476
R68499 VSS.n11034 VSS.n11032 0.00476
R68500 VSS.n11036 VSS.n11034 0.00476
R68501 VSS.n11072 VSS.n11071 0.00476
R68502 VSS.n11073 VSS.n11072 0.00476
R68503 VSS.n11074 VSS.n11073 0.00476
R68504 VSS.n2345 VSS.n2344 0.00475197
R68505 VSS.n17477 VSS.n17476 0.00475197
R68506 VSS.n11351 VSS.n11350 0.00475197
R68507 VSS.n13153 VSS.n13152 0.00475197
R68508 VSS.n12858 VSS.n12857 0.00475197
R68509 VSS.n12795 VSS.n12794 0.00475197
R68510 VSS.n12295 VSS.n12294 0.00475197
R68511 VSS.n11953 VSS.n11952 0.00475197
R68512 VSS.n11946 VSS.n11945 0.00475197
R68513 VSS.n11901 VSS.n11900 0.00475197
R68514 VSS.n11897 VSS.n11896 0.00475197
R68515 VSS.n2244 VSS.n2243 0.00475197
R68516 VSS.n2228 VSS.n2227 0.00475197
R68517 VSS.n15152 VSS.n15151 0.00475197
R68518 VSS.n2293 VSS.n2292 0.00475197
R68519 VSS.n20802 VSS.n20801 0.00475197
R68520 VSS.n17901 VSS.n17900 0.00475197
R68521 VSS.n2017 VSS.n2016 0.00475197
R68522 VSS.n21638 VSS.n21637 0.00475197
R68523 VSS.n21537 VSS.n21536 0.00475197
R68524 VSS.n21520 VSS.n21519 0.00475197
R68525 VSS.n21279 VSS.n21278 0.00475197
R68526 VSS.n7567 VSS.n7566 0.00475197
R68527 VSS.n3867 VSS.n3866 0.00475197
R68528 VSS.n4153 VSS.n4152 0.00475197
R68529 VSS.n4698 VSS.n4697 0.00475197
R68530 VSS.n11437 VSS.n11436 0.00475197
R68531 VSS.n11216 VSS.n11215 0.00475197
R68532 VSS.n555 VSS.n554 0.00475197
R68533 VSS.n496 VSS.n495 0.00475197
R68534 VSS.n10243 VSS.n10242 0.00475197
R68535 VSS.n9955 VSS.n9954 0.00475197
R68536 VSS.n9948 VSS.n9947 0.00475197
R68537 VSS.n9901 VSS.n9900 0.00475197
R68538 VSS.n9896 VSS.n9895 0.00475197
R68539 VSS.n7175 VSS.n7174 0.00474286
R68540 VSS.n7116 VSS.n7115 0.00474286
R68541 VSS.n18109 VSS.n2229 0.00473539
R68542 VSS.n2221 VSS.n2220 0.00473539
R68543 VSS.n2199 VSS.n2198 0.00473539
R68544 VSS.n2334 VSS.n2333 0.00473539
R68545 VSS.n13321 VSS.n13320 0.00473539
R68546 VSS.n13343 VSS.n13342 0.00473539
R68547 VSS.n17963 VSS.n17955 0.00473539
R68548 VSS.n17947 VSS.n17946 0.00473539
R68549 VSS.n13486 VSS.n13485 0.00473539
R68550 VSS.n18774 VSS.n18773 0.00472535
R68551 VSS.n18451 VSS.n18450 0.00472535
R68552 VSS.n18191 VSS.n18190 0.00472535
R68553 VSS.n18181 VSS.n18180 0.00472535
R68554 VSS.n16580 VSS.n16579 0.00472535
R68555 VSS.n14984 VSS.n14983 0.00472535
R68556 VSS.n14985 VSS.n14984 0.00472535
R68557 VSS.n15535 VSS.n15534 0.00472535
R68558 VSS.n8515 VSS.n8514 0.00472535
R68559 VSS.n19446 VSS.n19445 0.00472535
R68560 VSS.n19588 VSS.n19587 0.00472535
R68561 VSS.n19665 VSS.n19664 0.00472535
R68562 VSS.n19675 VSS.n19674 0.00472535
R68563 VSS.n788 VSS.n787 0.00472535
R68564 VSS.n820 VSS.n819 0.00472535
R68565 VSS.n821 VSS.n820 0.00472535
R68566 VSS.n1823 VSS.n1822 0.00472535
R68567 VSS.n8666 VSS.n8665 0.00472535
R68568 VSS.n3183 VSS.n3182 0.00467857
R68569 VSS.n2579 VSS.n2577 0.00467857
R68570 VSS.n4687 VSS.n4686 0.00467857
R68571 VSS.n4682 VSS.n4681 0.00467857
R68572 VSS.n17603 VSS.n2338 0.00467857
R68573 VSS.n17600 VSS.n17599 0.00467857
R68574 VSS.n20171 VSS.n20170 0.00467
R68575 VSS.n685 VSS.n684 0.00467
R68576 VSS.n20539 VSS.n20538 0.00467
R68577 VSS.n19692 VSS.n19691 0.00465899
R68578 VSS.n19718 VSS.n19717 0.00465899
R68579 VSS.n20370 VSS.n20369 0.00464
R68580 VSS.n9429 VSS.n9428 0.00464
R68581 VSS.n13248 VSS.n13247 0.00461744
R68582 VSS.n12996 VSS.n12995 0.00461744
R68583 VSS.n12897 VSS.n12896 0.00461744
R68584 VSS.n12884 VSS.n12883 0.00461744
R68585 VSS.n12830 VSS.n12829 0.00461744
R68586 VSS.n13215 VSS.n13214 0.00461744
R68587 VSS.n14401 VSS.n14400 0.00461744
R68588 VSS.n14422 VSS.n14421 0.00461744
R68589 VSS.n15075 VSS.n15074 0.00461744
R68590 VSS.n15108 VSS.n15107 0.00461744
R68591 VSS.n15178 VSS.n15177 0.00461744
R68592 VSS.n18988 VSS.n2165 0.00461744
R68593 VSS.n2210 VSS.n2209 0.00461744
R68594 VSS.n5714 VSS.n5639 0.00461744
R68595 VSS.n13365 VSS.n13364 0.00461744
R68596 VSS.n13416 VSS.n13415 0.00461744
R68597 VSS.n20687 VSS.n20686 0.00461744
R68598 VSS.n20738 VSS.n20737 0.00461744
R68599 VSS.n20830 VSS.n20829 0.00461744
R68600 VSS.n21734 VSS.n347 0.00461744
R68601 VSS.n13332 VSS.n13331 0.00461744
R68602 VSS.n21102 VSS.n21089 0.00461744
R68603 VSS.n13508 VSS.n13507 0.00461744
R68604 VSS.n20148 VSS.n20147 0.00461744
R68605 VSS.n2054 VSS.n2053 0.00461744
R68606 VSS.n2043 VSS.n2042 0.00461744
R68607 VSS.n884 VSS.n883 0.00461744
R68608 VSS.n17886 VSS.n17885 0.00461744
R68609 VSS.n13475 VSS.n13474 0.00461744
R68610 VSS.n592 VSS.n591 0.00461744
R68611 VSS.n579 VSS.n578 0.00461744
R68612 VSS.n529 VSS.n528 0.00461744
R68613 VSS.n21682 VSS.n21544 0.00461744
R68614 VSS.n2836 VSS.n2835 0.00461429
R68615 VSS.n18061 VSS.n18060 0.00461429
R68616 VSS.n14167 VSS.n14166 0.00459712
R68617 VSS.n16639 VSS.n16638 0.00459139
R68618 VSS.n759 VSS.n758 0.00459139
R68619 DVSS VSS.n7858 0.00458
R68620 VSS.n7861 DVSS 0.00458
R68621 VSS.n19055 VSS.n19054 0.00457827
R68622 VSS.n21770 VSS.n21769 0.00457827
R68623 VSS.n4011 VSS.n4010 0.0045748
R68624 VSS.n13036 VSS.n13035 0.0045748
R68625 VSS.n12527 VSS.n12526 0.0045748
R68626 VSS.n12306 VSS.n12305 0.0045748
R68627 VSS.n11954 VSS.n11953 0.0045748
R68628 VSS.n18882 VSS.n18881 0.0045748
R68629 VSS.n21809 VSS.n21808 0.0045748
R68630 VSS.n19094 VSS.n19093 0.0045748
R68631 VSS.n21580 VSS.n21579 0.0045748
R68632 VSS.n3813 VSS.n3812 0.0045748
R68633 VSS.n3258 VSS.n3257 0.0045748
R68634 VSS.n10472 VSS.n10471 0.0045748
R68635 VSS.n10254 VSS.n10253 0.0045748
R68636 VSS.n9956 VSS.n9955 0.0045748
R68637 VSS.n14236 VSS.n14235 0.00455714
R68638 VSS.n14235 VSS.n14234 0.00455714
R68639 VSS.n14234 VSS.n14233 0.00455714
R68640 VSS.n14233 VSS.n14232 0.00455714
R68641 VSS.n14232 VSS.n14231 0.00455714
R68642 VSS.n14211 VSS.n14210 0.00455714
R68643 VSS.n14212 VSS.n14211 0.00455714
R68644 VSS.n13940 VSS.n13939 0.00455714
R68645 VSS.n13939 VSS.n13938 0.00455714
R68646 VSS.n13938 VSS.n13937 0.00455714
R68647 VSS.n13937 VSS.n13936 0.00455714
R68648 VSS.n13936 VSS.n13935 0.00455714
R68649 VSS.n13935 VSS.n13934 0.00455714
R68650 VSS.n13934 VSS.n13933 0.00455714
R68651 VSS.n13933 VSS.n13932 0.00455714
R68652 VSS.n13932 VSS.n13931 0.00455714
R68653 VSS.n13931 VSS.n13930 0.00455714
R68654 VSS.n13930 VSS.n13929 0.00455714
R68655 VSS.n13929 VSS.n13928 0.00455714
R68656 VSS.n13928 VSS.n13927 0.00455714
R68657 VSS.n13927 VSS.n13926 0.00455714
R68658 VSS.n13926 VSS.n13925 0.00455714
R68659 VSS.n13925 VSS.n13924 0.00455714
R68660 VSS.n13924 VSS.n13923 0.00455714
R68661 VSS.n13923 VSS.n13922 0.00455714
R68662 VSS.n13922 VSS.n13921 0.00455714
R68663 VSS.n13921 VSS.n13920 0.00455714
R68664 VSS.n13920 VSS.n13919 0.00455714
R68665 VSS.n13919 VSS.n13918 0.00455714
R68666 VSS.n13918 VSS.n13917 0.00455714
R68667 VSS.n13917 VSS.n13916 0.00455714
R68668 VSS.n13916 VSS.n13915 0.00455714
R68669 VSS.n13915 VSS.n13914 0.00455714
R68670 VSS.n13914 VSS.n13913 0.00455714
R68671 VSS.n13913 VSS.n13912 0.00455714
R68672 VSS.n13912 VSS.n13911 0.00455714
R68673 VSS.n13911 VSS.n13910 0.00455714
R68674 VSS.n13910 VSS.n13909 0.00455714
R68675 VSS.n13909 VSS.n13908 0.00455714
R68676 VSS.n13908 VSS.n13907 0.00455714
R68677 VSS.n13907 VSS.n13906 0.00455714
R68678 VSS.n13906 VSS.n13905 0.00455714
R68679 VSS.n13905 VSS.n13904 0.00455714
R68680 VSS.n13904 VSS.n13903 0.00455714
R68681 VSS.n13903 VSS.n13902 0.00455714
R68682 VSS.n13902 VSS.n13901 0.00455714
R68683 VSS.n13901 VSS.n13900 0.00455714
R68684 VSS.n13900 VSS.n13899 0.00455714
R68685 VSS.n13899 VSS.n13898 0.00455714
R68686 VSS.n13898 VSS.n13897 0.00455714
R68687 VSS.n13897 VSS.n13896 0.00455714
R68688 VSS.n13896 VSS.n13895 0.00455714
R68689 VSS.n13895 VSS.n13894 0.00455714
R68690 VSS.n13894 VSS.n13893 0.00455714
R68691 VSS.n13893 VSS.n13892 0.00455714
R68692 VSS.n13892 VSS.n13891 0.00455714
R68693 VSS.n13891 VSS.n13890 0.00455714
R68694 VSS.n13890 VSS.n13889 0.00455714
R68695 VSS.n13889 VSS.n13888 0.00455714
R68696 VSS.n13888 VSS.n13887 0.00455714
R68697 VSS.n13887 VSS.n13886 0.00455714
R68698 VSS.n13886 VSS.n13885 0.00455714
R68699 VSS.n13885 VSS.n13884 0.00455714
R68700 VSS.n13884 VSS.n13883 0.00455714
R68701 VSS.n13883 VSS.n13882 0.00455714
R68702 VSS.n13882 VSS.n13881 0.00455714
R68703 VSS.n13881 VSS.n13880 0.00455714
R68704 VSS.n13880 VSS.n13879 0.00455714
R68705 VSS.n13879 VSS.n13878 0.00455714
R68706 VSS.n13878 VSS.n13877 0.00455714
R68707 VSS.n13877 VSS.n13876 0.00455714
R68708 VSS.n13876 VSS.n13875 0.00455714
R68709 VSS.n13875 VSS.n13874 0.00455714
R68710 VSS.n13874 VSS.n13873 0.00455714
R68711 VSS.n13873 VSS.n13872 0.00455714
R68712 VSS.n13872 VSS.n13871 0.00455714
R68713 VSS.n13871 VSS.n13870 0.00455714
R68714 VSS.n13870 VSS.n13869 0.00455714
R68715 VSS.n13869 VSS.n13868 0.00455714
R68716 VSS.n13868 VSS.n13867 0.00455714
R68717 VSS.n13867 VSS.n13866 0.00455714
R68718 VSS.n13866 VSS.n13865 0.00455714
R68719 VSS.n13865 VSS.n13864 0.00455714
R68720 VSS.n13864 VSS.n13863 0.00455714
R68721 VSS.n13863 VSS.n13862 0.00455714
R68722 VSS.n13862 VSS.n13861 0.00455714
R68723 VSS.n13861 VSS.n13860 0.00455714
R68724 VSS.n13860 VSS.n13859 0.00455714
R68725 VSS.n13859 VSS.n13858 0.00455714
R68726 VSS.n13858 VSS.n13857 0.00455714
R68727 VSS.n13857 VSS.n13856 0.00455714
R68728 VSS.n13856 VSS.n13855 0.00455714
R68729 VSS.n13855 VSS.n13854 0.00455714
R68730 VSS.n13854 VSS.n13853 0.00455714
R68731 VSS.n13853 VSS.n13852 0.00455714
R68732 VSS.n13663 VSS.n13662 0.00455714
R68733 VSS.n17606 VSS.n17605 0.00455714
R68734 VSS.n17607 VSS.n17606 0.00455714
R68735 VSS.n17608 VSS.n17607 0.00455714
R68736 VSS.n17609 VSS.n17608 0.00455714
R68737 VSS.n17610 VSS.n17609 0.00455714
R68738 VSS.n17611 VSS.n17610 0.00455714
R68739 VSS.n17612 VSS.n17611 0.00455714
R68740 VSS.n17613 VSS.n17612 0.00455714
R68741 VSS.n17614 VSS.n17613 0.00455714
R68742 VSS.n17615 VSS.n17614 0.00455714
R68743 VSS.n17616 VSS.n17615 0.00455714
R68744 VSS.n17617 VSS.n17616 0.00455714
R68745 VSS.n17618 VSS.n17617 0.00455714
R68746 VSS.n17619 VSS.n17618 0.00455714
R68747 VSS.n17620 VSS.n17619 0.00455714
R68748 VSS.n17621 VSS.n17620 0.00455714
R68749 VSS.n17622 VSS.n17621 0.00455714
R68750 VSS.n17623 VSS.n17622 0.00455714
R68751 VSS.n17624 VSS.n17623 0.00455714
R68752 VSS.n17625 VSS.n17624 0.00455714
R68753 VSS.n17626 VSS.n17625 0.00455714
R68754 VSS.n17627 VSS.n17626 0.00455714
R68755 VSS.n17628 VSS.n17627 0.00455714
R68756 VSS.n17629 VSS.n17628 0.00455714
R68757 VSS.n17630 VSS.n17629 0.00455714
R68758 VSS.n17631 VSS.n17630 0.00455714
R68759 VSS.n17632 VSS.n17631 0.00455714
R68760 VSS.n17633 VSS.n17632 0.00455714
R68761 VSS.n17634 VSS.n17633 0.00455714
R68762 VSS.n17635 VSS.n17634 0.00455714
R68763 VSS.n17636 VSS.n17635 0.00455714
R68764 VSS.n17637 VSS.n17636 0.00455714
R68765 VSS.n17638 VSS.n17637 0.00455714
R68766 VSS.n17639 VSS.n17638 0.00455714
R68767 VSS.n17640 VSS.n17639 0.00455714
R68768 VSS.n17641 VSS.n17640 0.00455714
R68769 VSS.n17642 VSS.n17641 0.00455714
R68770 VSS.n17643 VSS.n17642 0.00455714
R68771 VSS.n17644 VSS.n17643 0.00455714
R68772 VSS.n17645 VSS.n17644 0.00455714
R68773 VSS.n17646 VSS.n17645 0.00455714
R68774 VSS.n17647 VSS.n17646 0.00455714
R68775 VSS.n17648 VSS.n17647 0.00455714
R68776 VSS.n17649 VSS.n17648 0.00455714
R68777 VSS.n17650 VSS.n17649 0.00455714
R68778 VSS.n17651 VSS.n17650 0.00455714
R68779 VSS.n17652 VSS.n17651 0.00455714
R68780 VSS.n17653 VSS.n17652 0.00455714
R68781 VSS.n17654 VSS.n17653 0.00455714
R68782 VSS.n17655 VSS.n17654 0.00455714
R68783 VSS.n17656 VSS.n17655 0.00455714
R68784 VSS.n17657 VSS.n17656 0.00455714
R68785 VSS.n17658 VSS.n17657 0.00455714
R68786 VSS.n17659 VSS.n17658 0.00455714
R68787 VSS.n17660 VSS.n17659 0.00455714
R68788 VSS.n17661 VSS.n17660 0.00455714
R68789 VSS.n17662 VSS.n17661 0.00455714
R68790 VSS.n17663 VSS.n17662 0.00455714
R68791 VSS.n17664 VSS.n17663 0.00455714
R68792 VSS.n17665 VSS.n17664 0.00455714
R68793 VSS.n17666 VSS.n17665 0.00455714
R68794 VSS.n17667 VSS.n17666 0.00455714
R68795 VSS.n17668 VSS.n17667 0.00455714
R68796 VSS.n17669 VSS.n17668 0.00455714
R68797 VSS.n17670 VSS.n17669 0.00455714
R68798 VSS.n17671 VSS.n17670 0.00455714
R68799 VSS.n17672 VSS.n17671 0.00455714
R68800 VSS.n17673 VSS.n17672 0.00455714
R68801 VSS.n17674 VSS.n17673 0.00455714
R68802 VSS.n17675 VSS.n17674 0.00455714
R68803 VSS.n17676 VSS.n17675 0.00455714
R68804 VSS.n17677 VSS.n17676 0.00455714
R68805 VSS.n17678 VSS.n17677 0.00455714
R68806 VSS.n17679 VSS.n17678 0.00455714
R68807 VSS.n17680 VSS.n17679 0.00455714
R68808 VSS.n17681 VSS.n17680 0.00455714
R68809 VSS.n17682 VSS.n17681 0.00455714
R68810 VSS.n17683 VSS.n17682 0.00455714
R68811 VSS.n17684 VSS.n17683 0.00455714
R68812 VSS.n17685 VSS.n17684 0.00455714
R68813 VSS.n17686 VSS.n17685 0.00455714
R68814 VSS.n17687 VSS.n17686 0.00455714
R68815 VSS.n17688 VSS.n17687 0.00455714
R68816 VSS.n17689 VSS.n17688 0.00455714
R68817 VSS.n17690 VSS.n17689 0.00455714
R68818 VSS.n17691 VSS.n17690 0.00455714
R68819 VSS.n17692 VSS.n17691 0.00455714
R68820 VSS.n17693 VSS.n17692 0.00455714
R68821 VSS.n17694 VSS.n17693 0.00455714
R68822 VSS.n17695 VSS.n17694 0.00455714
R68823 VSS.n17696 VSS.n17695 0.00455714
R68824 VSS.n17697 VSS.n17696 0.00455714
R68825 VSS.n17698 VSS.n17697 0.00455714
R68826 VSS.n17699 VSS.n17698 0.00455714
R68827 VSS.n17700 VSS.n17699 0.00455714
R68828 VSS.n17701 VSS.n17700 0.00455714
R68829 VSS.n17712 VSS.n17711 0.00455714
R68830 VSS.n17711 VSS.n17710 0.00455714
R68831 VSS.n2539 VSS.n2538 0.00455714
R68832 VSS.n3180 VSS.n3179 0.00455714
R68833 VSS.n3179 VSS.n3178 0.00455714
R68834 VSS.n3178 VSS.n3177 0.00455714
R68835 VSS.n3177 VSS.n3176 0.00455714
R68836 VSS.n3176 VSS.n3175 0.00455714
R68837 VSS.n3175 VSS.n3174 0.00455714
R68838 VSS.n3174 VSS.n3173 0.00455714
R68839 VSS.n3173 VSS.n3172 0.00455714
R68840 VSS.n3172 VSS.n3171 0.00455714
R68841 VSS.n3171 VSS.n3170 0.00455714
R68842 VSS.n3170 VSS.n3169 0.00455714
R68843 VSS.n3169 VSS.n3168 0.00455714
R68844 VSS.n3168 VSS.n3167 0.00455714
R68845 VSS.n3167 VSS.n3166 0.00455714
R68846 VSS.n3166 VSS.n3165 0.00455714
R68847 VSS.n3165 VSS.n3164 0.00455714
R68848 VSS.n3164 VSS.n3163 0.00455714
R68849 VSS.n3163 VSS.n3162 0.00455714
R68850 VSS.n3162 VSS.n3161 0.00455714
R68851 VSS.n3161 VSS.n3160 0.00455714
R68852 VSS.n3160 VSS.n3159 0.00455714
R68853 VSS.n3159 VSS.n3158 0.00455714
R68854 VSS.n3158 VSS.n3157 0.00455714
R68855 VSS.n3157 VSS.n3156 0.00455714
R68856 VSS.n3156 VSS.n3155 0.00455714
R68857 VSS.n3155 VSS.n3154 0.00455714
R68858 VSS.n3154 VSS.n3153 0.00455714
R68859 VSS.n3153 VSS.n3152 0.00455714
R68860 VSS.n3152 VSS.n3151 0.00455714
R68861 VSS.n3151 VSS.n3150 0.00455714
R68862 VSS.n3150 VSS.n3149 0.00455714
R68863 VSS.n3149 VSS.n3148 0.00455714
R68864 VSS.n3148 VSS.n3147 0.00455714
R68865 VSS.n3147 VSS.n3146 0.00455714
R68866 VSS.n3146 VSS.n3145 0.00455714
R68867 VSS.n3145 VSS.n3144 0.00455714
R68868 VSS.n3144 VSS.n3143 0.00455714
R68869 VSS.n3143 VSS.n3142 0.00455714
R68870 VSS.n3142 VSS.n3141 0.00455714
R68871 VSS.n3141 VSS.n3140 0.00455714
R68872 VSS.n3140 VSS.n3139 0.00455714
R68873 VSS.n3139 VSS.n3138 0.00455714
R68874 VSS.n3138 VSS.n3137 0.00455714
R68875 VSS.n3137 VSS.n3136 0.00455714
R68876 VSS.n3136 VSS.n3135 0.00455714
R68877 VSS.n3135 VSS.n3134 0.00455714
R68878 VSS.n3134 VSS.n3133 0.00455714
R68879 VSS.n3133 VSS.n3132 0.00455714
R68880 VSS.n3132 VSS.n3131 0.00455714
R68881 VSS.n3131 VSS.n3130 0.00455714
R68882 VSS.n3130 VSS.n3129 0.00455714
R68883 VSS.n3129 VSS.n3128 0.00455714
R68884 VSS.n3128 VSS.n3127 0.00455714
R68885 VSS.n3127 VSS.n3126 0.00455714
R68886 VSS.n3126 VSS.n3125 0.00455714
R68887 VSS.n3125 VSS.n3124 0.00455714
R68888 VSS.n3124 VSS.n3123 0.00455714
R68889 VSS.n3123 VSS.n3122 0.00455714
R68890 VSS.n3122 VSS.n3121 0.00455714
R68891 VSS.n3121 VSS.n3120 0.00455714
R68892 VSS.n3120 VSS.n3119 0.00455714
R68893 VSS.n3119 VSS.n3118 0.00455714
R68894 VSS.n3118 VSS.n3117 0.00455714
R68895 VSS.n3117 VSS.n3116 0.00455714
R68896 VSS.n3116 VSS.n3115 0.00455714
R68897 VSS.n3115 VSS.n3114 0.00455714
R68898 VSS.n3114 VSS.n3113 0.00455714
R68899 VSS.n3113 VSS.n3112 0.00455714
R68900 VSS.n3112 VSS.n3111 0.00455714
R68901 VSS.n3111 VSS.n3110 0.00455714
R68902 VSS.n3110 VSS.n3109 0.00455714
R68903 VSS.n3109 VSS.n3108 0.00455714
R68904 VSS.n3108 VSS.n3107 0.00455714
R68905 VSS.n3107 VSS.n3106 0.00455714
R68906 VSS.n3106 VSS.n3105 0.00455714
R68907 VSS.n3105 VSS.n3104 0.00455714
R68908 VSS.n3104 VSS.n3103 0.00455714
R68909 VSS.n3103 VSS.n3102 0.00455714
R68910 VSS.n3102 VSS.n3101 0.00455714
R68911 VSS.n3101 VSS.n3100 0.00455714
R68912 VSS.n3100 VSS.n3099 0.00455714
R68913 VSS.n3099 VSS.n3098 0.00455714
R68914 VSS.n3098 VSS.n3097 0.00455714
R68915 VSS.n3097 VSS.n3096 0.00455714
R68916 VSS.n3096 VSS.n3095 0.00455714
R68917 VSS.n3095 VSS.n3094 0.00455714
R68918 VSS.n3094 VSS.n3093 0.00455714
R68919 VSS.n3093 VSS.n3092 0.00455714
R68920 VSS.n3092 VSS.n3091 0.00455714
R68921 VSS.n3091 VSS.n3090 0.00455714
R68922 VSS.n3090 VSS.n3089 0.00455714
R68923 VSS.n3089 VSS.n3088 0.00455714
R68924 VSS.n3088 VSS.n3087 0.00455714
R68925 VSS.n3087 VSS.n3086 0.00455714
R68926 VSS.n3086 VSS.n3085 0.00455714
R68927 VSS.n3085 VSS.n3084 0.00455714
R68928 VSS.n3084 VSS.n2575 0.00455714
R68929 VSS.n2552 VSS.n2551 0.00455714
R68930 VSS.n5409 VSS.n5408 0.00455714
R68931 VSS.n5408 VSS.n5407 0.00455714
R68932 VSS.n5407 VSS.n5406 0.00455714
R68933 VSS.n5406 VSS.n5405 0.00455714
R68934 VSS.n5405 VSS.n5404 0.00455714
R68935 VSS.n5404 VSS.n5403 0.00455714
R68936 VSS.n5403 VSS.n5402 0.00455714
R68937 VSS.n5402 VSS.n5401 0.00455714
R68938 VSS.n5401 VSS.n5400 0.00455714
R68939 VSS.n5400 VSS.n5399 0.00455714
R68940 VSS.n5399 VSS.n5398 0.00455714
R68941 VSS.n5398 VSS.n5397 0.00455714
R68942 VSS.n5397 VSS.n5396 0.00455714
R68943 VSS.n5396 VSS.n5395 0.00455714
R68944 VSS.n5395 VSS.n5394 0.00455714
R68945 VSS.n5394 VSS.n5393 0.00455714
R68946 VSS.n5393 VSS.n5392 0.00455714
R68947 VSS.n5392 VSS.n5391 0.00455714
R68948 VSS.n5391 VSS.n5390 0.00455714
R68949 VSS.n5390 VSS.n5389 0.00455714
R68950 VSS.n5389 VSS.n5388 0.00455714
R68951 VSS.n5388 VSS.n5387 0.00455714
R68952 VSS.n5387 VSS.n5386 0.00455714
R68953 VSS.n5386 VSS.n5385 0.00455714
R68954 VSS.n5385 VSS.n5384 0.00455714
R68955 VSS.n5384 VSS.n5383 0.00455714
R68956 VSS.n5383 VSS.n5382 0.00455714
R68957 VSS.n5382 VSS.n5381 0.00455714
R68958 VSS.n5381 VSS.n5380 0.00455714
R68959 VSS.n5380 VSS.n5379 0.00455714
R68960 VSS.n5379 VSS.n5378 0.00455714
R68961 VSS.n5378 VSS.n5377 0.00455714
R68962 VSS.n5377 VSS.n5376 0.00455714
R68963 VSS.n5376 VSS.n5375 0.00455714
R68964 VSS.n5375 VSS.n5374 0.00455714
R68965 VSS.n5374 VSS.n5373 0.00455714
R68966 VSS.n5373 VSS.n5372 0.00455714
R68967 VSS.n5372 VSS.n5371 0.00455714
R68968 VSS.n5371 VSS.n5370 0.00455714
R68969 VSS.n5370 VSS.n5369 0.00455714
R68970 VSS.n5369 VSS.n5368 0.00455714
R68971 VSS.n5368 VSS.n5367 0.00455714
R68972 VSS.n5367 VSS.n5366 0.00455714
R68973 VSS.n5366 VSS.n5365 0.00455714
R68974 VSS.n5365 VSS.n5364 0.00455714
R68975 VSS.n5364 VSS.n5363 0.00455714
R68976 VSS.n5363 VSS.n5362 0.00455714
R68977 VSS.n5362 VSS.n5361 0.00455714
R68978 VSS.n5361 VSS.n5360 0.00455714
R68979 VSS.n5360 VSS.n5359 0.00455714
R68980 VSS.n5359 VSS.n5358 0.00455714
R68981 VSS.n5358 VSS.n5357 0.00455714
R68982 VSS.n5357 VSS.n5356 0.00455714
R68983 VSS.n5356 VSS.n5355 0.00455714
R68984 VSS.n5355 VSS.n5354 0.00455714
R68985 VSS.n5354 VSS.n5353 0.00455714
R68986 VSS.n5353 VSS.n5352 0.00455714
R68987 VSS.n5352 VSS.n5351 0.00455714
R68988 VSS.n5351 VSS.n5350 0.00455714
R68989 VSS.n5350 VSS.n5349 0.00455714
R68990 VSS.n5349 VSS.n5348 0.00455714
R68991 VSS.n5348 VSS.n5347 0.00455714
R68992 VSS.n5347 VSS.n5346 0.00455714
R68993 VSS.n5346 VSS.n5345 0.00455714
R68994 VSS.n5345 VSS.n5344 0.00455714
R68995 VSS.n5344 VSS.n5343 0.00455714
R68996 VSS.n5343 VSS.n5342 0.00455714
R68997 VSS.n5342 VSS.n5341 0.00455714
R68998 VSS.n5341 VSS.n5340 0.00455714
R68999 VSS.n5340 VSS.n5339 0.00455714
R69000 VSS.n5339 VSS.n5338 0.00455714
R69001 VSS.n5338 VSS.n5337 0.00455714
R69002 VSS.n5337 VSS.n5336 0.00455714
R69003 VSS.n5336 VSS.n5335 0.00455714
R69004 VSS.n5335 VSS.n5334 0.00455714
R69005 VSS.n5334 VSS.n5333 0.00455714
R69006 VSS.n5333 VSS.n5332 0.00455714
R69007 VSS.n5332 VSS.n5331 0.00455714
R69008 VSS.n5331 VSS.n5330 0.00455714
R69009 VSS.n5330 VSS.n5329 0.00455714
R69010 VSS.n5329 VSS.n5328 0.00455714
R69011 VSS.n5328 VSS.n5327 0.00455714
R69012 VSS.n5327 VSS.n5326 0.00455714
R69013 VSS.n5326 VSS.n5325 0.00455714
R69014 VSS.n5325 VSS.n5324 0.00455714
R69015 VSS.n5324 VSS.n5323 0.00455714
R69016 VSS.n5323 VSS.n5322 0.00455714
R69017 VSS.n5322 VSS.n5321 0.00455714
R69018 VSS.n5321 VSS.n5320 0.00455714
R69019 VSS.n5320 VSS.n5319 0.00455714
R69020 VSS.n5319 VSS.n5318 0.00455714
R69021 VSS.n5318 VSS.n5317 0.00455714
R69022 VSS.n5317 VSS.n5316 0.00455714
R69023 VSS.n5316 VSS.n5315 0.00455714
R69024 VSS.n5315 VSS.n5314 0.00455714
R69025 VSS.n5314 VSS.n5313 0.00455714
R69026 VSS.n5313 VSS.n5312 0.00455714
R69027 VSS.n5312 VSS.n4973 0.00455714
R69028 VSS.n4954 VSS.n4953 0.00455714
R69029 VSS.n5918 VSS.n5917 0.00455714
R69030 VSS.n7422 VSS.n7421 0.00455714
R69031 VSS.n7423 VSS.n7422 0.00455714
R69032 VSS.n7424 VSS.n7423 0.00455714
R69033 VSS.n7425 VSS.n7424 0.00455714
R69034 VSS.n7426 VSS.n7425 0.00455714
R69035 VSS.n7427 VSS.n7426 0.00455714
R69036 VSS.n7428 VSS.n7427 0.00455714
R69037 VSS.n7429 VSS.n7428 0.00455714
R69038 VSS.n7430 VSS.n7429 0.00455714
R69039 VSS.n7431 VSS.n7430 0.00455714
R69040 VSS.n7432 VSS.n7431 0.00455714
R69041 VSS.n7433 VSS.n7432 0.00455714
R69042 VSS.n7434 VSS.n7433 0.00455714
R69043 VSS.n7435 VSS.n7434 0.00455714
R69044 VSS.n7436 VSS.n7435 0.00455714
R69045 VSS.n7437 VSS.n7436 0.00455714
R69046 VSS.n7438 VSS.n7437 0.00455714
R69047 VSS.n7439 VSS.n7438 0.00455714
R69048 VSS.n7440 VSS.n7439 0.00455714
R69049 VSS.n7441 VSS.n7440 0.00455714
R69050 VSS.n7442 VSS.n7441 0.00455714
R69051 VSS.n7443 VSS.n7442 0.00455714
R69052 VSS.n7444 VSS.n7443 0.00455714
R69053 VSS.n7445 VSS.n7444 0.00455714
R69054 VSS.n7446 VSS.n7445 0.00455714
R69055 VSS.n7447 VSS.n7446 0.00455714
R69056 VSS.n7448 VSS.n7447 0.00455714
R69057 VSS.n7449 VSS.n7448 0.00455714
R69058 VSS.n7450 VSS.n7449 0.00455714
R69059 VSS.n7451 VSS.n7450 0.00455714
R69060 VSS.n7452 VSS.n7451 0.00455714
R69061 VSS.n7453 VSS.n7452 0.00455714
R69062 VSS.n7454 VSS.n7453 0.00455714
R69063 VSS.n7455 VSS.n7454 0.00455714
R69064 VSS.n7456 VSS.n7455 0.00455714
R69065 VSS.n7457 VSS.n7456 0.00455714
R69066 VSS.n7458 VSS.n7457 0.00455714
R69067 VSS.n7459 VSS.n7458 0.00455714
R69068 VSS.n7460 VSS.n7459 0.00455714
R69069 VSS.n7461 VSS.n7460 0.00455714
R69070 VSS.n7462 VSS.n7461 0.00455714
R69071 VSS.n7463 VSS.n7462 0.00455714
R69072 VSS.n7464 VSS.n7463 0.00455714
R69073 VSS.n7465 VSS.n7464 0.00455714
R69074 VSS.n7466 VSS.n7465 0.00455714
R69075 VSS.n7467 VSS.n7466 0.00455714
R69076 VSS.n7468 VSS.n7467 0.00455714
R69077 VSS.n7469 VSS.n7468 0.00455714
R69078 VSS.n7470 VSS.n7469 0.00455714
R69079 VSS.n7471 VSS.n7470 0.00455714
R69080 VSS.n7472 VSS.n7471 0.00455714
R69081 VSS.n7473 VSS.n7472 0.00455714
R69082 VSS.n7474 VSS.n7473 0.00455714
R69083 VSS.n7475 VSS.n7474 0.00455714
R69084 VSS.n7476 VSS.n7475 0.00455714
R69085 VSS.n7477 VSS.n7476 0.00455714
R69086 VSS.n7478 VSS.n7477 0.00455714
R69087 VSS.n7479 VSS.n7478 0.00455714
R69088 VSS.n7480 VSS.n7479 0.00455714
R69089 VSS.n7481 VSS.n7480 0.00455714
R69090 VSS.n7482 VSS.n7481 0.00455714
R69091 VSS.n7483 VSS.n7482 0.00455714
R69092 VSS.n7484 VSS.n7483 0.00455714
R69093 VSS.n7485 VSS.n7484 0.00455714
R69094 VSS.n7486 VSS.n7485 0.00455714
R69095 VSS.n7487 VSS.n7486 0.00455714
R69096 VSS.n7488 VSS.n7487 0.00455714
R69097 VSS.n7489 VSS.n7488 0.00455714
R69098 VSS.n7490 VSS.n7489 0.00455714
R69099 VSS.n7491 VSS.n7490 0.00455714
R69100 VSS.n7492 VSS.n7491 0.00455714
R69101 VSS.n7493 VSS.n7492 0.00455714
R69102 VSS.n7494 VSS.n7493 0.00455714
R69103 VSS.n7495 VSS.n7494 0.00455714
R69104 VSS.n7496 VSS.n7495 0.00455714
R69105 VSS.n7497 VSS.n7496 0.00455714
R69106 VSS.n7498 VSS.n7497 0.00455714
R69107 VSS.n7499 VSS.n7498 0.00455714
R69108 VSS.n7500 VSS.n7499 0.00455714
R69109 VSS.n7501 VSS.n7500 0.00455714
R69110 VSS.n7502 VSS.n7501 0.00455714
R69111 VSS.n7503 VSS.n7502 0.00455714
R69112 VSS.n7504 VSS.n7503 0.00455714
R69113 VSS.n7505 VSS.n7504 0.00455714
R69114 VSS.n7506 VSS.n7505 0.00455714
R69115 VSS.n7507 VSS.n7506 0.00455714
R69116 VSS.n7508 VSS.n7507 0.00455714
R69117 VSS.n7509 VSS.n7508 0.00455714
R69118 VSS.n7510 VSS.n7509 0.00455714
R69119 VSS.n7511 VSS.n7510 0.00455714
R69120 VSS.n7512 VSS.n7511 0.00455714
R69121 VSS.n7513 VSS.n7512 0.00455714
R69122 VSS.n7514 VSS.n7513 0.00455714
R69123 VSS.n7515 VSS.n7514 0.00455714
R69124 VSS.n7516 VSS.n7515 0.00455714
R69125 VSS.n7518 VSS.n7517 0.00455714
R69126 VSS.n7537 VSS.n7536 0.00455714
R69127 VSS.n4214 VSS.n4213 0.00455714
R69128 VSS.n4215 VSS.n4214 0.00455714
R69129 VSS.n4216 VSS.n4215 0.00455714
R69130 VSS.n4217 VSS.n4216 0.00455714
R69131 VSS.n4218 VSS.n4217 0.00455714
R69132 VSS.n4219 VSS.n4218 0.00455714
R69133 VSS.n4220 VSS.n4219 0.00455714
R69134 VSS.n4221 VSS.n4220 0.00455714
R69135 VSS.n4222 VSS.n4221 0.00455714
R69136 VSS.n4223 VSS.n4222 0.00455714
R69137 VSS.n4224 VSS.n4223 0.00455714
R69138 VSS.n4225 VSS.n4224 0.00455714
R69139 VSS.n4226 VSS.n4225 0.00455714
R69140 VSS.n4227 VSS.n4226 0.00455714
R69141 VSS.n4228 VSS.n4227 0.00455714
R69142 VSS.n4229 VSS.n4228 0.00455714
R69143 VSS.n4230 VSS.n4229 0.00455714
R69144 VSS.n4231 VSS.n4230 0.00455714
R69145 VSS.n4232 VSS.n4231 0.00455714
R69146 VSS.n4233 VSS.n4232 0.00455714
R69147 VSS.n4234 VSS.n4233 0.00455714
R69148 VSS.n4235 VSS.n4234 0.00455714
R69149 VSS.n4236 VSS.n4235 0.00455714
R69150 VSS.n4237 VSS.n4236 0.00455714
R69151 VSS.n4238 VSS.n4237 0.00455714
R69152 VSS.n4239 VSS.n4238 0.00455714
R69153 VSS.n4240 VSS.n4239 0.00455714
R69154 VSS.n4241 VSS.n4240 0.00455714
R69155 VSS.n4242 VSS.n4241 0.00455714
R69156 VSS.n4243 VSS.n4242 0.00455714
R69157 VSS.n4244 VSS.n4243 0.00455714
R69158 VSS.n4245 VSS.n4244 0.00455714
R69159 VSS.n4246 VSS.n4245 0.00455714
R69160 VSS.n4247 VSS.n4246 0.00455714
R69161 VSS.n4248 VSS.n4247 0.00455714
R69162 VSS.n4249 VSS.n4248 0.00455714
R69163 VSS.n4250 VSS.n4249 0.00455714
R69164 VSS.n4251 VSS.n4250 0.00455714
R69165 VSS.n4252 VSS.n4251 0.00455714
R69166 VSS.n4253 VSS.n4252 0.00455714
R69167 VSS.n4254 VSS.n4253 0.00455714
R69168 VSS.n4255 VSS.n4254 0.00455714
R69169 VSS.n4256 VSS.n4255 0.00455714
R69170 VSS.n4257 VSS.n4256 0.00455714
R69171 VSS.n4258 VSS.n4257 0.00455714
R69172 VSS.n4259 VSS.n4258 0.00455714
R69173 VSS.n4260 VSS.n4259 0.00455714
R69174 VSS.n4261 VSS.n4260 0.00455714
R69175 VSS.n4262 VSS.n4261 0.00455714
R69176 VSS.n4263 VSS.n4262 0.00455714
R69177 VSS.n4264 VSS.n4263 0.00455714
R69178 VSS.n4265 VSS.n4264 0.00455714
R69179 VSS.n4266 VSS.n4265 0.00455714
R69180 VSS.n4267 VSS.n4266 0.00455714
R69181 VSS.n4268 VSS.n4267 0.00455714
R69182 VSS.n4269 VSS.n4268 0.00455714
R69183 VSS.n4270 VSS.n4269 0.00455714
R69184 VSS.n4271 VSS.n4270 0.00455714
R69185 VSS.n4272 VSS.n4271 0.00455714
R69186 VSS.n4273 VSS.n4272 0.00455714
R69187 VSS.n4274 VSS.n4273 0.00455714
R69188 VSS.n4275 VSS.n4274 0.00455714
R69189 VSS.n4276 VSS.n4275 0.00455714
R69190 VSS.n4277 VSS.n4276 0.00455714
R69191 VSS.n4278 VSS.n4277 0.00455714
R69192 VSS.n4279 VSS.n4278 0.00455714
R69193 VSS.n4280 VSS.n4279 0.00455714
R69194 VSS.n4281 VSS.n4280 0.00455714
R69195 VSS.n4282 VSS.n4281 0.00455714
R69196 VSS.n4283 VSS.n4282 0.00455714
R69197 VSS.n4284 VSS.n4283 0.00455714
R69198 VSS.n4285 VSS.n4284 0.00455714
R69199 VSS.n4286 VSS.n4285 0.00455714
R69200 VSS.n4287 VSS.n4286 0.00455714
R69201 VSS.n4288 VSS.n4287 0.00455714
R69202 VSS.n4289 VSS.n4288 0.00455714
R69203 VSS.n4290 VSS.n4289 0.00455714
R69204 VSS.n4291 VSS.n4290 0.00455714
R69205 VSS.n4292 VSS.n4291 0.00455714
R69206 VSS.n4293 VSS.n4292 0.00455714
R69207 VSS.n4294 VSS.n4293 0.00455714
R69208 VSS.n4295 VSS.n4294 0.00455714
R69209 VSS.n4296 VSS.n4295 0.00455714
R69210 VSS.n4297 VSS.n4296 0.00455714
R69211 VSS.n4298 VSS.n4297 0.00455714
R69212 VSS.n4299 VSS.n4298 0.00455714
R69213 VSS.n4300 VSS.n4299 0.00455714
R69214 VSS.n4301 VSS.n4300 0.00455714
R69215 VSS.n4302 VSS.n4301 0.00455714
R69216 VSS.n4303 VSS.n4302 0.00455714
R69217 VSS.n4304 VSS.n4303 0.00455714
R69218 VSS.n4305 VSS.n4304 0.00455714
R69219 VSS.n4306 VSS.n4305 0.00455714
R69220 VSS.n4307 VSS.n4306 0.00455714
R69221 VSS.n4308 VSS.n4307 0.00455714
R69222 VSS.n4309 VSS.n4308 0.00455714
R69223 VSS.n4322 VSS.n4309 0.00455714
R69224 VSS.n4321 VSS.n4311 0.00455714
R69225 VSS.n4311 VSS.n4310 0.00455714
R69226 VSS.n22010 VSS.n22009 0.00455714
R69227 VSS.n22011 VSS.n22010 0.00455714
R69228 VSS.n22012 VSS.n22011 0.00455714
R69229 VSS.n22013 VSS.n22012 0.00455714
R69230 VSS.n22014 VSS.n22013 0.00455714
R69231 VSS.n22015 VSS.n22014 0.00455714
R69232 VSS.n22016 VSS.n22015 0.00455714
R69233 VSS.n22017 VSS.n22016 0.00455714
R69234 VSS.n22018 VSS.n22017 0.00455714
R69235 VSS.n22019 VSS.n22018 0.00455714
R69236 VSS.n22020 VSS.n22019 0.00455714
R69237 VSS.n22021 VSS.n22020 0.00455714
R69238 VSS.n22022 VSS.n22021 0.00455714
R69239 VSS.n22023 VSS.n22022 0.00455714
R69240 VSS.n22024 VSS.n22023 0.00455714
R69241 VSS.n22025 VSS.n22024 0.00455714
R69242 VSS.n22026 VSS.n22025 0.00455714
R69243 VSS.n22027 VSS.n22026 0.00455714
R69244 VSS.n22028 VSS.n22027 0.00455714
R69245 VSS.n22029 VSS.n22028 0.00455714
R69246 VSS.n22030 VSS.n22029 0.00455714
R69247 VSS.n22031 VSS.n22030 0.00455714
R69248 VSS.n22032 VSS.n22031 0.00455714
R69249 VSS.n22033 VSS.n22032 0.00455714
R69250 VSS.n22034 VSS.n22033 0.00455714
R69251 VSS.n22035 VSS.n22034 0.00455714
R69252 VSS.n22036 VSS.n22035 0.00455714
R69253 VSS.n22037 VSS.n22036 0.00455714
R69254 VSS.n22038 VSS.n22037 0.00455714
R69255 VSS.n22039 VSS.n22038 0.00455714
R69256 VSS.n22040 VSS.n22039 0.00455714
R69257 VSS.n22041 VSS.n22040 0.00455714
R69258 VSS.n22042 VSS.n22041 0.00455714
R69259 VSS.n22043 VSS.n22042 0.00455714
R69260 VSS.n22044 VSS.n22043 0.00455714
R69261 VSS.n22045 VSS.n22044 0.00455714
R69262 VSS.n22046 VSS.n22045 0.00455714
R69263 VSS.n22047 VSS.n22046 0.00455714
R69264 VSS.n22048 VSS.n22047 0.00455714
R69265 VSS.n22049 VSS.n22048 0.00455714
R69266 VSS.n22050 VSS.n22049 0.00455714
R69267 VSS.n22051 VSS.n22050 0.00455714
R69268 VSS.n22052 VSS.n22051 0.00455714
R69269 VSS.n22053 VSS.n22052 0.00455714
R69270 VSS.n22054 VSS.n22053 0.00455714
R69271 VSS.n22055 VSS.n22054 0.00455714
R69272 VSS.n22056 VSS.n22055 0.00455714
R69273 VSS.n22057 VSS.n22056 0.00455714
R69274 VSS.n22058 VSS.n22057 0.00455714
R69275 VSS.n22059 VSS.n22058 0.00455714
R69276 VSS.n22060 VSS.n22059 0.00455714
R69277 VSS.n22061 VSS.n22060 0.00455714
R69278 VSS.n22062 VSS.n22061 0.00455714
R69279 VSS.n22063 VSS.n22062 0.00455714
R69280 VSS.n22064 VSS.n22063 0.00455714
R69281 VSS.n22065 VSS.n22064 0.00455714
R69282 VSS.n22066 VSS.n22065 0.00455714
R69283 VSS.n22067 VSS.n22066 0.00455714
R69284 VSS.n22068 VSS.n22067 0.00455714
R69285 VSS.n22069 VSS.n22068 0.00455714
R69286 VSS.n22070 VSS.n22069 0.00455714
R69287 VSS.n22071 VSS.n22070 0.00455714
R69288 VSS.n22072 VSS.n22071 0.00455714
R69289 VSS.n22073 VSS.n22072 0.00455714
R69290 VSS.n22074 VSS.n22073 0.00455714
R69291 VSS.n22075 VSS.n22074 0.00455714
R69292 VSS.n22076 VSS.n22075 0.00455714
R69293 VSS.n22077 VSS.n22076 0.00455714
R69294 VSS.n22078 VSS.n22077 0.00455714
R69295 VSS.n22079 VSS.n22078 0.00455714
R69296 VSS.n22080 VSS.n22079 0.00455714
R69297 VSS.n22081 VSS.n22080 0.00455714
R69298 VSS.n22082 VSS.n22081 0.00455714
R69299 VSS.n22083 VSS.n22082 0.00455714
R69300 VSS.n22084 VSS.n22083 0.00455714
R69301 VSS.n22085 VSS.n22084 0.00455714
R69302 VSS.n22086 VSS.n22085 0.00455714
R69303 VSS.n22087 VSS.n22086 0.00455714
R69304 VSS.n22088 VSS.n22087 0.00455714
R69305 VSS.n22089 VSS.n22088 0.00455714
R69306 VSS.n22090 VSS.n22089 0.00455714
R69307 VSS.n22091 VSS.n22090 0.00455714
R69308 VSS.n22092 VSS.n22091 0.00455714
R69309 VSS.n22093 VSS.n22092 0.00455714
R69310 VSS.n22094 VSS.n22093 0.00455714
R69311 VSS.n22095 VSS.n22094 0.00455714
R69312 VSS.n22096 VSS.n22095 0.00455714
R69313 VSS.n22097 VSS.n22096 0.00455714
R69314 VSS.n22098 VSS.n22097 0.00455714
R69315 VSS.n22099 VSS.n22098 0.00455714
R69316 VSS.n22100 VSS.n22099 0.00455714
R69317 VSS.n22101 VSS.n22100 0.00455714
R69318 VSS.n22102 VSS.n22101 0.00455714
R69319 VSS.n22103 VSS.n22102 0.00455714
R69320 VSS.n22104 VSS.n22103 0.00455714
R69321 VSS.n22105 VSS.n22104 0.00455714
R69322 VSS.n22262 VSS.n22105 0.00455714
R69323 VSS.n22262 VSS.n22261 0.00455714
R69324 VSS.n22261 VSS.n22260 0.00455714
R69325 VSS.n18366 VSS.n18363 0.00455
R69326 VSS.n16572 VSS.n16571 0.00455
R69327 VSS.n4669 VSS.n4666 0.00455
R69328 VSS.n13020 VSS.n13019 0.0045432
R69329 VSS.n21793 VSS.n21792 0.0045432
R69330 VSS.n19078 VSS.n19077 0.0045432
R69331 VSS.n10292 VSS.n10291 0.00453846
R69332 VSS.n10410 VSS.n10409 0.00453846
R69333 VSS.n10393 VSS.n10388 0.00453846
R69334 VSS.n10125 VSS.n10124 0.00453846
R69335 VSS.n10108 VSS.n10103 0.00453846
R69336 VSS.n8888 VSS.n8865 0.00453846
R69337 VSS.n12346 VSS.n12345 0.00453846
R69338 VSS.n12464 VSS.n12463 0.00453846
R69339 VSS.n12447 VSS.n12442 0.00453846
R69340 VSS.n12176 VSS.n12175 0.00453846
R69341 VSS.n12159 VSS.n12154 0.00453846
R69342 VSS.n12028 VSS.n12027 0.00453846
R69343 VSS.n12011 VSS.n11995 0.00453846
R69344 VSS.n9850 VSS.n9847 0.00453846
R69345 VSS.n12647 VSS.n12639 0.00453846
R69346 VSS.n20234 VSS.n20233 0.00452
R69347 VSS.n20229 VSS.n20228 0.00452
R69348 VSS.n10840 VSS.n10839 0.00452
R69349 VSS.n8747 VSS.n8746 0.00452
R69350 VSS.n8290 VSS.n8289 0.00452
R69351 VSS.n8285 VSS.n8284 0.00452
R69352 VSS.n8742 VSS.n8741 0.00452
R69353 VSS.n10844 VSS.n10843 0.00452
R69354 VSS.n15648 VSS.n15637 0.00451837
R69355 VSS.n15621 VSS.n15614 0.00451837
R69356 VSS.n15598 VSS.n15591 0.00451837
R69357 VSS.n15520 VSS.n15475 0.00451837
R69358 VSS.n1906 VSS.n1905 0.00451837
R69359 VSS.n1889 VSS.n1888 0.00451837
R69360 VSS.n1872 VSS.n1871 0.00451837
R69361 VSS.n1808 VSS.n1777 0.00451837
R69362 VSS.n1739 VSS.n1732 0.00451837
R69363 VSS.n18675 VSS.n18674 0.00451408
R69364 VSS.n18444 VSS.n18443 0.00451408
R69365 VSS.n18441 VSS.n18440 0.00451408
R69366 VSS.n18392 VSS.n18391 0.00451408
R69367 VSS.n17070 VSS.n17069 0.00451408
R69368 VSS.n17067 VSS.n17066 0.00451408
R69369 VSS.n17032 VSS.n17031 0.00451408
R69370 VSS.n16935 VSS.n16934 0.00451408
R69371 VSS.n16902 VSS.n16901 0.00451408
R69372 VSS.n16635 VSS.n16634 0.00451408
R69373 VSS.n16527 VSS.n16526 0.00451408
R69374 VSS.n15371 VSS.n15370 0.00451408
R69375 VSS.n8573 VSS.n8572 0.00451408
R69376 VSS.n8428 VSS.n8427 0.00451408
R69377 VSS.n19528 VSS.n19527 0.00451408
R69378 VSS.n19595 VSS.n19594 0.00451408
R69379 VSS.n19598 VSS.n19597 0.00451408
R69380 VSS.n19630 VSS.n19629 0.00451408
R69381 VSS.n19895 VSS.n19894 0.00451408
R69382 VSS.n19898 VSS.n19897 0.00451408
R69383 VSS.n19903 VSS.n19902 0.00451408
R69384 VSS.n19981 VSS.n19980 0.00451408
R69385 VSS.n20014 VSS.n20013 0.00451408
R69386 VSS.n763 VSS.n762 0.00451408
R69387 VSS.n811 VSS.n810 0.00451408
R69388 VSS.n1687 VSS.n1686 0.00451408
R69389 VSS.n8724 VSS.n8723 0.00451408
R69390 VSS.n8236 VSS.n8235 0.00451408
R69391 VSS.n13662 VSS 0.0045
R69392 VSS.n4187 VSS.n2450 0.00449949
R69393 VSS.n17344 VSS.n17343 0.00449949
R69394 VSS.n17333 VSS.n17332 0.00449949
R69395 VSS.n11522 VSS.n11521 0.00449949
R69396 VSS.n11324 VSS.n11323 0.00449949
R69397 VSS.n11319 VSS.n11318 0.00449949
R69398 VSS.n12833 VSS.n12832 0.00449949
R69399 VSS.n12887 VSS.n12886 0.00449949
R69400 VSS.n12900 VSS.n12899 0.00449949
R69401 VSS.n13001 VSS.n13000 0.00449949
R69402 VSS.n13245 VSS.n13244 0.00449949
R69403 VSS.n18986 VSS.n18979 0.00449949
R69404 VSS.n2213 VSS.n2212 0.00449949
R69405 VSS.n14398 VSS.n14397 0.00449949
R69406 VSS.n14425 VSS.n14424 0.00449949
R69407 VSS.n15072 VSS.n15071 0.00449949
R69408 VSS.n15105 VSS.n15104 0.00449949
R69409 VSS.n15175 VSS.n15174 0.00449949
R69410 VSS.n16314 VSS.n16313 0.00449949
R69411 VSS.n16279 VSS.n16278 0.00449949
R69412 VSS.n16359 VSS.n16358 0.00449949
R69413 VSS.n5717 VSS.n5716 0.00449949
R69414 VSS.n21743 VSS.n21742 0.00449949
R69415 VSS.n13329 VSS.n13328 0.00449949
R69416 VSS.n13362 VSS.n13361 0.00449949
R69417 VSS.n13413 VSS.n13412 0.00449949
R69418 VSS.n20684 VSS.n20683 0.00449949
R69419 VSS.n20735 VSS.n20734 0.00449949
R69420 VSS.n20827 VSS.n20826 0.00449949
R69421 VSS.n21105 VSS.n21104 0.00449949
R69422 VSS.n19028 VSS.n19027 0.00449949
R69423 VSS.n20145 VSS.n20144 0.00449949
R69424 VSS.n13505 VSS.n13504 0.00449949
R69425 VSS.n881 VSS.n880 0.00449949
R69426 VSS.n2046 VSS.n2045 0.00449949
R69427 VSS.n2051 VSS.n2050 0.00449949
R69428 VSS.n4163 VSS.n4140 0.00449949
R69429 VSS.n582 VSS.n581 0.00449949
R69430 VSS.n595 VSS.n594 0.00449949
R69431 VSS.n532 VSS.n531 0.00449949
R69432 VSS.n15344 VSS.n15343 0.00448591
R69433 VSS.n1660 VSS.n1659 0.00448591
R69434 VSS.n2531 VSS.n2530 0.00448571
R69435 VSS.n2883 VSS.n2882 0.00448571
R69436 VSS.n2921 VSS.n2920 0.00448571
R69437 VSS.n2985 VSS.n2984 0.00448571
R69438 VSS.n3033 VSS.n3032 0.00448571
R69439 VSS.n2441 VSS.n2440 0.00448571
R69440 VSS.n4742 VSS.n4741 0.00448571
R69441 VSS.n18017 VSS.n18016 0.00448571
R69442 VSS.n17982 VSS.n17979 0.00448571
R69443 VSS.n17828 VSS.n17825 0.00448571
R69444 VSS.n17783 VSS.n17780 0.00448571
R69445 VSS.n4954 DVSS 0.00447143
R69446 VSS.n3242 VSS.n3241 0.00444366
R69447 VSS.n3325 VSS.n3324 0.00444366
R69448 VSS.n3379 VSS.n3378 0.00444366
R69449 VSS.n3441 VSS.n3440 0.00444366
R69450 VSS.n2562 VSS.n2561 0.00442143
R69451 VSS.n4671 VSS.n4669 0.00442143
R69452 VSS.n4328 VSS.n4327 0.00442143
R69453 VSS.n17720 VSS.n17719 0.00442143
R69454 VSS.n5840 VSS.n5839 0.00439764
R69455 VSS.n9498 VSS.n9497 0.00439764
R69456 VSS.n11892 VSS.n11891 0.00439764
R69457 VSS.n11875 VSS.n11874 0.00439764
R69458 VSS.n11796 VSS.n11795 0.00439764
R69459 VSS.n16201 VSS.n16200 0.00439764
R69460 VSS.n9615 VSS.n9614 0.00439764
R69461 VSS.n21143 VSS.n21142 0.00439764
R69462 VSS.n6929 VSS.n6928 0.00439764
R69463 VSS.n1272 VSS.n1271 0.00439764
R69464 VSS.n6806 VSS.n6805 0.00439764
R69465 VSS.n8983 VSS.n8982 0.00439764
R69466 VSS.n8899 VSS.n8898 0.00439764
R69467 VSS.n18709 VSS.n18708 0.00437965
R69468 VSS.n19191 VSS.n19190 0.00437965
R69469 VSS.n15651 VSS.n15650 0.00437774
R69470 VSS.n15624 VSS.n15623 0.00437774
R69471 VSS.n15601 VSS.n15600 0.00437774
R69472 VSS.n1909 VSS.n1908 0.00437774
R69473 VSS.n1892 VSS.n1891 0.00437774
R69474 VSS.n1875 VSS.n1874 0.00437774
R69475 VSS.n19513 VSS.n19512 0.00437774
R69476 VSS.n18840 VSS.n18690 0.00437774
R69477 VSS.n3533 VSS.n3532 0.00437324
R69478 VSS.n3592 VSS.n3591 0.00437324
R69479 VSS.n3635 VSS.n3634 0.00437324
R69480 VSS.n14201 VSS.n14200 0.00437247
R69481 VSS.n14155 VSS.n14154 0.00437247
R69482 VSS.n19255 VSS.n19252 0.004325
R69483 VSS.n19264 VSS.n19263 0.004325
R69484 VSS.n16983 VSS.n16982 0.004325
R69485 VSS.n16977 VSS.n16975 0.004325
R69486 VSS.n11714 VSS.n11713 0.00431
R69487 VSS.n18811 VSS.n18810 0.00430282
R69488 VSS.n18825 VSS.n18824 0.00430282
R69489 VSS.n17077 VSS.n17076 0.00430282
R69490 VSS.n16919 VSS.n16918 0.00430282
R69491 VSS.n8461 VSS.n8460 0.00430282
R69492 VSS.n8543 VSS.n8542 0.00430282
R69493 VSS.n8309 VSS.n8308 0.00430282
R69494 VSS.n8398 VSS.n8397 0.00430282
R69495 VSS.n8379 VSS.n8378 0.00430282
R69496 VSS.n19483 VSS.n19482 0.00430282
R69497 VSS.n19497 VSS.n19496 0.00430282
R69498 VSS.n19888 VSS.n19887 0.00430282
R69499 VSS.n19997 VSS.n19996 0.00430282
R69500 VSS.n8612 VSS.n8611 0.00430282
R69501 VSS.n8694 VSS.n8693 0.00430282
R69502 VSS.n8105 VSS.n8104 0.00430282
R69503 VSS.n8206 VSS.n8205 0.00430282
R69504 VSS.n8187 VSS.n8186 0.00430282
R69505 VSS.n13097 VSS.n13096 0.00427756
R69506 VSS.n21870 VSS.n21869 0.00427756
R69507 VSS.n19155 VSS.n19154 0.00427756
R69508 VSS.n21234 VSS.n21233 0.00426578
R69509 VSS.n330 VSS.n329 0.00426578
R69510 VSS.n3466 VSS.n3465 0.00423239
R69511 VSS.n2699 VSS.n2694 0.00422857
R69512 VSS.n2752 VSS.n2738 0.00422857
R69513 VSS.n2802 VSS.n2798 0.00422857
R69514 VSS.n17531 VSS.n17530 0.00422857
R69515 VSS.n18097 VSS.n18096 0.00422857
R69516 VSS.n4002 VSS.n4001 0.00422047
R69517 VSS.n17456 VSS.n17455 0.00422047
R69518 VSS.n13027 VSS.n13026 0.00422047
R69519 VSS.n12542 VSS.n12541 0.00422047
R69520 VSS.n12541 VSS.n12540 0.00422047
R69521 VSS.n11972 VSS.n11971 0.00422047
R69522 VSS.n11945 VSS.n11944 0.00422047
R69523 VSS.n11873 VSS.n11872 0.00422047
R69524 VSS.n18873 VSS.n18872 0.00422047
R69525 VSS.n2207 VSS.n2206 0.00422047
R69526 VSS.n21800 VSS.n21799 0.00422047
R69527 VSS.n19085 VSS.n19084 0.00422047
R69528 VSS.n21571 VSS.n21570 0.00422047
R69529 VSS.n21676 VSS.n21675 0.00422047
R69530 VSS.n21453 VSS.n21452 0.00422047
R69531 VSS.n3804 VSS.n3803 0.00422047
R69532 VSS.n4137 VSS.n4136 0.00422047
R69533 VSS.n4782 VSS.n4781 0.00422047
R69534 VSS.n3282 VSS.n3281 0.00422047
R69535 VSS.n10487 VSS.n10486 0.00422047
R69536 VSS.n10486 VSS.n10485 0.00422047
R69537 VSS.n9975 VSS.n9974 0.00422047
R69538 VSS.n9947 VSS.n9946 0.00422047
R69539 VSS.n8788 VSS.n8787 0.00422047
R69540 VSS.n20521 VSS.n20520 0.00422
R69541 VSS.n14982 VSS.n14981 0.00416802
R69542 VSS.n818 VSS.n817 0.00416802
R69543 VSS.n14902 VSS.n14901 0.00416734
R69544 VSS.n19973 VSS.n19972 0.00416734
R69545 VSS.n4976 VSS.n4975 0.00416429
R69546 VSS.n5006 VSS.n5005 0.00416429
R69547 VSS.n5036 VSS.n5035 0.00416429
R69548 VSS.n5082 VSS.n5081 0.00416429
R69549 VSS.n7419 VSS.n7418 0.00416429
R69550 VSS.n7390 VSS.n7388 0.00416429
R69551 VSS.n4620 VSS.n4618 0.00416429
R69552 VSS.n4574 VSS.n4572 0.00416429
R69553 VSS.n10322 VSS.n10321 0.00415385
R69554 VSS.n10440 VSS.n10439 0.00415385
R69555 VSS.n10348 VSS.n10347 0.00415385
R69556 VSS.n10155 VSS.n10154 0.00415385
R69557 VSS.n10063 VSS.n10062 0.00415385
R69558 VSS.n10022 VSS.n10017 0.00415385
R69559 VSS.n12376 VSS.n12375 0.00415385
R69560 VSS.n12494 VSS.n12493 0.00415385
R69561 VSS.n12402 VSS.n12401 0.00415385
R69562 VSS.n12206 VSS.n12205 0.00415385
R69563 VSS.n12114 VSS.n12113 0.00415385
R69564 VSS.n12073 VSS.n12068 0.00415385
R69565 VSS.n5900 VSS.n5899 0.00414027
R69566 VSS.n5899 VSS.n5898 0.00414027
R69567 VSS.n18482 VSS.n2162 0.0041
R69568 VSS.n18375 VSS.n18374 0.0041
R69569 VSS.n14964 VSS.n14963 0.0041
R69570 VSS.n14764 VSS.n14379 0.0041
R69571 VSS.n14659 VSS.n14658 0.0041
R69572 VSS.n14933 VSS.n14932 0.0041
R69573 VSS.n16565 VSS.n16564 0.0041
R69574 VSS.n16424 VSS.n16423 0.0041
R69575 VSS.n5126 VSS.n5125 0.0041
R69576 VSS.n7367 VSS.n7366 0.0041
R69577 VSS.n7313 VSS.n7312 0.0041
R69578 DVSS VSS.n4321 0.0041
R69579 VSS.n4529 VSS.n4528 0.0041
R69580 VSS.n15899 VSS.n15898 0.0041
R69581 VSS.n186 VSS.n174 0.00409785
R69582 VSS.n5897 VSS.n5894 0.00409785
R69583 VSS.n18740 VSS.n18739 0.00409155
R69584 VSS.n18808 VSS.n18807 0.00409155
R69585 VSS.n18408 VSS.n18407 0.00409155
R69586 VSS.n14858 VSS.n14857 0.00409155
R69587 VSS.n14884 VSS.n14883 0.00409155
R69588 VSS.n14893 VSS.n14892 0.00409155
R69589 VSS.n16900 VSS.n16899 0.00409155
R69590 VSS.n16588 VSS.n16587 0.00409155
R69591 VSS.n15352 VSS.n15351 0.00409155
R69592 VSS.n8472 VSS.n8471 0.00409155
R69593 VSS.n8554 VSS.n8553 0.00409155
R69594 VSS.n8320 VSS.n8319 0.00409155
R69595 VSS.n8409 VSS.n8408 0.00409155
R69596 VSS.n8368 VSS.n8367 0.00409155
R69597 VSS.n19222 VSS.n19221 0.00409155
R69598 VSS.n19480 VSS.n19479 0.00409155
R69599 VSS.n19614 VSS.n19613 0.00409155
R69600 VSS.n19929 VSS.n19928 0.00409155
R69601 VSS.n19955 VSS.n19954 0.00409155
R69602 VSS.n19964 VSS.n19963 0.00409155
R69603 VSS.n20016 VSS.n20015 0.00409155
R69604 VSS.n780 VSS.n779 0.00409155
R69605 VSS.n1668 VSS.n1667 0.00409155
R69606 VSS.n8623 VSS.n8622 0.00409155
R69607 VSS.n8705 VSS.n8704 0.00409155
R69608 VSS.n8116 VSS.n8115 0.00409155
R69609 VSS.n8217 VSS.n8216 0.00409155
R69610 VSS.n8176 VSS.n8175 0.00409155
R69611 VSS.n17479 VSS.n17478 0.00406877
R69612 VSS.n17470 VSS.n17469 0.00406877
R69613 VSS.n17439 VSS.n17438 0.00406877
R69614 VSS.n13195 VSS.n13194 0.00406877
R69615 VSS.n13204 VSS.n13203 0.00406877
R69616 VSS.n13226 VSS.n13225 0.00406877
R69617 VSS.n13234 VSS.n13233 0.00406877
R69618 VSS.n17448 VSS.n17447 0.00406877
R69619 VSS.n2190 VSS.n2189 0.00406877
R69620 VSS.n13351 VSS.n13350 0.00406877
R69621 VSS.n13494 VSS.n13493 0.00406877
R69622 VSS.n14989 VSS.n14988 0.00406336
R69623 VSS.n15386 VSS.n15385 0.00406336
R69624 VSS.n825 VSS.n824 0.00406336
R69625 VSS.n1702 VSS.n1701 0.00406336
R69626 VSS.n14896 VSS.n14895 0.00406318
R69627 VSS.n19967 VSS.n19966 0.00406318
R69628 VSS.n4208 VSS.n4207 0.00404331
R69629 VSS.n2377 VSS.n2376 0.00404331
R69630 VSS.n11346 VSS.n11345 0.00404331
R69631 VSS.n5851 VSS.n5850 0.00404331
R69632 VSS.n13147 VSS.n13146 0.00404331
R69633 VSS.n13189 VSS.n13188 0.00404331
R69634 VSS.n12863 VSS.n12862 0.00404331
R69635 VSS.n12800 VSS.n12799 0.00404331
R69636 VSS.n12677 VSS.n12676 0.00404331
R69637 VSS.n12587 VSS.n12586 0.00404331
R69638 VSS.n11836 VSS.n11835 0.00404331
R69639 VSS.n2238 VSS.n2237 0.00404331
R69640 VSS.n2276 VSS.n2275 0.00404331
R69641 VSS.n15147 VSS.n15146 0.00404331
R69642 VSS.n16212 VSS.n16211 0.00404331
R69643 VSS.n2287 VSS.n2286 0.00404331
R69644 VSS.n2329 VSS.n2328 0.00404331
R69645 VSS.n20797 VSS.n20796 0.00404331
R69646 VSS.n21154 VSS.n21153 0.00404331
R69647 VSS.n17895 VSS.n17894 0.00404331
R69648 VSS.n17937 VSS.n17936 0.00404331
R69649 VSS.n2022 VSS.n2021 0.00404331
R69650 VSS.n1283 VSS.n1282 0.00404331
R69651 VSS.n21484 VSS.n21483 0.00404331
R69652 VSS.n21284 VSS.n21283 0.00404331
R69653 VSS.n7545 VSS.n7544 0.00404331
R69654 VSS.n7562 VSS.n7561 0.00404331
R69655 VSS.n3852 VSS.n3851 0.00404331
R69656 VSS.n4730 VSS.n4729 0.00404331
R69657 VSS.n11442 VSS.n11441 0.00404331
R69658 VSS.n11221 VSS.n11220 0.00404331
R69659 VSS.n560 VSS.n559 0.00404331
R69660 VSS.n501 VSS.n500 0.00404331
R69661 VSS.n10545 VSS.n10544 0.00404331
R69662 VSS.n10522 VSS.n10521 0.00404331
R69663 VSS.n8909 VSS.n8908 0.00404331
R69664 VSS.n7906 VSS.n7905 0.00404
R69665 VSS.n7999 VSS.n7998 0.00404
R69666 VSS.n11030 VSS.n11028 0.00404
R69667 VSS.n2847 VSS.n2846 0.00403571
R69668 VSS.n7165 VSS.n7164 0.00403571
R69669 VSS.n7106 VSS.n7105 0.00403571
R69670 VSS.n18050 VSS.n18049 0.00403571
R69671 VSS.n15393 VSS.n15392 0.0040341
R69672 VSS.n1709 VSS.n1708 0.0040341
R69673 VSS.n151 VSS.n149 0.00401955
R69674 VSS.n127 VSS.n126 0.00401955
R69675 VSS.n119 VSS.n118 0.00401955
R69676 VSS.n96 VSS.n95 0.00401955
R69677 VSS.n88 VSS.n86 0.00401955
R69678 VSS.n64 VSS.n63 0.00401955
R69679 VSS.n229 VSS.n228 0.00401955
R69680 VSS.n254 VSS.n251 0.00401955
R69681 VSS.n261 VSS.n260 0.00401955
R69682 VSS.n286 VSS.n283 0.00401955
R69683 VSS.n293 VSS.n292 0.00401955
R69684 VSS.n317 VSS.n315 0.00401955
R69685 VSS.n3973 VSS.n3972 0.00397904
R69686 VSS.n2607 VSS.n2606 0.00397904
R69687 VSS.n2516 VSS.n2515 0.00397222
R69688 VSS.n4119 VSS.n3941 0.00397222
R69689 VSS.n17591 VSS.n17589 0.00397143
R69690 VSS.n1634 VSS.n1633 0.0039558
R69691 VSS.n1635 VSS.n1634 0.0039558
R69692 VSS.n8533 VSS.n8532 0.0039558
R69693 VSS.n8388 VSS.n8387 0.0039558
R69694 VSS.n8389 VSS.n8388 0.0039558
R69695 VSS.n8534 VSS.n8533 0.0039558
R69696 VSS.n8684 VSS.n8683 0.0039558
R69697 VSS.n8196 VSS.n8195 0.0039558
R69698 VSS.n8685 VSS.n8684 0.0039558
R69699 VSS.n8197 VSS.n8196 0.0039558
R69700 VSS.n4199 VSS.n4198 0.00395082
R69701 VSS.n5837 VSS.n5749 0.00395082
R69702 VSS.n17347 VSS.n17346 0.00395082
R69703 VSS.n17330 VSS.n17329 0.00395082
R69704 VSS.n11519 VSS.n11518 0.00395082
R69705 VSS.n11327 VSS.n11326 0.00395082
R69706 VSS.n11316 VSS.n11315 0.00395082
R69707 VSS.n16356 VSS.n16327 0.00395082
R69708 VSS.n16311 VSS.n16292 0.00395082
R69709 VSS.n16276 VSS.n16256 0.00395082
R69710 VSS.n1437 VSS.n1408 0.00395082
R69711 VSS.n1392 VSS.n1373 0.00395082
R69712 VSS.n1357 VSS.n1337 0.00395082
R69713 VSS.n1269 VSS.n1189 0.00395082
R69714 VSS.n1152 VSS.n1141 0.00395082
R69715 VSS.n3218 VSS.n3217 0.0039507
R69716 VSS.n13237 VSS.n13236 0.00392323
R69717 VSS.n13354 VSS.n13353 0.00392323
R69718 VSS.n13497 VSS.n13496 0.00392323
R69719 VSS.n14157 VSS.n14156 0.0039231
R69720 VSS.n14199 VSS.n14198 0.0039231
R69721 VSS.n20517 DVSS 0.00392
R69722 VSS.n20552 DVSS 0.00392
R69723 VSS.n11077 DVSS 0.00392
R69724 DVSS VSS.n11074 0.00392
R69725 VSS.n3677 DVSS 0.00391158
R69726 VSS.n2673 VSS.n2672 0.00390714
R69727 VSS.n2717 VSS.n2716 0.00390714
R69728 VSS.n2777 VSS.n2776 0.00390714
R69729 VSS.n2872 VSS.n2871 0.00390714
R69730 VSS.n5147 VSS.n5146 0.00390714
R69731 VSS.n4508 VSS.n4507 0.00390714
R69732 VSS.n17552 VSS.n17551 0.00390714
R69733 VSS.n17494 VSS.n17493 0.00390714
R69734 VSS.n18027 VSS.n18026 0.00390714
R69735 VSS.n11852 VSS.n11851 0.00389099
R69736 VSS.n12268 VSS.n12267 0.00389055
R69737 VSS.n18800 VSS.n18799 0.00388028
R69738 VSS.n18475 VSS.n18474 0.00388028
R69739 VSS.n18400 VSS.n18399 0.00388028
R69740 VSS.n18162 VSS.n18161 0.00388028
R69741 VSS.n14573 VSS.n14572 0.00388028
R69742 VSS.n14822 VSS.n14821 0.00388028
R69743 VSS.n14866 VSS.n14865 0.00388028
R69744 VSS.n16895 VSS.n16894 0.00388028
R69745 VSS.n16697 VSS.n16696 0.00388028
R69746 VSS.n16535 VSS.n16534 0.00388028
R69747 VSS.n16446 VSS.n16445 0.00388028
R69748 VSS.n15863 VSS.n15862 0.00388028
R69749 VSS.n8521 VSS.n8520 0.00388028
R69750 VSS.n8339 VSS.n8338 0.00388028
R69751 VSS.n19472 VSS.n19471 0.00388028
R69752 VSS.n19564 VSS.n19563 0.00388028
R69753 VSS.n19622 VSS.n19621 0.00388028
R69754 VSS.n19694 VSS.n19693 0.00388028
R69755 VSS.n19755 VSS.n19754 0.00388028
R69756 VSS.n19845 VSS.n19844 0.00388028
R69757 VSS.n19937 VSS.n19936 0.00388028
R69758 VSS.n20021 VSS.n20020 0.00388028
R69759 VSS.n2099 VSS.n2098 0.00388028
R69760 VSS.n803 VSS.n802 0.00388028
R69761 VSS.n843 VSS.n842 0.00388028
R69762 VSS.n1937 VSS.n1936 0.00388028
R69763 VSS.n8672 VSS.n8671 0.00388028
R69764 VSS.n8135 VSS.n8134 0.00388028
R69765 VSS.n19239 VSS.n19238 0.003875
R69766 VSS.n18658 VSS.n18657 0.003875
R69767 VSS.n16857 VSS.n16856 0.003875
R69768 VSS.n19773 VSS.n19772 0.003875
R69769 VSS.n14462 VSS.n14461 0.003875
R69770 VSS.n17133 VSS.n17132 0.003875
R69771 VSS.n17106 VSS.n17105 0.003875
R69772 VSS.n17055 VSS.n17053 0.003875
R69773 VSS.n16956 VSS.n16955 0.003875
R69774 VSS.n14918 VSS.n14915 0.003875
R69775 VSS.n16668 VSS.n16667 0.003875
R69776 VSS.n15707 VSS.n15706 0.003875
R69777 VSS.n3961 VSS.n3960 0.00386614
R69778 VSS.n11527 VSS.n11526 0.00386614
R69779 VSS.n5596 VSS.n5595 0.00386614
R69780 VSS.n9592 VSS.n9591 0.00386614
R69781 VSS.n9155 VSS.n9154 0.00386614
R69782 VSS.n12977 VSS.n12976 0.00386614
R69783 VSS.n12759 VSS.n12758 0.00386614
R69784 VSS.n12687 VSS.n12686 0.00386614
R69785 VSS.n12234 VSS.n12233 0.00386614
R69786 VSS.n11970 VSS.n11969 0.00386614
R69787 VSS.n11891 VSS.n11890 0.00386614
R69788 VSS.n11855 VSS.n11854 0.00386614
R69789 VSS.n18964 VSS.n18963 0.00386614
R69790 VSS.n15001 VSS.n15000 0.00386614
R69791 VSS.n16112 VSS.n16111 0.00386614
R69792 VSS.n9709 VSS.n9708 0.00386614
R69793 VSS.n9318 VSS.n9317 0.00386614
R69794 VSS.n20607 VSS.n20606 0.00386614
R69795 VSS.n21046 VSS.n21045 0.00386614
R69796 VSS.n7004 VSS.n7003 0.00386614
R69797 VSS.n6644 VSS.n6643 0.00386614
R69798 VSS.n20142 VSS.n20141 0.00386614
R69799 VSS.n1092 VSS.n1091 0.00386614
R69800 VSS.n6902 VSS.n6901 0.00386614
R69801 VSS.n6494 VSS.n6493 0.00386614
R69802 VSS.n21626 VSS.n21625 0.00386614
R69803 VSS.n21646 VSS.n21645 0.00386614
R69804 VSS.n21529 VSS.n21528 0.00386614
R69805 VSS.n21394 VSS.n21393 0.00386614
R69806 VSS.n7603 VSS.n7602 0.00386614
R69807 VSS.n7691 VSS.n7690 0.00386614
R69808 VSS.n7848 VSS.n7847 0.00386614
R69809 VSS.n3854 VSS.n3853 0.00386614
R69810 VSS.n3875 VSS.n3874 0.00386614
R69811 VSS.n4146 VSS.n4145 0.00386614
R69812 VSS.n11708 VSS.n11707 0.00386614
R69813 VSS.n6151 VSS.n6150 0.00386614
R69814 VSS.n6070 VSS.n6069 0.00386614
R69815 VSS.n5989 VSS.n5988 0.00386614
R69816 VSS.n2595 VSS.n2594 0.00386614
R69817 VSS.n665 VSS.n664 0.00386614
R69818 VSS.n10623 VSS.n10622 0.00386614
R69819 VSS.n10555 VSS.n10554 0.00386614
R69820 VSS.n10182 VSS.n10181 0.00386614
R69821 VSS.n9973 VSS.n9972 0.00386614
R69822 VSS.n8982 VSS.n8981 0.00386614
R69823 VSS.n8795 VSS.n8794 0.00386614
R69824 VSS.n5691 VSS.n5689 0.00385106
R69825 VSS.n5670 VSS.n5669 0.00385106
R69826 VSS.n16013 VSS.n16012 0.00385106
R69827 VSS.n16025 VSS.n16020 0.00385106
R69828 VSS.n994 VSS.n993 0.00385106
R69829 VSS.n985 VSS.n984 0.00385106
R69830 VSS.n20939 VSS.n20938 0.00385106
R69831 VSS.n20960 VSS.n20958 0.00385106
R69832 VSS.n5771 VSS.n5770 0.00385106
R69833 VSS.n5823 VSS.n5822 0.00385106
R69834 VSS.n5812 VSS.n5811 0.00385106
R69835 VSS.n15482 VSS.n15479 0.00385106
R69836 VSS.n1195 VSS.n1194 0.00385106
R69837 VSS.n1253 VSS.n1252 0.00385106
R69838 VSS.n1223 VSS.n1222 0.00385106
R69839 VSS.n18818 VSS.n18817 0.00385031
R69840 VSS.n16888 VSS.n16887 0.00385031
R69841 VSS.n15361 VSS.n15360 0.00385031
R69842 VSS.n8563 VSS.n8562 0.00385031
R69843 VSS.n8330 VSS.n8329 0.00385031
R69844 VSS.n8418 VSS.n8417 0.00385031
R69845 VSS.n16546 VSS.n16545 0.00385031
R69846 VSS.n16887 VSS.n16886 0.00385031
R69847 VSS.n8419 VSS.n8418 0.00385031
R69848 VSS.n8564 VSS.n8563 0.00385031
R69849 VSS.n8329 VSS.n8328 0.00385031
R69850 VSS.n15362 VSS.n15361 0.00385031
R69851 VSS.n19491 VSS.n19490 0.00385031
R69852 VSS.n20028 VSS.n20027 0.00385031
R69853 VSS.n1678 VSS.n1677 0.00385031
R69854 VSS.n8714 VSS.n8713 0.00385031
R69855 VSS.n8126 VSS.n8125 0.00385031
R69856 VSS.n8226 VSS.n8225 0.00385031
R69857 VSS.n8715 VSS.n8714 0.00385031
R69858 VSS.n8227 VSS.n8226 0.00385031
R69859 VSS.n8125 VSS.n8124 0.00385031
R69860 VSS.n1677 VSS.n1676 0.00385031
R69861 VSS.n792 VSS.n791 0.00385031
R69862 VSS.n20029 VSS.n20028 0.00385031
R69863 VSS.n19490 VSS.n19489 0.00385031
R69864 VSS.n18819 VSS.n18818 0.00385031
R69865 VSS.n2947 VSS.n2946 0.00384286
R69866 VSS.n3012 VSS.n3011 0.00384286
R69867 VSS.n3060 VSS.n3059 0.00384286
R69868 VSS.n17577 VSS.n17576 0.00384286
R69869 VSS.n17863 VSS.n17862 0.00384286
R69870 VSS.n17802 VSS.n17801 0.00384286
R69871 VSS.n17757 VSS.n17756 0.00384286
R69872 VSS.n13101 VSS.n13100 0.00383286
R69873 VSS.n13212 VSS.n13211 0.00383286
R69874 VSS.n21873 VSS.n21776 0.00383286
R69875 VSS.n19158 VSS.n19061 0.00383286
R69876 VSS.n1440 VSS.n1439 0.00383286
R69877 VSS.n1395 VSS.n1394 0.00383286
R69878 VSS.n1360 VSS.n1359 0.00383286
R69879 VSS.n1155 VSS.n1154 0.00383286
R69880 VSS.n2614 VSS.n2613 0.00383286
R69881 VSS.n4073 VSS.n3979 0.00383286
R69882 VSS.n18945 VSS.n18944 0.00383286
R69883 VSS.n12237 VSS.n12236 0.00380239
R69884 VSS.n10167 VSS.n10166 0.00380234
R69885 VSS.n11823 VSS.n11822 0.00380214
R69886 VSS.n4780 VSS.n4779 0.00380206
R69887 VSS.n10885 VSS.n10884 0.0038
R69888 VSS.n10880 VSS.n10879 0.0038
R69889 VSS.n6784 VSS.n6783 0.0038
R69890 VSS.n8100 VSS.n8099 0.0038
R69891 VSS.n10910 VSS.n10905 0.0038
R69892 VSS.n20261 VSS.n20260 0.00377
R69893 VSS.n9876 VSS.n9875 0.00376923
R69894 VSS.n9883 VSS.n9878 0.00376923
R69895 VSS.n10378 VSS.n10377 0.00376923
R69896 VSS.n10369 VSS.n10364 0.00376923
R69897 VSS.n10093 VSS.n10092 0.00376923
R69898 VSS.n10084 VSS.n10079 0.00376923
R69899 VSS.n10001 VSS.n10000 0.00376923
R69900 VSS.n9992 VSS.n9987 0.00376923
R69901 VSS.n11777 VSS.n11776 0.00376923
R69902 VSS.n11784 VSS.n11779 0.00376923
R69903 VSS.n12432 VSS.n12431 0.00376923
R69904 VSS.n12423 VSS.n12418 0.00376923
R69905 VSS.n12144 VSS.n12143 0.00376923
R69906 VSS.n12135 VSS.n12130 0.00376923
R69907 VSS.n12052 VSS.n12051 0.00376923
R69908 VSS.n12043 VSS.n12038 0.00376923
R69909 VSS.n13207 VSS.n13206 0.00374606
R69910 VSS.n13324 VSS.n13323 0.00374606
R69911 VSS.n17944 VSS.n17943 0.00374606
R69912 VSS.n5566 VSS.n5565 0.00374577
R69913 VSS.n16082 VSS.n16081 0.00374577
R69914 VSS.n21015 VSS.n21014 0.00374577
R69915 VSS.n1061 VSS.n1060 0.00374577
R69916 VSS.n18466 VSS.n18465 0.0037448
R69917 VSS.n18143 VSS.n18142 0.0037448
R69918 VSS.n15544 VSS.n15543 0.0037448
R69919 VSS.n8358 VSS.n8357 0.0037448
R69920 VSS.n18467 VSS.n18466 0.0037448
R69921 VSS.n14903 VSS.n14902 0.0037448
R69922 VSS.n18142 VSS.n18141 0.0037448
R69923 VSS.n15545 VSS.n15544 0.0037448
R69924 VSS.n8359 VSS.n8358 0.0037448
R69925 VSS.n19573 VSS.n19572 0.0037448
R69926 VSS.n19713 VSS.n19712 0.0037448
R69927 VSS.n19974 VSS.n19973 0.0037448
R69928 VSS.n1833 VSS.n1832 0.0037448
R69929 VSS.n8166 VSS.n8165 0.0037448
R69930 VSS.n8167 VSS.n8166 0.0037448
R69931 VSS.n19572 VSS.n19571 0.0037448
R69932 VSS.n19714 VSS.n19713 0.0037448
R69933 VSS.n1832 VSS.n1831 0.0037448
R69934 VSS.n15311 VSS.n15306 0.00374324
R69935 VSS.n15315 VSS.n15313 0.00374324
R69936 VSS.n1629 VSS.n1624 0.00374324
R69937 VSS.n1618 VSS.n1616 0.00374324
R69938 VSS.n20203 VSS.n20202 0.00371
R69939 VSS.n14187 VSS.n14186 0.00369838
R69940 VSS.n4056 VSS.n4055 0.00368898
R69941 VSS.n4070 VSS.n4069 0.00368898
R69942 VSS.n11555 VSS.n11554 0.00368898
R69943 VSS.n11571 VSS.n11570 0.00368898
R69944 VSS.n9564 VSS.n9563 0.00368898
R69945 VSS.n9018 VSS.n9017 0.00368898
R69946 VSS.n9127 VSS.n9126 0.00368898
R69947 VSS.n9111 VSS.n9110 0.00368898
R69948 VSS.n13085 VSS.n13084 0.00368898
R69949 VSS.n12947 VSS.n12946 0.00368898
R69950 VSS.n12928 VSS.n12927 0.00368898
R69951 VSS.n12729 VSS.n12728 0.00368898
R69952 VSS.n12711 VSS.n12710 0.00368898
R69953 VSS.n12679 VSS.n12678 0.00368898
R69954 VSS.n12528 VSS.n12527 0.00368898
R69955 VSS.n12255 VSS.n12254 0.00368898
R69956 VSS.n11879 VSS.n11878 0.00368898
R69957 VSS.n11845 VSS.n11844 0.00368898
R69958 VSS.n18927 VSS.n18926 0.00368898
R69959 VSS.n18941 VSS.n18940 0.00368898
R69960 VSS.n15029 VSS.n15028 0.00368898
R69961 VSS.n15046 VSS.n15045 0.00368898
R69962 VSS.n16049 VSS.n16048 0.00368898
R69963 VSS.n9681 VSS.n9680 0.00368898
R69964 VSS.n9161 VSS.n9160 0.00368898
R69965 VSS.n9290 VSS.n9289 0.00368898
R69966 VSS.n9274 VSS.n9273 0.00368898
R69967 VSS.n21858 VSS.n21857 0.00368898
R69968 VSS.n20637 VSS.n20636 0.00368898
R69969 VSS.n20656 VSS.n20655 0.00368898
R69970 VSS.n6908 VSS.n6907 0.00368898
R69971 VSS.n6974 VSS.n6973 0.00368898
R69972 VSS.n6649 VSS.n6648 0.00368898
R69973 VSS.n6614 VSS.n6613 0.00368898
R69974 VSS.n6595 VSS.n6594 0.00368898
R69975 VSS.n19143 VSS.n19142 0.00368898
R69976 VSS.n20112 VSS.n20111 0.00368898
R69977 VSS.n20093 VSS.n20092 0.00368898
R69978 VSS.n6872 VSS.n6871 0.00368898
R69979 VSS.n6499 VSS.n6498 0.00368898
R69980 VSS.n6464 VSS.n6463 0.00368898
R69981 VSS.n6445 VSS.n6444 0.00368898
R69982 VSS.n21440 VSS.n21439 0.00368898
R69983 VSS.n21439 VSS.n21438 0.00368898
R69984 VSS.n21364 VSS.n21363 0.00368898
R69985 VSS.n21345 VSS.n21344 0.00368898
R69986 VSS.n7633 VSS.n7632 0.00368898
R69987 VSS.n7652 VSS.n7651 0.00368898
R69988 VSS.n7721 VSS.n7720 0.00368898
R69989 VSS.n7740 VSS.n7739 0.00368898
R69990 VSS.n7818 VSS.n7817 0.00368898
R69991 VSS.n7799 VSS.n7798 0.00368898
R69992 VSS.n4769 VSS.n4768 0.00368898
R69993 VSS.n4795 VSS.n4794 0.00368898
R69994 VSS.n4796 VSS.n4795 0.00368898
R69995 VSS.n11680 VSS.n11679 0.00368898
R69996 VSS.n11663 VSS.n11662 0.00368898
R69997 VSS.n6123 VSS.n6122 0.00368898
R69998 VSS.n6107 VSS.n6106 0.00368898
R69999 VSS.n6042 VSS.n6041 0.00368898
R70000 VSS.n6026 VSS.n6025 0.00368898
R70001 VSS.n5961 VSS.n5960 0.00368898
R70002 VSS.n5945 VSS.n5944 0.00368898
R70003 VSS.n2632 VSS.n2631 0.00368898
R70004 VSS.n2618 VSS.n2617 0.00368898
R70005 VSS.n637 VSS.n636 0.00368898
R70006 VSS.n621 VSS.n620 0.00368898
R70007 VSS.n10595 VSS.n10594 0.00368898
R70008 VSS.n10579 VSS.n10578 0.00368898
R70009 VSS.n10547 VSS.n10546 0.00368898
R70010 VSS.n10473 VSS.n10472 0.00368898
R70011 VSS.n10203 VSS.n10202 0.00368898
R70012 VSS.n8941 VSS.n8940 0.00368898
R70013 VSS.n9004 VSS.n9003 0.00368898
R70014 VSS.n174 VSS.n171 0.00368083
R70015 VSS.n5898 VSS.n5897 0.00368083
R70016 VSS.n3213 VSS.n3197 0.00366901
R70017 VSS.n3301 VSS.n3300 0.00366901
R70018 VSS.n3339 VSS.n3338 0.00366901
R70019 VSS.n3393 VSS.n3392 0.00366901
R70020 VSS.n3520 VSS.n3519 0.00366901
R70021 VSS.n3579 VSS.n3578 0.00366901
R70022 VSS.n3622 VSS.n3621 0.00366901
R70023 VSS.n18724 VSS.n18723 0.00366901
R70024 VSS.n18669 VSS.n18668 0.00366901
R70025 VSS.n18459 VSS.n18458 0.00366901
R70026 VSS.n18424 VSS.n18423 0.00366901
R70027 VSS.n14459 VSS.n14458 0.00366901
R70028 VSS.n14673 VSS.n14672 0.00366901
R70029 VSS.n17163 VSS.n17162 0.00366901
R70030 VSS.n17076 VSS.n17075 0.00366901
R70031 VSS.n17023 VSS.n17022 0.00366901
R70032 VSS.n17022 VSS.n17021 0.00366901
R70033 VSS.n16926 VSS.n16925 0.00366901
R70034 VSS.n16871 VSS.n16870 0.00366901
R70035 VSS.n16682 VSS.n16681 0.00366901
R70036 VSS.n16533 VSS.n16532 0.00366901
R70037 VSS.n15704 VSS.n15703 0.00366901
R70038 VSS.n15463 VSS.n15462 0.00366901
R70039 VSS.n19206 VSS.n19205 0.00366901
R70040 VSS.n19534 VSS.n19533 0.00366901
R70041 VSS.n19580 VSS.n19579 0.00366901
R70042 VSS.n19605 VSS.n19604 0.00366901
R70043 VSS.n19725 VSS.n19724 0.00366901
R70044 VSS.n19770 VSS.n19769 0.00366901
R70045 VSS.n19860 VSS.n19859 0.00366901
R70046 VSS.n19889 VSS.n19888 0.00366901
R70047 VSS.n19912 VSS.n19911 0.00366901
R70048 VSS.n19913 VSS.n19912 0.00366901
R70049 VSS.n19990 VSS.n19989 0.00366901
R70050 VSS.n2129 VSS.n2128 0.00366901
R70051 VSS.n750 VSS.n749 0.00366901
R70052 VSS.n805 VSS.n804 0.00366901
R70053 VSS.n1967 VSS.n1966 0.00366901
R70054 VSS.n1765 VSS.n1764 0.00366901
R70055 VSS.n19402 VSS.n19400 0.00365
R70056 VSS.n18264 VSS.n18263 0.00365
R70057 VSS.n18250 VSS.n18249 0.00365
R70058 VSS.n18247 VSS.n18246 0.00365
R70059 VSS.n16660 VSS.n16658 0.00365
R70060 VSS.n16618 VSS.n16617 0.00365
R70061 VSS.n3182 VSS.n2544 0.00365
R70062 VSS.n20524 VSS.n20523 0.00365
R70063 VSS.n4686 VSS.n4684 0.00365
R70064 VSS.n17603 VSS.n17602 0.00365
R70065 VSS.n8444 VSS.n8443 0.00365
R70066 VSS.n8776 VSS.n8775 0.00365
R70067 VSS.n10805 VSS.n10804 0.00365
R70068 VSS.n7517 DVSS 0.00364286
R70069 VSS.n16938 VSS.n16937 0.00364043
R70070 VSS.n19978 VSS.n19977 0.00364043
R70071 VSS.n16525 VSS.n16524 0.00363995
R70072 VSS.n813 VSS.n812 0.00363995
R70073 VSS.n18697 VSS.n18696 0.0036393
R70074 VSS.n18460 VSS.n18459 0.0036393
R70075 VSS.n18155 VSS.n18154 0.0036393
R70076 VSS.n15632 VSS.n15631 0.0036393
R70077 VSS.n15609 VSS.n15608 0.0036393
R70078 VSS.n15586 VSS.n15585 0.0036393
R70079 VSS.n15453 VSS.n15452 0.0036393
R70080 VSS.n15411 VSS.n15410 0.0036393
R70081 VSS.n15454 VSS.n15453 0.0036393
R70082 VSS.n15587 VSS.n15586 0.0036393
R70083 VSS.n15610 VSS.n15609 0.0036393
R70084 VSS.n15633 VSS.n15632 0.0036393
R70085 VSS.n14882 VSS.n14881 0.0036393
R70086 VSS.n18698 VSS.n18697 0.0036393
R70087 VSS.n15412 VSS.n15411 0.0036393
R70088 VSS.n19180 VSS.n19179 0.0036393
R70089 VSS.n19579 VSS.n19578 0.0036393
R70090 VSS.n19701 VSS.n19700 0.0036393
R70091 VSS.n1900 VSS.n1899 0.0036393
R70092 VSS.n1883 VSS.n1882 0.0036393
R70093 VSS.n1866 VSS.n1865 0.0036393
R70094 VSS.n1755 VSS.n1754 0.0036393
R70095 VSS.n1727 VSS.n1726 0.0036393
R70096 VSS.n1756 VSS.n1755 0.0036393
R70097 VSS.n19953 VSS.n19952 0.0036393
R70098 VSS.n1901 VSS.n1900 0.0036393
R70099 VSS.n1884 VSS.n1883 0.0036393
R70100 VSS.n1867 VSS.n1866 0.0036393
R70101 VSS.n19179 VSS.n19178 0.0036393
R70102 VSS.n1728 VSS.n1727 0.0036393
R70103 VSS.n18156 VSS.n18155 0.0036393
R70104 VSS.n19578 VSS.n19577 0.0036393
R70105 VSS.n18461 VSS.n18460 0.0036393
R70106 VSS.n19700 VSS.n19699 0.0036393
R70107 VSS.n1229 VSS.n1228 0.00363144
R70108 VSS.n1230 VSS.n1229 0.00363144
R70109 VSS.n21564 VSS.n21563 0.00362543
R70110 VSS.n3665 VSS.n3664 0.00359859
R70111 VSS.n10787 VSS.n10786 0.00356
R70112 VSS.n10782 VSS.n10781 0.00356
R70113 VSS.n10771 VSS.n10770 0.00356
R70114 VSS.n8453 VSS.n8452 0.00356
R70115 VSS.n8785 VSS.n8784 0.00356
R70116 VSS.n10791 VSS.n10790 0.00356
R70117 VSS.n21696 VSS.n21692 0.00355556
R70118 VSS.n441 VSS.n437 0.00355556
R70119 VSS.n424 VSS.n420 0.00355556
R70120 VSS.n407 VSS.n403 0.00355556
R70121 VSS.n14289 VSS.n14288 0.00355556
R70122 VSS.n389 VSS.n385 0.00355556
R70123 VSS.n363 VSS.n359 0.00355556
R70124 VSS.n21930 VSS.n21924 0.00355556
R70125 VSS.n16532 VSS.n16531 0.0035352
R70126 VSS.n806 VSS.n805 0.0035352
R70127 VSS.n18752 VSS.n18751 0.00353378
R70128 VSS.n18821 VSS.n18820 0.00353378
R70129 VSS.n18831 VSS.n18830 0.00353378
R70130 VSS.n18682 VSS.n18681 0.00353378
R70131 VSS.n18673 VSS.n18672 0.00353378
R70132 VSS.n18462 VSS.n18461 0.00353378
R70133 VSS.n18157 VSS.n18156 0.00353378
R70134 VSS.n15656 VSS.n15655 0.00353378
R70135 VSS.n15629 VSS.n15628 0.00353378
R70136 VSS.n15606 VSS.n15605 0.00353378
R70137 VSS.n15445 VSS.n15444 0.00353378
R70138 VSS.n8355 VSS.n8354 0.00353378
R70139 VSS.n16913 VSS.n16912 0.00353378
R70140 VSS.n15657 VSS.n15656 0.00353378
R70141 VSS.n15630 VSS.n15629 0.00353378
R70142 VSS.n15607 VSS.n15606 0.00353378
R70143 VSS.n18158 VSS.n18157 0.00353378
R70144 VSS.n18463 VSS.n18462 0.00353378
R70145 VSS.n18751 VSS.n18750 0.00353378
R70146 VSS.n15446 VSS.n15445 0.00353378
R70147 VSS.n19234 VSS.n19233 0.00353378
R70148 VSS.n19493 VSS.n19492 0.00353378
R70149 VSS.n19503 VSS.n19502 0.00353378
R70150 VSS.n19521 VSS.n19520 0.00353378
R70151 VSS.n19530 VSS.n19529 0.00353378
R70152 VSS.n19577 VSS.n19576 0.00353378
R70153 VSS.n19699 VSS.n19698 0.00353378
R70154 VSS.n1914 VSS.n1913 0.00353378
R70155 VSS.n1897 VSS.n1896 0.00353378
R70156 VSS.n1880 VSS.n1879 0.00353378
R70157 VSS.n1747 VSS.n1746 0.00353378
R70158 VSS.n8162 VSS.n8161 0.00353378
R70159 VSS.n8163 VSS.n8162 0.00353378
R70160 VSS.n1748 VSS.n1747 0.00353378
R70161 VSS.n20003 VSS.n20002 0.00353378
R70162 VSS.n1915 VSS.n1914 0.00353378
R70163 VSS.n1898 VSS.n1897 0.00353378
R70164 VSS.n1881 VSS.n1880 0.00353378
R70165 VSS.n19698 VSS.n19697 0.00353378
R70166 VSS.n19576 VSS.n19575 0.00353378
R70167 VSS.n19233 VSS.n19232 0.00353378
R70168 VSS.n19520 VSS.n19519 0.00353378
R70169 VSS.n18683 VSS.n18682 0.00353378
R70170 VSS.n18830 VSS.n18829 0.00353378
R70171 VSS.n19492 VSS.n19491 0.00353378
R70172 VSS.n18820 VSS.n18819 0.00353378
R70173 VSS.n19502 VSS.n19501 0.00353378
R70174 VSS.n19529 VSS.n19528 0.00353378
R70175 VSS.n18674 VSS.n18673 0.00353378
R70176 VSS.n8354 VSS.n8353 0.00353378
R70177 VSS.n8257 VSS.n8256 0.00353
R70178 VSS.n8594 VSS.n8593 0.00353
R70179 VSS.n10896 VSS.n10875 0.00353
R70180 VSS.n3300 VSS.n3298 0.00352817
R70181 VSS.n3338 VSS.n3336 0.00352817
R70182 VSS.n3392 VSS.n3390 0.00352817
R70183 VSS.n152 VSS.n151 0.00351676
R70184 VSS.n126 VSS.n123 0.00351676
R70185 VSS.n120 VSS.n119 0.00351676
R70186 VSS.n95 VSS.n92 0.00351676
R70187 VSS.n89 VSS.n88 0.00351676
R70188 VSS.n63 VSS.n60 0.00351676
R70189 VSS.n228 VSS.n226 0.00351676
R70190 VSS.n255 VSS.n254 0.00351676
R70191 VSS.n260 VSS.n258 0.00351676
R70192 VSS.n287 VSS.n286 0.00351676
R70193 VSS.n292 VSS.n290 0.00351676
R70194 VSS.n318 VSS.n317 0.00351676
R70195 VSS.n11544 VSS.n11543 0.00351181
R70196 VSS.n11582 VSS.n11581 0.00351181
R70197 VSS.n5579 VSS.n5578 0.00351181
R70198 VSS.n9488 VSS.n9487 0.00351181
R70199 VSS.n9575 VSS.n9574 0.00351181
R70200 VSS.n9029 VSS.n9028 0.00351181
R70201 VSS.n9138 VSS.n9137 0.00351181
R70202 VSS.n9100 VSS.n9099 0.00351181
R70203 VSS.n12958 VSS.n12957 0.00351181
R70204 VSS.n12917 VSS.n12916 0.00351181
R70205 VSS.n12740 VSS.n12739 0.00351181
R70206 VSS.n12700 VSS.n12699 0.00351181
R70207 VSS.n12578 VSS.n12577 0.00351181
R70208 VSS.n12520 VSS.n12519 0.00351181
R70209 VSS.n12293 VSS.n12292 0.00351181
R70210 VSS.n12264 VSS.n12263 0.00351181
R70211 VSS.n12246 VSS.n12245 0.00351181
R70212 VSS.n11910 VSS.n11909 0.00351181
R70213 VSS.n11827 VSS.n11826 0.00351181
R70214 VSS.n15018 VSS.n15017 0.00351181
R70215 VSS.n15057 VSS.n15056 0.00351181
R70216 VSS.n16095 VSS.n16094 0.00351181
R70217 VSS.n9605 VSS.n9604 0.00351181
R70218 VSS.n9692 VSS.n9691 0.00351181
R70219 VSS.n9172 VSS.n9171 0.00351181
R70220 VSS.n9301 VSS.n9300 0.00351181
R70221 VSS.n9263 VSS.n9262 0.00351181
R70222 VSS.n20626 VSS.n20625 0.00351181
R70223 VSS.n20667 VSS.n20666 0.00351181
R70224 VSS.n21027 VSS.n21026 0.00351181
R70225 VSS.n6919 VSS.n6918 0.00351181
R70226 VSS.n6985 VSS.n6984 0.00351181
R70227 VSS.n6660 VSS.n6659 0.00351181
R70228 VSS.n6625 VSS.n6624 0.00351181
R70229 VSS.n6584 VSS.n6583 0.00351181
R70230 VSS.n20123 VSS.n20122 0.00351181
R70231 VSS.n20082 VSS.n20081 0.00351181
R70232 VSS.n1073 VSS.n1072 0.00351181
R70233 VSS.n6796 VSS.n6795 0.00351181
R70234 VSS.n6883 VSS.n6882 0.00351181
R70235 VSS.n6510 VSS.n6509 0.00351181
R70236 VSS.n6475 VSS.n6474 0.00351181
R70237 VSS.n6434 VSS.n6433 0.00351181
R70238 VSS.n21375 VSS.n21374 0.00351181
R70239 VSS.n21334 VSS.n21333 0.00351181
R70240 VSS.n7622 VSS.n7621 0.00351181
R70241 VSS.n7663 VSS.n7662 0.00351181
R70242 VSS.n7710 VSS.n7709 0.00351181
R70243 VSS.n7751 VSS.n7750 0.00351181
R70244 VSS.n7829 VSS.n7828 0.00351181
R70245 VSS.n7788 VSS.n7787 0.00351181
R70246 VSS.n11691 VSS.n11690 0.00351181
R70247 VSS.n11652 VSS.n11651 0.00351181
R70248 VSS.n6134 VSS.n6133 0.00351181
R70249 VSS.n6096 VSS.n6095 0.00351181
R70250 VSS.n6053 VSS.n6052 0.00351181
R70251 VSS.n6015 VSS.n6014 0.00351181
R70252 VSS.n5972 VSS.n5971 0.00351181
R70253 VSS.n5934 VSS.n5933 0.00351181
R70254 VSS.n648 VSS.n647 0.00351181
R70255 VSS.n610 VSS.n609 0.00351181
R70256 VSS.n10606 VSS.n10605 0.00351181
R70257 VSS.n10568 VSS.n10567 0.00351181
R70258 VSS.n10513 VSS.n10512 0.00351181
R70259 VSS.n10465 VSS.n10464 0.00351181
R70260 VSS.n10241 VSS.n10240 0.00351181
R70261 VSS.n10212 VSS.n10211 0.00351181
R70262 VSS.n10195 VSS.n10194 0.00351181
R70263 VSS.n9911 VSS.n9910 0.00351181
R70264 VSS.n8987 VSS.n8986 0.00351181
R70265 VSS.n11563 VSS.n11562 0.00347895
R70266 VSS.n12937 VSS.n12936 0.00347895
R70267 VSS.n12938 VSS.n12937 0.00347895
R70268 VSS.n15038 VSS.n15037 0.00347895
R70269 VSS.n15037 VSS.n15036 0.00347895
R70270 VSS.n20647 VSS.n20646 0.00347895
R70271 VSS.n20991 VSS.n20990 0.00347895
R70272 VSS.n6964 VSS.n6963 0.00347895
R70273 VSS.n6604 VSS.n6603 0.00347895
R70274 VSS.n20646 VSS.n20645 0.00347895
R70275 VSS.n20102 VSS.n20101 0.00347895
R70276 VSS.n1033 VSS.n1032 0.00347895
R70277 VSS.n6862 VSS.n6861 0.00347895
R70278 VSS.n6454 VSS.n6453 0.00347895
R70279 VSS.n20103 VSS.n20102 0.00347895
R70280 VSS.n21354 VSS.n21353 0.00347895
R70281 VSS.n7643 VSS.n7642 0.00347895
R70282 VSS.n7731 VSS.n7730 0.00347895
R70283 VSS.n7808 VSS.n7807 0.00347895
R70284 VSS.n21355 VSS.n21354 0.00347895
R70285 VSS.n9282 VSS.n9281 0.00347895
R70286 VSS.n7809 VSS.n7808 0.00347895
R70287 VSS.n9119 VSS.n9118 0.00347895
R70288 VSS.n6605 VSS.n6604 0.00347895
R70289 VSS.n6455 VSS.n6454 0.00347895
R70290 VSS.n9673 VSS.n9672 0.00347895
R70291 VSS.n7730 VSS.n7729 0.00347895
R70292 VSS.n9556 VSS.n9555 0.00347895
R70293 VSS.n6965 VSS.n6964 0.00347895
R70294 VSS.n6863 VSS.n6862 0.00347895
R70295 VSS.n5547 VSS.n5546 0.00347895
R70296 VSS.n7642 VSS.n7641 0.00347895
R70297 VSS.n16057 VSS.n16056 0.00347895
R70298 VSS.n1032 VSS.n1031 0.00347895
R70299 VSS.n20990 VSS.n20989 0.00347895
R70300 VSS.n11671 VSS.n11670 0.00347895
R70301 VSS.n11672 VSS.n11671 0.00347895
R70302 VSS.n6115 VSS.n6114 0.00347895
R70303 VSS.n6034 VSS.n6033 0.00347895
R70304 VSS.n5953 VSS.n5952 0.00347895
R70305 VSS.n10587 VSS.n10586 0.00347895
R70306 VSS.n629 VSS.n628 0.00347895
R70307 VSS.n14142 VSS.n14141 0.00347364
R70308 VSS.n20385 VSS.n20383 0.00347
R70309 VSS.n20354 VSS.n20353 0.00347
R70310 VSS.n20308 VSS.n20306 0.00347
R70311 VSS.n8829 VSS.n8828 0.00347
R70312 VSS.n9442 VSS.n9441 0.00347
R70313 VSS.n9817 VSS.n9816 0.00347
R70314 VSS.n18748 VSS.n18747 0.00345775
R70315 VSS.n18783 VSS.n18782 0.00345775
R70316 VSS.n18179 VSS.n18178 0.00345775
R70317 VSS.n18177 VSS.n18176 0.00345775
R70318 VSS.n17128 VSS.n17127 0.00345775
R70319 VSS.n16929 VSS.n16928 0.00345775
R70320 VSS.n16642 VSS.n16641 0.00345775
R70321 VSS.n16595 VSS.n16594 0.00345775
R70322 VSS.n14993 VSS.n14992 0.00345775
R70323 VSS.n19230 VSS.n19229 0.00345775
R70324 VSS.n19455 VSS.n19454 0.00345775
R70325 VSS.n19677 VSS.n19676 0.00345775
R70326 VSS.n19679 VSS.n19678 0.00345775
R70327 VSS.n19867 VSS.n19866 0.00345775
R70328 VSS.n19987 VSS.n19986 0.00345775
R70329 VSS.n756 VSS.n755 0.00345775
R70330 VSS.n773 VSS.n772 0.00345775
R70331 VSS.n829 VSS.n828 0.00345775
R70332 VSS.n10500 VSS.n10499 0.00344838
R70333 VSS.n18687 VSS.n18686 0.00342827
R70334 VSS.n19517 VSS.n19516 0.00342827
R70335 VSS.n18688 VSS.n18687 0.00342827
R70336 VSS.n19516 VSS.n19515 0.00342827
R70337 VSS.n19437 DVSS 0.003425
R70338 VSS.n18564 DVSS 0.003425
R70339 VSS.n18302 DVSS 0.003425
R70340 VSS.n16763 DVSS 0.003425
R70341 VSS.n14807 DVSS 0.003425
R70342 DVSS VSS.n14587 0.003425
R70343 VSS.n17155 VSS.n17154 0.003425
R70344 VSS.n17154 VSS.n17152 0.003425
R70345 VSS.n16999 VSS.n16998 0.003425
R70346 VSS.n16998 VSS.n16996 0.003425
R70347 VSS.n16992 DVSS 0.003425
R70348 VSS.n16510 DVSS 0.003425
R70349 DVSS VSS.n15813 0.003425
R70350 VSS.n390 VSS.n389 0.00340612
R70351 VSS.n14289 VSS.n14282 0.00340612
R70352 VSS.n408 VSS.n407 0.00340612
R70353 VSS.n425 VSS.n424 0.00340612
R70354 VSS.n442 VSS.n441 0.00340612
R70355 VSS.n2543 VSS.n2542 0.00339286
R70356 VSS.n7354 VSS.n7352 0.00339286
R70357 VSS.n7300 VSS.n7298 0.00339286
R70358 VSS.n7178 VSS.n7177 0.00339286
R70359 VSS.n7119 VSS.n7118 0.00339286
R70360 VSS.n4690 VSS.n4689 0.00339286
R70361 VSS.n4753 VSS.n4752 0.00339286
R70362 VSS.n5604 VSS.n5603 0.00339173
R70363 VSS.n16120 VSS.n16119 0.00339173
R70364 VSS.n21054 VSS.n21053 0.00339173
R70365 VSS.n1100 VSS.n1099 0.00339173
R70366 VSS.n6946 VSS.n6945 0.00339144
R70367 VSS.n6844 VSS.n6843 0.00339144
R70368 VSS.n6933 VSS.n6932 0.00339064
R70369 VSS.n6810 VSS.n6809 0.00339064
R70370 VSS.n4050 VSS.n4049 0.00339046
R70371 VSS.n11590 VSS.n11589 0.00339046
R70372 VSS.n9037 VSS.n9036 0.00339046
R70373 VSS.n11536 VSS.n11535 0.00339046
R70374 VSS.n4049 VSS.n4048 0.00339046
R70375 VSS.n13079 VSS.n13078 0.00339046
R70376 VSS.n12967 VSS.n12966 0.00339046
R70377 VSS.n12908 VSS.n12907 0.00339046
R70378 VSS.n12749 VSS.n12748 0.00339046
R70379 VSS.n12907 VSS.n12906 0.00339046
R70380 VSS.n12968 VSS.n12967 0.00339046
R70381 VSS.n13078 VSS.n13077 0.00339046
R70382 VSS.n18921 VSS.n18920 0.00339046
R70383 VSS.n15065 VSS.n15064 0.00339046
R70384 VSS.n9180 VSS.n9179 0.00339046
R70385 VSS.n15010 VSS.n15009 0.00339046
R70386 VSS.n18920 VSS.n18919 0.00339046
R70387 VSS.n21852 VSS.n21851 0.00339046
R70388 VSS.n20617 VSS.n20616 0.00339046
R70389 VSS.n20676 VSS.n20675 0.00339046
R70390 VSS.n21036 VSS.n21035 0.00339046
R70391 VSS.n6994 VSS.n6993 0.00339046
R70392 VSS.n6670 VSS.n6669 0.00339046
R70393 VSS.n6634 VSS.n6633 0.00339046
R70394 VSS.n20616 VSS.n20615 0.00339046
R70395 VSS.n20677 VSS.n20676 0.00339046
R70396 VSS.n21851 VSS.n21850 0.00339046
R70397 VSS.n19137 VSS.n19136 0.00339046
R70398 VSS.n20132 VSS.n20131 0.00339046
R70399 VSS.n20073 VSS.n20072 0.00339046
R70400 VSS.n1082 VSS.n1081 0.00339046
R70401 VSS.n6892 VSS.n6891 0.00339046
R70402 VSS.n6520 VSS.n6519 0.00339046
R70403 VSS.n6484 VSS.n6483 0.00339046
R70404 VSS.n20133 VSS.n20132 0.00339046
R70405 VSS.n20072 VSS.n20071 0.00339046
R70406 VSS.n19136 VSS.n19135 0.00339046
R70407 VSS.n21384 VSS.n21383 0.00339046
R70408 VSS.n21325 VSS.n21324 0.00339046
R70409 VSS.n7613 VSS.n7612 0.00339046
R70410 VSS.n7673 VSS.n7672 0.00339046
R70411 VSS.n7701 VSS.n7700 0.00339046
R70412 VSS.n7761 VSS.n7760 0.00339046
R70413 VSS.n7838 VSS.n7837 0.00339046
R70414 VSS.n7779 VSS.n7778 0.00339046
R70415 VSS.n21324 VSS.n21323 0.00339046
R70416 VSS.n21385 VSS.n21384 0.00339046
R70417 VSS.n9309 VSS.n9308 0.00339046
R70418 VSS.n7839 VSS.n7838 0.00339046
R70419 VSS.n9146 VSS.n9145 0.00339046
R70420 VSS.n6635 VSS.n6634 0.00339046
R70421 VSS.n6485 VSS.n6484 0.00339046
R70422 VSS.n7778 VSS.n7777 0.00339046
R70423 VSS.n9700 VSS.n9699 0.00339046
R70424 VSS.n7700 VSS.n7699 0.00339046
R70425 VSS.n9583 VSS.n9582 0.00339046
R70426 VSS.n7760 VSS.n7759 0.00339046
R70427 VSS.n6669 VSS.n6668 0.00339046
R70428 VSS.n6519 VSS.n6518 0.00339046
R70429 VSS.n6995 VSS.n6994 0.00339046
R70430 VSS.n6893 VSS.n6892 0.00339046
R70431 VSS.n7672 VSS.n7671 0.00339046
R70432 VSS.n7612 VSS.n7611 0.00339046
R70433 VSS.n12750 VSS.n12749 0.00339046
R70434 VSS.n16103 VSS.n16102 0.00339046
R70435 VSS.n5587 VSS.n5586 0.00339046
R70436 VSS.n21037 VSS.n21036 0.00339046
R70437 VSS.n1083 VSS.n1082 0.00339046
R70438 VSS.n11644 VSS.n11643 0.00339046
R70439 VSS.n6088 VSS.n6087 0.00339046
R70440 VSS.n6007 VSS.n6006 0.00339046
R70441 VSS.n5926 VSS.n5925 0.00339046
R70442 VSS.n11699 VSS.n11698 0.00339046
R70443 VSS.n6142 VSS.n6141 0.00339046
R70444 VSS.n6061 VSS.n6060 0.00339046
R70445 VSS.n5980 VSS.n5979 0.00339046
R70446 VSS.n3972 VSS.n3971 0.00339046
R70447 VSS.n2638 VSS.n2637 0.00339046
R70448 VSS.n2606 VSS.n2605 0.00339046
R70449 VSS.n2639 VSS.n2638 0.00339046
R70450 VSS.n10614 VSS.n10613 0.00339046
R70451 VSS.n602 VSS.n601 0.00339046
R70452 VSS.n656 VSS.n655 0.00339046
R70453 VSS.n10313 VSS.n10308 0.00338462
R70454 VSS.n10431 VSS.n10426 0.00338462
R70455 VSS.n10339 VSS.n10334 0.00338462
R70456 VSS.n10146 VSS.n10141 0.00338462
R70457 VSS.n10054 VSS.n10049 0.00338462
R70458 VSS.n10031 VSS.n10030 0.00338462
R70459 VSS.n12367 VSS.n12362 0.00338462
R70460 VSS.n12485 VSS.n12480 0.00338462
R70461 VSS.n12393 VSS.n12388 0.00338462
R70462 VSS.n12197 VSS.n12192 0.00338462
R70463 VSS.n12105 VSS.n12100 0.00338462
R70464 VSS.n12082 VSS.n12081 0.00338462
R70465 VSS.n718 VSS.n717 0.00338
R70466 VSS.n20578 VSS.n20577 0.00338
R70467 VSS.n20556 VSS.n20555 0.00338
R70468 VSS.n7866 VSS.n7865 0.00338
R70469 VSS.n7959 VSS.n7958 0.00338
R70470 VSS.n11071 VSS.n11069 0.00338
R70471 VSS.n21771 VSS.n21770 0.00337808
R70472 VSS.n19056 VSS.n19055 0.00337808
R70473 VSS.n5692 VSS.n5691 0.00337234
R70474 VSS.n5669 VSS.n5667 0.00337234
R70475 VSS.n16012 VSS.n16010 0.00337234
R70476 VSS.n16025 VSS.n16023 0.00337234
R70477 VSS.n993 VSS.n991 0.00337234
R70478 VSS.n984 VSS.n982 0.00337234
R70479 VSS.n20938 VSS.n20936 0.00337234
R70480 VSS.n20961 VSS.n20960 0.00337234
R70481 VSS.n1246 VSS.n1245 0.00337234
R70482 VSS.n11907 VSS.n11906 0.00335985
R70483 VSS.n11940 VSS.n11939 0.00335984
R70484 VSS.n3994 VSS.n3993 0.00333465
R70485 VSS.n4039 VSS.n4038 0.00333465
R70486 VSS.n17436 VSS.n17435 0.00333465
R70487 VSS.n17318 VSS.n17317 0.00333465
R70488 VSS.n9545 VSS.n9544 0.00333465
R70489 VSS.n9046 VSS.n9045 0.00333465
R70490 VSS.n13068 VSS.n13067 0.00333465
R70491 VSS.n12986 VSS.n12985 0.00333465
R70492 VSS.n12768 VSS.n12767 0.00333465
R70493 VSS.n12604 VSS.n12603 0.00333465
R70494 VSS.n12313 VSS.n12312 0.00333465
R70495 VSS.n12274 VSS.n12273 0.00333465
R70496 VSS.n11966 VSS.n11965 0.00333465
R70497 VSS.n11929 VSS.n11928 0.00333465
R70498 VSS.n11918 VSS.n11917 0.00333465
R70499 VSS.n11798 VSS.n11797 0.00333465
R70500 VSS.n18865 VSS.n18864 0.00333465
R70501 VSS.n18910 VSS.n18909 0.00333465
R70502 VSS.n2187 VSS.n2186 0.00333465
R70503 VSS.n14410 VSS.n14409 0.00333465
R70504 VSS.n9662 VSS.n9661 0.00333465
R70505 VSS.n9189 VSS.n9188 0.00333465
R70506 VSS.n21841 VSS.n21840 0.00333465
R70507 VSS.n20598 VSS.n20597 0.00333465
R70508 VSS.n6952 VSS.n6951 0.00333465
R70509 VSS.n6679 VSS.n6678 0.00333465
R70510 VSS.n19126 VSS.n19125 0.00333465
R70511 VSS.n20160 VSS.n20159 0.00333465
R70512 VSS.n6850 VSS.n6849 0.00333465
R70513 VSS.n6529 VSS.n6528 0.00333465
R70514 VSS.n21612 VSS.n21611 0.00333465
R70515 VSS.n21538 VSS.n21537 0.00333465
R70516 VSS.n21403 VSS.n21402 0.00333465
R70517 VSS.n7594 VSS.n7593 0.00333465
R70518 VSS.n7682 VSS.n7681 0.00333465
R70519 VSS.n7770 VSS.n7769 0.00333465
R70520 VSS.n3841 VSS.n3840 0.00333465
R70521 VSS.n4154 VSS.n4153 0.00333465
R70522 VSS.n11728 VSS.n11727 0.00333465
R70523 VSS.n11191 VSS.n11190 0.00333465
R70524 VSS.n6079 VSS.n6078 0.00333465
R70525 VSS.n5998 VSS.n5997 0.00333465
R70526 VSS.n3274 VSS.n3273 0.00333465
R70527 VSS.n2656 VSS.n2655 0.00333465
R70528 VSS.n674 VSS.n673 0.00333465
R70529 VSS.n471 VSS.n470 0.00333465
R70530 VSS.n10538 VSS.n10537 0.00333465
R70531 VSS.n10260 VSS.n10259 0.00333465
R70532 VSS.n10223 VSS.n10222 0.00333465
R70533 VSS.n9969 VSS.n9968 0.00333465
R70534 VSS.n9930 VSS.n9929 0.00333465
R70535 VSS.n9919 VSS.n9918 0.00333465
R70536 VSS.n8901 VSS.n8900 0.00333465
R70537 VSS.n2683 VSS.n2682 0.00332857
R70538 VSS.n2728 VSS.n2727 0.00332857
R70539 VSS.n2788 VSS.n2787 0.00332857
R70540 VSS.n2569 VSS.n2568 0.00332857
R70541 VSS.n4335 VSS.n4334 0.00332857
R70542 VSS.n17542 VSS.n17541 0.00332857
R70543 VSS.n17484 VSS.n17483 0.00332857
R70544 VSS.n17727 VSS.n17726 0.00332857
R70545 VSS.n18693 VSS.n18692 0.00332274
R70546 VSS.n18694 VSS.n18693 0.00332274
R70547 VSS.n19175 VSS.n19174 0.00332274
R70548 VSS.n19176 VSS.n19175 0.00332274
R70549 VSS.n15457 VSS.n15456 0.00332274
R70550 VSS.n15458 VSS.n15457 0.00332274
R70551 VSS.n1759 VSS.n1758 0.00332274
R70552 VSS.n1760 VSS.n1759 0.00332274
R70553 VSS.n10649 VSS.n10648 0.00332
R70554 VSS.n9410 VSS.n9409 0.00332
R70555 VSS.n9802 VSS.n9801 0.00332
R70556 VSS.n10656 VSS.n10654 0.00332
R70557 VSS.n18684 VSS.n18683 0.00330302
R70558 VSS.n3948 VSS.n3947 0.00330197
R70559 VSS.n2368 VSS.n2367 0.00330197
R70560 VSS.n11337 VSS.n11336 0.00330197
R70561 VSS.n9091 VSS.n9090 0.00330197
R70562 VSS.n3949 VSS.n3948 0.00330197
R70563 VSS.n4031 VSS.n4030 0.00330197
R70564 VSS.n5860 VSS.n5859 0.00330197
R70565 VSS.n13059 VSS.n13058 0.00330197
R70566 VSS.n13132 VSS.n13131 0.00330197
R70567 VSS.n13179 VSS.n13178 0.00330197
R70568 VSS.n12872 VSS.n12871 0.00330197
R70569 VSS.n12809 VSS.n12808 0.00330197
R70570 VSS.n12505 VSS.n12504 0.00330197
R70571 VSS.n12267 VSS.n12266 0.00330197
R70572 VSS.n11922 VSS.n11921 0.00330197
R70573 VSS.n13131 VSS.n13130 0.00330197
R70574 VSS.n12873 VSS.n12872 0.00330197
R70575 VSS.n13058 VSS.n13057 0.00330197
R70576 VSS.n12810 VSS.n12809 0.00330197
R70577 VSS.n13180 VSS.n13179 0.00330197
R70578 VSS.n18977 VSS.n18976 0.00330197
R70579 VSS.n15138 VSS.n15137 0.00330197
R70580 VSS.n16221 VSS.n16220 0.00330197
R70581 VSS.n9255 VSS.n9254 0.00330197
R70582 VSS.n18976 VSS.n18975 0.00330197
R70583 VSS.n18902 VSS.n18901 0.00330197
R70584 VSS.n2267 VSS.n2266 0.00330197
R70585 VSS.n21832 VSS.n21831 0.00330197
R70586 VSS.n21746 VSS.n21745 0.00330197
R70587 VSS.n2319 VSS.n2318 0.00330197
R70588 VSS.n20788 VSS.n20787 0.00330197
R70589 VSS.n21164 VSS.n21163 0.00330197
R70590 VSS.n6574 VSS.n6573 0.00330197
R70591 VSS.n21747 VSS.n21746 0.00330197
R70592 VSS.n20787 VSS.n20786 0.00330197
R70593 VSS.n21831 VSS.n21830 0.00330197
R70594 VSS.n2320 VSS.n2319 0.00330197
R70595 VSS.n21163 VSS.n21162 0.00330197
R70596 VSS.n19117 VSS.n19116 0.00330197
R70597 VSS.n19031 VSS.n19030 0.00330197
R70598 VSS.n17927 VSS.n17926 0.00330197
R70599 VSS.n2031 VSS.n2030 0.00330197
R70600 VSS.n1293 VSS.n1292 0.00330197
R70601 VSS.n6424 VSS.n6423 0.00330197
R70602 VSS.n19032 VSS.n19031 0.00330197
R70603 VSS.n2032 VSS.n2031 0.00330197
R70604 VSS.n19116 VSS.n19115 0.00330197
R70605 VSS.n17928 VSS.n17927 0.00330197
R70606 VSS.n1292 VSS.n1291 0.00330197
R70607 VSS.n21603 VSS.n21602 0.00330197
R70608 VSS.n21494 VSS.n21493 0.00330197
R70609 VSS.n21293 VSS.n21292 0.00330197
R70610 VSS.n7553 VSS.n7552 0.00330197
R70611 VSS.n21294 VSS.n21293 0.00330197
R70612 VSS.n21602 VSS.n21601 0.00330197
R70613 VSS.n21493 VSS.n21492 0.00330197
R70614 VSS.n7552 VSS.n7551 0.00330197
R70615 VSS.n6575 VSS.n6574 0.00330197
R70616 VSS.n6425 VSS.n6424 0.00330197
R70617 VSS.n11923 VSS.n11922 0.00330197
R70618 VSS.n9092 VSS.n9091 0.00330197
R70619 VSS.n12506 VSS.n12505 0.00330197
R70620 VSS.n4721 VSS.n4720 0.00330197
R70621 VSS.n11451 VSS.n11450 0.00330197
R70622 VSS.n11230 VSS.n11229 0.00330197
R70623 VSS.n3833 VSS.n3832 0.00330197
R70624 VSS.n2648 VSS.n2647 0.00330197
R70625 VSS.n569 VSS.n568 0.00330197
R70626 VSS.n510 VSS.n509 0.00330197
R70627 VSS.n10451 VSS.n10450 0.00330197
R70628 VSS.n10215 VSS.n10214 0.00330197
R70629 VSS.n9923 VSS.n9922 0.00330197
R70630 VSS.n10452 VSS.n10451 0.00330197
R70631 VSS.n10216 VSS.n10215 0.00330197
R70632 VSS.n9924 VSS.n9923 0.00330197
R70633 VSS.n4165 VSS.n2521 0.00327778
R70634 VSS.n21707 VSS.n21705 0.00327778
R70635 VSS.n17401 VSS.n17399 0.00327778
R70636 VSS.n375 VSS.n372 0.00327778
R70637 VSS.n4114 VSS.n4113 0.00327778
R70638 VSS.n21910 VSS.n21909 0.00327778
R70639 VSS.n10228 VSS.n10227 0.00327131
R70640 VSS.n10266 VSS.n10265 0.00327102
R70641 VSS.n2937 VSS.n2936 0.00326429
R70642 VSS.n3001 VSS.n3000 0.00326429
R70643 VSS.n3049 VSS.n3048 0.00326429
R70644 VSS.n7355 VSS.n7354 0.00326429
R70645 VSS.n7301 VSS.n7300 0.00326429
R70646 VSS.n17872 VSS.n17871 0.00326429
R70647 VSS.n17811 VSS.n17810 0.00326429
R70648 VSS.n17766 VSS.n17765 0.00326429
R70649 VSS.n18706 VSS.n18705 0.00324648
R70650 VSS.n18784 VSS.n18783 0.00324648
R70651 VSS.n18199 VSS.n18198 0.00324648
R70652 VSS.n18196 VSS.n18195 0.00324648
R70653 VSS.n18194 VSS.n18193 0.00324648
R70654 VSS.n17131 VSS.n17130 0.00324648
R70655 VSS.n14869 VSS.n14868 0.00324648
R70656 VSS.n16936 VSS.n16935 0.00324648
R70657 VSS.n15397 VSS.n15396 0.00324648
R70658 VSS.n15378 VSS.n15377 0.00324648
R70659 VSS.n19188 VSS.n19187 0.00324648
R70660 VSS.n19456 VSS.n19455 0.00324648
R70661 VSS.n19657 VSS.n19656 0.00324648
R70662 VSS.n19660 VSS.n19659 0.00324648
R70663 VSS.n19662 VSS.n19661 0.00324648
R70664 VSS.n19864 VSS.n19863 0.00324648
R70665 VSS.n19940 VSS.n19939 0.00324648
R70666 VSS.n19980 VSS.n19979 0.00324648
R70667 VSS.n1713 VSS.n1712 0.00324648
R70668 VSS.n1694 VSS.n1693 0.00324648
R70669 VSS.n18793 VSS.n18792 0.00321722
R70670 VSS.n18470 VSS.n18469 0.00321722
R70671 VSS.n18202 VSS.n18201 0.00321722
R70672 VSS.n18149 VSS.n18148 0.00321722
R70673 VSS.n15549 VSS.n15548 0.00321722
R70674 VSS.n15408 VSS.n15407 0.00321722
R70675 VSS.n8334 VSS.n8333 0.00321722
R70676 VSS.n16924 VSS.n16923 0.00321722
R70677 VSS.n18203 VSS.n18202 0.00321722
R70678 VSS.n18471 VSS.n18470 0.00321722
R70679 VSS.n18792 VSS.n18791 0.00321722
R70680 VSS.n18150 VSS.n18149 0.00321722
R70681 VSS.n15548 VSS.n15547 0.00321722
R70682 VSS.n15392 VSS.n15391 0.00321722
R70683 VSS.n8333 VSS.n8332 0.00321722
R70684 VSS.n15409 VSS.n15408 0.00321722
R70685 VSS.n19465 VSS.n19464 0.00321722
R70686 VSS.n19569 VSS.n19568 0.00321722
R70687 VSS.n19654 VSS.n19653 0.00321722
R70688 VSS.n19707 VSS.n19706 0.00321722
R70689 VSS.n1837 VSS.n1836 0.00321722
R70690 VSS.n1724 VSS.n1723 0.00321722
R70691 VSS.n8130 VSS.n8129 0.00321722
R70692 VSS.n8129 VSS.n8128 0.00321722
R70693 VSS.n1725 VSS.n1724 0.00321722
R70694 VSS.n1708 VSS.n1707 0.00321722
R70695 VSS.n19992 VSS.n19991 0.00321722
R70696 VSS.n19568 VSS.n19567 0.00321722
R70697 VSS.n19464 VSS.n19463 0.00321722
R70698 VSS.n19653 VSS.n19652 0.00321722
R70699 VSS.n19706 VSS.n19705 0.00321722
R70700 VSS.n1836 VSS.n1835 0.00321722
R70701 VSS.n2357 VSS.n2356 0.00321348
R70702 VSS.n3985 VSS.n3984 0.00321348
R70703 VSS.n12844 VSS.n12843 0.00321348
R70704 VSS.n12845 VSS.n12844 0.00321348
R70705 VSS.n20816 VSS.n20815 0.00321348
R70706 VSS.n20815 VSS.n20814 0.00321348
R70707 VSS.n21265 VSS.n21264 0.00321348
R70708 VSS.n21266 VSS.n21265 0.00321348
R70709 VSS.n17459 VSS.n17458 0.00321348
R70710 VSS.n11363 VSS.n11362 0.00321348
R70711 VSS.n5730 VSS.n5729 0.00321348
R70712 VSS.n5634 VSS.n5633 0.00321348
R70713 VSS.n9502 VSS.n9501 0.00321348
R70714 VSS.n13010 VSS.n13009 0.00321348
R70715 VSS.n13138 VSS.n13137 0.00321348
R70716 VSS.n13167 VSS.n13166 0.00321348
R70717 VSS.n12781 VSS.n12780 0.00321348
R70718 VSS.n13166 VSS.n13165 0.00321348
R70719 VSS.n12782 VSS.n12781 0.00321348
R70720 VSS.n13011 VSS.n13010 0.00321348
R70721 VSS.n15164 VSS.n15163 0.00321348
R70722 VSS.n16322 VSS.n16321 0.00321348
R70723 VSS.n16287 VSS.n16286 0.00321348
R70724 VSS.n16251 VSS.n16250 0.00321348
R70725 VSS.n16198 VSS.n16197 0.00321348
R70726 VSS.n16178 VSS.n16177 0.00321348
R70727 VSS.n16162 VSS.n16161 0.00321348
R70728 VSS.n16156 VSS.n16155 0.00321348
R70729 VSS.n9619 VSS.n9618 0.00321348
R70730 VSS.n16323 VSS.n16322 0.00321348
R70731 VSS.n16288 VSS.n16287 0.00321348
R70732 VSS.n16252 VSS.n16251 0.00321348
R70733 VSS.n2256 VSS.n2255 0.00321348
R70734 VSS.n18856 VSS.n18855 0.00321348
R70735 VSS.n16157 VSS.n16156 0.00321348
R70736 VSS.n5635 VSS.n5634 0.00321348
R70737 VSS.n16163 VSS.n16162 0.00321348
R70738 VSS.n16199 VSS.n16198 0.00321348
R70739 VSS.n21783 VSS.n21782 0.00321348
R70740 VSS.n2307 VSS.n2306 0.00321348
R70741 VSS.n21140 VSS.n21139 0.00321348
R70742 VSS.n21118 VSS.n21117 0.00321348
R70743 VSS.n21084 VSS.n21083 0.00321348
R70744 VSS.n2306 VSS.n2305 0.00321348
R70745 VSS.n21119 VSS.n21118 0.00321348
R70746 VSS.n21784 VSS.n21783 0.00321348
R70747 VSS.n21141 VSS.n21140 0.00321348
R70748 VSS.n21085 VSS.n21084 0.00321348
R70749 VSS.n19068 VSS.n19067 0.00321348
R70750 VSS.n17915 VSS.n17914 0.00321348
R70751 VSS.n2003 VSS.n2002 0.00321348
R70752 VSS.n1403 VSS.n1402 0.00321348
R70753 VSS.n1368 VSS.n1367 0.00321348
R70754 VSS.n1332 VSS.n1331 0.00321348
R70755 VSS.n1168 VSS.n1167 0.00321348
R70756 VSS.n1136 VSS.n1135 0.00321348
R70757 VSS.n17914 VSS.n17913 0.00321348
R70758 VSS.n1137 VSS.n1136 0.00321348
R70759 VSS.n1169 VSS.n1168 0.00321348
R70760 VSS.n2004 VSS.n2003 0.00321348
R70761 VSS.n1333 VSS.n1332 0.00321348
R70762 VSS.n1369 VSS.n1368 0.00321348
R70763 VSS.n1404 VSS.n1403 0.00321348
R70764 VSS.n19069 VSS.n19068 0.00321348
R70765 VSS.n21551 VSS.n21550 0.00321348
R70766 VSS.n21506 VSS.n21505 0.00321348
R70767 VSS.n7581 VSS.n7580 0.00321348
R70768 VSS.n21507 VSS.n21506 0.00321348
R70769 VSS.n7580 VSS.n7579 0.00321348
R70770 VSS.n21552 VSS.n21551 0.00321348
R70771 VSS.n3785 VSS.n3784 0.00321348
R70772 VSS.n4161 VSS.n4160 0.00321348
R70773 VSS.n4710 VSS.n4709 0.00321348
R70774 VSS.n11425 VSS.n11424 0.00321348
R70775 VSS.n11204 VSS.n11203 0.00321348
R70776 VSS.n4162 VSS.n4161 0.00321348
R70777 VSS.n3265 VSS.n3264 0.00321348
R70778 VSS.n543 VSS.n542 0.00321348
R70779 VSS.n484 VSS.n483 0.00321348
R70780 VSS.n6932 VSS.n6931 0.00321348
R70781 VSS.n6809 VSS.n6808 0.00321348
R70782 VSS.n9618 VSS.n9617 0.00321348
R70783 VSS.n9501 VSS.n9500 0.00321348
R70784 VSS.n21426 VSS.n21425 0.00321348
R70785 VSS.n21415 VSS.n21414 0.00321348
R70786 VSS.n21316 VSS.n21315 0.00321348
R70787 VSS.n21305 VSS.n21304 0.00321348
R70788 VSS.n21253 VSS.n21252 0.00321348
R70789 VSS.n13137 VSS.n13136 0.00321348
R70790 VSS.n17460 VSS.n17459 0.00321348
R70791 VSS.n4779 VSS.n4778 0.00321348
R70792 VSS.n19403 VSS.n19402 0.0032
R70793 VSS.n18263 VSS.n18261 0.0032
R70794 VSS.n18249 VSS.n18247 0.0032
R70795 VSS.n16661 VSS.n16660 0.0032
R70796 VSS.n16617 VSS.n16616 0.0032
R70797 VSS.n16511 VSS.n16510 0.0032
R70798 VSS.n2932 VSS.n2931 0.0032
R70799 VSS.n2996 VSS.n2995 0.0032
R70800 VSS.n3044 VSS.n3043 0.0032
R70801 VSS.n17970 VSS.n17969 0.0032
R70802 VSS.n17816 VSS.n17815 0.0032
R70803 VSS.n17771 VSS.n17770 0.0032
R70804 VSS.n21635 VSS.n21634 0.0031825
R70805 VSS.n21245 VSS.n21244 0.00317666
R70806 VSS.n11139 VSS.n6295 0.00316667
R70807 VSS.n11114 VSS.n6345 0.00316667
R70808 VSS.n6245 VSS.n6205 0.00316667
R70809 VSS.n6295 VSS.n6270 0.00316667
R70810 VSS.n6345 VSS.n6320 0.00316667
R70811 VSS.n11089 VSS.n6346 0.00316667
R70812 VSS.n7009 VSS.n6346 0.00316667
R70813 VSS.n11164 VSS.n6245 0.00316667
R70814 VSS.n18139 VSS.n18138 0.00316244
R70815 VSS.n18172 VSS.n18171 0.00316244
R70816 VSS.n18165 VSS.n18164 0.00316244
R70817 VSS.n18147 VSS.n18146 0.00316244
R70818 VSS.n19684 VSS.n19683 0.00316244
R70819 VSS.n19709 VSS.n19708 0.00316244
R70820 VSS.n4200 VSS.n4199 0.00315748
R70821 VSS.n2349 VSS.n2348 0.00315748
R70822 VSS.n17468 VSS.n17467 0.00315748
R70823 VSS.n11355 VSS.n11354 0.00315748
R70824 VSS.n5738 VSS.n5737 0.00315748
R70825 VSS.n13139 VSS.n13138 0.00315748
R70826 VSS.n13157 VSS.n13156 0.00315748
R70827 VSS.n12854 VSS.n12853 0.00315748
R70828 VSS.n12791 VSS.n12790 0.00315748
R70829 VSS.n12518 VSS.n12517 0.00315748
R70830 VSS.n12305 VSS.n12304 0.00315748
R70831 VSS.n12224 VSS.n12223 0.00315748
R70832 VSS.n11962 VSS.n11961 0.00315748
R70833 VSS.n11882 VSS.n11881 0.00315748
R70834 VSS.n11864 VSS.n11863 0.00315748
R70835 VSS.n11817 VSS.n11816 0.00315748
R70836 VSS.n2230 VSS.n2165 0.00315748
R70837 VSS.n2248 VSS.n2247 0.00315748
R70838 VSS.n2219 VSS.n2218 0.00315748
R70839 VSS.n15156 VSS.n15155 0.00315748
R70840 VSS.n16186 VSS.n16185 0.00315748
R70841 VSS.n2279 VSS.n347 0.00315748
R70842 VSS.n2297 VSS.n2296 0.00315748
R70843 VSS.n20806 VSS.n20805 0.00315748
R70844 VSS.n21128 VSS.n21127 0.00315748
R70845 VSS.n17887 VSS.n17886 0.00315748
R70846 VSS.n17905 VSS.n17904 0.00315748
R70847 VSS.n2013 VSS.n2012 0.00315748
R70848 VSS.n1178 VSS.n1177 0.00315748
R70849 VSS.n21674 VSS.n21673 0.00315748
R70850 VSS.n21544 VSS.n21543 0.00315748
R70851 VSS.n21527 VSS.n21526 0.00315748
R70852 VSS.n21516 VSS.n21515 0.00315748
R70853 VSS.n21464 VSS.n21463 0.00315748
R70854 VSS.n21275 VSS.n21274 0.00315748
R70855 VSS.n7571 VSS.n7570 0.00315748
R70856 VSS.n4135 VSS.n4134 0.00315748
R70857 VSS.n4160 VSS.n4159 0.00315748
R70858 VSS.n4144 VSS.n4143 0.00315748
R70859 VSS.n4702 VSS.n4701 0.00315748
R70860 VSS.n4771 VSS.n4770 0.00315748
R70861 VSS.n11433 VSS.n11432 0.00315748
R70862 VSS.n11212 VSS.n11211 0.00315748
R70863 VSS.n551 VSS.n550 0.00315748
R70864 VSS.n492 VSS.n491 0.00315748
R70865 VSS.n10463 VSS.n10462 0.00315748
R70866 VSS.n10253 VSS.n10252 0.00315748
R70867 VSS.n10172 VSS.n10171 0.00315748
R70868 VSS.n9965 VSS.n9964 0.00315748
R70869 VSS.n8944 VSS.n8943 0.00315748
R70870 VSS.n8975 VSS.n8974 0.00315748
R70871 VSS.n8832 VSS.n8831 0.00315748
R70872 VSS.n15513 VSS.n15512 0.00315322
R70873 VSS.n1783 VSS.n1782 0.00315322
R70874 VSS.n15512 VSS.n15511 0.00315322
R70875 VSS.n1782 VSS.n1781 0.00315322
R70876 VSS.n9772 VSS.n9771 0.00314496
R70877 VSS.n20178 VSS.n20176 0.00314
R70878 VSS.n693 VSS.n691 0.00314
R70879 VSS.n20573 VSS.n20572 0.00314
R70880 VSS.n7860 VSS.n7008 0.00314
R70881 VSS.n4023 VSS.n4022 0.00312498
R70882 VSS.n4052 VSS.n4051 0.00312498
R70883 VSS.n4063 VSS.n4062 0.00312498
R70884 VSS.n3970 VSS.n3969 0.00312498
R70885 VSS.n3959 VSS.n3958 0.00312498
R70886 VSS.n17461 VSS.n17460 0.00312498
R70887 VSS.n5722 VSS.n5721 0.00312498
R70888 VSS.n9085 VSS.n9084 0.00312498
R70889 VSS.n17462 VSS.n17461 0.00312498
R70890 VSS.n13050 VSS.n13049 0.00312498
R70891 VSS.n13081 VSS.n13080 0.00312498
R70892 VSS.n13091 VSS.n13090 0.00312498
R70893 VSS.n13110 VSS.n13109 0.00312498
R70894 VSS.n13121 VSS.n13120 0.00312498
R70895 VSS.n13136 VSS.n13135 0.00312498
R70896 VSS.n12575 VSS.n12574 0.00312498
R70897 VSS.n13135 VSS.n13134 0.00312498
R70898 VSS.n13049 VSS.n13048 0.00312498
R70899 VSS.n18923 VSS.n18922 0.00312498
R70900 VSS.n18934 VSS.n18933 0.00312498
R70901 VSS.n18955 VSS.n18954 0.00312498
R70902 VSS.n18966 VSS.n18965 0.00312498
R70903 VSS.n16364 VSS.n16363 0.00312498
R70904 VSS.n16319 VSS.n16318 0.00312498
R70905 VSS.n16284 VSS.n16283 0.00312498
R70906 VSS.n16170 VSS.n16169 0.00312498
R70907 VSS.n16164 VSS.n16163 0.00312498
R70908 VSS.n9249 VSS.n9248 0.00312498
R70909 VSS.n16365 VSS.n16364 0.00312498
R70910 VSS.n16320 VSS.n16319 0.00312498
R70911 VSS.n16285 VSS.n16284 0.00312498
R70912 VSS.n18894 VSS.n18893 0.00312498
R70913 VSS.n16165 VSS.n16164 0.00312498
R70914 VSS.n16171 VSS.n16170 0.00312498
R70915 VSS.n5723 VSS.n5722 0.00312498
R70916 VSS.n21823 VSS.n21822 0.00312498
R70917 VSS.n21854 VSS.n21853 0.00312498
R70918 VSS.n21864 VSS.n21863 0.00312498
R70919 VSS.n21768 VSS.n21767 0.00312498
R70920 VSS.n21757 VSS.n21756 0.00312498
R70921 VSS.n21110 VSS.n21109 0.00312498
R70922 VSS.n6570 VSS.n6569 0.00312498
R70923 VSS.n21111 VSS.n21110 0.00312498
R70924 VSS.n21822 VSS.n21821 0.00312498
R70925 VSS.n19108 VSS.n19107 0.00312498
R70926 VSS.n19139 VSS.n19138 0.00312498
R70927 VSS.n19149 VSS.n19148 0.00312498
R70928 VSS.n19053 VSS.n19052 0.00312498
R70929 VSS.n19042 VSS.n19041 0.00312498
R70930 VSS.n1445 VSS.n1444 0.00312498
R70931 VSS.n1400 VSS.n1399 0.00312498
R70932 VSS.n1365 VSS.n1364 0.00312498
R70933 VSS.n1160 VSS.n1159 0.00312498
R70934 VSS.n6419 VSS.n6418 0.00312498
R70935 VSS.n1161 VSS.n1160 0.00312498
R70936 VSS.n1446 VSS.n1445 0.00312498
R70937 VSS.n1401 VSS.n1400 0.00312498
R70938 VSS.n1366 VSS.n1365 0.00312498
R70939 VSS.n19107 VSS.n19106 0.00312498
R70940 VSS.n21594 VSS.n21593 0.00312498
R70941 VSS.n21681 VSS.n21680 0.00312498
R70942 VSS.n21457 VSS.n21456 0.00312498
R70943 VSS.n21254 VSS.n21253 0.00312498
R70944 VSS.n21306 VSS.n21305 0.00312498
R70945 VSS.n21317 VSS.n21316 0.00312498
R70946 VSS.n21416 VSS.n21415 0.00312498
R70947 VSS.n21427 VSS.n21426 0.00312498
R70948 VSS.n21458 VSS.n21457 0.00312498
R70949 VSS.n21680 VSS.n21679 0.00312498
R70950 VSS.n21593 VSS.n21592 0.00312498
R70951 VSS.n11824 VSS.n11823 0.00312498
R70952 VSS.n9086 VSS.n9085 0.00312498
R70953 VSS.n9250 VSS.n9249 0.00312498
R70954 VSS.n6420 VSS.n6419 0.00312498
R70955 VSS.n12576 VSS.n12575 0.00312498
R70956 VSS.n3825 VSS.n3824 0.00312498
R70957 VSS.n4778 VSS.n4777 0.00312498
R70958 VSS.n17247 VSS.n17246 0.00312498
R70959 VSS.n11741 VSS.n11740 0.00312498
R70960 VSS.n4925 VSS.n4924 0.00312498
R70961 VSS.n11462 VSS.n11461 0.00312498
R70962 VSS.n11243 VSS.n11242 0.00312498
R70963 VSS.n4777 VSS.n4776 0.00312498
R70964 VSS.n18965 VSS.n18964 0.00312498
R70965 VSS.n3960 VSS.n3959 0.00312498
R70966 VSS.n19054 VSS.n19053 0.00312498
R70967 VSS.n18954 VSS.n18953 0.00312498
R70968 VSS.n18933 VSS.n18932 0.00312498
R70969 VSS.n4062 VSS.n4061 0.00312498
R70970 VSS.n13090 VSS.n13089 0.00312498
R70971 VSS.n21863 VSS.n21862 0.00312498
R70972 VSS.n18922 VSS.n18921 0.00312498
R70973 VSS.n21853 VSS.n21852 0.00312498
R70974 VSS.n13120 VSS.n13119 0.00312498
R70975 VSS.n13109 VSS.n13108 0.00312498
R70976 VSS.n21758 VSS.n21757 0.00312498
R70977 VSS.n21769 VSS.n21768 0.00312498
R70978 VSS.n13080 VSS.n13079 0.00312498
R70979 VSS.n4051 VSS.n4050 0.00312498
R70980 VSS.n19138 VSS.n19137 0.00312498
R70981 VSS.n19148 VSS.n19147 0.00312498
R70982 VSS.n3971 VSS.n3970 0.00312498
R70983 VSS.n19043 VSS.n19042 0.00312498
R70984 VSS.n3246 VSS.n3245 0.00312498
R70985 VSS.n2636 VSS.n2635 0.00312498
R70986 VSS.n2625 VSS.n2624 0.00312498
R70987 VSS.n2604 VSS.n2603 0.00312498
R70988 VSS.n2593 VSS.n2592 0.00312498
R70989 VSS.n2594 VSS.n2593 0.00312498
R70990 VSS.n2626 VSS.n2625 0.00312498
R70991 VSS.n2637 VSS.n2636 0.00312498
R70992 VSS.n2605 VSS.n2604 0.00312498
R70993 VSS.n10510 VSS.n10509 0.00312498
R70994 VSS.n8936 VSS.n8933 0.00312498
R70995 VSS.n10511 VSS.n10510 0.00312498
R70996 VSS.n8936 VSS.n8935 0.00312498
R70997 VSS.n6569 VSS.n6568 0.00312498
R70998 VSS.n1770 VSS.n1769 0.00311264
R70999 VSS.n15468 VSS.n15467 0.00311264
R71000 VSS.n16597 VSS.n16596 0.00311219
R71001 VSS.n771 VSS.n770 0.00311219
R71002 VSS.n17013 VSS.n17012 0.00311168
R71003 VSS.n16891 VSS.n16890 0.00311168
R71004 VSS.n15671 VSS.n15670 0.00311168
R71005 VSS.n15357 VSS.n15356 0.00311168
R71006 VSS.n8478 VSS.n8477 0.00311168
R71007 VSS.n8559 VSS.n8558 0.00311168
R71008 VSS.n8326 VSS.n8325 0.00311168
R71009 VSS.n8414 VSS.n8413 0.00311168
R71010 VSS.n8363 VSS.n8362 0.00311168
R71011 VSS.n16892 VSS.n16891 0.00311168
R71012 VSS.n14871 VSS.n14870 0.00311168
R71013 VSS.n17014 VSS.n17013 0.00311168
R71014 VSS.n14981 VSS.n14973 0.00311168
R71015 VSS.n8415 VSS.n8414 0.00311168
R71016 VSS.n8362 VSS.n8361 0.00311168
R71017 VSS.n8325 VSS.n8324 0.00311168
R71018 VSS.n8560 VSS.n8559 0.00311168
R71019 VSS.n8477 VSS.n8476 0.00311168
R71020 VSS.n15358 VSS.n15357 0.00311168
R71021 VSS.n19922 VSS.n19921 0.00311168
R71022 VSS.n19942 VSS.n19941 0.00311168
R71023 VSS.n20025 VSS.n20024 0.00311168
R71024 VSS.n817 VSS.n816 0.00311168
R71025 VSS.n1928 VSS.n1927 0.00311168
R71026 VSS.n1673 VSS.n1672 0.00311168
R71027 VSS.n8628 VSS.n8627 0.00311168
R71028 VSS.n8710 VSS.n8709 0.00311168
R71029 VSS.n8122 VSS.n8121 0.00311168
R71030 VSS.n8222 VSS.n8221 0.00311168
R71031 VSS.n8171 VSS.n8170 0.00311168
R71032 VSS.n8629 VSS.n8628 0.00311168
R71033 VSS.n8121 VSS.n8120 0.00311168
R71034 VSS.n8711 VSS.n8710 0.00311168
R71035 VSS.n8223 VSS.n8222 0.00311168
R71036 VSS.n1674 VSS.n1673 0.00311168
R71037 VSS.n19921 VSS.n19920 0.00311168
R71038 VSS.n20024 VSS.n20023 0.00311168
R71039 VSS.n1929 VSS.n1928 0.00311168
R71040 VSS.n8170 VSS.n8169 0.00311168
R71041 VSS.n15670 VSS.n15669 0.00311168
R71042 VSS.n10459 VSS.n10458 0.00309404
R71043 VSS.n15428 VSS.n15427 0.00309215
R71044 VSS.n14565 VSS.n14564 0.00309215
R71045 VSS.n19763 VSS.n19762 0.00309215
R71046 VSS.n14830 VSS.n14829 0.00309215
R71047 VSS.n19853 VSS.n19852 0.00309215
R71048 VSS.n16878 VSS.n16877 0.00309215
R71049 VSS.n20038 VSS.n20037 0.00309215
R71050 VSS.n16689 VSS.n16688 0.00309215
R71051 VSS.n2091 VSS.n2090 0.00309215
R71052 VSS.n16438 VSS.n16437 0.00309215
R71053 VSS.n851 VSS.n850 0.00309215
R71054 VSS.n2689 VSS.n2687 0.00307143
R71055 VSS.n2733 VSS.n2732 0.00307143
R71056 VSS.n2793 VSS.n2792 0.00307143
R71057 VSS.n17537 VSS.n17536 0.00307143
R71058 VSS.n18103 VSS.n18102 0.00307143
R71059 VSS.n20394 VSS.n20393 0.00305
R71060 VSS.n20364 VSS.n20363 0.00305
R71061 VSS.n20333 VSS.n20332 0.00305
R71062 VSS.n20287 VSS.n20286 0.00305
R71063 VSS.n8820 VSS.n8818 0.00305
R71064 VSS.n9433 VSS.n9431 0.00305
R71065 VSS.n9808 VSS.n9806 0.00305
R71066 VSS.n3976 VSS.n3975 0.00303648
R71067 VSS.n4020 VSS.n4019 0.00303648
R71068 VSS.n13046 VSS.n13045 0.00303648
R71069 VSS.n13105 VSS.n13104 0.00303648
R71070 VSS.n13045 VSS.n13044 0.00303648
R71071 VSS.n18949 VSS.n18948 0.00303648
R71072 VSS.n18891 VSS.n18890 0.00303648
R71073 VSS.n21819 VSS.n21818 0.00303648
R71074 VSS.n21773 VSS.n21772 0.00303648
R71075 VSS.n21818 VSS.n21817 0.00303648
R71076 VSS.n19104 VSS.n19103 0.00303648
R71077 VSS.n19058 VSS.n19057 0.00303648
R71078 VSS.n19103 VSS.n19102 0.00303648
R71079 VSS.n21590 VSS.n21589 0.00303648
R71080 VSS.n21642 VSS.n21641 0.00303648
R71081 VSS.n21589 VSS.n21588 0.00303648
R71082 VSS.n3871 VSS.n3870 0.00303648
R71083 VSS.n3822 VSS.n3821 0.00303648
R71084 VSS.n3870 VSS.n3869 0.00303648
R71085 VSS.n3977 VSS.n3976 0.00303648
R71086 VSS.n18948 VSS.n18947 0.00303648
R71087 VSS.n19059 VSS.n19058 0.00303648
R71088 VSS.n21774 VSS.n21773 0.00303648
R71089 VSS.n13104 VSS.n13103 0.00303648
R71090 VSS.n21641 VSS.n21640 0.00303648
R71091 VSS.n3249 VSS.n3248 0.00303648
R71092 VSS.n2610 VSS.n2609 0.00303648
R71093 VSS.n2611 VSS.n2610 0.00303648
R71094 VSS.n18743 VSS.n18742 0.00303521
R71095 VSS.n18782 VSS.n18781 0.00303521
R71096 VSS.n18425 VSS.n18424 0.00303521
R71097 VSS.n18197 VSS.n18196 0.00303521
R71098 VSS.n18178 VSS.n18177 0.00303521
R71099 VSS.n18163 VSS.n18162 0.00303521
R71100 VSS.n16911 VSS.n16910 0.00303521
R71101 VSS.n16908 VSS.n16907 0.00303521
R71102 VSS.n16643 VSS.n16642 0.00303521
R71103 VSS.n16585 VSS.n16584 0.00303521
R71104 VSS.n14990 VSS.n14989 0.00303521
R71105 VSS.n14992 VSS.n14991 0.00303521
R71106 VSS.n15533 VSS.n15532 0.00303521
R71107 VSS.n15448 VSS.n15447 0.00303521
R71108 VSS.n15377 VSS.n15376 0.00303521
R71109 VSS.n19225 VSS.n19224 0.00303521
R71110 VSS.n19454 VSS.n19453 0.00303521
R71111 VSS.n19604 VSS.n19603 0.00303521
R71112 VSS.n19659 VSS.n19658 0.00303521
R71113 VSS.n19678 VSS.n19677 0.00303521
R71114 VSS.n19693 VSS.n19692 0.00303521
R71115 VSS.n20005 VSS.n20004 0.00303521
R71116 VSS.n20008 VSS.n20007 0.00303521
R71117 VSS.n755 VSS.n754 0.00303521
R71118 VSS.n783 VSS.n782 0.00303521
R71119 VSS.n826 VSS.n825 0.00303521
R71120 VSS.n828 VSS.n827 0.00303521
R71121 VSS.n1821 VSS.n1820 0.00303521
R71122 VSS.n1750 VSS.n1749 0.00303521
R71123 VSS.n1693 VSS.n1692 0.00303521
R71124 VSS.n16439 VSS.n16438 0.00302184
R71125 VSS.n14566 VSS.n14565 0.00302184
R71126 VSS.n14829 VSS.n14828 0.00302184
R71127 VSS.n16879 VSS.n16878 0.00302184
R71128 VSS.n16690 VSS.n16689 0.00302184
R71129 VSS.n1741 VSS.n1740 0.00302184
R71130 VSS.n19852 VSS.n19851 0.00302184
R71131 VSS.n19762 VSS.n19761 0.00302184
R71132 VSS.n850 VSS.n849 0.00302184
R71133 VSS.n2092 VSS.n2091 0.00302184
R71134 VSS.n20037 VSS.n20036 0.00302184
R71135 VSS.n15439 VSS.n15428 0.00302184
R71136 VSS.n9409 VSS.n9408 0.00302
R71137 VSS.n9356 VSS.n9354 0.00302
R71138 VSS.n9801 VSS.n9799 0.00302
R71139 VSS.n9747 VSS.n9745 0.00302
R71140 VSS.n10657 VSS.n10656 0.00302
R71141 VSS.n10719 VSS.n10718 0.00302
R71142 VSS.n16899 VSS.n16898 0.00300702
R71143 VSS.n20017 VSS.n20016 0.00300702
R71144 VSS.n18837 VSS.n18836 0.00300615
R71145 VSS.n18677 VSS.n18676 0.00300615
R71146 VSS.n15322 VSS.n15321 0.00300615
R71147 VSS.n8456 VSS.n8455 0.00300615
R71148 VSS.n8537 VSS.n8536 0.00300615
R71149 VSS.n8529 VSS.n8528 0.00300615
R71150 VSS.n8392 VSS.n8391 0.00300615
R71151 VSS.n8384 VSS.n8383 0.00300615
R71152 VSS.n17034 VSS.n17033 0.00300615
R71153 VSS.n16583 VSS.n16582 0.00300615
R71154 VSS.n16524 VSS.n16523 0.00300615
R71155 VSS.n18836 VSS.n18835 0.00300615
R71156 VSS.n18678 VSS.n18677 0.00300615
R71157 VSS.n8393 VSS.n8392 0.00300615
R71158 VSS.n8385 VSS.n8384 0.00300615
R71159 VSS.n8538 VSS.n8537 0.00300615
R71160 VSS.n8530 VSS.n8529 0.00300615
R71161 VSS.n15323 VSS.n15322 0.00300615
R71162 VSS.n19509 VSS.n19508 0.00300615
R71163 VSS.n19526 VSS.n19525 0.00300615
R71164 VSS.n785 VSS.n784 0.00300615
R71165 VSS.n814 VSS.n813 0.00300615
R71166 VSS.n1638 VSS.n1637 0.00300615
R71167 VSS.n8688 VSS.n8687 0.00300615
R71168 VSS.n8680 VSS.n8679 0.00300615
R71169 VSS.n8200 VSS.n8199 0.00300615
R71170 VSS.n8192 VSS.n8191 0.00300615
R71171 VSS.n8689 VSS.n8688 0.00300615
R71172 VSS.n8201 VSS.n8200 0.00300615
R71173 VSS.n8681 VSS.n8680 0.00300615
R71174 VSS.n8193 VSS.n8192 0.00300615
R71175 VSS.n1631 VSS.n1630 0.00300615
R71176 VSS.n19901 VSS.n19900 0.00300615
R71177 VSS.n19508 VSS.n19507 0.00300615
R71178 VSS.n19525 VSS.n19524 0.00300615
R71179 VSS.n1639 VSS.n1638 0.00300615
R71180 VSS.n4764 VSS.n4763 0.00300558
R71181 VSS.n10283 VSS.n10278 0.003
R71182 VSS.n10284 VSS.n10283 0.003
R71183 VSS.n10402 VSS.n10401 0.003
R71184 VSS.n10401 VSS.n10396 0.003
R71185 VSS.n10117 VSS.n10116 0.003
R71186 VSS.n10116 VSS.n10111 0.003
R71187 VSS.n8962 VSS.n8955 0.003
R71188 VSS.n8964 VSS.n8962 0.003
R71189 VSS.n21699 VSS.n21698 0.003
R71190 VSS.n21697 VSS.n21696 0.003
R71191 VSS.n366 VSS.n365 0.003
R71192 VSS.n364 VSS.n363 0.003
R71193 VSS.n12337 VSS.n12332 0.003
R71194 VSS.n12338 VSS.n12337 0.003
R71195 VSS.n12456 VSS.n12455 0.003
R71196 VSS.n12455 VSS.n12450 0.003
R71197 VSS.n12168 VSS.n12167 0.003
R71198 VSS.n12167 VSS.n12162 0.003
R71199 VSS.n12020 VSS.n12019 0.003
R71200 VSS.n12019 VSS.n12014 0.003
R71201 VSS.n21917 VSS.n21916 0.003
R71202 VSS.n21924 VSS.n21918 0.003
R71203 VSS.n9829 VSS.n9828 0.003
R71204 VSS.n9830 VSS.n9829 0.003
R71205 VSS.n12654 VSS.n12653 0.003
R71206 VSS.n12653 VSS.n12652 0.003
R71207 VSS.n4015 VSS.n4014 0.00298032
R71208 VSS.n13040 VSS.n13039 0.00298032
R71209 VSS.n18886 VSS.n18885 0.00298032
R71210 VSS.n21813 VSS.n21812 0.00298032
R71211 VSS.n19098 VSS.n19097 0.00298032
R71212 VSS.n21584 VSS.n21583 0.00298032
R71213 VSS.n3817 VSS.n3816 0.00298032
R71214 VSS.n3254 VSS.n3253 0.00298032
R71215 VSS.n19241 VSS.n19239 0.002975
R71216 VSS.n18660 VSS.n18658 0.002975
R71217 VSS.n16859 VSS.n16857 0.002975
R71218 VSS.n19775 VSS.n19773 0.002975
R71219 VSS.n14464 VSS.n14462 0.002975
R71220 VSS.n17135 VSS.n17133 0.002975
R71221 VSS.n17105 VSS.n17104 0.002975
R71222 VSS.n17056 VSS.n17055 0.002975
R71223 VSS.n16957 VSS.n16956 0.002975
R71224 VSS.n14919 VSS.n14918 0.002975
R71225 VSS.n16670 VSS.n16668 0.002975
R71226 VSS.n15709 VSS.n15707 0.002975
R71227 VSS.n3982 VSS.n3981 0.00294798
R71228 VSS.n2354 VSS.n2353 0.00294798
R71229 VSS.n5733 VSS.n5732 0.00294798
R71230 VSS.n11360 VSS.n11359 0.00294798
R71231 VSS.n13007 VSS.n13006 0.00294798
R71232 VSS.n13163 VSS.n13162 0.00294798
R71233 VSS.n12848 VSS.n12847 0.00294798
R71234 VSS.n12785 VSS.n12784 0.00294798
R71235 VSS.n12786 VSS.n12785 0.00294798
R71236 VSS.n12849 VSS.n12848 0.00294798
R71237 VSS.n13006 VSS.n13005 0.00294798
R71238 VSS.n13162 VSS.n13161 0.00294798
R71239 VSS.n15161 VSS.n15160 0.00294798
R71240 VSS.n16181 VSS.n16180 0.00294798
R71241 VSS.n2253 VSS.n2252 0.00294798
R71242 VSS.n18853 VSS.n18852 0.00294798
R71243 VSS.n21780 VSS.n21779 0.00294798
R71244 VSS.n2303 VSS.n2302 0.00294798
R71245 VSS.n20812 VSS.n20811 0.00294798
R71246 VSS.n21122 VSS.n21121 0.00294798
R71247 VSS.n21123 VSS.n21122 0.00294798
R71248 VSS.n20811 VSS.n20810 0.00294798
R71249 VSS.n21779 VSS.n21778 0.00294798
R71250 VSS.n2302 VSS.n2301 0.00294798
R71251 VSS.n19065 VSS.n19064 0.00294798
R71252 VSS.n17911 VSS.n17910 0.00294798
R71253 VSS.n2007 VSS.n2006 0.00294798
R71254 VSS.n1172 VSS.n1171 0.00294798
R71255 VSS.n1173 VSS.n1172 0.00294798
R71256 VSS.n2008 VSS.n2007 0.00294798
R71257 VSS.n19064 VSS.n19063 0.00294798
R71258 VSS.n17910 VSS.n17909 0.00294798
R71259 VSS.n21548 VSS.n21547 0.00294798
R71260 VSS.n21510 VSS.n21509 0.00294798
R71261 VSS.n21269 VSS.n21268 0.00294798
R71262 VSS.n7577 VSS.n7576 0.00294798
R71263 VSS.n7576 VSS.n7575 0.00294798
R71264 VSS.n21270 VSS.n21269 0.00294798
R71265 VSS.n21511 VSS.n21510 0.00294798
R71266 VSS.n21547 VSS.n21546 0.00294798
R71267 VSS.n4707 VSS.n4706 0.00294798
R71268 VSS.n11428 VSS.n11427 0.00294798
R71269 VSS.n11207 VSS.n11206 0.00294798
R71270 VSS.n3782 VSS.n3781 0.00294798
R71271 VSS.n3262 VSS.n3261 0.00294798
R71272 VSS.n487 VSS.n486 0.00294798
R71273 VSS.n546 VSS.n545 0.00294798
R71274 VSS.n2575 DVSS 0.00292857
R71275 VSS.n15402 VSS.n15401 0.00290105
R71276 VSS.n1718 VSS.n1717 0.00290105
R71277 VSS.n18829 VSS.n18828 0.00290061
R71278 VSS.n17027 VSS.n17026 0.00290061
R71279 VSS.n15365 VSS.n15364 0.00290061
R71280 VSS.n8567 VSS.n8566 0.00290061
R71281 VSS.n8422 VSS.n8421 0.00290061
R71282 VSS.n17028 VSS.n17027 0.00290061
R71283 VSS.n17073 VSS.n17072 0.00290061
R71284 VSS.n18828 VSS.n18827 0.00290061
R71285 VSS.n8423 VSS.n8422 0.00290061
R71286 VSS.n8568 VSS.n8567 0.00290061
R71287 VSS.n15366 VSS.n15365 0.00290061
R71288 VSS.n19500 VSS.n19499 0.00290061
R71289 VSS.n19908 VSS.n19907 0.00290061
R71290 VSS.n1682 VSS.n1681 0.00290061
R71291 VSS.n8718 VSS.n8717 0.00290061
R71292 VSS.n8230 VSS.n8229 0.00290061
R71293 VSS.n8719 VSS.n8718 0.00290061
R71294 VSS.n8231 VSS.n8230 0.00290061
R71295 VSS.n1681 VSS.n1680 0.00290061
R71296 VSS.n19892 VSS.n19891 0.00290061
R71297 VSS.n19907 VSS.n19906 0.00290061
R71298 VSS.n19501 VSS.n19500 0.00290061
R71299 VSS.n6746 VSS.n6745 0.0029
R71300 VSS.n8062 VSS.n8061 0.0029
R71301 VSS.n8002 VSS.n8001 0.0029
R71302 VSS.n10957 VSS.n10954 0.0029
R71303 VSS.n11027 VSS.n11021 0.0029
R71304 VSS.n2200 VSS.n2199 0.00286739
R71305 VSS.n18109 VSS.n18108 0.00286739
R71306 VSS.n2222 VSS.n2221 0.00286739
R71307 VSS.n2335 VSS.n2334 0.00286739
R71308 VSS.n13320 VSS.n13319 0.00286739
R71309 VSS.n13342 VSS.n13341 0.00286739
R71310 VSS.n17948 VSS.n17947 0.00286739
R71311 VSS.n17964 VSS.n17963 0.00286739
R71312 VSS.n13485 VSS.n13484 0.00286739
R71313 VSS.n2510 VSS.n2509 0.00286111
R71314 VSS.n2514 VSS.n2513 0.00286111
R71315 VSS.n2424 VSS.n2423 0.00286111
R71316 VSS.n2428 VSS.n2427 0.00286111
R71317 VSS.n3936 VSS.n3935 0.00286111
R71318 VSS.n3940 VSS.n3939 0.00286111
R71319 VSS.n4034 VSS.n4033 0.00285947
R71320 VSS.n3953 VSS.n3952 0.00285947
R71321 VSS.n17451 VSS.n17450 0.00285947
R71322 VSS.n17324 VSS.n17323 0.00285947
R71323 VSS.n11334 VSS.n11333 0.00285947
R71324 VSS.n5863 VSS.n5862 0.00285947
R71325 VSS.n5631 VSS.n5630 0.00285947
R71326 VSS.n5615 VSS.n5614 0.00285947
R71327 VSS.n9041 VSS.n9040 0.00285947
R71328 VSS.n3952 VSS.n3951 0.00285947
R71329 VSS.n17323 VSS.n17322 0.00285947
R71330 VSS.n13063 VSS.n13062 0.00285947
R71331 VSS.n13128 VSS.n13127 0.00285947
R71332 VSS.n13175 VSS.n13174 0.00285947
R71333 VSS.n13219 VSS.n13218 0.00285947
R71334 VSS.n13223 VSS.n13222 0.00285947
R71335 VSS.n12991 VSS.n12990 0.00285947
R71336 VSS.n12876 VSS.n12875 0.00285947
R71337 VSS.n12813 VSS.n12812 0.00285947
R71338 VSS.n12773 VSS.n12772 0.00285947
R71339 VSS.n12537 VSS.n12536 0.00285947
R71340 VSS.n12217 VSS.n12216 0.00285947
R71341 VSS.n12814 VSS.n12813 0.00285947
R71342 VSS.n12877 VSS.n12876 0.00285947
R71343 VSS.n12992 VSS.n12991 0.00285947
R71344 VSS.n13062 VSS.n13061 0.00285947
R71345 VSS.n13127 VSS.n13126 0.00285947
R71346 VSS.n2365 VSS.n2364 0.00285947
R71347 VSS.n13218 VSS.n13217 0.00285947
R71348 VSS.n13176 VSS.n13175 0.00285947
R71349 VSS.n13222 VSS.n13221 0.00285947
R71350 VSS.n17452 VSS.n17451 0.00285947
R71351 VSS.n18905 VSS.n18904 0.00285947
R71352 VSS.n18973 VSS.n18972 0.00285947
R71353 VSS.n2202 VSS.n2201 0.00285947
R71354 VSS.n14415 VSS.n14414 0.00285947
R71355 VSS.n15135 VSS.n15134 0.00285947
R71356 VSS.n16153 VSS.n16152 0.00285947
R71357 VSS.n16131 VSS.n16130 0.00285947
R71358 VSS.n9184 VSS.n9183 0.00285947
R71359 VSS.n2203 VSS.n2202 0.00285947
R71360 VSS.n16224 VSS.n16223 0.00285947
R71361 VSS.n14416 VSS.n14415 0.00285947
R71362 VSS.n18972 VSS.n18971 0.00285947
R71363 VSS.n2264 VSS.n2263 0.00285947
R71364 VSS.n16132 VSS.n16131 0.00285947
R71365 VSS.n5616 VSS.n5615 0.00285947
R71366 VSS.n21836 VSS.n21835 0.00285947
R71367 VSS.n21750 VSS.n21749 0.00285947
R71368 VSS.n2315 VSS.n2314 0.00285947
R71369 VSS.n13336 VSS.n13335 0.00285947
R71370 VSS.n13340 VSS.n13339 0.00285947
R71371 VSS.n20593 VSS.n20592 0.00285947
R71372 VSS.n20784 VSS.n20783 0.00285947
R71373 VSS.n21168 VSS.n21167 0.00285947
R71374 VSS.n21081 VSS.n21080 0.00285947
R71375 VSS.n21065 VSS.n21064 0.00285947
R71376 VSS.n6674 VSS.n6673 0.00285947
R71377 VSS.n21066 VSS.n21065 0.00285947
R71378 VSS.n20783 VSS.n20782 0.00285947
R71379 VSS.n20592 VSS.n20591 0.00285947
R71380 VSS.n13335 VSS.n13334 0.00285947
R71381 VSS.n21835 VSS.n21834 0.00285947
R71382 VSS.n21751 VSS.n21750 0.00285947
R71383 VSS.n2316 VSS.n2315 0.00285947
R71384 VSS.n13339 VSS.n13338 0.00285947
R71385 VSS.n21167 VSS.n21166 0.00285947
R71386 VSS.n19121 VSS.n19120 0.00285947
R71387 VSS.n19035 VSS.n19034 0.00285947
R71388 VSS.n17923 VSS.n17922 0.00285947
R71389 VSS.n13479 VSS.n13478 0.00285947
R71390 VSS.n13483 VSS.n13482 0.00285947
R71391 VSS.n20155 VSS.n20154 0.00285947
R71392 VSS.n2035 VSS.n2034 0.00285947
R71393 VSS.n1297 VSS.n1296 0.00285947
R71394 VSS.n1133 VSS.n1132 0.00285947
R71395 VSS.n1111 VSS.n1110 0.00285947
R71396 VSS.n6524 VSS.n6523 0.00285947
R71397 VSS.n1112 VSS.n1111 0.00285947
R71398 VSS.n20154 VSS.n20153 0.00285947
R71399 VSS.n2036 VSS.n2035 0.00285947
R71400 VSS.n13478 VSS.n13477 0.00285947
R71401 VSS.n19120 VSS.n19119 0.00285947
R71402 VSS.n19036 VSS.n19035 0.00285947
R71403 VSS.n17924 VSS.n17923 0.00285947
R71404 VSS.n13482 VSS.n13481 0.00285947
R71405 VSS.n1296 VSS.n1295 0.00285947
R71406 VSS.n21607 VSS.n21606 0.00285947
R71407 VSS.n21497 VSS.n21496 0.00285947
R71408 VSS.n21448 VSS.n21447 0.00285947
R71409 VSS.n21408 VSS.n21407 0.00285947
R71410 VSS.n21297 VSS.n21296 0.00285947
R71411 VSS.n7549 VSS.n7548 0.00285947
R71412 VSS.n7589 VSS.n7588 0.00285947
R71413 VSS.n7677 VSS.n7676 0.00285947
R71414 VSS.n7765 VSS.n7764 0.00285947
R71415 VSS.n7548 VSS.n7547 0.00285947
R71416 VSS.n21298 VSS.n21297 0.00285947
R71417 VSS.n21409 VSS.n21408 0.00285947
R71418 VSS.n21449 VSS.n21448 0.00285947
R71419 VSS.n21606 VSS.n21605 0.00285947
R71420 VSS.n21498 VSS.n21497 0.00285947
R71421 VSS.n7764 VSS.n7763 0.00285947
R71422 VSS.n12218 VSS.n12217 0.00285947
R71423 VSS.n6673 VSS.n6672 0.00285947
R71424 VSS.n6523 VSS.n6522 0.00285947
R71425 VSS.n9183 VSS.n9182 0.00285947
R71426 VSS.n9040 VSS.n9039 0.00285947
R71427 VSS.n12536 VSS.n12535 0.00285947
R71428 VSS.n7676 VSS.n7675 0.00285947
R71429 VSS.n7588 VSS.n7587 0.00285947
R71430 VSS.n12774 VSS.n12773 0.00285947
R71431 VSS.n21082 VSS.n21081 0.00285947
R71432 VSS.n1134 VSS.n1133 0.00285947
R71433 VSS.n16154 VSS.n16153 0.00285947
R71434 VSS.n5632 VSS.n5631 0.00285947
R71435 VSS.n3836 VSS.n3835 0.00285947
R71436 VSS.n4786 VSS.n4785 0.00285947
R71437 VSS.n11733 VSS.n11732 0.00285947
R71438 VSS.n11196 VSS.n11195 0.00285947
R71439 VSS.n6084 VSS.n6083 0.00285947
R71440 VSS.n6003 VSS.n6002 0.00285947
R71441 VSS.n4718 VSS.n4717 0.00285947
R71442 VSS.n11454 VSS.n11453 0.00285947
R71443 VSS.n11233 VSS.n11232 0.00285947
R71444 VSS.n6004 VSS.n6003 0.00285947
R71445 VSS.n11734 VSS.n11733 0.00285947
R71446 VSS.n11197 VSS.n11196 0.00285947
R71447 VSS.n4787 VSS.n4786 0.00285947
R71448 VSS.n6085 VSS.n6084 0.00285947
R71449 VSS.n2651 VSS.n2650 0.00285947
R71450 VSS.n669 VSS.n668 0.00285947
R71451 VSS.n476 VSS.n475 0.00285947
R71452 VSS.n10482 VSS.n10481 0.00285947
R71453 VSS.n10166 VSS.n10165 0.00285947
R71454 VSS.n10481 VSS.n10480 0.00285947
R71455 VSS.n513 VSS.n512 0.00285947
R71456 VSS.n572 VSS.n571 0.00285947
R71457 VSS.n668 VSS.n667 0.00285947
R71458 VSS.n477 VSS.n476 0.00285947
R71459 VSS.n19717 VSS.n19716 0.0028295
R71460 VSS.n19691 VSS.n19690 0.0028295
R71461 VSS.n11959 VSS.n11958 0.00282847
R71462 VSS.n11886 VSS.n11885 0.0028284
R71463 VSS.n18725 VSS.n18724 0.00282394
R71464 VSS.n18745 VSS.n18744 0.00282394
R71465 VSS.n18668 VSS.n18667 0.00282394
R71466 VSS.n18456 VSS.n18455 0.00282394
R71467 VSS.n14457 VSS.n14456 0.00282394
R71468 VSS.n14460 VSS.n14459 0.00282394
R71469 VSS.n14674 VSS.n14673 0.00282394
R71470 VSS.n17162 VSS.n17161 0.00282394
R71471 VSS.n17075 VSS.n17074 0.00282394
R71472 VSS.n17024 VSS.n17023 0.00282394
R71473 VSS.n16909 VSS.n16908 0.00282394
R71474 VSS.n16870 VSS.n16869 0.00282394
R71475 VSS.n16681 VSS.n16680 0.00282394
R71476 VSS.n16596 VSS.n16595 0.00282394
R71477 VSS.n16586 VSS.n16585 0.00282394
R71478 VSS.n16544 VSS.n16543 0.00282394
R71479 VSS.n15705 VSS.n15704 0.00282394
R71480 VSS.n15539 VSS.n15538 0.00282394
R71481 VSS.n15345 VSS.n15344 0.00282394
R71482 VSS.n19207 VSS.n19206 0.00282394
R71483 VSS.n19227 VSS.n19226 0.00282394
R71484 VSS.n19535 VSS.n19534 0.00282394
R71485 VSS.n19583 VSS.n19582 0.00282394
R71486 VSS.n19723 VSS.n19722 0.00282394
R71487 VSS.n19726 VSS.n19725 0.00282394
R71488 VSS.n19771 VSS.n19770 0.00282394
R71489 VSS.n19861 VSS.n19860 0.00282394
R71490 VSS.n19890 VSS.n19889 0.00282394
R71491 VSS.n19911 VSS.n19910 0.00282394
R71492 VSS.n20007 VSS.n20006 0.00282394
R71493 VSS.n2128 VSS.n2127 0.00282394
R71494 VSS.n751 VSS.n750 0.00282394
R71495 VSS.n772 VSS.n771 0.00282394
R71496 VSS.n782 VSS.n781 0.00282394
R71497 VSS.n794 VSS.n793 0.00282394
R71498 VSS.n1966 VSS.n1965 0.00282394
R71499 VSS.n1827 VSS.n1826 0.00282394
R71500 VSS.n1661 VSS.n1660 0.00282394
R71501 VSS.n2926 VSS.n2925 0.0028235
R71502 VSS.n13660 VSS.n13659 0.00282169
R71503 VSS.n17582 VSS.n17580 0.00281429
R71504 VSS.n11719 VSS.n11718 0.00281
R71505 VSS.n20376 VSS.n20375 0.00281
R71506 VSS.n20345 VSS.n20344 0.00281
R71507 VSS.n20299 VSS.n20298 0.00281
R71508 VSS.n20252 VSS.n20251 0.00281
R71509 VSS.n20212 VSS.n20211 0.00281
R71510 VSS.n727 VSS.n726 0.00281
R71511 VSS.n20583 VSS.n20582 0.00281
R71512 VSS.n20562 VSS.n20561 0.00281
R71513 VSS.n20533 VSS.n20532 0.00281
R71514 VSS.n8807 VSS.n8806 0.00281
R71515 VSS.n7036 VSS.n7035 0.00281
R71516 VSS.n9420 VSS.n9419 0.00281
R71517 VSS.n6162 VSS.n6161 0.00281
R71518 VSS.n13214 VSS.n13213 0.00280842
R71519 VSS.n2211 VSS.n2210 0.00280842
R71520 VSS.n5715 VSS.n5714 0.00280842
R71521 VSS.n21103 VSS.n21102 0.00280842
R71522 VSS.n21456 VSS.n21455 0.00280842
R71523 VSS.n21682 VSS.n21681 0.00280842
R71524 VSS.n17246 VSS.n17245 0.00280842
R71525 VSS.n11740 VSS.n11739 0.00280842
R71526 VSS.n4926 VSS.n4925 0.00280842
R71527 VSS.n11461 VSS.n11460 0.00280842
R71528 VSS.n11244 VSS.n11243 0.00280842
R71529 VSS.n14400 VSS.n14399 0.00280842
R71530 VSS.n13507 VSS.n13506 0.00280842
R71531 VSS.n13364 VSS.n13363 0.00280842
R71532 VSS.n13247 VSS.n13246 0.00280842
R71533 VSS.n14423 VSS.n14422 0.00280842
R71534 VSS.n20147 VSS.n20146 0.00280842
R71535 VSS.n13415 VSS.n13414 0.00280842
R71536 VSS.n12995 VSS.n12994 0.00280842
R71537 VSS.n593 VSS.n592 0.00280842
R71538 VSS.n15074 VSS.n15073 0.00280842
R71539 VSS.n2053 VSS.n2052 0.00280842
R71540 VSS.n20686 VSS.n20685 0.00280842
R71541 VSS.n12898 VSS.n12897 0.00280842
R71542 VSS.n580 VSS.n579 0.00280842
R71543 VSS.n15107 VSS.n15106 0.00280842
R71544 VSS.n2044 VSS.n2043 0.00280842
R71545 VSS.n20737 VSS.n20736 0.00280842
R71546 VSS.n12885 VSS.n12884 0.00280842
R71547 VSS.n530 VSS.n529 0.00280842
R71548 VSS.n15177 VSS.n15176 0.00280842
R71549 VSS.n883 VSS.n882 0.00280842
R71550 VSS.n20829 VSS.n20828 0.00280842
R71551 VSS.n12831 VSS.n12830 0.00280842
R71552 VSS.n13331 VSS.n13330 0.00280842
R71553 VSS.n13474 VSS.n13473 0.00280842
R71554 VSS.n21735 VSS.n21734 0.00280842
R71555 VSS.n17885 VSS.n2161 0.00280842
R71556 VSS.n18988 VSS.n18987 0.00280842
R71557 VSS.n21915 VSS.n21914 0.00280483
R71558 VSS.n21702 VSS.n21700 0.00280483
R71559 VSS.n369 VSS.n367 0.00280483
R71560 VSS.n3992 VSS.n3991 0.00280315
R71561 VSS.n5621 VSS.n5620 0.00280315
R71562 VSS.n5611 VSS.n5610 0.00280315
R71563 VSS.n9539 VSS.n9538 0.00280315
R71564 VSS.n13018 VSS.n13017 0.00280315
R71565 VSS.n12561 VSS.n12560 0.00280315
R71566 VSS.n12552 VSS.n12551 0.00280315
R71567 VSS.n12551 VSS.n12550 0.00280315
R71568 VSS.n12315 VSS.n12314 0.00280315
R71569 VSS.n12284 VSS.n12283 0.00280315
R71570 VSS.n12283 VSS.n12282 0.00280315
R71571 VSS.n12226 VSS.n12225 0.00280315
R71572 VSS.n11961 VSS.n11960 0.00280315
R71573 VSS.n11957 VSS.n11956 0.00280315
R71574 VSS.n11937 VSS.n11936 0.00280315
R71575 VSS.n11936 VSS.n11935 0.00280315
R71576 VSS.n11888 VSS.n11887 0.00280315
R71577 VSS.n11884 VSS.n11883 0.00280315
R71578 VSS.n11808 VSS.n11807 0.00280315
R71579 VSS.n11807 VSS.n11806 0.00280315
R71580 VSS.n18863 VSS.n18862 0.00280315
R71581 VSS.n16137 VSS.n16136 0.00280315
R71582 VSS.n16127 VSS.n16126 0.00280315
R71583 VSS.n9656 VSS.n9655 0.00280315
R71584 VSS.n21791 VSS.n21790 0.00280315
R71585 VSS.n21071 VSS.n21070 0.00280315
R71586 VSS.n21061 VSS.n21060 0.00280315
R71587 VSS.n19076 VSS.n19075 0.00280315
R71588 VSS.n1117 VSS.n1116 0.00280315
R71589 VSS.n1107 VSS.n1106 0.00280315
R71590 VSS.n21479 VSS.n21478 0.00280315
R71591 VSS.n4758 VSS.n4757 0.00280315
R71592 VSS.n3272 VSS.n3271 0.00280315
R71593 VSS.n10505 VSS.n10504 0.00280315
R71594 VSS.n10497 VSS.n10496 0.00280315
R71595 VSS.n10496 VSS.n10495 0.00280315
R71596 VSS.n10262 VSS.n10261 0.00280315
R71597 VSS.n10232 VSS.n10231 0.00280315
R71598 VSS.n10231 VSS.n10230 0.00280315
R71599 VSS.n10174 VSS.n10173 0.00280315
R71600 VSS.n9964 VSS.n9963 0.00280315
R71601 VSS.n9959 VSS.n9958 0.00280315
R71602 VSS.n9938 VSS.n9937 0.00280315
R71603 VSS.n9937 VSS.n9936 0.00280315
R71604 VSS.n8950 VSS.n8949 0.00280315
R71605 VSS.n8946 VSS.n8945 0.00280315
R71606 VSS.n8953 VSS.n8952 0.00280315
R71607 VSS.n8965 VSS.n8953 0.00280315
R71608 VSS.n14145 VSS.n14144 0.00279928
R71609 VSS.n14183 VSS.n14182 0.00279928
R71610 VSS.n14182 VSS.n14181 0.00279928
R71611 VSS.n14144 VSS.n14143 0.00279928
R71612 VSS.n18779 VSS.n18778 0.00279506
R71613 VSS.n18457 VSS.n18456 0.00279506
R71614 VSS.n18188 VSS.n18187 0.00279506
R71615 VSS.n14456 VSS.n14455 0.00279506
R71616 VSS.n15540 VSS.n15539 0.00279506
R71617 VSS.n18458 VSS.n18457 0.00279506
R71618 VSS.n14455 VSS.n14454 0.00279506
R71619 VSS.n18778 VSS.n18777 0.00279506
R71620 VSS.n18189 VSS.n18188 0.00279506
R71621 VSS.n15541 VSS.n15540 0.00279506
R71622 VSS.n19451 VSS.n19450 0.00279506
R71623 VSS.n19582 VSS.n19581 0.00279506
R71624 VSS.n19668 VSS.n19667 0.00279506
R71625 VSS.n19722 VSS.n19721 0.00279506
R71626 VSS.n1828 VSS.n1827 0.00279506
R71627 VSS.n19581 VSS.n19580 0.00279506
R71628 VSS.n19721 VSS.n19720 0.00279506
R71629 VSS.n19450 VSS.n19449 0.00279506
R71630 VSS.n19667 VSS.n19666 0.00279506
R71631 VSS.n1829 VSS.n1828 0.00279506
R71632 VSS.n3990 VSS.n3989 0.00277159
R71633 VSS.n13016 VSS.n13015 0.00277159
R71634 VSS.n18861 VSS.n18860 0.00277159
R71635 VSS.n21789 VSS.n21788 0.00277159
R71636 VSS.n19074 VSS.n19073 0.00277159
R71637 VSS.n3270 VSS.n3269 0.00277159
R71638 VSS.n11539 VSS.n11538 0.00277096
R71639 VSS.n11587 VSS.n11586 0.00277096
R71640 VSS.n5877 VSS.n5876 0.00277096
R71641 VSS.n5584 VSS.n5583 0.00277096
R71642 VSS.n9494 VSS.n9493 0.00277096
R71643 VSS.n9580 VSS.n9579 0.00277096
R71644 VSS.n9143 VSS.n9142 0.00277096
R71645 VSS.n9094 VSS.n9093 0.00277096
R71646 VSS.n12964 VSS.n12963 0.00277096
R71647 VSS.n12911 VSS.n12910 0.00277096
R71648 VSS.n12817 VSS.n12816 0.00277096
R71649 VSS.n12745 VSS.n12744 0.00277096
R71650 VSS.n12694 VSS.n12693 0.00277096
R71651 VSS.n12236 VSS.n12235 0.00277096
R71652 VSS.n12912 VSS.n12911 0.00277096
R71653 VSS.n12963 VSS.n12962 0.00277096
R71654 VSS.n16378 VSS.n16377 0.00277096
R71655 VSS.n16100 VSS.n16099 0.00277096
R71656 VSS.n9611 VSS.n9610 0.00277096
R71657 VSS.n9697 VSS.n9696 0.00277096
R71658 VSS.n9306 VSS.n9305 0.00277096
R71659 VSS.n9258 VSS.n9257 0.00277096
R71660 VSS.n15013 VSS.n15012 0.00277096
R71661 VSS.n15062 VSS.n15061 0.00277096
R71662 VSS.n20620 VSS.n20619 0.00277096
R71663 VSS.n20673 VSS.n20672 0.00277096
R71664 VSS.n21186 VSS.n21185 0.00277096
R71665 VSS.n21032 VSS.n21031 0.00277096
R71666 VSS.n6925 VSS.n6924 0.00277096
R71667 VSS.n6990 VSS.n6989 0.00277096
R71668 VSS.n6666 VSS.n6665 0.00277096
R71669 VSS.n6630 VSS.n6629 0.00277096
R71670 VSS.n6578 VSS.n6577 0.00277096
R71671 VSS.n20621 VSS.n20620 0.00277096
R71672 VSS.n20672 VSS.n20671 0.00277096
R71673 VSS.n20129 VSS.n20128 0.00277096
R71674 VSS.n20076 VSS.n20075 0.00277096
R71675 VSS.n1461 VSS.n1460 0.00277096
R71676 VSS.n1078 VSS.n1077 0.00277096
R71677 VSS.n6802 VSS.n6801 0.00277096
R71678 VSS.n6888 VSS.n6887 0.00277096
R71679 VSS.n6516 VSS.n6515 0.00277096
R71680 VSS.n6480 VSS.n6479 0.00277096
R71681 VSS.n6428 VSS.n6427 0.00277096
R71682 VSS.n20128 VSS.n20127 0.00277096
R71683 VSS.n20077 VSS.n20076 0.00277096
R71684 VSS.n1462 VSS.n1461 0.00277096
R71685 VSS.n12818 VSS.n12817 0.00277096
R71686 VSS.n21187 VSS.n21186 0.00277096
R71687 VSS.n21624 VSS.n21623 0.00277096
R71688 VSS.n21381 VSS.n21380 0.00277096
R71689 VSS.n21328 VSS.n21327 0.00277096
R71690 VSS.n7617 VSS.n7616 0.00277096
R71691 VSS.n7669 VSS.n7668 0.00277096
R71692 VSS.n7705 VSS.n7704 0.00277096
R71693 VSS.n7757 VSS.n7756 0.00277096
R71694 VSS.n7834 VSS.n7833 0.00277096
R71695 VSS.n7782 VSS.n7781 0.00277096
R71696 VSS.n21329 VSS.n21328 0.00277096
R71697 VSS.n21380 VSS.n21379 0.00277096
R71698 VSS.n7835 VSS.n7834 0.00277096
R71699 VSS.n6631 VSS.n6630 0.00277096
R71700 VSS.n6481 VSS.n6480 0.00277096
R71701 VSS.n7783 VSS.n7782 0.00277096
R71702 VSS.n6429 VSS.n6428 0.00277096
R71703 VSS.n6579 VSS.n6578 0.00277096
R71704 VSS.n9095 VSS.n9094 0.00277096
R71705 VSS.n9177 VSS.n9176 0.00277096
R71706 VSS.n7756 VSS.n7755 0.00277096
R71707 VSS.n9034 VSS.n9033 0.00277096
R71708 VSS.n7704 VSS.n7703 0.00277096
R71709 VSS.n6991 VSS.n6990 0.00277096
R71710 VSS.n6889 VSS.n6888 0.00277096
R71711 VSS.n6665 VSS.n6664 0.00277096
R71712 VSS.n6515 VSS.n6514 0.00277096
R71713 VSS.n6801 VSS.n6800 0.00277096
R71714 VSS.n6924 VSS.n6923 0.00277096
R71715 VSS.n12695 VSS.n12694 0.00277096
R71716 VSS.n7668 VSS.n7667 0.00277096
R71717 VSS.n7616 VSS.n7615 0.00277096
R71718 VSS.n12746 VSS.n12745 0.00277096
R71719 VSS.n21033 VSS.n21032 0.00277096
R71720 VSS.n1079 VSS.n1078 0.00277096
R71721 VSS.n9610 VSS.n9609 0.00277096
R71722 VSS.n9493 VSS.n9492 0.00277096
R71723 VSS.n16379 VSS.n16378 0.00277096
R71724 VSS.n5878 VSS.n5877 0.00277096
R71725 VSS.n11236 VSS.n11235 0.00277096
R71726 VSS.n6139 VSS.n6138 0.00277096
R71727 VSS.n6058 VSS.n6057 0.00277096
R71728 VSS.n5977 VSS.n5976 0.00277096
R71729 VSS.n11696 VSS.n11695 0.00277096
R71730 VSS.n11647 VSS.n11646 0.00277096
R71731 VSS.n11237 VSS.n11236 0.00277096
R71732 VSS.n6091 VSS.n6090 0.00277096
R71733 VSS.n6010 VSS.n6009 0.00277096
R71734 VSS.n5929 VSS.n5928 0.00277096
R71735 VSS.n21623 VSS.n21622 0.00277096
R71736 VSS.n516 VSS.n515 0.00277096
R71737 VSS.n10611 VSS.n10610 0.00277096
R71738 VSS.n10562 VSS.n10561 0.00277096
R71739 VSS.n10184 VSS.n10183 0.00277096
R71740 VSS.n10185 VSS.n10184 0.00277096
R71741 VSS.n517 VSS.n516 0.00277096
R71742 VSS.n605 VSS.n604 0.00277096
R71743 VSS.n653 VSS.n652 0.00277096
R71744 VSS.n10563 VSS.n10562 0.00277096
R71745 VSS.n15649 VSS.n15648 0.00275919
R71746 VSS.n15622 VSS.n15621 0.00275919
R71747 VSS.n15599 VSS.n15598 0.00275919
R71748 VSS.n15521 VSS.n15520 0.00275919
R71749 VSS.n1740 VSS.n1739 0.00275919
R71750 VSS.n1809 VSS.n1808 0.00275919
R71751 VSS.n1907 VSS.n1906 0.00275919
R71752 VSS.n1890 VSS.n1889 0.00275919
R71753 VSS.n1873 VSS.n1872 0.00275919
R71754 VSS.n18484 VSS.n18482 0.00275
R71755 VSS.n18374 VSS.n18371 0.00275
R71756 VSS.n14963 VSS.n14962 0.00275
R71757 VSS.n14765 VSS.n14764 0.00275
R71758 VSS.n14658 VSS.n14657 0.00275
R71759 VSS.n14932 VSS.n14931 0.00275
R71760 VSS.n16566 VSS.n16565 0.00275
R71761 VSS.n16423 VSS.n16422 0.00275
R71762 DVSS VSS.n7952 0.00275
R71763 VSS.n15898 VSS.n15897 0.00275
R71764 VSS.n5716 VSS.n5715 0.00274945
R71765 VSS.n13246 VSS.n13245 0.00274945
R71766 VSS.n12899 VSS.n12898 0.00274945
R71767 VSS.n12886 VSS.n12885 0.00274945
R71768 VSS.n12832 VSS.n12831 0.00274945
R71769 VSS.n14399 VSS.n14398 0.00274945
R71770 VSS.n14424 VSS.n14423 0.00274945
R71771 VSS.n15073 VSS.n15072 0.00274945
R71772 VSS.n15106 VSS.n15105 0.00274945
R71773 VSS.n15176 VSS.n15175 0.00274945
R71774 VSS.n16358 VSS.n16357 0.00274945
R71775 VSS.n16313 VSS.n16312 0.00274945
R71776 VSS.n16278 VSS.n16277 0.00274945
R71777 VSS.n13363 VSS.n13362 0.00274945
R71778 VSS.n13414 VSS.n13413 0.00274945
R71779 VSS.n20685 VSS.n20684 0.00274945
R71780 VSS.n20736 VSS.n20735 0.00274945
R71781 VSS.n20828 VSS.n20827 0.00274945
R71782 VSS.n21104 VSS.n21103 0.00274945
R71783 VSS.n13506 VSS.n13505 0.00274945
R71784 VSS.n20146 VSS.n20145 0.00274945
R71785 VSS.n2052 VSS.n2051 0.00274945
R71786 VSS.n2045 VSS.n2044 0.00274945
R71787 VSS.n882 VSS.n881 0.00274945
R71788 VSS.n594 VSS.n593 0.00274945
R71789 VSS.n581 VSS.n580 0.00274945
R71790 VSS.n531 VSS.n530 0.00274945
R71791 VSS.n17345 VSS.n17344 0.00274945
R71792 VSS.n17332 VSS.n17331 0.00274945
R71793 VSS.n11521 VSS.n11520 0.00274945
R71794 VSS.n11325 VSS.n11324 0.00274945
R71795 VSS.n11318 VSS.n11317 0.00274945
R71796 VSS.n13330 VSS.n13329 0.00274945
R71797 VSS.n13473 VSS.n13472 0.00274945
R71798 VSS.n21742 VSS.n21735 0.00274945
R71799 VSS.n19027 VSS.n2161 0.00274945
R71800 VSS.n18987 VSS.n18986 0.00274945
R71801 VSS.n4188 VSS.n4187 0.00274945
R71802 VSS.n4163 VSS.n4162 0.00274945
R71803 VSS.n2212 VSS.n2211 0.00274945
R71804 VSS.n5474 VSS.n5473 0.00273544
R71805 VSS.n4919 VSS.n4918 0.00273544
R71806 VSS.n4855 VSS.n4854 0.00273544
R71807 VSS.n14294 VSS.n14293 0.00273544
R71808 VSS.n17307 VSS.n17306 0.00273544
R71809 VSS.n17394 VSS.n2429 0.00273544
R71810 VSS.n5473 VSS.n5472 0.00273544
R71811 VSS.n4918 VSS.n4917 0.00273544
R71812 VSS.n4854 VSS.n4853 0.00273544
R71813 VSS.n14295 VSS.n14294 0.00273544
R71814 VSS.n17306 VSS.n17305 0.00273544
R71815 VSS.n9389 VSS.n9388 0.00272496
R71816 VSS.n9335 VSS.n9334 0.00272496
R71817 VSS.n2508 VSS.n2507 0.00271192
R71818 VSS.n5471 VSS.n5470 0.00271192
R71819 VSS.n4916 VSS.n4915 0.00271192
R71820 VSS.n4852 VSS.n4851 0.00271192
R71821 VSS.n14303 VSS.n14302 0.00271192
R71822 VSS.n17304 VSS.n17303 0.00271192
R71823 VSS.n2422 VSS.n2421 0.00271192
R71824 VSS.n3934 VSS.n3933 0.00271192
R71825 DVSS VSS.n17701 0.0027
R71826 VSS.n15450 VSS.n15449 0.00268951
R71827 VSS.n15449 VSS.n15448 0.00268951
R71828 VSS.n18396 VSS.n18395 0.00268951
R71829 VSS.n15526 VSS.n15525 0.00268951
R71830 VSS.n18397 VSS.n18396 0.00268951
R71831 VSS.n18708 VSS.n18707 0.00268951
R71832 VSS.n15527 VSS.n15526 0.00268951
R71833 VSS.n19626 VSS.n19625 0.00268951
R71834 VSS.n1814 VSS.n1813 0.00268951
R71835 VSS.n1751 VSS.n1750 0.00268951
R71836 VSS.n19625 VSS.n19624 0.00268951
R71837 VSS.n1752 VSS.n1751 0.00268951
R71838 VSS.n19190 VSS.n19189 0.00268951
R71839 VSS.n1815 VSS.n1814 0.00268951
R71840 VSS.n18840 VSS.n18839 0.00268887
R71841 VSS.n15650 VSS.n15649 0.00268887
R71842 VSS.n15623 VSS.n15622 0.00268887
R71843 VSS.n15600 VSS.n15599 0.00268887
R71844 VSS.n19512 VSS.n19511 0.00268887
R71845 VSS.n1908 VSS.n1907 0.00268887
R71846 VSS.n1891 VSS.n1890 0.00268887
R71847 VSS.n1874 VSS.n1873 0.00268887
R71848 VSS.n17583 VSS.n17582 0.00268571
R71849 VSS.n13087 VSS.n13086 0.00268307
R71850 VSS.n21860 VSS.n21859 0.00268307
R71851 VSS.n19145 VSS.n19144 0.00268307
R71852 VSS.n3965 VSS.n3964 0.00268244
R71853 VSS.n11561 VSS.n11560 0.00268244
R71854 VSS.n11566 VSS.n11565 0.00268244
R71855 VSS.n5544 VSS.n5543 0.00268244
R71856 VSS.n9553 VSS.n9552 0.00268244
R71857 VSS.n9116 VSS.n9115 0.00268244
R71858 VSS.n11560 VSS.n11559 0.00268244
R71859 VSS.n3966 VSS.n3965 0.00268244
R71860 VSS.n13115 VSS.n13114 0.00268244
R71861 VSS.n13118 VSS.n13117 0.00268244
R71862 VSS.n12941 VSS.n12940 0.00268244
R71863 VSS.n12933 VSS.n12932 0.00268244
R71864 VSS.n12723 VSS.n12722 0.00268244
R71865 VSS.n12717 VSS.n12716 0.00268244
R71866 VSS.n12318 VSS.n12317 0.00268244
R71867 VSS.n11868 VSS.n11867 0.00268244
R71868 VSS.n12942 VSS.n12941 0.00268244
R71869 VSS.n12934 VSS.n12933 0.00268244
R71870 VSS.n13119 VSS.n13118 0.00268244
R71871 VSS.n13114 VSS.n13113 0.00268244
R71872 VSS.n18960 VSS.n18959 0.00268244
R71873 VSS.n15041 VSS.n15040 0.00268244
R71874 VSS.n9670 VSS.n9669 0.00268244
R71875 VSS.n9279 VSS.n9278 0.00268244
R71876 VSS.n15034 VSS.n15033 0.00268244
R71877 VSS.n15040 VSS.n15039 0.00268244
R71878 VSS.n18959 VSS.n18958 0.00268244
R71879 VSS.n21763 VSS.n21762 0.00268244
R71880 VSS.n21760 VSS.n21759 0.00268244
R71881 VSS.n20643 VSS.n20642 0.00268244
R71882 VSS.n20651 VSS.n20650 0.00268244
R71883 VSS.n20994 VSS.n20993 0.00268244
R71884 VSS.n20987 VSS.n20986 0.00268244
R71885 VSS.n6968 VSS.n6967 0.00268244
R71886 VSS.n6960 VSS.n6959 0.00268244
R71887 VSS.n6608 VSS.n6607 0.00268244
R71888 VSS.n6600 VSS.n6599 0.00268244
R71889 VSS.n20642 VSS.n20641 0.00268244
R71890 VSS.n20650 VSS.n20649 0.00268244
R71891 VSS.n21759 VSS.n21758 0.00268244
R71892 VSS.n21764 VSS.n21763 0.00268244
R71893 VSS.n19048 VSS.n19047 0.00268244
R71894 VSS.n19045 VSS.n19044 0.00268244
R71895 VSS.n20106 VSS.n20105 0.00268244
R71896 VSS.n20098 VSS.n20097 0.00268244
R71897 VSS.n1037 VSS.n1036 0.00268244
R71898 VSS.n1029 VSS.n1028 0.00268244
R71899 VSS.n6866 VSS.n6865 0.00268244
R71900 VSS.n6858 VSS.n6857 0.00268244
R71901 VSS.n6458 VSS.n6457 0.00268244
R71902 VSS.n6450 VSS.n6449 0.00268244
R71903 VSS.n20107 VSS.n20106 0.00268244
R71904 VSS.n20099 VSS.n20098 0.00268244
R71905 VSS.n19044 VSS.n19043 0.00268244
R71906 VSS.n19049 VSS.n19048 0.00268244
R71907 VSS.n21358 VSS.n21357 0.00268244
R71908 VSS.n21350 VSS.n21349 0.00268244
R71909 VSS.n7639 VSS.n7638 0.00268244
R71910 VSS.n7646 VSS.n7645 0.00268244
R71911 VSS.n7727 VSS.n7726 0.00268244
R71912 VSS.n7735 VSS.n7734 0.00268244
R71913 VSS.n7812 VSS.n7811 0.00268244
R71914 VSS.n7804 VSS.n7803 0.00268244
R71915 VSS.n21359 VSS.n21358 0.00268244
R71916 VSS.n21351 VSS.n21350 0.00268244
R71917 VSS.n9285 VSS.n9284 0.00268244
R71918 VSS.n11869 VSS.n11868 0.00268244
R71919 VSS.n7813 VSS.n7812 0.00268244
R71920 VSS.n9122 VSS.n9121 0.00268244
R71921 VSS.n7805 VSS.n7804 0.00268244
R71922 VSS.n11853 VSS.n11852 0.00268244
R71923 VSS.n6601 VSS.n6600 0.00268244
R71924 VSS.n6451 VSS.n6450 0.00268244
R71925 VSS.n6609 VSS.n6608 0.00268244
R71926 VSS.n6459 VSS.n6458 0.00268244
R71927 VSS.n9676 VSS.n9675 0.00268244
R71928 VSS.n7726 VSS.n7725 0.00268244
R71929 VSS.n9559 VSS.n9558 0.00268244
R71930 VSS.n12319 VSS.n12318 0.00268244
R71931 VSS.n7734 VSS.n7733 0.00268244
R71932 VSS.n6961 VSS.n6960 0.00268244
R71933 VSS.n6859 VSS.n6858 0.00268244
R71934 VSS.n6969 VSS.n6968 0.00268244
R71935 VSS.n6867 VSS.n6866 0.00268244
R71936 VSS.n5550 VSS.n5549 0.00268244
R71937 VSS.n20986 VSS.n20985 0.00268244
R71938 VSS.n20995 VSS.n20994 0.00268244
R71939 VSS.n12724 VSS.n12723 0.00268244
R71940 VSS.n12716 VSS.n12715 0.00268244
R71941 VSS.n7647 VSS.n7646 0.00268244
R71942 VSS.n16054 VSS.n16053 0.00268244
R71943 VSS.n1028 VSS.n1027 0.00268244
R71944 VSS.n7638 VSS.n7637 0.00268244
R71945 VSS.n16060 VSS.n16059 0.00268244
R71946 VSS.n1036 VSS.n1035 0.00268244
R71947 VSS.n11668 VSS.n11667 0.00268244
R71948 VSS.n6112 VSS.n6111 0.00268244
R71949 VSS.n6031 VSS.n6030 0.00268244
R71950 VSS.n5950 VSS.n5949 0.00268244
R71951 VSS.n11675 VSS.n11674 0.00268244
R71952 VSS.n6118 VSS.n6117 0.00268244
R71953 VSS.n6037 VSS.n6036 0.00268244
R71954 VSS.n5956 VSS.n5955 0.00268244
R71955 VSS.n11669 VSS.n11668 0.00268244
R71956 VSS.n2599 VSS.n2598 0.00268244
R71957 VSS.n2600 VSS.n2599 0.00268244
R71958 VSS.n626 VSS.n625 0.00268244
R71959 VSS.n10584 VSS.n10583 0.00268244
R71960 VSS.n10265 VSS.n10264 0.00268244
R71961 VSS.n8792 VSS.n8791 0.00268244
R71962 VSS.n10590 VSS.n10589 0.00268244
R71963 VSS.n8797 VSS.n8796 0.00268244
R71964 VSS.n632 VSS.n631 0.00268244
R71965 VSS.n1243 VSS.n1242 0.00267491
R71966 VSS.n1245 VSS.n1243 0.00267491
R71967 VSS.n6770 VSS.n6769 0.00266496
R71968 VSS.n6710 VSS.n6709 0.00266496
R71969 VSS.n20398 VSS.n20397 0.00263
R71970 VSS.n20367 VSS.n20366 0.00263
R71971 VSS.n20337 VSS.n20336 0.00263
R71972 VSS.n20291 VSS.n20290 0.00263
R71973 VSS.n8815 VSS.n8814 0.00263
R71974 VSS.n9427 VSS.n9426 0.00263
R71975 VSS.n9803 VSS.n6163 0.00263
R71976 VSS.n2362 VSS.n2361 0.00262598
R71977 VSS.n17469 VSS.n17468 0.00262598
R71978 VSS.n11368 VSS.n11367 0.00262598
R71979 VSS.n5849 VSS.n5848 0.00262598
R71980 VSS.n5725 VSS.n5724 0.00262598
R71981 VSS.n5626 VSS.n5625 0.00262598
R71982 VSS.n5603 VSS.n5602 0.00262598
R71983 VSS.n13172 VSS.n13171 0.00262598
R71984 VSS.n12839 VSS.n12838 0.00262598
R71985 VSS.n12776 VSS.n12775 0.00262598
R71986 VSS.n12691 VSS.n12690 0.00262598
R71987 VSS.n12603 VSS.n12602 0.00262598
R71988 VSS.n12585 VSS.n12584 0.00262598
R71989 VSS.n12580 VSS.n12579 0.00262598
R71990 VSS.n12324 VSS.n12323 0.00262598
R71991 VSS.n11862 VSS.n11861 0.00262598
R71992 VSS.n11829 VSS.n11828 0.00262598
R71993 VSS.n2261 VSS.n2260 0.00262598
R71994 VSS.n2220 VSS.n2219 0.00262598
R71995 VSS.n15169 VSS.n15168 0.00262598
R71996 VSS.n16210 VSS.n16209 0.00262598
R71997 VSS.n16173 VSS.n16172 0.00262598
R71998 VSS.n16148 VSS.n16147 0.00262598
R71999 VSS.n16119 VSS.n16118 0.00262598
R72000 VSS.n2312 VSS.n2311 0.00262598
R72001 VSS.n20821 VSS.n20820 0.00262598
R72002 VSS.n21152 VSS.n21151 0.00262598
R72003 VSS.n21113 VSS.n21112 0.00262598
R72004 VSS.n21076 VSS.n21075 0.00262598
R72005 VSS.n21053 VSS.n21052 0.00262598
R72006 VSS.n17920 VSS.n17919 0.00262598
R72007 VSS.n1998 VSS.n1997 0.00262598
R72008 VSS.n1281 VSS.n1280 0.00262598
R72009 VSS.n1163 VSS.n1162 0.00262598
R72010 VSS.n1128 VSS.n1127 0.00262598
R72011 VSS.n1099 VSS.n1098 0.00262598
R72012 VSS.n21664 VSS.n21663 0.00262598
R72013 VSS.n21501 VSS.n21500 0.00262598
R72014 VSS.n21433 VSS.n21432 0.00262598
R72015 VSS.n21260 VSS.n21259 0.00262598
R72016 VSS.n7586 VSS.n7585 0.00262598
R72017 VSS.n4125 VSS.n4124 0.00262598
R72018 VSS.n4715 VSS.n4714 0.00262598
R72019 VSS.n17389 VSS.n17388 0.00262598
R72020 VSS.n11420 VSS.n11419 0.00262598
R72021 VSS.n11199 VSS.n11198 0.00262598
R72022 VSS.n538 VSS.n537 0.00262598
R72023 VSS.n479 VSS.n478 0.00262598
R72024 VSS.n10559 VSS.n10558 0.00262598
R72025 VSS.n10537 VSS.n10536 0.00262598
R72026 VSS.n10520 VSS.n10519 0.00262598
R72027 VSS.n10515 VSS.n10514 0.00262598
R72028 VSS.n10270 VSS.n10269 0.00262598
R72029 VSS.n8977 VSS.n8976 0.00262598
R72030 VSS.n8989 VSS.n8988 0.00262598
R72031 VSS.n10314 VSS.n10313 0.00261538
R72032 VSS.n10432 VSS.n10431 0.00261538
R72033 VSS.n10340 VSS.n10339 0.00261538
R72034 VSS.n10147 VSS.n10146 0.00261538
R72035 VSS.n10055 VSS.n10054 0.00261538
R72036 VSS.n10030 VSS.n10025 0.00261538
R72037 VSS.n12368 VSS.n12367 0.00261538
R72038 VSS.n12486 VSS.n12485 0.00261538
R72039 VSS.n12394 VSS.n12393 0.00261538
R72040 VSS.n12198 VSS.n12197 0.00261538
R72041 VSS.n12106 VSS.n12105 0.00261538
R72042 VSS.n12081 VSS.n12076 0.00261538
R72043 VSS.n18476 VSS.n18475 0.00261268
R72044 VSS.n18402 VSS.n18401 0.00261268
R72045 VSS.n18401 VSS.n18400 0.00261268
R72046 VSS.n14574 VSS.n14573 0.00261268
R72047 VSS.n14821 VSS.n14820 0.00261268
R72048 VSS.n17122 VSS.n17121 0.00261268
R72049 VSS.n17118 VSS.n17117 0.00261268
R72050 VSS.n17072 VSS.n17071 0.00261268
R72051 VSS.n14867 VSS.n14866 0.00261268
R72052 VSS.n14887 VSS.n14886 0.00261268
R72053 VSS.n16896 VSS.n16895 0.00261268
R72054 VSS.n16698 VSS.n16697 0.00261268
R72055 VSS.n16536 VSS.n16535 0.00261268
R72056 VSS.n16447 VSS.n16446 0.00261268
R72057 VSS.n15862 VSS.n15861 0.00261268
R72058 VSS.n15531 VSS.n15530 0.00261268
R72059 VSS.n15473 VSS.n15472 0.00261268
R72060 VSS.n15398 VSS.n15397 0.00261268
R72061 VSS.n15367 VSS.n15366 0.00261268
R72062 VSS.n15333 VSS.n15332 0.00261268
R72063 VSS.n8569 VSS.n8568 0.00261268
R72064 VSS.n8424 VSS.n8423 0.00261268
R72065 VSS.n19563 VSS.n19562 0.00261268
R72066 VSS.n19620 VSS.n19619 0.00261268
R72067 VSS.n19621 VSS.n19620 0.00261268
R72068 VSS.n19754 VSS.n19753 0.00261268
R72069 VSS.n19844 VSS.n19843 0.00261268
R72070 VSS.n19873 VSS.n19872 0.00261268
R72071 VSS.n19877 VSS.n19876 0.00261268
R72072 VSS.n19893 VSS.n19892 0.00261268
R72073 VSS.n19938 VSS.n19937 0.00261268
R72074 VSS.n19958 VSS.n19957 0.00261268
R72075 VSS.n20020 VSS.n20019 0.00261268
R72076 VSS.n2100 VSS.n2099 0.00261268
R72077 VSS.n802 VSS.n801 0.00261268
R72078 VSS.n842 VSS.n841 0.00261268
R72079 VSS.n1938 VSS.n1937 0.00261268
R72080 VSS.n1819 VSS.n1818 0.00261268
R72081 VSS.n1775 VSS.n1774 0.00261268
R72082 VSS.n1714 VSS.n1713 0.00261268
R72083 VSS.n1683 VSS.n1682 0.00261268
R72084 VSS.n1649 VSS.n1648 0.00261268
R72085 VSS.n8720 VSS.n8719 0.00261268
R72086 VSS.n8232 VSS.n8231 0.00261268
R72087 VSS.n9777 VSS.n9776 0.00260496
R72088 VSS.n9723 VSS.n9722 0.00260496
R72089 VSS.n20167 VSS.n733 0.0026
R72090 VSS.n20590 VSS.n20589 0.0026
R72091 VSS.n20567 VSS.n20566 0.0026
R72092 VSS.n20544 VSS.n20543 0.0026
R72093 VSS.n7851 VSS.n7045 0.0026
R72094 VSS.n5846 VSS.n5845 0.00259448
R72095 VSS.n16207 VSS.n16206 0.00259448
R72096 VSS.n21149 VSS.n21148 0.00259448
R72097 VSS.n1278 VSS.n1277 0.00259448
R72098 VSS.n21018 VSS.n21017 0.00259404
R72099 VSS.n1064 VSS.n1063 0.00259404
R72100 VSS.n4061 VSS.n4060 0.00259392
R72101 VSS.n11533 VSS.n11532 0.00259392
R72102 VSS.n5590 VSS.n5589 0.00259392
R72103 VSS.n9586 VSS.n9585 0.00259392
R72104 VSS.n9149 VSS.n9148 0.00259392
R72105 VSS.n11532 VSS.n11531 0.00259392
R72106 VSS.n4060 VSS.n4059 0.00259392
R72107 VSS.n13089 VSS.n13088 0.00259392
R72108 VSS.n12971 VSS.n12970 0.00259392
R72109 VSS.n12753 VSS.n12752 0.00259392
R72110 VSS.n12532 VSS.n12531 0.00259392
R72111 VSS.n12260 VSS.n12259 0.00259392
R72112 VSS.n12972 VSS.n12971 0.00259392
R72113 VSS.n13088 VSS.n13087 0.00259392
R72114 VSS.n18932 VSS.n18931 0.00259392
R72115 VSS.n15007 VSS.n15006 0.00259392
R72116 VSS.n16106 VSS.n16105 0.00259392
R72117 VSS.n9703 VSS.n9702 0.00259392
R72118 VSS.n9312 VSS.n9311 0.00259392
R72119 VSS.n15006 VSS.n15005 0.00259392
R72120 VSS.n18931 VSS.n18930 0.00259392
R72121 VSS.n21862 VSS.n21861 0.00259392
R72122 VSS.n20613 VSS.n20612 0.00259392
R72123 VSS.n21040 VSS.n21039 0.00259392
R72124 VSS.n6998 VSS.n6997 0.00259392
R72125 VSS.n6638 VSS.n6637 0.00259392
R72126 VSS.n20612 VSS.n20611 0.00259392
R72127 VSS.n21861 VSS.n21860 0.00259392
R72128 VSS.n19147 VSS.n19146 0.00259392
R72129 VSS.n20136 VSS.n20135 0.00259392
R72130 VSS.n1086 VSS.n1085 0.00259392
R72131 VSS.n6896 VSS.n6895 0.00259392
R72132 VSS.n6488 VSS.n6487 0.00259392
R72133 VSS.n20137 VSS.n20136 0.00259392
R72134 VSS.n19146 VSS.n19145 0.00259392
R72135 VSS.n21636 VSS.n21635 0.00259392
R72136 VSS.n21660 VSS.n21659 0.00259392
R72137 VSS.n21466 VSS.n21465 0.00259392
R72138 VSS.n21444 VSS.n21443 0.00259392
R72139 VSS.n21388 VSS.n21387 0.00259392
R72140 VSS.n7609 VSS.n7608 0.00259392
R72141 VSS.n7697 VSS.n7696 0.00259392
R72142 VSS.n7842 VSS.n7841 0.00259392
R72143 VSS.n21389 VSS.n21388 0.00259392
R72144 VSS.n21445 VSS.n21444 0.00259392
R72145 VSS.n21467 VSS.n21466 0.00259392
R72146 VSS.n9313 VSS.n9312 0.00259392
R72147 VSS.n7843 VSS.n7842 0.00259392
R72148 VSS.n9150 VSS.n9149 0.00259392
R72149 VSS.n6639 VSS.n6638 0.00259392
R72150 VSS.n6489 VSS.n6488 0.00259392
R72151 VSS.n9704 VSS.n9703 0.00259392
R72152 VSS.n7696 VSS.n7695 0.00259392
R72153 VSS.n12533 VSS.n12532 0.00259392
R72154 VSS.n12261 VSS.n12260 0.00259392
R72155 VSS.n9587 VSS.n9586 0.00259392
R72156 VSS.n6897 VSS.n6896 0.00259392
R72157 VSS.n6999 VSS.n6998 0.00259392
R72158 VSS.n7608 VSS.n7607 0.00259392
R72159 VSS.n12754 VSS.n12753 0.00259392
R72160 VSS.n16107 VSS.n16106 0.00259392
R72161 VSS.n5591 VSS.n5590 0.00259392
R72162 VSS.n21041 VSS.n21040 0.00259392
R72163 VSS.n1087 VSS.n1086 0.00259392
R72164 VSS.n3865 VSS.n3864 0.00259392
R72165 VSS.n4121 VSS.n4120 0.00259392
R72166 VSS.n4791 VSS.n4790 0.00259392
R72167 VSS.n11702 VSS.n11701 0.00259392
R72168 VSS.n6145 VSS.n6144 0.00259392
R72169 VSS.n6064 VSS.n6063 0.00259392
R72170 VSS.n5983 VSS.n5982 0.00259392
R72171 VSS.n3864 VSS.n3863 0.00259392
R72172 VSS.n11703 VSS.n11702 0.00259392
R72173 VSS.n6146 VSS.n6145 0.00259392
R72174 VSS.n6065 VSS.n6064 0.00259392
R72175 VSS.n5984 VSS.n5983 0.00259392
R72176 VSS.n4790 VSS.n4789 0.00259392
R72177 VSS.n21659 VSS.n21658 0.00259392
R72178 VSS.n4120 VSS.n3887 0.00259392
R72179 VSS.n2627 VSS.n2626 0.00259392
R72180 VSS.n2628 VSS.n2627 0.00259392
R72181 VSS.n659 VSS.n658 0.00259392
R72182 VSS.n10617 VSS.n10616 0.00259392
R72183 VSS.n10477 VSS.n10476 0.00259392
R72184 VSS.n10208 VSS.n10207 0.00259392
R72185 VSS.n10478 VSS.n10477 0.00259392
R72186 VSS.n10209 VSS.n10208 0.00259392
R72187 VSS.n10618 VSS.n10617 0.00259392
R72188 VSS.n660 VSS.n659 0.00259392
R72189 VSS.n14857 VSS.n14856 0.00258439
R72190 VSS.n19928 VSS.n19927 0.00258439
R72191 VSS.n18799 VSS.n18798 0.00258431
R72192 VSS.n19471 VSS.n19470 0.00258431
R72193 VSS.n17019 VSS.n17018 0.00258395
R72194 VSS.n16538 VSS.n16537 0.00258395
R72195 VSS.n19916 VSS.n19915 0.00258395
R72196 VSS.n800 VSS.n799 0.00258395
R72197 VSS.n14170 VSS.n14169 0.00257445
R72198 VSS.n14133 VSS.n14132 0.00257445
R72199 VSS.n20168 VSS.n20167 0.00257
R72200 VSS.n20590 VSS.n460 0.00257
R72201 VSS.n20568 VSS.n20567 0.00257
R72202 VSS.n20545 VSS.n20544 0.00257
R72203 VSS.n7852 VSS.n7851 0.00257
R72204 VSS.n7949 VSS.n7948 0.00257
R72205 VSS.n6375 VSS.n6374 0.00257
R72206 VSS.n10258 VSS.n10257 0.00256281
R72207 VSS.n17449 VSS.n17448 0.00253439
R72208 VSS.n17440 VSS.n17439 0.00253439
R72209 VSS.n17480 VSS.n17479 0.00253439
R72210 VSS.n17471 VSS.n17470 0.00253439
R72211 VSS.n13233 VSS.n13232 0.00253439
R72212 VSS.n13225 VSS.n13224 0.00253439
R72213 VSS.n13194 VSS.n13193 0.00253439
R72214 VSS.n13203 VSS.n13202 0.00253439
R72215 VSS.n2191 VSS.n2190 0.00253439
R72216 VSS.n13350 VSS.n13349 0.00253439
R72217 VSS.n13493 VSS.n13492 0.00253439
R72218 VSS.n19256 VSS.n19255 0.002525
R72219 VSS.n19263 VSS.n19260 0.002525
R72220 VSS.n16982 VSS.n16981 0.002525
R72221 VSS.n16978 VSS.n16977 0.002525
R72222 VSS.n170 VSS.n169 0.00251117
R72223 VSS.n57 VSS.n56 0.00251117
R72224 VSS.n40 VSS.n37 0.00251117
R72225 VSS.n205 VSS.n203 0.00251117
R72226 VSS.n223 VSS.n222 0.00251117
R72227 VSS.n333 VSS.n332 0.00251117
R72228 VSS.n20397 VSS.n20396 0.00251
R72229 VSS.n20366 VSS.n20365 0.00251
R72230 VSS.n20336 VSS.n20335 0.00251
R72231 VSS.n20290 VSS.n20289 0.00251
R72232 VSS.n8817 VSS.n8815 0.00251
R72233 VSS.n8848 VSS.n8847 0.00251
R72234 VSS.n9430 VSS.n9427 0.00251
R72235 VSS.n9451 VSS.n9450 0.00251
R72236 VSS.n9805 VSS.n9803 0.00251
R72237 VSS.n9825 VSS.n9824 0.00251
R72238 VSS.n13117 VSS.n13116 0.0025059
R72239 VSS.n21761 VSS.n21760 0.0025059
R72240 VSS.n19046 VSS.n19045 0.0025059
R72241 VSS.n4028 VSS.n4027 0.0025054
R72242 VSS.n4202 VSS.n4201 0.0025054
R72243 VSS.n2372 VSS.n2371 0.0025054
R72244 VSS.n11340 VSS.n11339 0.0025054
R72245 VSS.n5857 VSS.n5856 0.0025054
R72246 VSS.n4201 VSS.n4200 0.0025054
R72247 VSS.n11341 VSS.n11340 0.0025054
R72248 VSS.n4027 VSS.n4026 0.0025054
R72249 VSS.n5856 VSS.n5855 0.0025054
R72250 VSS.n13055 VSS.n13054 0.0025054
R72251 VSS.n13141 VSS.n13140 0.0025054
R72252 VSS.n13184 VSS.n13183 0.0025054
R72253 VSS.n12868 VSS.n12867 0.0025054
R72254 VSS.n12805 VSS.n12804 0.0025054
R72255 VSS.n13140 VSS.n13139 0.0025054
R72256 VSS.n12869 VSS.n12868 0.0025054
R72257 VSS.n13054 VSS.n13053 0.0025054
R72258 VSS.n12806 VSS.n12805 0.0025054
R72259 VSS.n2371 VSS.n2370 0.0025054
R72260 VSS.n13183 VSS.n13182 0.0025054
R72261 VSS.n18899 VSS.n18898 0.0025054
R72262 VSS.n2232 VSS.n2231 0.0025054
R72263 VSS.n2271 VSS.n2270 0.0025054
R72264 VSS.n15142 VSS.n15141 0.0025054
R72265 VSS.n16217 VSS.n16216 0.0025054
R72266 VSS.n2231 VSS.n2230 0.0025054
R72267 VSS.n15141 VSS.n15140 0.0025054
R72268 VSS.n2270 VSS.n2269 0.0025054
R72269 VSS.n18898 VSS.n18897 0.0025054
R72270 VSS.n16218 VSS.n16217 0.0025054
R72271 VSS.n21828 VSS.n21827 0.0025054
R72272 VSS.n2281 VSS.n2280 0.0025054
R72273 VSS.n2324 VSS.n2323 0.0025054
R72274 VSS.n20792 VSS.n20791 0.0025054
R72275 VSS.n21159 VSS.n21158 0.0025054
R72276 VSS.n2280 VSS.n2279 0.0025054
R72277 VSS.n20791 VSS.n20790 0.0025054
R72278 VSS.n21827 VSS.n21826 0.0025054
R72279 VSS.n2323 VSS.n2322 0.0025054
R72280 VSS.n21160 VSS.n21159 0.0025054
R72281 VSS.n19113 VSS.n19112 0.0025054
R72282 VSS.n17889 VSS.n17888 0.0025054
R72283 VSS.n17932 VSS.n17931 0.0025054
R72284 VSS.n2027 VSS.n2026 0.0025054
R72285 VSS.n1288 VSS.n1287 0.0025054
R72286 VSS.n17888 VSS.n17887 0.0025054
R72287 VSS.n2028 VSS.n2027 0.0025054
R72288 VSS.n19112 VSS.n19111 0.0025054
R72289 VSS.n17931 VSS.n17930 0.0025054
R72290 VSS.n1289 VSS.n1288 0.0025054
R72291 VSS.n21599 VSS.n21598 0.0025054
R72292 VSS.n21655 VSS.n21654 0.0025054
R72293 VSS.n21489 VSS.n21488 0.0025054
R72294 VSS.n21289 VSS.n21288 0.0025054
R72295 VSS.n7557 VSS.n7556 0.0025054
R72296 VSS.n21290 VSS.n21289 0.0025054
R72297 VSS.n21654 VSS.n21653 0.0025054
R72298 VSS.n21598 VSS.n21597 0.0025054
R72299 VSS.n21490 VSS.n21489 0.0025054
R72300 VSS.n7556 VSS.n7555 0.0025054
R72301 VSS.n3830 VSS.n3829 0.0025054
R72302 VSS.n3884 VSS.n3883 0.0025054
R72303 VSS.n4725 VSS.n4724 0.0025054
R72304 VSS.n11447 VSS.n11446 0.0025054
R72305 VSS.n11226 VSS.n11225 0.0025054
R72306 VSS.n3829 VSS.n3828 0.0025054
R72307 VSS.n3883 VSS.n3882 0.0025054
R72308 VSS.n11448 VSS.n11447 0.0025054
R72309 VSS.n4724 VSS.n4723 0.0025054
R72310 VSS.n11227 VSS.n11226 0.0025054
R72311 VSS.n2645 VSS.n2644 0.0025054
R72312 VSS.n2644 VSS.n2643 0.0025054
R72313 VSS.n565 VSS.n564 0.0025054
R72314 VSS.n506 VSS.n505 0.0025054
R72315 VSS.n566 VSS.n565 0.0025054
R72316 VSS.n507 VSS.n506 0.0025054
R72317 VSS.n2509 VSS.n2508 0.00248147
R72318 VSS.n3935 VSS.n3934 0.00248147
R72319 VSS.n5472 VSS.n5471 0.00248147
R72320 VSS.n4917 VSS.n4916 0.00248147
R72321 VSS.n4853 VSS.n4852 0.00248147
R72322 VSS.n14303 VSS.n14295 0.00248147
R72323 VSS.n17305 VSS.n17304 0.00248147
R72324 VSS.n2423 VSS.n2422 0.00248147
R72325 VSS.n7875 VSS.n7874 0.00248
R72326 VSS.n7968 VSS.n7967 0.00248
R72327 VSS.n11061 VSS.n11060 0.00248
R72328 VSS.n18423 VSS.n18422 0.00247852
R72329 VSS.n19606 VSS.n19605 0.00247852
R72330 VSS.n18738 VSS.n18737 0.00247839
R72331 VSS.n8510 VSS.n8509 0.00247839
R72332 VSS.n16905 VSS.n16904 0.00247839
R72333 VSS.n16598 VSS.n16597 0.00247839
R72334 VSS.n18737 VSS.n18736 0.00247839
R72335 VSS.n19220 VSS.n19219 0.00247839
R72336 VSS.n770 VSS.n769 0.00247839
R72337 VSS.n8661 VSS.n8660 0.00247839
R72338 VSS.n20011 VSS.n20010 0.00247839
R72339 VSS.n19219 VSS.n19218 0.00247839
R72340 VSS.n8511 VSS.n8510 0.00247839
R72341 VSS.n8662 VSS.n8661 0.00247839
R72342 VSS.n17346 VSS.n17345 0.00247541
R72343 VSS.n17331 VSS.n17330 0.00247541
R72344 VSS.n11520 VSS.n11519 0.00247541
R72345 VSS.n11326 VSS.n11325 0.00247541
R72346 VSS.n11317 VSS.n11316 0.00247541
R72347 VSS.n4198 VSS.n4188 0.00247541
R72348 VSS.n16357 VSS.n16356 0.00247541
R72349 VSS.n16312 VSS.n16311 0.00247541
R72350 VSS.n16277 VSS.n16276 0.00247541
R72351 VSS.n5838 VSS.n5837 0.00247541
R72352 VSS.n1438 VSS.n1437 0.00247541
R72353 VSS.n1393 VSS.n1392 0.00247541
R72354 VSS.n1358 VSS.n1357 0.00247541
R72355 VSS.n1270 VSS.n1269 0.00247541
R72356 VSS.n1153 VSS.n1152 0.00247541
R72357 VSS.n3676 DVSS 0.00247183
R72358 VSS.n3675 DVSS 0.00247183
R72359 VSS.n4026 VSS.n4025 0.00244882
R72360 VSS.n4203 VSS.n4202 0.00244882
R72361 VSS.n2373 VSS.n2372 0.00244882
R72362 VSS.n17433 VSS.n17432 0.00244882
R72363 VSS.n11342 VSS.n11341 0.00244882
R72364 VSS.n5855 VSS.n5854 0.00244882
R72365 VSS.n5572 VSS.n5571 0.00244882
R72366 VSS.n13053 VSS.n13052 0.00244882
R72367 VSS.n13142 VSS.n13141 0.00244882
R72368 VSS.n13185 VSS.n13184 0.00244882
R72369 VSS.n13239 VSS.n13238 0.00244882
R72370 VSS.n12867 VSS.n12866 0.00244882
R72371 VSS.n12804 VSS.n12803 0.00244882
R72372 VSS.n12517 VSS.n12516 0.00244882
R72373 VSS.n12316 VSS.n12315 0.00244882
R72374 VSS.n12225 VSS.n12224 0.00244882
R72375 VSS.n11963 VSS.n11962 0.00244882
R72376 VSS.n11883 VSS.n11882 0.00244882
R72377 VSS.n11863 VSS.n11862 0.00244882
R72378 VSS.n18897 VSS.n18896 0.00244882
R72379 VSS.n2233 VSS.n2232 0.00244882
R72380 VSS.n2272 VSS.n2271 0.00244882
R72381 VSS.n2184 VSS.n2183 0.00244882
R72382 VSS.n15143 VSS.n15142 0.00244882
R72383 VSS.n16216 VSS.n16215 0.00244882
R72384 VSS.n16088 VSS.n16087 0.00244882
R72385 VSS.n21826 VSS.n21825 0.00244882
R72386 VSS.n2282 VSS.n2281 0.00244882
R72387 VSS.n2325 VSS.n2324 0.00244882
R72388 VSS.n13356 VSS.n13355 0.00244882
R72389 VSS.n20793 VSS.n20792 0.00244882
R72390 VSS.n21158 VSS.n21157 0.00244882
R72391 VSS.n21020 VSS.n21019 0.00244882
R72392 VSS.n19111 VSS.n19110 0.00244882
R72393 VSS.n17890 VSS.n17889 0.00244882
R72394 VSS.n17933 VSS.n17932 0.00244882
R72395 VSS.n13499 VSS.n13498 0.00244882
R72396 VSS.n2026 VSS.n2025 0.00244882
R72397 VSS.n1287 VSS.n1286 0.00244882
R72398 VSS.n1066 VSS.n1065 0.00244882
R72399 VSS.n21597 VSS.n21596 0.00244882
R72400 VSS.n21539 VSS.n21538 0.00244882
R72401 VSS.n21488 VSS.n21487 0.00244882
R72402 VSS.n21475 VSS.n21474 0.00244882
R72403 VSS.n21288 VSS.n21287 0.00244882
R72404 VSS.n7558 VSS.n7557 0.00244882
R72405 VSS.n3828 VSS.n3827 0.00244882
R72406 VSS.n4155 VSS.n4154 0.00244882
R72407 VSS.n4726 VSS.n4725 0.00244882
R72408 VSS.n4762 VSS.n4761 0.00244882
R72409 VSS.n11446 VSS.n11445 0.00244882
R72410 VSS.n11225 VSS.n11224 0.00244882
R72411 VSS.n2643 VSS.n2642 0.00244882
R72412 VSS.n564 VSS.n563 0.00244882
R72413 VSS.n505 VSS.n504 0.00244882
R72414 VSS.n10462 VSS.n10461 0.00244882
R72415 VSS.n10263 VSS.n10262 0.00244882
R72416 VSS.n10173 VSS.n10172 0.00244882
R72417 VSS.n9966 VSS.n9965 0.00244882
R72418 VSS.n8945 VSS.n8944 0.00244882
R72419 VSS.n8976 VSS.n8975 0.00244882
R72420 VSS.n15484 VSS.n15483 0.00243571
R72421 VSS.n1220 VSS.n1219 0.00243571
R72422 VSS.n15483 VSS.n15482 0.00243571
R72423 VSS.n1222 VSS.n1220 0.00243571
R72424 VSS.n5767 VSS.n5766 0.00243571
R72425 VSS.n5819 VSS.n5818 0.00243571
R72426 VSS.n5813 VSS.n5812 0.00243571
R72427 VSS.n1191 VSS.n1190 0.00243571
R72428 VSS.n1251 VSS.n1250 0.00243571
R72429 VSS.n5814 VSS.n5813 0.00243571
R72430 VSS.n5822 VSS.n5819 0.00243571
R72431 VSS.n5770 VSS.n5767 0.00243571
R72432 VSS.n1252 VSS.n1251 0.00243571
R72433 VSS.n1194 VSS.n1191 0.00243571
R72434 VSS.n2690 VSS.n2689 0.00242857
R72435 VSS.n2734 VSS.n2733 0.00242857
R72436 VSS.n2794 VSS.n2793 0.00242857
R72437 VSS.n17536 VSS.n17535 0.00242857
R72438 VSS.n18102 VSS.n18101 0.00242857
R72439 VSS.n8434 VSS.n8433 0.00242
R72440 VSS.n7899 VSS.n7897 0.00242
R72441 VSS.n8766 VSS.n8765 0.00242
R72442 VSS.n7992 VSS.n7990 0.00242
R72443 VSS.n10817 VSS.n10816 0.00242
R72444 VSS.n11037 VSS.n11036 0.00242
R72445 VSS.n5843 VSS.n5842 0.00241688
R72446 VSS.n5570 VSS.n5569 0.00241688
R72447 VSS.n13171 VSS.n13170 0.00241688
R72448 VSS.n12840 VSS.n12839 0.00241688
R72449 VSS.n12581 VSS.n12580 0.00241688
R72450 VSS.n12515 VSS.n12514 0.00241688
R72451 VSS.n11860 VSS.n11859 0.00241688
R72452 VSS.n11830 VSS.n11829 0.00241688
R72453 VSS.n13170 VSS.n13169 0.00241688
R72454 VSS.n12841 VSS.n12840 0.00241688
R72455 VSS.n2260 VSS.n2259 0.00241688
R72456 VSS.n15168 VSS.n15167 0.00241688
R72457 VSS.n16204 VSS.n16203 0.00241688
R72458 VSS.n16086 VSS.n16085 0.00241688
R72459 VSS.n2259 VSS.n2258 0.00241688
R72460 VSS.n15167 VSS.n15166 0.00241688
R72461 VSS.n5844 VSS.n5843 0.00241688
R72462 VSS.n16205 VSS.n16204 0.00241688
R72463 VSS.n2311 VSS.n2310 0.00241688
R72464 VSS.n20820 VSS.n20819 0.00241688
R72465 VSS.n21146 VSS.n21145 0.00241688
R72466 VSS.n2310 VSS.n2309 0.00241688
R72467 VSS.n20819 VSS.n20818 0.00241688
R72468 VSS.n21147 VSS.n21146 0.00241688
R72469 VSS.n17919 VSS.n17918 0.00241688
R72470 VSS.n1999 VSS.n1998 0.00241688
R72471 VSS.n1275 VSS.n1274 0.00241688
R72472 VSS.n1164 VSS.n1163 0.00241688
R72473 VSS.n17918 VSS.n17917 0.00241688
R72474 VSS.n2000 VSS.n1999 0.00241688
R72475 VSS.n1276 VSS.n1275 0.00241688
R72476 VSS.n1165 VSS.n1164 0.00241688
R72477 VSS.n21542 VSS.n21541 0.00241688
R72478 VSS.n21502 VSS.n21501 0.00241688
R72479 VSS.n21434 VSS.n21433 0.00241688
R72480 VSS.n21261 VSS.n21260 0.00241688
R72481 VSS.n21435 VSS.n21434 0.00241688
R72482 VSS.n21543 VSS.n21542 0.00241688
R72483 VSS.n21503 VSS.n21502 0.00241688
R72484 VSS.n21262 VSS.n21261 0.00241688
R72485 VSS.n21563 VSS.n21562 0.00241688
R72486 VSS.n11831 VSS.n11830 0.00241688
R72487 VSS.n11861 VSS.n11860 0.00241688
R72488 VSS.n12582 VSS.n12581 0.00241688
R72489 VSS.n12514 VSS.n12513 0.00241688
R72490 VSS.n5571 VSS.n5570 0.00241688
R72491 VSS.n16087 VSS.n16086 0.00241688
R72492 VSS.n21019 VSS.n21018 0.00241688
R72493 VSS.n1065 VSS.n1064 0.00241688
R72494 VSS.n3796 VSS.n3795 0.00241688
R72495 VSS.n4158 VSS.n4157 0.00241688
R72496 VSS.n4714 VSS.n4713 0.00241688
R72497 VSS.n17390 VSS.n17389 0.00241688
R72498 VSS.n11421 VSS.n11420 0.00241688
R72499 VSS.n11200 VSS.n11199 0.00241688
R72500 VSS.n4159 VSS.n4158 0.00241688
R72501 VSS.n4713 VSS.n4712 0.00241688
R72502 VSS.n11422 VSS.n11421 0.00241688
R72503 VSS.n11201 VSS.n11200 0.00241688
R72504 VSS.n17391 VSS.n17390 0.00241688
R72505 VSS.n3795 VSS.n3794 0.00241688
R72506 VSS.n480 VSS.n479 0.00241688
R72507 VSS.n10516 VSS.n10515 0.00241688
R72508 VSS.n10460 VSS.n10459 0.00241688
R72509 VSS.n8979 VSS.n8978 0.00241688
R72510 VSS.n8991 VSS.n8989 0.00241688
R72511 VSS.n10517 VSS.n10516 0.00241688
R72512 VSS.n8991 VSS.n8990 0.00241688
R72513 VSS.n8979 VSS.n8977 0.00241688
R72514 VSS.n481 VSS.n480 0.00241688
R72515 VSS.n2361 VSS.n2360 0.00241688
R72516 VSS.n11366 VSS.n11365 0.00241688
R72517 VSS.n5727 VSS.n5726 0.00241688
R72518 VSS.n2360 VSS.n2359 0.00241688
R72519 VSS.n5726 VSS.n5725 0.00241688
R72520 VSS.n11367 VSS.n11366 0.00241688
R72521 VSS.n12777 VSS.n12776 0.00241688
R72522 VSS.n12778 VSS.n12777 0.00241688
R72523 VSS.n16174 VSS.n16173 0.00241688
R72524 VSS.n16175 VSS.n16174 0.00241688
R72525 VSS.n21115 VSS.n21114 0.00241688
R72526 VSS.n21114 VSS.n21113 0.00241688
R72527 VSS.n7585 VSS.n7584 0.00241688
R72528 VSS.n7584 VSS.n7583 0.00241688
R72529 VSS.n540 VSS.n539 0.00241688
R72530 VSS.n539 VSS.n538 0.00241688
R72531 VSS.n4073 VSS.n4072 0.00241643
R72532 VSS.n13213 VSS.n13212 0.00241643
R72533 VSS.n18944 VSS.n18943 0.00241643
R72534 VSS.n1439 VSS.n1438 0.00241643
R72535 VSS.n1394 VSS.n1393 0.00241643
R72536 VSS.n1359 VSS.n1358 0.00241643
R72537 VSS.n1154 VSS.n1153 0.00241643
R72538 VSS.n13100 VSS.n13099 0.00241643
R72539 VSS.n21873 VSS.n21872 0.00241643
R72540 VSS.n19158 VSS.n19157 0.00241643
R72541 VSS.n2615 VSS.n2614 0.00241643
R72542 VSS.n15290 VSS.n15287 0.00241489
R72543 VSS.n15297 VSS.n15295 0.00241489
R72544 VSS.n1610 VSS.n1608 0.00241489
R72545 VSS.n1607 VSS.n1605 0.00241489
R72546 VSS.n15511 VSS.n15510 0.00241489
R72547 VSS.n1781 VSS.n1778 0.00241489
R72548 VSS.n3526 VSS.n3525 0.00240141
R72549 VSS.n3585 VSS.n3584 0.00240141
R72550 VSS.n3628 VSS.n3627 0.00240141
R72551 VSS.n3205 VSS.n3204 0.00240141
R72552 VSS.n3528 VSS.n3527 0.00240141
R72553 VSS.n3587 VSS.n3586 0.00240141
R72554 VSS.n3630 VSS.n3629 0.00240141
R72555 VSS.n3663 VSS.n3662 0.00240141
R72556 VSS.n18736 VSS.n18735 0.00240141
R72557 VSS.n18741 VSS.n18740 0.00240141
R72558 VSS.n18746 VSS.n18745 0.00240141
R72559 VSS.n18801 VSS.n18800 0.00240141
R72560 VSS.n18835 VSS.n18834 0.00240141
R72561 VSS.n18676 VSS.n18675 0.00240141
R72562 VSS.n14892 VSS.n14891 0.00240141
R72563 VSS.n14894 VSS.n14893 0.00240141
R72564 VSS.n14895 VSS.n14894 0.00240141
R72565 VSS.n16937 VSS.n16936 0.00240141
R72566 VSS.n16582 VSS.n16581 0.00240141
R72567 VSS.n16541 VSS.n16540 0.00240141
R72568 VSS.n15472 VSS.n15471 0.00240141
R72569 VSS.n15465 VSS.n15464 0.00240141
R72570 VSS.n15340 VSS.n15339 0.00240141
R72571 VSS.n15324 VSS.n15323 0.00240141
R72572 VSS.n8457 VSS.n8456 0.00240141
R72573 VSS.n8539 VSS.n8538 0.00240141
R72574 VSS.n8528 VSS.n8527 0.00240141
R72575 VSS.n8394 VSS.n8393 0.00240141
R72576 VSS.n8383 VSS.n8382 0.00240141
R72577 VSS.n19218 VSS.n19217 0.00240141
R72578 VSS.n19223 VSS.n19222 0.00240141
R72579 VSS.n19228 VSS.n19227 0.00240141
R72580 VSS.n19473 VSS.n19472 0.00240141
R72581 VSS.n19507 VSS.n19506 0.00240141
R72582 VSS.n19527 VSS.n19526 0.00240141
R72583 VSS.n19963 VSS.n19962 0.00240141
R72584 VSS.n19965 VSS.n19964 0.00240141
R72585 VSS.n19966 VSS.n19965 0.00240141
R72586 VSS.n19979 VSS.n19978 0.00240141
R72587 VSS.n786 VSS.n785 0.00240141
R72588 VSS.n797 VSS.n796 0.00240141
R72589 VSS.n1774 VSS.n1773 0.00240141
R72590 VSS.n1767 VSS.n1766 0.00240141
R72591 VSS.n1656 VSS.n1655 0.00240141
R72592 VSS.n1640 VSS.n1639 0.00240141
R72593 VSS.n8608 VSS.n8607 0.00240141
R72594 VSS.n8690 VSS.n8689 0.00240141
R72595 VSS.n8679 VSS.n8678 0.00240141
R72596 VSS.n8202 VSS.n8201 0.00240141
R72597 VSS.n8191 VSS.n8190 0.00240141
R72598 VSS.n20401 VSS.n461 0.00239333
R72599 VSS.n20402 VSS.n20401 0.00239333
R72600 VSS.n20403 VSS.n20402 0.00239333
R72601 VSS.n20404 VSS.n20403 0.00239333
R72602 VSS.n20405 VSS.n20404 0.00239333
R72603 VSS.n20406 VSS.n20405 0.00239333
R72604 VSS.n20407 VSS.n20406 0.00239333
R72605 VSS.n20408 VSS.n20407 0.00239333
R72606 VSS.n20409 VSS.n20408 0.00239333
R72607 VSS.n20410 VSS.n20409 0.00239333
R72608 VSS.n20411 VSS.n20410 0.00239333
R72609 VSS.n20412 VSS.n20411 0.00239333
R72610 VSS.n20413 VSS.n20412 0.00239333
R72611 VSS.n20414 VSS.n20413 0.00239333
R72612 VSS.n20415 VSS.n20414 0.00239333
R72613 VSS.n20416 VSS.n20415 0.00239333
R72614 VSS.n20417 VSS.n20416 0.00239333
R72615 VSS.n20418 VSS.n20417 0.00239333
R72616 VSS.n20419 VSS.n20418 0.00239333
R72617 VSS.n20420 VSS.n20419 0.00239333
R72618 VSS.n20421 VSS.n20420 0.00239333
R72619 VSS.n20422 VSS.n20421 0.00239333
R72620 VSS.n20423 VSS.n20422 0.00239333
R72621 VSS.n20424 VSS.n20423 0.00239333
R72622 VSS.n20425 VSS.n20424 0.00239333
R72623 VSS.n20426 VSS.n20425 0.00239333
R72624 VSS.n20427 VSS.n20426 0.00239333
R72625 VSS.n20428 VSS.n20427 0.00239333
R72626 VSS.n20429 VSS.n20428 0.00239333
R72627 VSS.n20430 VSS.n20429 0.00239333
R72628 VSS.n20431 VSS.n20430 0.00239333
R72629 VSS.n20432 VSS.n20431 0.00239333
R72630 VSS.n20433 VSS.n20432 0.00239333
R72631 VSS.n20434 VSS.n20433 0.00239333
R72632 VSS.n20435 VSS.n20434 0.00239333
R72633 VSS.n20436 VSS.n20435 0.00239333
R72634 VSS.n20437 VSS.n20436 0.00239333
R72635 VSS.n20438 VSS.n20437 0.00239333
R72636 VSS.n20439 VSS.n20438 0.00239333
R72637 VSS.n20440 VSS.n20439 0.00239333
R72638 VSS.n20441 VSS.n20440 0.00239333
R72639 VSS.n20442 VSS.n20441 0.00239333
R72640 VSS.n20443 VSS.n20442 0.00239333
R72641 VSS.n20444 VSS.n20443 0.00239333
R72642 VSS.n20445 VSS.n20444 0.00239333
R72643 VSS.n20446 VSS.n20445 0.00239333
R72644 VSS.n20447 VSS.n20446 0.00239333
R72645 VSS.n20448 VSS.n20447 0.00239333
R72646 VSS.n20449 VSS.n20448 0.00239333
R72647 VSS.n20450 VSS.n20449 0.00239333
R72648 VSS.n20451 VSS.n20450 0.00239333
R72649 VSS.n20452 VSS.n20451 0.00239333
R72650 VSS.n20453 VSS.n20452 0.00239333
R72651 VSS.n20454 VSS.n20453 0.00239333
R72652 VSS.n20455 VSS.n20454 0.00239333
R72653 VSS.n20456 VSS.n20455 0.00239333
R72654 VSS.n20457 VSS.n20456 0.00239333
R72655 VSS.n20458 VSS.n20457 0.00239333
R72656 VSS.n20459 VSS.n20458 0.00239333
R72657 VSS.n20460 VSS.n20459 0.00239333
R72658 VSS.n20461 VSS.n20460 0.00239333
R72659 VSS.n20462 VSS.n20461 0.00239333
R72660 VSS.n20463 VSS.n20462 0.00239333
R72661 VSS.n20464 VSS.n20463 0.00239333
R72662 VSS.n20465 VSS.n20464 0.00239333
R72663 VSS.n20466 VSS.n20465 0.00239333
R72664 VSS.n20467 VSS.n20466 0.00239333
R72665 VSS.n20468 VSS.n20467 0.00239333
R72666 VSS.n20469 VSS.n20468 0.00239333
R72667 VSS.n20470 VSS.n20469 0.00239333
R72668 VSS.n20471 VSS.n20470 0.00239333
R72669 VSS.n20472 VSS.n20471 0.00239333
R72670 VSS.n20473 VSS.n20472 0.00239333
R72671 VSS.n20474 VSS.n20473 0.00239333
R72672 VSS.n20475 VSS.n20474 0.00239333
R72673 VSS.n20476 VSS.n20475 0.00239333
R72674 VSS.n20477 VSS.n20476 0.00239333
R72675 VSS.n20478 VSS.n20477 0.00239333
R72676 VSS.n20479 VSS.n20478 0.00239333
R72677 VSS.n20480 VSS.n20479 0.00239333
R72678 VSS.n20481 VSS.n20480 0.00239333
R72679 VSS.n20482 VSS.n20481 0.00239333
R72680 VSS.n20483 VSS.n20482 0.00239333
R72681 VSS.n20484 VSS.n20483 0.00239333
R72682 VSS.n20488 VSS.n20484 0.00239333
R72683 VSS.n20490 VSS.n20488 0.00239333
R72684 VSS.n20492 VSS.n20490 0.00239333
R72685 VSS.n20494 VSS.n20492 0.00239333
R72686 VSS.n20496 VSS.n20494 0.00239333
R72687 VSS.n20498 VSS.n20496 0.00239333
R72688 VSS.n20502 VSS.n20498 0.00239333
R72689 VSS.n20506 VSS.n20502 0.00239333
R72690 VSS.n20510 VSS.n20506 0.00239333
R72691 VSS.n20512 VSS.n20510 0.00239333
R72692 VSS.n20514 VSS.n20512 0.00239333
R72693 VSS.n20516 VSS.n20514 0.00239333
R72694 VSS.n20518 VSS.n20516 0.00239333
R72695 VSS.n20549 VSS.n20518 0.00239333
R72696 VSS.n20549 VSS.n20548 0.00239333
R72697 VSS.n20526 VSS.n20525 0.00239333
R72698 VSS.n6167 VSS.n6166 0.00239333
R72699 VSS.n6168 VSS.n6167 0.00239333
R72700 VSS.n6169 VSS.n6168 0.00239333
R72701 VSS.n6170 VSS.n6169 0.00239333
R72702 VSS.n6171 VSS.n6170 0.00239333
R72703 VSS.n6172 VSS.n6171 0.00239333
R72704 VSS.n6173 VSS.n6172 0.00239333
R72705 VSS.n6174 VSS.n6173 0.00239333
R72706 VSS.n6175 VSS.n6174 0.00239333
R72707 VSS.n6176 VSS.n6175 0.00239333
R72708 VSS.n6177 VSS.n6176 0.00239333
R72709 VSS.n6178 VSS.n6177 0.00239333
R72710 VSS.n6179 VSS.n6178 0.00239333
R72711 VSS.n6180 VSS.n6179 0.00239333
R72712 VSS.n6204 VSS.n6203 0.00239333
R72713 VSS.n6203 VSS.n6202 0.00239333
R72714 VSS.n6202 VSS.n6201 0.00239333
R72715 VSS.n6201 VSS.n6200 0.00239333
R72716 VSS.n6200 VSS.n6199 0.00239333
R72717 VSS.n6199 VSS.n6198 0.00239333
R72718 VSS.n6198 VSS.n6197 0.00239333
R72719 VSS.n6197 VSS.n6196 0.00239333
R72720 VSS.n6196 VSS.n6195 0.00239333
R72721 VSS.n6195 VSS.n6194 0.00239333
R72722 VSS.n6194 VSS.n6193 0.00239333
R72723 VSS.n6193 VSS.n6192 0.00239333
R72724 VSS.n6192 VSS.n6191 0.00239333
R72725 VSS.n6191 VSS.n6190 0.00239333
R72726 VSS.n6190 VSS.n6189 0.00239333
R72727 VSS.n6189 VSS.n6188 0.00239333
R72728 VSS.n6188 VSS.n6187 0.00239333
R72729 VSS.n6187 VSS.n6186 0.00239333
R72730 VSS.n6186 VSS.n6185 0.00239333
R72731 VSS.n6185 VSS.n6184 0.00239333
R72732 VSS.n6184 VSS.n6183 0.00239333
R72733 VSS.n6183 VSS.n6182 0.00239333
R72734 VSS.n6182 VSS.n6181 0.00239333
R72735 VSS.n6269 VSS.n6268 0.00239333
R72736 VSS.n6268 VSS.n6267 0.00239333
R72737 VSS.n6267 VSS.n6266 0.00239333
R72738 VSS.n6266 VSS.n6265 0.00239333
R72739 VSS.n6265 VSS.n6264 0.00239333
R72740 VSS.n6264 VSS.n6263 0.00239333
R72741 VSS.n6263 VSS.n6262 0.00239333
R72742 VSS.n6262 VSS.n6261 0.00239333
R72743 VSS.n6261 VSS.n6260 0.00239333
R72744 VSS.n6260 VSS.n6259 0.00239333
R72745 VSS.n6259 VSS.n6258 0.00239333
R72746 VSS.n6258 VSS.n6257 0.00239333
R72747 VSS.n6257 VSS.n6256 0.00239333
R72748 VSS.n6256 VSS.n6255 0.00239333
R72749 VSS.n6255 VSS.n6254 0.00239333
R72750 VSS.n6254 VSS.n6253 0.00239333
R72751 VSS.n6253 VSS.n6252 0.00239333
R72752 VSS.n6252 VSS.n6251 0.00239333
R72753 VSS.n6251 VSS.n6250 0.00239333
R72754 VSS.n6250 VSS.n6249 0.00239333
R72755 VSS.n6249 VSS.n6248 0.00239333
R72756 VSS.n6248 VSS.n6247 0.00239333
R72757 VSS.n6247 VSS.n6246 0.00239333
R72758 VSS.n6319 VSS.n6318 0.00239333
R72759 VSS.n6318 VSS.n6317 0.00239333
R72760 VSS.n6317 VSS.n6316 0.00239333
R72761 VSS.n6316 VSS.n6315 0.00239333
R72762 VSS.n6315 VSS.n6314 0.00239333
R72763 VSS.n6314 VSS.n6313 0.00239333
R72764 VSS.n6313 VSS.n6312 0.00239333
R72765 VSS.n6312 VSS.n6311 0.00239333
R72766 VSS.n6311 VSS.n6310 0.00239333
R72767 VSS.n6310 VSS.n6309 0.00239333
R72768 VSS.n6309 VSS.n6308 0.00239333
R72769 VSS.n6308 VSS.n6307 0.00239333
R72770 VSS.n6307 VSS.n6306 0.00239333
R72771 VSS.n6306 VSS.n6305 0.00239333
R72772 VSS.n6305 VSS.n6304 0.00239333
R72773 VSS.n6304 VSS.n6303 0.00239333
R72774 VSS.n6303 VSS.n6302 0.00239333
R72775 VSS.n6302 VSS.n6301 0.00239333
R72776 VSS.n6301 VSS.n6300 0.00239333
R72777 VSS.n6300 VSS.n6299 0.00239333
R72778 VSS.n6299 VSS.n6298 0.00239333
R72779 VSS.n6298 VSS.n6297 0.00239333
R72780 VSS.n6297 VSS.n6296 0.00239333
R72781 VSS.n7011 VSS.n7010 0.00239333
R72782 VSS.n7012 VSS.n7011 0.00239333
R72783 VSS.n7013 VSS.n7012 0.00239333
R72784 VSS.n7014 VSS.n7013 0.00239333
R72785 VSS.n7015 VSS.n7014 0.00239333
R72786 VSS.n7016 VSS.n7015 0.00239333
R72787 VSS.n7017 VSS.n7016 0.00239333
R72788 VSS.n7019 VSS.n7017 0.00239333
R72789 VSS.n7021 VSS.n7019 0.00239333
R72790 VSS.n7857 VSS.n7021 0.00239333
R72791 VSS.n7856 VSS.n7855 0.00239333
R72792 VSS.n7042 VSS.n7041 0.00239333
R72793 VSS.n6207 VSS.n6206 0.00239333
R72794 VSS.n6208 VSS.n6207 0.00239333
R72795 VSS.n6209 VSS.n6208 0.00239333
R72796 VSS.n6210 VSS.n6209 0.00239333
R72797 VSS.n6211 VSS.n6210 0.00239333
R72798 VSS.n6212 VSS.n6211 0.00239333
R72799 VSS.n6213 VSS.n6212 0.00239333
R72800 VSS.n6214 VSS.n6213 0.00239333
R72801 VSS.n6215 VSS.n6214 0.00239333
R72802 VSS.n6216 VSS.n6215 0.00239333
R72803 VSS.n6217 VSS.n6216 0.00239333
R72804 VSS.n6218 VSS.n6217 0.00239333
R72805 VSS.n6219 VSS.n6218 0.00239333
R72806 VSS.n6220 VSS.n6219 0.00239333
R72807 VSS.n6244 VSS.n6243 0.00239333
R72808 VSS.n6243 VSS.n6242 0.00239333
R72809 VSS.n6242 VSS.n6241 0.00239333
R72810 VSS.n6241 VSS.n6240 0.00239333
R72811 VSS.n6240 VSS.n6239 0.00239333
R72812 VSS.n6239 VSS.n6238 0.00239333
R72813 VSS.n6238 VSS.n6237 0.00239333
R72814 VSS.n6237 VSS.n6236 0.00239333
R72815 VSS.n6236 VSS.n6235 0.00239333
R72816 VSS.n6235 VSS.n6234 0.00239333
R72817 VSS.n6234 VSS.n6233 0.00239333
R72818 VSS.n6233 VSS.n6232 0.00239333
R72819 VSS.n6232 VSS.n6231 0.00239333
R72820 VSS.n6231 VSS.n6230 0.00239333
R72821 VSS.n6230 VSS.n6229 0.00239333
R72822 VSS.n6229 VSS.n6228 0.00239333
R72823 VSS.n6228 VSS.n6227 0.00239333
R72824 VSS.n6227 VSS.n6226 0.00239333
R72825 VSS.n6226 VSS.n6225 0.00239333
R72826 VSS.n6225 VSS.n6224 0.00239333
R72827 VSS.n6224 VSS.n6223 0.00239333
R72828 VSS.n6223 VSS.n6222 0.00239333
R72829 VSS.n6222 VSS.n6221 0.00239333
R72830 VSS.n6294 VSS.n6293 0.00239333
R72831 VSS.n6293 VSS.n6292 0.00239333
R72832 VSS.n6292 VSS.n6291 0.00239333
R72833 VSS.n6291 VSS.n6290 0.00239333
R72834 VSS.n6290 VSS.n6289 0.00239333
R72835 VSS.n6289 VSS.n6288 0.00239333
R72836 VSS.n6288 VSS.n6287 0.00239333
R72837 VSS.n6287 VSS.n6286 0.00239333
R72838 VSS.n6286 VSS.n6285 0.00239333
R72839 VSS.n6285 VSS.n6284 0.00239333
R72840 VSS.n6284 VSS.n6283 0.00239333
R72841 VSS.n6283 VSS.n6282 0.00239333
R72842 VSS.n6282 VSS.n6281 0.00239333
R72843 VSS.n6281 VSS.n6280 0.00239333
R72844 VSS.n6280 VSS.n6279 0.00239333
R72845 VSS.n6279 VSS.n6278 0.00239333
R72846 VSS.n6278 VSS.n6277 0.00239333
R72847 VSS.n6277 VSS.n6276 0.00239333
R72848 VSS.n6276 VSS.n6275 0.00239333
R72849 VSS.n6275 VSS.n6274 0.00239333
R72850 VSS.n6274 VSS.n6273 0.00239333
R72851 VSS.n6273 VSS.n6272 0.00239333
R72852 VSS.n6272 VSS.n6271 0.00239333
R72853 VSS.n6344 VSS.n6343 0.00239333
R72854 VSS.n6343 VSS.n6342 0.00239333
R72855 VSS.n6342 VSS.n6341 0.00239333
R72856 VSS.n6341 VSS.n6340 0.00239333
R72857 VSS.n6340 VSS.n6339 0.00239333
R72858 VSS.n6339 VSS.n6338 0.00239333
R72859 VSS.n6338 VSS.n6337 0.00239333
R72860 VSS.n6337 VSS.n6336 0.00239333
R72861 VSS.n6336 VSS.n6335 0.00239333
R72862 VSS.n6335 VSS.n6334 0.00239333
R72863 VSS.n6334 VSS.n6333 0.00239333
R72864 VSS.n6333 VSS.n6332 0.00239333
R72865 VSS.n6332 VSS.n6331 0.00239333
R72866 VSS.n6331 VSS.n6330 0.00239333
R72867 VSS.n6330 VSS.n6329 0.00239333
R72868 VSS.n6329 VSS.n6328 0.00239333
R72869 VSS.n6328 VSS.n6327 0.00239333
R72870 VSS.n6327 VSS.n6326 0.00239333
R72871 VSS.n6326 VSS.n6325 0.00239333
R72872 VSS.n6325 VSS.n6324 0.00239333
R72873 VSS.n6324 VSS.n6323 0.00239333
R72874 VSS.n6323 VSS.n6322 0.00239333
R72875 VSS.n6322 VSS.n6321 0.00239333
R72876 VSS.n7909 VSS.n7908 0.00239333
R72877 VSS.n7910 VSS.n7909 0.00239333
R72878 VSS.n7911 VSS.n7910 0.00239333
R72879 VSS.n7912 VSS.n7911 0.00239333
R72880 VSS.n7913 VSS.n7912 0.00239333
R72881 VSS.n7914 VSS.n7913 0.00239333
R72882 VSS.n7915 VSS.n7914 0.00239333
R72883 VSS.n7916 VSS.n7915 0.00239333
R72884 VSS.n7917 VSS.n7916 0.00239333
R72885 VSS.n7919 VSS.n7918 0.00239333
R72886 VSS.n7940 VSS.n7919 0.00239333
R72887 VSS.n7940 VSS.n7939 0.00239333
R72888 VSS.n7939 VSS.n7930 0.00239333
R72889 VSS.n11178 VSS.n6165 0.00239333
R72890 VSS.n11178 VSS.n11177 0.00239333
R72891 VSS.n11177 VSS.n11176 0.00239333
R72892 VSS.n11176 VSS.n11175 0.00239333
R72893 VSS.n11175 VSS.n11174 0.00239333
R72894 VSS.n11174 VSS.n11173 0.00239333
R72895 VSS.n11173 VSS.n11172 0.00239333
R72896 VSS.n11172 VSS.n11171 0.00239333
R72897 VSS.n11171 VSS.n11170 0.00239333
R72898 VSS.n11170 VSS.n11169 0.00239333
R72899 VSS.n11169 VSS.n11168 0.00239333
R72900 VSS.n11168 VSS.n11167 0.00239333
R72901 VSS.n11167 VSS.n11166 0.00239333
R72902 VSS.n11166 VSS.n11165 0.00239333
R72903 VSS.n11163 VSS.n11162 0.00239333
R72904 VSS.n11162 VSS.n11161 0.00239333
R72905 VSS.n11161 VSS.n11160 0.00239333
R72906 VSS.n11160 VSS.n11159 0.00239333
R72907 VSS.n11159 VSS.n11158 0.00239333
R72908 VSS.n11158 VSS.n11157 0.00239333
R72909 VSS.n11157 VSS.n11156 0.00239333
R72910 VSS.n11156 VSS.n11155 0.00239333
R72911 VSS.n11155 VSS.n11154 0.00239333
R72912 VSS.n11154 VSS.n11153 0.00239333
R72913 VSS.n11153 VSS.n11152 0.00239333
R72914 VSS.n11152 VSS.n11151 0.00239333
R72915 VSS.n11151 VSS.n11150 0.00239333
R72916 VSS.n11150 VSS.n11149 0.00239333
R72917 VSS.n11149 VSS.n11148 0.00239333
R72918 VSS.n11148 VSS.n11147 0.00239333
R72919 VSS.n11147 VSS.n11146 0.00239333
R72920 VSS.n11146 VSS.n11145 0.00239333
R72921 VSS.n11145 VSS.n11144 0.00239333
R72922 VSS.n11144 VSS.n11143 0.00239333
R72923 VSS.n11143 VSS.n11142 0.00239333
R72924 VSS.n11142 VSS.n11141 0.00239333
R72925 VSS.n11141 VSS.n11140 0.00239333
R72926 VSS.n11138 VSS.n11137 0.00239333
R72927 VSS.n11137 VSS.n11136 0.00239333
R72928 VSS.n11136 VSS.n11135 0.00239333
R72929 VSS.n11135 VSS.n11134 0.00239333
R72930 VSS.n11134 VSS.n11133 0.00239333
R72931 VSS.n11133 VSS.n11132 0.00239333
R72932 VSS.n11132 VSS.n11131 0.00239333
R72933 VSS.n11131 VSS.n11130 0.00239333
R72934 VSS.n11130 VSS.n11129 0.00239333
R72935 VSS.n11129 VSS.n11128 0.00239333
R72936 VSS.n11128 VSS.n11127 0.00239333
R72937 VSS.n11127 VSS.n11126 0.00239333
R72938 VSS.n11126 VSS.n11125 0.00239333
R72939 VSS.n11125 VSS.n11124 0.00239333
R72940 VSS.n11124 VSS.n11123 0.00239333
R72941 VSS.n11123 VSS.n11122 0.00239333
R72942 VSS.n11122 VSS.n11121 0.00239333
R72943 VSS.n11121 VSS.n11120 0.00239333
R72944 VSS.n11120 VSS.n11119 0.00239333
R72945 VSS.n11119 VSS.n11118 0.00239333
R72946 VSS.n11118 VSS.n11117 0.00239333
R72947 VSS.n11117 VSS.n11116 0.00239333
R72948 VSS.n11116 VSS.n11115 0.00239333
R72949 VSS.n11113 VSS.n11112 0.00239333
R72950 VSS.n11112 VSS.n11111 0.00239333
R72951 VSS.n11111 VSS.n11110 0.00239333
R72952 VSS.n11110 VSS.n11109 0.00239333
R72953 VSS.n11109 VSS.n11108 0.00239333
R72954 VSS.n11108 VSS.n11107 0.00239333
R72955 VSS.n11107 VSS.n11106 0.00239333
R72956 VSS.n11106 VSS.n11105 0.00239333
R72957 VSS.n11105 VSS.n11104 0.00239333
R72958 VSS.n11104 VSS.n11103 0.00239333
R72959 VSS.n11103 VSS.n11102 0.00239333
R72960 VSS.n11102 VSS.n11101 0.00239333
R72961 VSS.n11101 VSS.n11100 0.00239333
R72962 VSS.n11100 VSS.n11099 0.00239333
R72963 VSS.n11099 VSS.n11098 0.00239333
R72964 VSS.n11098 VSS.n11097 0.00239333
R72965 VSS.n11097 VSS.n11096 0.00239333
R72966 VSS.n11096 VSS.n11095 0.00239333
R72967 VSS.n11095 VSS.n11094 0.00239333
R72968 VSS.n11094 VSS.n11093 0.00239333
R72969 VSS.n11093 VSS.n11092 0.00239333
R72970 VSS.n11092 VSS.n11091 0.00239333
R72971 VSS.n11091 VSS.n11090 0.00239333
R72972 VSS.n11088 VSS.n11087 0.00239333
R72973 VSS.n11087 VSS.n11086 0.00239333
R72974 VSS.n11086 VSS.n11085 0.00239333
R72975 VSS.n11085 VSS.n11084 0.00239333
R72976 VSS.n11084 VSS.n11083 0.00239333
R72977 VSS.n11083 VSS.n11082 0.00239333
R72978 VSS.n11082 VSS.n11081 0.00239333
R72979 VSS.n11081 VSS.n11080 0.00239333
R72980 VSS.n11079 VSS.n6347 0.00239333
R72981 VSS.n6379 VSS.n6347 0.00239333
R72982 VSS.n6379 VSS.n6378 0.00239333
R72983 VSS.n6378 VSS.n6368 0.00239333
R72984 VSS.n6368 VSS.n6359 0.00239333
R72985 VSS.n10201 VSS.n10200 0.00238571
R72986 VSS.n18702 VSS.n18701 0.00237282
R72987 VSS.n18787 VSS.n18786 0.00237282
R72988 VSS.n15667 VSS.n15666 0.00237282
R72989 VSS.n15665 VSS.n15664 0.00237282
R72990 VSS.n15661 VSS.n15660 0.00237282
R72991 VSS.n15659 VSS.n15658 0.00237282
R72992 VSS.n15584 VSS.n15583 0.00237282
R72993 VSS.n15573 VSS.n15572 0.00237282
R72994 VSS.n15569 VSS.n15568 0.00237282
R72995 VSS.n15567 VSS.n15566 0.00237282
R72996 VSS.n15564 VSS.n15563 0.00237282
R72997 VSS.n15562 VSS.n15557 0.00237282
R72998 VSS.n15554 VSS.n15553 0.00237282
R72999 VSS.n15552 VSS.n15551 0.00237282
R73000 VSS.n15461 VSS.n15460 0.00237282
R73001 VSS.n15338 VSS.n15337 0.00237282
R73002 VSS.n15462 VSS.n15461 0.00237282
R73003 VSS.n15568 VSS.n15567 0.00237282
R73004 VSS.n15583 VSS.n15574 0.00237282
R73005 VSS.n15574 VSS.n15573 0.00237282
R73006 VSS.n15660 VSS.n15659 0.00237282
R73007 VSS.n15666 VSS.n15665 0.00237282
R73008 VSS.n16939 VSS.n16938 0.00237282
R73009 VSS.n15570 VSS.n15569 0.00237282
R73010 VSS.n15662 VSS.n15661 0.00237282
R73011 VSS.n15668 VSS.n15667 0.00237282
R73012 VSS.n15339 VSS.n15338 0.00237282
R73013 VSS.n15555 VSS.n15554 0.00237282
R73014 VSS.n15553 VSS.n15552 0.00237282
R73015 VSS.n15565 VSS.n15564 0.00237282
R73016 VSS.n15563 VSS.n15562 0.00237282
R73017 VSS.n15375 VSS.n15374 0.00237282
R73018 VSS.n19184 VSS.n19183 0.00237282
R73019 VSS.n1925 VSS.n1924 0.00237282
R73020 VSS.n1923 VSS.n1922 0.00237282
R73021 VSS.n1919 VSS.n1918 0.00237282
R73022 VSS.n1917 VSS.n1916 0.00237282
R73023 VSS.n1863 VSS.n1862 0.00237282
R73024 VSS.n1861 VSS.n1860 0.00237282
R73025 VSS.n1857 VSS.n1856 0.00237282
R73026 VSS.n1856 VSS.n1855 0.00237282
R73027 VSS.n1852 VSS.n1851 0.00237282
R73028 VSS.n1850 VSS.n1845 0.00237282
R73029 VSS.n1842 VSS.n1841 0.00237282
R73030 VSS.n1840 VSS.n1839 0.00237282
R73031 VSS.n1763 VSS.n1762 0.00237282
R73032 VSS.n1654 VSS.n1653 0.00237282
R73033 VSS.n1655 VSS.n1654 0.00237282
R73034 VSS.n1691 VSS.n1690 0.00237282
R73035 VSS.n1764 VSS.n1763 0.00237282
R73036 VSS.n1843 VSS.n1842 0.00237282
R73037 VSS.n1841 VSS.n1840 0.00237282
R73038 VSS.n1853 VSS.n1852 0.00237282
R73039 VSS.n19977 VSS.n19976 0.00237282
R73040 VSS.n1924 VSS.n1923 0.00237282
R73041 VSS.n1918 VSS.n1917 0.00237282
R73042 VSS.n1862 VSS.n1861 0.00237282
R73043 VSS.n1858 VSS.n1857 0.00237282
R73044 VSS.n1920 VSS.n1919 0.00237282
R73045 VSS.n1864 VSS.n1863 0.00237282
R73046 VSS.n1926 VSS.n1925 0.00237282
R73047 VSS.n1855 VSS.n1854 0.00237282
R73048 VSS.n1851 VSS.n1850 0.00237282
R73049 VSS.n19459 VSS.n19458 0.00237282
R73050 VSS.n19183 VSS.n19182 0.00237282
R73051 VSS.n18701 VSS.n18700 0.00237282
R73052 VSS.n20526 DVSS 0.00236667
R73053 VSS.n8268 VSS.n8267 0.00236
R73054 VSS.n6780 VSS.n6779 0.00236
R73055 VSS.n6721 VSS.n6719 0.00236
R73056 VSS.n7888 VSS.n7887 0.00236
R73057 VSS.n8605 VSS.n8604 0.00236
R73058 VSS.n8096 VSS.n8095 0.00236
R73059 VSS.n8037 VSS.n8035 0.00236
R73060 VSS.n7981 VSS.n7980 0.00236
R73061 VSS.n10863 VSS.n10862 0.00236
R73062 VSS.n10914 VSS.n10913 0.00236
R73063 VSS.n10981 VSS.n10980 0.00236
R73064 VSS.n11047 VSS.n11046 0.00236
R73065 VSS.n17712 DVSS 0.00235714
R73066 VSS.n14197 VSS.n14196 0.0023496
R73067 VSS.n14159 VSS.n14158 0.0023496
R73068 VSS.n3212 VSS.n3211 0.00233099
R73069 VSS.n3214 VSS.n3213 0.00233099
R73070 VSS.n3518 VSS.n3515 0.00233099
R73071 VSS.n3577 VSS.n3574 0.00233099
R73072 VSS.n3620 VSS.n3617 0.00233099
R73073 VSS.n3670 VSS.n3669 0.00233099
R73074 VSS.n3666 VSS.n3665 0.00233099
R73075 VSS.n12301 VSS.n12300 0.00232835
R73076 VSS.n21668 VSS.n21667 0.00232835
R73077 VSS.n21667 VSS.n21666 0.00232835
R73078 VSS.n12300 VSS.n12299 0.00232835
R73079 VSS.n4129 VSS.n4128 0.00232835
R73080 VSS.n4128 VSS.n4127 0.00232835
R73081 VSS.n10249 VSS.n10248 0.00232835
R73082 VSS.n10248 VSS.n10247 0.00232835
R73083 VSS.n9385 VSS.n9383 0.00230496
R73084 VSS.n9331 VSS.n9329 0.00230496
R73085 VSS.n9722 VSS.n9720 0.00230496
R73086 VSS.n13851 VSS 0.0023
R73087 VSS.n13850 VSS 0.0023
R73088 VSS.n18367 VSS.n18366 0.0023
R73089 DVSS VSS.n16991 0.0023
R73090 VSS.n16571 VSS.n16569 0.0023
R73091 VSS.n3083 DVSS 0.0023
R73092 VSS.n3082 DVSS 0.0023
R73093 VSS.n5311 DVSS 0.0023
R73094 VSS.n5310 DVSS 0.0023
R73095 DVSS VSS.n7054 0.0023
R73096 VSS.n7053 DVSS 0.0023
R73097 DVSS VSS.n4346 0.0023
R73098 VSS.n4345 DVSS 0.0023
R73099 VSS.n17737 DVSS 0.0023
R73100 DVSS VSS.n17738 0.0023
R73101 VSS.n8995 VSS.n8993 0.0023
R73102 VSS.n9008 VSS.n9006 0.0023
R73103 VSS.n9465 VSS.n9463 0.0023
R73104 VSS.n9470 VSS.n9468 0.0023
R73105 VSS.n10638 VSS.n10636 0.0023
R73106 VSS.n10643 VSS.n10641 0.0023
R73107 VSS.n22264 VSS 0.0023
R73108 VSS VSS.n22265 0.0023
R73109 VSS.n4148 VSS.n4147 0.00229713
R73110 VSS.n7918 DVSS 0.00227333
R73111 VSS.n11531 VSS.n11530 0.00227165
R73112 VSS.n5847 VSS.n5846 0.00227165
R73113 VSS.n5747 VSS.n5746 0.00227165
R73114 VSS.n5622 VSS.n5621 0.00227165
R73115 VSS.n5592 VSS.n5591 0.00227165
R73116 VSS.n5560 VSS.n5559 0.00227165
R73117 VSS.n9588 VSS.n9587 0.00227165
R73118 VSS.n9151 VSS.n9150 0.00227165
R73119 VSS.n12973 VSS.n12972 0.00227165
R73120 VSS.n12755 VSS.n12754 0.00227165
R73121 VSS.n12549 VSS.n12548 0.00227165
R73122 VSS.n12511 VSS.n12510 0.00227165
R73123 VSS.n12508 VSS.n12507 0.00227165
R73124 VSS.n12262 VSS.n12261 0.00227165
R73125 VSS.n11934 VSS.n11933 0.00227165
R73126 VSS.n11933 VSS.n11932 0.00227165
R73127 VSS.n11915 VSS.n11914 0.00227165
R73128 VSS.n11913 VSS.n11912 0.00227165
R73129 VSS.n11844 VSS.n11843 0.00227165
R73130 VSS.n11834 VSS.n11833 0.00227165
R73131 VSS.n15005 VSS.n15004 0.00227165
R73132 VSS.n16208 VSS.n16207 0.00227165
R73133 VSS.n16195 VSS.n16194 0.00227165
R73134 VSS.n16138 VSS.n16137 0.00227165
R73135 VSS.n16108 VSS.n16107 0.00227165
R73136 VSS.n16070 VSS.n16069 0.00227165
R73137 VSS.n9705 VSS.n9704 0.00227165
R73138 VSS.n9314 VSS.n9313 0.00227165
R73139 VSS.n20611 VSS.n20610 0.00227165
R73140 VSS.n21150 VSS.n21149 0.00227165
R73141 VSS.n21137 VSS.n21136 0.00227165
R73142 VSS.n21072 VSS.n21071 0.00227165
R73143 VSS.n21042 VSS.n21041 0.00227165
R73144 VSS.n21009 VSS.n21008 0.00227165
R73145 VSS.n7000 VSS.n6999 0.00227165
R73146 VSS.n6640 VSS.n6639 0.00227165
R73147 VSS.n20138 VSS.n20137 0.00227165
R73148 VSS.n1279 VSS.n1278 0.00227165
R73149 VSS.n1187 VSS.n1186 0.00227165
R73150 VSS.n1118 VSS.n1117 0.00227165
R73151 VSS.n1088 VSS.n1087 0.00227165
R73152 VSS.n1055 VSS.n1054 0.00227165
R73153 VSS.n6898 VSS.n6897 0.00227165
R73154 VSS.n6490 VSS.n6489 0.00227165
R73155 VSS.n21390 VSS.n21389 0.00227165
R73156 VSS.n7607 VSS.n7606 0.00227165
R73157 VSS.n7695 VSS.n7694 0.00227165
R73158 VSS.n7844 VSS.n7843 0.00227165
R73159 VSS.n11704 VSS.n11703 0.00227165
R73160 VSS.n6147 VSS.n6146 0.00227165
R73161 VSS.n6066 VSS.n6065 0.00227165
R73162 VSS.n5985 VSS.n5984 0.00227165
R73163 VSS.n661 VSS.n660 0.00227165
R73164 VSS.n10619 VSS.n10618 0.00227165
R73165 VSS.n10494 VSS.n10493 0.00227165
R73166 VSS.n10457 VSS.n10456 0.00227165
R73167 VSS.n10454 VSS.n10453 0.00227165
R73168 VSS.n10210 VSS.n10209 0.00227165
R73169 VSS.n9935 VSS.n9934 0.00227165
R73170 VSS.n9934 VSS.n9933 0.00227165
R73171 VSS.n9916 VSS.n9915 0.00227165
R73172 VSS.n9914 VSS.n9913 0.00227165
R73173 VSS.n9003 VSS.n9002 0.00227165
R73174 VSS.n8907 VSS.n8906 0.00227165
R73175 VSS.n18422 VSS.n18421 0.00226725
R73176 VSS.n18160 VSS.n18159 0.00226725
R73177 VSS.n17120 VSS.n17119 0.00226725
R73178 VSS.n15381 VSS.n15380 0.00226725
R73179 VSS.n15326 VSS.n15325 0.00226725
R73180 VSS.n8520 VSS.n8519 0.00226725
R73181 VSS.n8338 VSS.n8337 0.00226725
R73182 VSS.n17121 VSS.n17120 0.00226725
R73183 VSS.n18161 VSS.n18160 0.00226725
R73184 VSS.n15327 VSS.n15326 0.00226725
R73185 VSS.n15382 VSS.n15381 0.00226725
R73186 VSS.n8337 VSS.n8336 0.00226725
R73187 VSS.n8519 VSS.n8518 0.00226725
R73188 VSS.n15403 VSS.n15402 0.00226725
R73189 VSS.n19607 VSS.n19606 0.00226725
R73190 VSS.n19696 VSS.n19695 0.00226725
R73191 VSS.n19875 VSS.n19874 0.00226725
R73192 VSS.n1697 VSS.n1696 0.00226725
R73193 VSS.n1643 VSS.n1642 0.00226725
R73194 VSS.n8671 VSS.n8670 0.00226725
R73195 VSS.n8134 VSS.n8133 0.00226725
R73196 VSS.n8133 VSS.n8132 0.00226725
R73197 VSS.n8670 VSS.n8669 0.00226725
R73198 VSS.n1719 VSS.n1718 0.00226725
R73199 VSS.n19874 VSS.n19873 0.00226725
R73200 VSS.n19695 VSS.n19694 0.00226725
R73201 VSS.n1698 VSS.n1697 0.00226725
R73202 VSS.n1642 VSS.n1641 0.00226725
R73203 VSS.n3456 VSS.n3455 0.00226056
R73204 VSS.n9381 VSS.n9380 0.00224
R73205 VSS.n9327 VSS.n9326 0.00224
R73206 VSS.n9718 VSS.n9717 0.00224
R73207 VSS.n10694 VSS.n10692 0.00224
R73208 VSS.n10757 VSS.n10754 0.00224
R73209 VSS.n4017 VSS.n4016 0.00223982
R73210 VSS.n9535 VSS.n9534 0.00223982
R73211 VSS.n4016 VSS.n4015 0.00223982
R73212 VSS.n13042 VSS.n13041 0.00223982
R73213 VSS.n12547 VSS.n12546 0.00223982
R73214 VSS.n12228 VSS.n12227 0.00223982
R73215 VSS.n11803 VSS.n11802 0.00223982
R73216 VSS.n13041 VSS.n13040 0.00223982
R73217 VSS.n18888 VSS.n18887 0.00223982
R73218 VSS.n9652 VSS.n9651 0.00223982
R73219 VSS.n18887 VSS.n18886 0.00223982
R73220 VSS.n21815 VSS.n21814 0.00223982
R73221 VSS.n6941 VSS.n6940 0.00223982
R73222 VSS.n21814 VSS.n21813 0.00223982
R73223 VSS.n19100 VSS.n19099 0.00223982
R73224 VSS.n6839 VSS.n6838 0.00223982
R73225 VSS.n19099 VSS.n19098 0.00223982
R73226 VSS.n21586 VSS.n21585 0.00223982
R73227 VSS.n21663 VSS.n21662 0.00223982
R73228 VSS.n21585 VSS.n21584 0.00223982
R73229 VSS.n21662 VSS.n21661 0.00223982
R73230 VSS.n11887 VSS.n11886 0.00223982
R73231 VSS.n11804 VSS.n11803 0.00223982
R73232 VSS.n12229 VSS.n12228 0.00223982
R73233 VSS.n12548 VSS.n12547 0.00223982
R73234 VSS.n3819 VSS.n3818 0.00223982
R73235 VSS.n4124 VSS.n4123 0.00223982
R73236 VSS.n3818 VSS.n3817 0.00223982
R73237 VSS.n4123 VSS.n4122 0.00223982
R73238 VSS.n3252 VSS.n3251 0.00223982
R73239 VSS.n3253 VSS.n3252 0.00223982
R73240 VSS.n10492 VSS.n10491 0.00223982
R73241 VSS.n10176 VSS.n10175 0.00223982
R73242 VSS.n8951 VSS.n8948 0.00223982
R73243 VSS.n8969 VSS.n8968 0.00223982
R73244 VSS.n10177 VSS.n10176 0.00223982
R73245 VSS.n8951 VSS.n8950 0.00223982
R73246 VSS.n10493 VSS.n10492 0.00223982
R73247 VSS.n8969 VSS.n8967 0.00223982
R73248 VSS.n9534 VSS.n9533 0.00223982
R73249 VSS.n9651 VSS.n9650 0.00223982
R73250 VSS.n6940 VSS.n6939 0.00223982
R73251 VSS.n6838 VSS.n6837 0.00223982
R73252 VSS.n14254 VSS.n13564 0.00223571
R73253 VSS.n14254 VSS.n14241 0.00223571
R73254 VSS.n13676 VSS.n13673 0.00223571
R73255 VSS.n13658 VSS.n13623 0.00223571
R73256 VSS.n2939 VSS.n2938 0.00223571
R73257 VSS.n3004 VSS.n3003 0.00223571
R73258 VSS.n3052 VSS.n3051 0.00223571
R73259 VSS.n2553 VSS.n2550 0.00223571
R73260 VSS.n2567 VSS.n2566 0.00223571
R73261 VSS.n5201 VSS.n5200 0.00223571
R73262 VSS.n5252 VSS.n5251 0.00223571
R73263 VSS.n5287 VSS.n5286 0.00223571
R73264 VSS.n4964 VSS.n4952 0.00223571
R73265 VSS.n5192 VSS.n5191 0.00223571
R73266 VSS.n5203 VSS.n5202 0.00223571
R73267 VSS.n5243 VSS.n5242 0.00223571
R73268 VSS.n5254 VSS.n5253 0.00223571
R73269 VSS.n5278 VSS.n5277 0.00223571
R73270 VSS.n5289 VSS.n5288 0.00223571
R73271 VSS.n4963 VSS.n4962 0.00223571
R73272 VSS.n7172 VSS.n7171 0.00223571
R73273 VSS.n7113 VSS.n7112 0.00223571
R73274 VSS.n7073 VSS.n7072 0.00223571
R73275 VSS.n7538 VSS.n7535 0.00223571
R73276 VSS.n7173 VSS.n7169 0.00223571
R73277 VSS.n7114 VSS.n7110 0.00223571
R73278 VSS.n7083 VSS.n7082 0.00223571
R73279 VSS.n7074 VSS.n7071 0.00223571
R73280 VSS.n7051 VSS.n7046 0.00223571
R73281 VSS.n7539 VSS.n7533 0.00223571
R73282 VSS.n4453 VSS.n4452 0.00223571
R73283 VSS.n4402 VSS.n4401 0.00223571
R73284 VSS.n4367 VSS.n4366 0.00223571
R73285 VSS.n4317 VSS.n4316 0.00223571
R73286 VSS.n4463 VSS.n4462 0.00223571
R73287 VSS.n4454 VSS.n4451 0.00223571
R73288 VSS.n4412 VSS.n4411 0.00223571
R73289 VSS.n4403 VSS.n4400 0.00223571
R73290 VSS.n4377 VSS.n4376 0.00223571
R73291 VSS.n4368 VSS.n4365 0.00223571
R73292 VSS.n4333 VSS.n4332 0.00223571
R73293 VSS.n17580 VSS.n17579 0.00223571
R73294 VSS.n17725 VSS.n17724 0.00223571
R73295 VSS.n17869 VSS.n17868 0.00223571
R73296 VSS.n17808 VSS.n17807 0.00223571
R73297 VSS.n17763 VSS.n17762 0.00223571
R73298 VSS.n17707 VSS.n17706 0.00223571
R73299 VSS.n21987 VSS.n3 0.00223571
R73300 VSS.n21988 VSS.n21987 0.00223571
R73301 VSS.n14124 VSS.n14123 0.00223571
R73302 VSS.n22255 VSS.n22254 0.00223571
R73303 VSS.n14126 VSS.n14125 0.00223571
R73304 VSS.n9875 VSS.n9870 0.00223077
R73305 VSS.n9884 VSS.n9883 0.00223077
R73306 VSS.n10377 VSS.n10372 0.00223077
R73307 VSS.n10370 VSS.n10369 0.00223077
R73308 VSS.n10092 VSS.n10087 0.00223077
R73309 VSS.n10085 VSS.n10084 0.00223077
R73310 VSS.n10000 VSS.n9995 0.00223077
R73311 VSS.n9993 VSS.n9992 0.00223077
R73312 VSS.n11776 VSS.n11771 0.00223077
R73313 VSS.n11785 VSS.n11784 0.00223077
R73314 VSS.n12431 VSS.n12426 0.00223077
R73315 VSS.n12424 VSS.n12423 0.00223077
R73316 VSS.n12143 VSS.n12138 0.00223077
R73317 VSS.n12136 VSS.n12135 0.00223077
R73318 VSS.n12051 VSS.n12046 0.00223077
R73319 VSS.n12044 VSS.n12043 0.00223077
R73320 VSS.n20396 VSS.n20394 0.00221
R73321 VSS.n20365 VSS.n20364 0.00221
R73322 VSS.n20335 VSS.n20333 0.00221
R73323 VSS.n20289 VSS.n20287 0.00221
R73324 VSS.n8818 VSS.n8817 0.00221
R73325 VSS.n9431 VSS.n9430 0.00221
R73326 VSS.n9806 VSS.n9805 0.00221
R73327 VSS.n10524 VSS.n10523 0.0022086
R73328 VSS.n8912 VSS.n8910 0.00220857
R73329 VSS.n443 VSS.n442 0.00220306
R73330 VSS.n426 VSS.n425 0.00220306
R73331 VSS.n409 VSS.n408 0.00220306
R73332 VSS.n14282 VSS.n14281 0.00220306
R73333 VSS.n391 VSS.n390 0.00220306
R73334 VSS.n3775 VSS.n3198 0.00219014
R73335 VSS.n3777 VSS.n3776 0.00219014
R73336 VSS.n3294 VSS.n3291 0.00219014
R73337 VSS.n3298 VSS.n3297 0.00219014
R73338 VSS.n3332 VSS.n3329 0.00219014
R73339 VSS.n3336 VSS.n3335 0.00219014
R73340 VSS.n3386 VSS.n3383 0.00219014
R73341 VSS.n3390 VSS.n3389 0.00219014
R73342 VSS.n3521 VSS.n3520 0.00219014
R73343 VSS.n3580 VSS.n3579 0.00219014
R73344 VSS.n3623 VSS.n3622 0.00219014
R73345 VSS.n18407 VSS.n18406 0.00219014
R73346 VSS.n17065 VSS.n17034 0.00219014
R73347 VSS.n17029 VSS.n17028 0.00219014
R73348 VSS.n14872 VSS.n14871 0.00219014
R73349 VSS.n14886 VSS.n14885 0.00219014
R73350 VSS.n16893 VSS.n16892 0.00219014
R73351 VSS.n16641 VSS.n16640 0.00219014
R73352 VSS.n16542 VSS.n16541 0.00219014
R73353 VSS.n15530 VSS.n15529 0.00219014
R73354 VSS.n15404 VSS.n15403 0.00219014
R73355 VSS.n15385 VSS.n15384 0.00219014
R73356 VSS.n15356 VSS.n15355 0.00219014
R73357 VSS.n15332 VSS.n15331 0.00219014
R73358 VSS.n15328 VSS.n15327 0.00219014
R73359 VSS.n8476 VSS.n8475 0.00219014
R73360 VSS.n8516 VSS.n8515 0.00219014
R73361 VSS.n8558 VSS.n8557 0.00219014
R73362 VSS.n8324 VSS.n8323 0.00219014
R73363 VSS.n8413 VSS.n8412 0.00219014
R73364 VSS.n8364 VSS.n8363 0.00219014
R73365 VSS.n19615 VSS.n19614 0.00219014
R73366 VSS.n19900 VSS.n19899 0.00219014
R73367 VSS.n19906 VSS.n19905 0.00219014
R73368 VSS.n19943 VSS.n19942 0.00219014
R73369 VSS.n19957 VSS.n19956 0.00219014
R73370 VSS.n20023 VSS.n20022 0.00219014
R73371 VSS.n757 VSS.n756 0.00219014
R73372 VSS.n796 VSS.n795 0.00219014
R73373 VSS.n1818 VSS.n1817 0.00219014
R73374 VSS.n1720 VSS.n1719 0.00219014
R73375 VSS.n1701 VSS.n1700 0.00219014
R73376 VSS.n1672 VSS.n1671 0.00219014
R73377 VSS.n1648 VSS.n1647 0.00219014
R73378 VSS.n1644 VSS.n1643 0.00219014
R73379 VSS.n8627 VSS.n8626 0.00219014
R73380 VSS.n8667 VSS.n8666 0.00219014
R73381 VSS.n8709 VSS.n8708 0.00219014
R73382 VSS.n8120 VSS.n8119 0.00219014
R73383 VSS.n8221 VSS.n8220 0.00219014
R73384 VSS.n8172 VSS.n8171 0.00219014
R73385 VSS.n20243 VSS.n20242 0.00218
R73386 VSS.n2574 VSS.n2545 0.00217143
R73387 VSS.n3184 VSS.n2543 0.00217143
R73388 VSS.n2922 VSS.n2921 0.00217143
R73389 VSS.n2930 VSS.n2926 0.00217143
R73390 VSS.n2941 VSS.n2940 0.00217143
R73391 VSS.n2943 VSS.n2942 0.00217143
R73392 VSS.n2986 VSS.n2985 0.00217143
R73393 VSS.n2994 VSS.n2990 0.00217143
R73394 VSS.n3006 VSS.n3005 0.00217143
R73395 VSS.n3034 VSS.n3033 0.00217143
R73396 VSS.n3042 VSS.n3038 0.00217143
R73397 VSS.n3054 VSS.n3053 0.00217143
R73398 VSS.n2573 VSS.n2556 0.00217143
R73399 VSS.n2570 VSS.n2569 0.00217143
R73400 VSS.n4972 VSS.n4947 0.00217143
R73401 VSS.n5196 VSS.n5192 0.00217143
R73402 VSS.n5204 VSS.n5203 0.00217143
R73403 VSS.n5247 VSS.n5243 0.00217143
R73404 VSS.n5255 VSS.n5254 0.00217143
R73405 VSS.n5281 VSS.n5278 0.00217143
R73406 VSS.n5290 VSS.n5289 0.00217143
R73407 VSS.n4971 VSS.n4967 0.00217143
R73408 VSS.n4962 VSS.n4961 0.00217143
R73409 VSS.n7181 VSS.n7179 0.00217143
R73410 VSS.n7122 VSS.n7120 0.00217143
R73411 VSS.n7519 VSS.n7047 0.00217143
R73412 VSS.n7183 VSS.n7182 0.00217143
R73413 VSS.n7124 VSS.n7123 0.00217143
R73414 VSS.n7082 VSS.n7081 0.00217143
R73415 VSS.n7071 VSS.n7070 0.00217143
R73416 VSS.n7520 VSS.n7046 0.00217143
R73417 VSS.n7533 VSS.n7532 0.00217143
R73418 VSS.n4320 VSS.n4212 0.00217143
R73419 VSS.n4689 VSS.n4688 0.00217143
R73420 VSS.n4462 VSS.n4461 0.00217143
R73421 VSS.n4451 VSS.n4450 0.00217143
R73422 VSS.n4411 VSS.n4410 0.00217143
R73423 VSS.n4400 VSS.n4399 0.00217143
R73424 VSS.n4376 VSS.n4375 0.00217143
R73425 VSS.n4365 VSS.n4364 0.00217143
R73426 VSS.n4340 VSS.n4339 0.00217143
R73427 VSS.n4336 VSS.n4335 0.00217143
R73428 VSS.n4754 VSS.n4753 0.00217143
R73429 VSS.n17979 VSS.n17978 0.00217143
R73430 VSS.n17975 VSS.n17974 0.00217143
R73431 VSS.n17870 VSS.n17867 0.00217143
R73432 VSS.n17866 VSS.n17865 0.00217143
R73433 VSS.n17825 VSS.n17824 0.00217143
R73434 VSS.n17821 VSS.n17820 0.00217143
R73435 VSS.n17809 VSS.n17806 0.00217143
R73436 VSS.n17805 VSS.n17804 0.00217143
R73437 VSS.n17780 VSS.n17779 0.00217143
R73438 VSS.n17776 VSS.n17775 0.00217143
R73439 VSS.n17764 VSS.n17761 0.00217143
R73440 VSS.n17760 VSS.n17759 0.00217143
R73441 VSS.n17732 VSS.n17731 0.00217143
R73442 VSS.n17728 VSS.n17727 0.00217143
R73443 VSS.n17714 VSS.n17713 0.00217143
R73444 VSS.n14454 VSS.n14453 0.00216167
R73445 VSS.n15353 VSS.n15352 0.00216167
R73446 VSS.n8474 VSS.n8473 0.00216167
R73447 VSS.n8555 VSS.n8554 0.00216167
R73448 VSS.n8322 VSS.n8321 0.00216167
R73449 VSS.n8410 VSS.n8409 0.00216167
R73450 VSS.n8366 VSS.n8365 0.00216167
R73451 VSS.n14453 VSS.n2182 0.00216167
R73452 VSS.n8367 VSS.n8366 0.00216167
R73453 VSS.n8411 VSS.n8410 0.00216167
R73454 VSS.n8321 VSS.n8320 0.00216167
R73455 VSS.n8556 VSS.n8555 0.00216167
R73456 VSS.n8473 VSS.n8472 0.00216167
R73457 VSS.n15354 VSS.n15353 0.00216167
R73458 VSS.n19720 VSS.n19719 0.00216167
R73459 VSS.n1669 VSS.n1668 0.00216167
R73460 VSS.n8625 VSS.n8624 0.00216167
R73461 VSS.n8706 VSS.n8705 0.00216167
R73462 VSS.n8118 VSS.n8117 0.00216167
R73463 VSS.n8218 VSS.n8217 0.00216167
R73464 VSS.n8174 VSS.n8173 0.00216167
R73465 VSS.n8117 VSS.n8116 0.00216167
R73466 VSS.n8175 VSS.n8174 0.00216167
R73467 VSS.n8707 VSS.n8706 0.00216167
R73468 VSS.n8219 VSS.n8218 0.00216167
R73469 VSS.n1670 VSS.n1669 0.00216167
R73470 VSS.n19719 VSS.n19718 0.00216167
R73471 VSS.n8624 VSS.n8623 0.00216167
R73472 VSS.n5744 VSS.n5743 0.00215157
R73473 VSS.n13220 VSS.n13219 0.00215157
R73474 VSS.n16192 VSS.n16191 0.00215157
R73475 VSS.n13337 VSS.n13336 0.00215157
R73476 VSS.n21134 VSS.n21133 0.00215157
R73477 VSS.n13480 VSS.n13479 0.00215157
R73478 VSS.n1184 VSS.n1183 0.00215157
R73479 VSS.n3988 VSS.n3987 0.00215128
R73480 VSS.n2350 VSS.n2349 0.00215128
R73481 VSS.n11357 VSS.n11356 0.00215128
R73482 VSS.n5874 VSS.n5873 0.00215128
R73483 VSS.n5872 VSS.n5871 0.00215128
R73484 VSS.n5868 VSS.n5867 0.00215128
R73485 VSS.n5866 VSS.n5865 0.00215128
R73486 VSS.n5736 VSS.n5735 0.00215128
R73487 VSS.n5600 VSS.n5599 0.00215128
R73488 VSS.n5565 VSS.n5564 0.00215128
R73489 VSS.n2351 VSS.n2350 0.00215128
R73490 VSS.n5737 VSS.n5736 0.00215128
R73491 VSS.n11356 VSS.n11355 0.00215128
R73492 VSS.n3989 VSS.n3988 0.00215128
R73493 VSS.n13015 VSS.n13014 0.00215128
R73494 VSS.n13159 VSS.n13158 0.00215128
R73495 VSS.n12852 VSS.n12851 0.00215128
R73496 VSS.n12789 VSS.n12788 0.00215128
R73497 VSS.n12554 VSS.n12553 0.00215128
R73498 VSS.n12230 VSS.n12229 0.00215128
R73499 VSS.n12790 VSS.n12789 0.00215128
R73500 VSS.n12853 VSS.n12852 0.00215128
R73501 VSS.n13158 VSS.n13157 0.00215128
R73502 VSS.n18860 VSS.n18859 0.00215128
R73503 VSS.n2250 VSS.n2249 0.00215128
R73504 VSS.n15158 VSS.n15157 0.00215128
R73505 VSS.n16375 VSS.n16374 0.00215128
R73506 VSS.n16373 VSS.n16372 0.00215128
R73507 VSS.n16369 VSS.n16368 0.00215128
R73508 VSS.n16367 VSS.n16366 0.00215128
R73509 VSS.n16248 VSS.n16247 0.00215128
R73510 VSS.n16246 VSS.n16245 0.00215128
R73511 VSS.n16240 VSS.n16239 0.00215128
R73512 VSS.n16238 VSS.n16237 0.00215128
R73513 VSS.n16235 VSS.n16234 0.00215128
R73514 VSS.n16233 VSS.n16232 0.00215128
R73515 VSS.n16229 VSS.n16228 0.00215128
R73516 VSS.n16227 VSS.n16226 0.00215128
R73517 VSS.n16184 VSS.n16183 0.00215128
R73518 VSS.n16116 VSS.n16115 0.00215128
R73519 VSS.n16081 VSS.n16080 0.00215128
R73520 VSS.n15157 VSS.n15156 0.00215128
R73521 VSS.n16374 VSS.n16373 0.00215128
R73522 VSS.n16368 VSS.n16367 0.00215128
R73523 VSS.n16247 VSS.n16246 0.00215128
R73524 VSS.n16239 VSS.n16238 0.00215128
R73525 VSS.n16185 VSS.n16184 0.00215128
R73526 VSS.n16241 VSS.n16240 0.00215128
R73527 VSS.n16370 VSS.n16369 0.00215128
R73528 VSS.n16249 VSS.n16248 0.00215128
R73529 VSS.n16376 VSS.n16375 0.00215128
R73530 VSS.n2249 VSS.n2248 0.00215128
R73531 VSS.n16234 VSS.n16233 0.00215128
R73532 VSS.n16228 VSS.n16227 0.00215128
R73533 VSS.n5867 VSS.n5866 0.00215128
R73534 VSS.n5873 VSS.n5872 0.00215128
R73535 VSS.n16230 VSS.n16229 0.00215128
R73536 VSS.n5869 VSS.n5868 0.00215128
R73537 VSS.n16236 VSS.n16235 0.00215128
R73538 VSS.n5875 VSS.n5874 0.00215128
R73539 VSS.n21788 VSS.n21787 0.00215128
R73540 VSS.n2299 VSS.n2298 0.00215128
R73541 VSS.n20808 VSS.n20807 0.00215128
R73542 VSS.n21183 VSS.n21182 0.00215128
R73543 VSS.n21182 VSS.n21181 0.00215128
R73544 VSS.n21173 VSS.n21172 0.00215128
R73545 VSS.n21171 VSS.n21170 0.00215128
R73546 VSS.n21126 VSS.n21125 0.00215128
R73547 VSS.n21050 VSS.n21049 0.00215128
R73548 VSS.n21014 VSS.n21013 0.00215128
R73549 VSS.n21127 VSS.n21126 0.00215128
R73550 VSS.n20807 VSS.n20806 0.00215128
R73551 VSS.n21174 VSS.n21173 0.00215128
R73552 VSS.n21184 VSS.n21183 0.00215128
R73553 VSS.n21181 VSS.n21176 0.00215128
R73554 VSS.n21172 VSS.n21171 0.00215128
R73555 VSS.n2298 VSS.n2297 0.00215128
R73556 VSS.n19073 VSS.n19072 0.00215128
R73557 VSS.n17907 VSS.n17906 0.00215128
R73558 VSS.n2011 VSS.n2010 0.00215128
R73559 VSS.n1458 VSS.n1457 0.00215128
R73560 VSS.n1457 VSS.n1456 0.00215128
R73561 VSS.n1450 VSS.n1449 0.00215128
R73562 VSS.n1448 VSS.n1447 0.00215128
R73563 VSS.n1329 VSS.n1328 0.00215128
R73564 VSS.n1327 VSS.n1326 0.00215128
R73565 VSS.n1323 VSS.n1322 0.00215128
R73566 VSS.n1322 VSS.n1321 0.00215128
R73567 VSS.n1316 VSS.n1315 0.00215128
R73568 VSS.n1315 VSS.n1314 0.00215128
R73569 VSS.n1309 VSS.n1308 0.00215128
R73570 VSS.n1300 VSS.n1299 0.00215128
R73571 VSS.n1176 VSS.n1175 0.00215128
R73572 VSS.n1096 VSS.n1095 0.00215128
R73573 VSS.n1060 VSS.n1059 0.00215128
R73574 VSS.n1177 VSS.n1176 0.00215128
R73575 VSS.n1308 VSS.n1301 0.00215128
R73576 VSS.n1301 VSS.n1300 0.00215128
R73577 VSS.n1317 VSS.n1316 0.00215128
R73578 VSS.n1324 VSS.n1323 0.00215128
R73579 VSS.n1328 VSS.n1327 0.00215128
R73580 VSS.n1449 VSS.n1448 0.00215128
R73581 VSS.n1451 VSS.n1450 0.00215128
R73582 VSS.n1330 VSS.n1329 0.00215128
R73583 VSS.n1459 VSS.n1458 0.00215128
R73584 VSS.n1456 VSS.n1453 0.00215128
R73585 VSS.n2012 VSS.n2011 0.00215128
R73586 VSS.n1321 VSS.n1318 0.00215128
R73587 VSS.n1314 VSS.n1311 0.00215128
R73588 VSS.n17906 VSS.n17905 0.00215128
R73589 VSS.n21556 VSS.n21555 0.00215128
R73590 VSS.n21561 VSS.n21560 0.00215128
R73591 VSS.n21514 VSS.n21513 0.00215128
R73592 VSS.n21471 VSS.n21470 0.00215128
R73593 VSS.n21273 VSS.n21272 0.00215128
R73594 VSS.n7573 VSS.n7572 0.00215128
R73595 VSS.n7572 VSS.n7571 0.00215128
R73596 VSS.n21274 VSS.n21273 0.00215128
R73597 VSS.n21515 VSS.n21514 0.00215128
R73598 VSS.n21560 VSS.n21559 0.00215128
R73599 VSS.n21472 VSS.n21471 0.00215128
R73600 VSS.n12231 VSS.n12230 0.00215128
R73601 VSS.n12555 VSS.n12554 0.00215128
R73602 VSS.n16117 VSS.n16116 0.00215128
R73603 VSS.n1097 VSS.n1096 0.00215128
R73604 VSS.n21051 VSS.n21050 0.00215128
R73605 VSS.n5601 VSS.n5600 0.00215128
R73606 VSS.n3789 VSS.n3788 0.00215128
R73607 VSS.n3793 VSS.n3792 0.00215128
R73608 VSS.n4704 VSS.n4703 0.00215128
R73609 VSS.n4765 VSS.n4764 0.00215128
R73610 VSS.n11431 VSS.n11430 0.00215128
R73611 VSS.n11210 VSS.n11209 0.00215128
R73612 VSS.n4703 VSS.n4702 0.00215128
R73613 VSS.n11432 VSS.n11431 0.00215128
R73614 VSS.n11211 VSS.n11210 0.00215128
R73615 VSS.n3792 VSS.n3791 0.00215128
R73616 VSS.n3269 VSS.n3268 0.00215128
R73617 VSS.n549 VSS.n548 0.00215128
R73618 VSS.n490 VSS.n489 0.00215128
R73619 VSS.n10499 VSS.n10498 0.00215128
R73620 VSS.n10178 VSS.n10177 0.00215128
R73621 VSS.n10179 VSS.n10178 0.00215128
R73622 VSS.n491 VSS.n490 0.00215128
R73623 VSS.n550 VSS.n549 0.00215128
R73624 VSS.n6945 VSS.n6944 0.00215128
R73625 VSS.n6843 VSS.n6842 0.00215128
R73626 VSS.n3788 VSS.n3787 0.00215128
R73627 VSS.n21555 VSS.n21554 0.00215128
R73628 VSS.n13014 VSS.n13013 0.00215128
R73629 VSS.n21787 VSS.n21786 0.00215128
R73630 VSS.n19072 VSS.n19071 0.00215128
R73631 VSS.n3268 VSS.n3267 0.00215128
R73632 VSS.n18859 VSS.n18858 0.00215128
R73633 VSS.n8299 VSS.n8298 0.00215
R73634 VSS.n8756 VSS.n8755 0.00215
R73635 VSS.n10828 VSS.n10827 0.00215
R73636 VSS.n2552 DVSS 0.00212857
R73637 VSS.n5654 VSS.n5653 0.00212162
R73638 VSS.n5538 VSS.n5536 0.00212162
R73639 VSS.n16028 VSS.n16026 0.00212162
R73640 VSS.n16042 VSS.n16041 0.00212162
R73641 VSS.n1003 VSS.n1001 0.00212162
R73642 VSS.n1022 VSS.n1020 0.00212162
R73643 VSS.n20910 VSS.n20908 0.00212162
R73644 VSS.n20921 VSS.n20920 0.00212162
R73645 VSS.n8996 VSS.n8995 0.00212
R73646 VSS.n9466 VSS.n9465 0.00212
R73647 VSS.n10639 VSS.n10638 0.00212
R73648 VSS.n3429 VSS.n3428 0.00211972
R73649 VSS.n3431 VSS.n3430 0.00211972
R73650 VSS.n3458 VSS.n3457 0.00211972
R73651 VSS.n2863 VSS.n2862 0.00210714
R73652 VSS.n2677 VSS.n2676 0.00210714
R73653 VSS.n2721 VSS.n2720 0.00210714
R73654 VSS.n2781 VSS.n2780 0.00210714
R73655 VSS.n2946 VSS.n2945 0.00210714
R73656 VSS.n3011 VSS.n3010 0.00210714
R73657 VSS.n3059 VSS.n3058 0.00210714
R73658 VSS.n5139 VSS.n5138 0.00210714
R73659 VSS.n5413 VSS.n5412 0.00210714
R73660 VSS.n4998 VSS.n4997 0.00210714
R73661 VSS.n5028 VSS.n5027 0.00210714
R73662 VSS.n5074 VSS.n5073 0.00210714
R73663 VSS.n7238 VSS.n7237 0.00210714
R73664 VSS.n5915 VSS.n5914 0.00210714
R73665 VSS.n7397 VSS.n7396 0.00210714
R73666 VSS.n7239 VSS.n7236 0.00210714
R73667 VSS.n4515 VSS.n4514 0.00210714
R73668 VSS.n4627 VSS.n4626 0.00210714
R73669 VSS.n4581 VSS.n4580 0.00210714
R73670 VSS.n17549 VSS.n17548 0.00210714
R73671 VSS.n17491 VSS.n17490 0.00210714
R73672 VSS.n17864 VSS.n17863 0.00210714
R73673 VSS.n17803 VSS.n17802 0.00210714
R73674 VSS.n17758 VSS.n17757 0.00210714
R73675 VSS.n18034 VSS.n18033 0.00210714
R73676 VSS.n4059 VSS.n4058 0.00209449
R73677 VSS.n4067 VSS.n4066 0.00209449
R73678 VSS.n11559 VSS.n11558 0.00209449
R73679 VSS.n11567 VSS.n11566 0.00209449
R73680 VSS.n5746 VSS.n5745 0.00209449
R73681 VSS.n5740 VSS.n5739 0.00209449
R73682 VSS.n5551 VSS.n5550 0.00209449
R73683 VSS.n5543 VSS.n5542 0.00209449
R73684 VSS.n9560 VSS.n9559 0.00209449
R73685 VSS.n9552 VSS.n9551 0.00209449
R73686 VSS.n9123 VSS.n9122 0.00209449
R73687 VSS.n9115 VSS.n9114 0.00209449
R73688 VSS.n13095 VSS.n13094 0.00209449
R73689 VSS.n12943 VSS.n12942 0.00209449
R73690 VSS.n12932 VSS.n12931 0.00209449
R73691 VSS.n12725 VSS.n12724 0.00209449
R73692 VSS.n12715 VSS.n12714 0.00209449
R73693 VSS.n12584 VSS.n12583 0.00209449
R73694 VSS.n12579 VSS.n12578 0.00209449
R73695 VSS.n12509 VSS.n12508 0.00209449
R73696 VSS.n12304 VSS.n12303 0.00209449
R73697 VSS.n12286 VSS.n12285 0.00209449
R73698 VSS.n12263 VSS.n12262 0.00209449
R73699 VSS.n12258 VSS.n12257 0.00209449
R73700 VSS.n12257 VSS.n12256 0.00209449
R73701 VSS.n12247 VSS.n12246 0.00209449
R73702 VSS.n11916 VSS.n11915 0.00209449
R73703 VSS.n11911 VSS.n11910 0.00209449
R73704 VSS.n11833 VSS.n11832 0.00209449
R73705 VSS.n11828 VSS.n11827 0.00209449
R73706 VSS.n18930 VSS.n18929 0.00209449
R73707 VSS.n18938 VSS.n18937 0.00209449
R73708 VSS.n15033 VSS.n15032 0.00209449
R73709 VSS.n15042 VSS.n15041 0.00209449
R73710 VSS.n16194 VSS.n16193 0.00209449
R73711 VSS.n16188 VSS.n16187 0.00209449
R73712 VSS.n16061 VSS.n16060 0.00209449
R73713 VSS.n16053 VSS.n16052 0.00209449
R73714 VSS.n9677 VSS.n9676 0.00209449
R73715 VSS.n9669 VSS.n9668 0.00209449
R73716 VSS.n9286 VSS.n9285 0.00209449
R73717 VSS.n9278 VSS.n9277 0.00209449
R73718 VSS.n21868 VSS.n21867 0.00209449
R73719 VSS.n20641 VSS.n20640 0.00209449
R73720 VSS.n20652 VSS.n20651 0.00209449
R73721 VSS.n21136 VSS.n21135 0.00209449
R73722 VSS.n21130 VSS.n21129 0.00209449
R73723 VSS.n20996 VSS.n20995 0.00209449
R73724 VSS.n20985 VSS.n20984 0.00209449
R73725 VSS.n6970 VSS.n6969 0.00209449
R73726 VSS.n6959 VSS.n6958 0.00209449
R73727 VSS.n6610 VSS.n6609 0.00209449
R73728 VSS.n6599 VSS.n6598 0.00209449
R73729 VSS.n19153 VSS.n19152 0.00209449
R73730 VSS.n20108 VSS.n20107 0.00209449
R73731 VSS.n20097 VSS.n20096 0.00209449
R73732 VSS.n1186 VSS.n1185 0.00209449
R73733 VSS.n1180 VSS.n1179 0.00209449
R73734 VSS.n1038 VSS.n1037 0.00209449
R73735 VSS.n1027 VSS.n1026 0.00209449
R73736 VSS.n6868 VSS.n6867 0.00209449
R73737 VSS.n6857 VSS.n6856 0.00209449
R73738 VSS.n6460 VSS.n6459 0.00209449
R73739 VSS.n6449 VSS.n6448 0.00209449
R73740 VSS.n21633 VSS.n21632 0.00209449
R73741 VSS.n21637 VSS.n21636 0.00209449
R73742 VSS.n21360 VSS.n21359 0.00209449
R73743 VSS.n21349 VSS.n21348 0.00209449
R73744 VSS.n7637 VSS.n7636 0.00209449
R73745 VSS.n7648 VSS.n7647 0.00209449
R73746 VSS.n7725 VSS.n7724 0.00209449
R73747 VSS.n7736 VSS.n7735 0.00209449
R73748 VSS.n7814 VSS.n7813 0.00209449
R73749 VSS.n7803 VSS.n7802 0.00209449
R73750 VSS.n3861 VSS.n3860 0.00209449
R73751 VSS.n3866 VSS.n3865 0.00209449
R73752 VSS.n11676 VSS.n11675 0.00209449
R73753 VSS.n11667 VSS.n11666 0.00209449
R73754 VSS.n6119 VSS.n6118 0.00209449
R73755 VSS.n6111 VSS.n6110 0.00209449
R73756 VSS.n6038 VSS.n6037 0.00209449
R73757 VSS.n6030 VSS.n6029 0.00209449
R73758 VSS.n5957 VSS.n5956 0.00209449
R73759 VSS.n5949 VSS.n5948 0.00209449
R73760 VSS.n2629 VSS.n2628 0.00209449
R73761 VSS.n2621 VSS.n2620 0.00209449
R73762 VSS.n633 VSS.n632 0.00209449
R73763 VSS.n625 VSS.n624 0.00209449
R73764 VSS.n10591 VSS.n10590 0.00209449
R73765 VSS.n10583 VSS.n10582 0.00209449
R73766 VSS.n10519 VSS.n10518 0.00209449
R73767 VSS.n10514 VSS.n10513 0.00209449
R73768 VSS.n10455 VSS.n10454 0.00209449
R73769 VSS.n10252 VSS.n10251 0.00209449
R73770 VSS.n10234 VSS.n10233 0.00209449
R73771 VSS.n10211 VSS.n10210 0.00209449
R73772 VSS.n10206 VSS.n10205 0.00209449
R73773 VSS.n10205 VSS.n10204 0.00209449
R73774 VSS.n10196 VSS.n10195 0.00209449
R73775 VSS.n9917 VSS.n9916 0.00209449
R73776 VSS.n9912 VSS.n9911 0.00209449
R73777 VSS.n8906 VSS.n8905 0.00209449
R73778 VSS.n8988 VSS.n8987 0.00209449
R73779 VSS.n20221 VSS.n20220 0.00209
R73780 VSS.n9399 VSS.n9398 0.00209
R73781 VSS.n9345 VSS.n9344 0.00209
R73782 VSS.n8278 VSS.n8277 0.00209
R73783 VSS.n9790 VSS.n9789 0.00209
R73784 VSS.n9736 VSS.n9735 0.00209
R73785 VSS.n8735 VSS.n8734 0.00209
R73786 VSS.n10669 VSS.n10668 0.00209
R73787 VSS.n10731 VSS.n10730 0.00209
R73788 VSS.n10853 VSS.n10852 0.00209
R73789 VSS.n18427 VSS.n18426 0.002075
R73790 VSS.n18431 VSS.n18430 0.002075
R73791 VSS.n17101 VSS.n17100 0.002075
R73792 VSS.n17060 VSS.n17059 0.002075
R73793 VSS.n16961 VSS.n16960 0.002075
R73794 VSS.n14926 VSS.n14923 0.002075
R73795 VSS.n7010 VSS.n7009 0.00207333
R73796 VSS.n7908 VSS.n6346 0.00207333
R73797 VSS.n11089 VSS.n11088 0.00207333
R73798 VSS.n4038 VSS.n4037 0.00206274
R73799 VSS.n17464 VSS.n17463 0.00206274
R73800 VSS.n17320 VSS.n17319 0.00206274
R73801 VSS.n5606 VSS.n5605 0.00206274
R73802 VSS.n5554 VSS.n5553 0.00206274
R73803 VSS.n9045 VSS.n9044 0.00206274
R73804 VSS.n17319 VSS.n17318 0.00206274
R73805 VSS.n4037 VSS.n4036 0.00206274
R73806 VSS.n13067 VSS.n13066 0.00206274
R73807 VSS.n13206 VSS.n13205 0.00206274
R73808 VSS.n13210 VSS.n13209 0.00206274
R73809 VSS.n12987 VSS.n12986 0.00206274
R73810 VSS.n12769 VSS.n12768 0.00206274
R73811 VSS.n12605 VSS.n12604 0.00206274
R73812 VSS.n12287 VSS.n12286 0.00206274
R73813 VSS.n11958 VSS.n11957 0.00206274
R73814 VSS.n11859 VSS.n11858 0.00206274
R73815 VSS.n12988 VSS.n12987 0.00206274
R73816 VSS.n13066 VSS.n13065 0.00206274
R73817 VSS.n13205 VSS.n13204 0.00206274
R73818 VSS.n13209 VSS.n13208 0.00206274
R73819 VSS.n17465 VSS.n17464 0.00206274
R73820 VSS.n5553 VSS.n5552 0.00206274
R73821 VSS.n18909 VSS.n18908 0.00206274
R73822 VSS.n2215 VSS.n2214 0.00206274
R73823 VSS.n14411 VSS.n14410 0.00206274
R73824 VSS.n16122 VSS.n16121 0.00206274
R73825 VSS.n16064 VSS.n16063 0.00206274
R73826 VSS.n9661 VSS.n9660 0.00206274
R73827 VSS.n9188 VSS.n9187 0.00206274
R73828 VSS.n2216 VSS.n2215 0.00206274
R73829 VSS.n14412 VSS.n14411 0.00206274
R73830 VSS.n18908 VSS.n18907 0.00206274
R73831 VSS.n16063 VSS.n16062 0.00206274
R73832 VSS.n16123 VSS.n16122 0.00206274
R73833 VSS.n5607 VSS.n5606 0.00206274
R73834 VSS.n21840 VSS.n21839 0.00206274
R73835 VSS.n13323 VSS.n13322 0.00206274
R73836 VSS.n13327 VSS.n13326 0.00206274
R73837 VSS.n20597 VSS.n20596 0.00206274
R73838 VSS.n21056 VSS.n21055 0.00206274
R73839 VSS.n21002 VSS.n20997 0.00206274
R73840 VSS.n6950 VSS.n6949 0.00206274
R73841 VSS.n6678 VSS.n6677 0.00206274
R73842 VSS.n21057 VSS.n21056 0.00206274
R73843 VSS.n20596 VSS.n20595 0.00206274
R73844 VSS.n13322 VSS.n13321 0.00206274
R73845 VSS.n21839 VSS.n21838 0.00206274
R73846 VSS.n13326 VSS.n13325 0.00206274
R73847 VSS.n21003 VSS.n21002 0.00206274
R73848 VSS.n19125 VSS.n19124 0.00206274
R73849 VSS.n17946 VSS.n17945 0.00206274
R73850 VSS.n17941 VSS.n17940 0.00206274
R73851 VSS.n20159 VSS.n20158 0.00206274
R73852 VSS.n1102 VSS.n1101 0.00206274
R73853 VSS.n1049 VSS.n1048 0.00206274
R73854 VSS.n6849 VSS.n6848 0.00206274
R73855 VSS.n6528 VSS.n6527 0.00206274
R73856 VSS.n1103 VSS.n1102 0.00206274
R73857 VSS.n20158 VSS.n20157 0.00206274
R73858 VSS.n19124 VSS.n19123 0.00206274
R73859 VSS.n17942 VSS.n17941 0.00206274
R73860 VSS.n17945 VSS.n17944 0.00206274
R73861 VSS.n1048 VSS.n1039 0.00206274
R73862 VSS.n21611 VSS.n21610 0.00206274
R73863 VSS.n21404 VSS.n21403 0.00206274
R73864 VSS.n7593 VSS.n7592 0.00206274
R73865 VSS.n7681 VSS.n7680 0.00206274
R73866 VSS.n7769 VSS.n7768 0.00206274
R73867 VSS.n21405 VSS.n21404 0.00206274
R73868 VSS.n21610 VSS.n21609 0.00206274
R73869 VSS.n11941 VSS.n11940 0.00206274
R73870 VSS.n7768 VSS.n7767 0.00206274
R73871 VSS.n6677 VSS.n6676 0.00206274
R73872 VSS.n6527 VSS.n6526 0.00206274
R73873 VSS.n9187 VSS.n9186 0.00206274
R73874 VSS.n9044 VSS.n9043 0.00206274
R73875 VSS.n11858 VSS.n11857 0.00206274
R73876 VSS.n12288 VSS.n12287 0.00206274
R73877 VSS.n9544 VSS.n9543 0.00206274
R73878 VSS.n12606 VSS.n12605 0.00206274
R73879 VSS.n7680 VSS.n7679 0.00206274
R73880 VSS.n6848 VSS.n6847 0.00206274
R73881 VSS.n6951 VSS.n6950 0.00206274
R73882 VSS.n12770 VSS.n12769 0.00206274
R73883 VSS.n7592 VSS.n7591 0.00206274
R73884 VSS.n3840 VSS.n3839 0.00206274
R73885 VSS.n11729 VSS.n11728 0.00206274
R73886 VSS.n11192 VSS.n11191 0.00206274
R73887 VSS.n6080 VSS.n6079 0.00206274
R73888 VSS.n5999 VSS.n5998 0.00206274
R73889 VSS.n6000 VSS.n5999 0.00206274
R73890 VSS.n6081 VSS.n6080 0.00206274
R73891 VSS.n11730 VSS.n11729 0.00206274
R73892 VSS.n3839 VSS.n3838 0.00206274
R73893 VSS.n11193 VSS.n11192 0.00206274
R73894 VSS.n2655 VSS.n2654 0.00206274
R73895 VSS.n2654 VSS.n2653 0.00206274
R73896 VSS.n673 VSS.n672 0.00206274
R73897 VSS.n472 VSS.n471 0.00206274
R73898 VSS.n10539 VSS.n10538 0.00206274
R73899 VSS.n10235 VSS.n10234 0.00206274
R73900 VSS.n9960 VSS.n9959 0.00206274
R73901 VSS.n9942 VSS.n9941 0.00206274
R73902 VSS.n10236 VSS.n10235 0.00206274
R73903 VSS.n9943 VSS.n9942 0.00206274
R73904 VSS.n9961 VSS.n9960 0.00206274
R73905 VSS.n8916 VSS.n8915 0.00206274
R73906 VSS.n10540 VSS.n10539 0.00206274
R73907 VSS.n672 VSS.n671 0.00206274
R73908 VSS.n473 VSS.n472 0.00206274
R73909 VSS.n6757 VSS.n6756 0.00206
R73910 VSS.n6697 VSS.n6696 0.00206
R73911 VSS.n8073 VSS.n8072 0.00206
R73912 VSS.n8013 VSS.n8012 0.00206
R73913 VSS.n10942 VSS.n10941 0.00206
R73914 VSS.n11010 VSS.n11009 0.00206
R73915 VSS.n8611 VSS.n8610 0.00205609
R73916 VSS.n8610 VSS.n8609 0.00205609
R73917 VSS.n18827 VSS.n18826 0.00205609
R73918 VSS.n18405 VSS.n18404 0.00205609
R73919 VSS.n14889 VSS.n14888 0.00205609
R73920 VSS.n16930 VSS.n16929 0.00205609
R73921 VSS.n8460 VSS.n8459 0.00205609
R73922 VSS.n8541 VSS.n8540 0.00205609
R73923 VSS.n8308 VSS.n8307 0.00205609
R73924 VSS.n8396 VSS.n8395 0.00205609
R73925 VSS.n8380 VSS.n8379 0.00205609
R73926 VSS.n14888 VSS.n14887 0.00205609
R73927 VSS.n16931 VSS.n16930 0.00205609
R73928 VSS.n14863 VSS.n14862 0.00205609
R73929 VSS.n17078 VSS.n17077 0.00205609
R73930 VSS.n18826 VSS.n18825 0.00205609
R73931 VSS.n8397 VSS.n8396 0.00205609
R73932 VSS.n8381 VSS.n8380 0.00205609
R73933 VSS.n8542 VSS.n8541 0.00205609
R73934 VSS.n8307 VSS.n8306 0.00205609
R73935 VSS.n8459 VSS.n8458 0.00205609
R73936 VSS.n19499 VSS.n19498 0.00205609
R73937 VSS.n19617 VSS.n19616 0.00205609
R73938 VSS.n19960 VSS.n19959 0.00205609
R73939 VSS.n19986 VSS.n19985 0.00205609
R73940 VSS.n8692 VSS.n8691 0.00205609
R73941 VSS.n8104 VSS.n8103 0.00205609
R73942 VSS.n8204 VSS.n8203 0.00205609
R73943 VSS.n8188 VSS.n8187 0.00205609
R73944 VSS.n8693 VSS.n8692 0.00205609
R73945 VSS.n8205 VSS.n8204 0.00205609
R73946 VSS.n8103 VSS.n8102 0.00205609
R73947 VSS.n8189 VSS.n8188 0.00205609
R73948 VSS.n19985 VSS.n19984 0.00205609
R73949 VSS.n19934 VSS.n19933 0.00205609
R73950 VSS.n19887 VSS.n19886 0.00205609
R73951 VSS.n19959 VSS.n19958 0.00205609
R73952 VSS.n19498 VSS.n19497 0.00205609
R73953 VSS.n3529 VSS.n3528 0.0020493
R73954 VSS.n3532 VSS.n3531 0.0020493
R73955 VSS.n3588 VSS.n3587 0.0020493
R73956 VSS.n3591 VSS.n3590 0.0020493
R73957 VSS.n3631 VSS.n3630 0.0020493
R73958 VSS.n3634 VSS.n3633 0.0020493
R73959 VSS.n2540 VSS.n2536 0.00204286
R73960 VSS.n2541 VSS.n2535 0.00204286
R73961 VSS.n2674 VSS.n2673 0.00204286
R73962 VSS.n2718 VSS.n2717 0.00204286
R73963 VSS.n2778 VSS.n2777 0.00204286
R73964 VSS.n2867 VSS.n2866 0.00204286
R73965 VSS.n2871 VSS.n2870 0.00204286
R73966 VSS.n5410 VSS.n4944 0.00204286
R73967 VSS.n5412 VSS.n5411 0.00204286
R73968 VSS.n5001 VSS.n4998 0.00204286
R73969 VSS.n5031 VSS.n5028 0.00204286
R73970 VSS.n5077 VSS.n5074 0.00204286
R73971 VSS.n5143 VSS.n5142 0.00204286
R73972 VSS.n5146 VSS.n5145 0.00204286
R73973 VSS.n5920 VSS.n5916 0.00204286
R73974 VSS.n5921 VSS.n5915 0.00204286
R73975 VSS.n7396 VSS.n7395 0.00204286
R73976 VSS.n7362 VSS.n7361 0.00204286
R73977 VSS.n7356 VSS.n7355 0.00204286
R73978 VSS.n7308 VSS.n7307 0.00204286
R73979 VSS.n7302 VSS.n7301 0.00204286
R73980 VSS.n7177 VSS.n7176 0.00204286
R73981 VSS.n7118 VSS.n7117 0.00204286
R73982 VSS.n2445 VSS.n2443 0.00204286
R73983 VSS.n4692 VSS.n4691 0.00204286
R73984 VSS.n4626 VSS.n4625 0.00204286
R73985 VSS.n4580 VSS.n4579 0.00204286
R73986 VSS.n4512 VSS.n4511 0.00204286
R73987 VSS.n4509 VSS.n4508 0.00204286
R73988 VSS.n4751 VSS.n4746 0.00204286
R73989 VSS.n17551 VSS.n17550 0.00204286
R73990 VSS.n17493 VSS.n17492 0.00204286
R73991 VSS.n18031 VSS.n18030 0.00204286
R73992 VSS.n18028 VSS.n18027 0.00204286
R73993 VSS.n4750 VSS.n4747 0.00204286
R73994 VSS.n8887 VSS.n8878 0.00203846
R73995 VSS.n11994 VSS.n11993 0.00203846
R73996 VSS.n9852 VSS.n9831 0.00203846
R73997 VSS.n12656 VSS.n12655 0.00203846
R73998 VSS.n158 VSS.n155 0.00200838
R73999 VSS.n324 VSS.n321 0.00200838
R74000 VSS.n8927 VSS.n8926 0.002
R74001 VSS.n9461 VSS.n9460 0.002
R74002 VSS.n10634 VSS.n10633 0.002
R74003 VSS.n3243 VSS.n3242 0.00197887
R74004 VSS.n3291 VSS.n3290 0.00197887
R74005 VSS.n3326 VSS.n3325 0.00197887
R74006 VSS.n3329 VSS.n3328 0.00197887
R74007 VSS.n3380 VSS.n3379 0.00197887
R74008 VSS.n3383 VSS.n3382 0.00197887
R74009 VSS.n3478 VSS.n3475 0.00197887
R74010 VSS.n18703 VSS.n18702 0.00197887
R74011 VSS.n18716 VSS.n18715 0.00197887
R74012 VSS.n18777 VSS.n18776 0.00197887
R74013 VSS.n18472 VSS.n18471 0.00197887
R74014 VSS.n18445 VSS.n18444 0.00197887
R74015 VSS.n18187 VSS.n18186 0.00197887
R74016 VSS.n18180 VSS.n18179 0.00197887
R74017 VSS.n18151 VSS.n18150 0.00197887
R74018 VSS.n17129 VSS.n17128 0.00197887
R74019 VSS.n17127 VSS.n17126 0.00197887
R74020 VSS.n17126 VSS.n17125 0.00197887
R74021 VSS.n17071 VSS.n17070 0.00197887
R74022 VSS.n17068 VSS.n17067 0.00197887
R74023 VSS.n14859 VSS.n14858 0.00197887
R74024 VSS.n16934 VSS.n16933 0.00197887
R74025 VSS.n16927 VSS.n16926 0.00197887
R74026 VSS.n16903 VSS.n16902 0.00197887
R74027 VSS.n16640 VSS.n16639 0.00197887
R74028 VSS.n16543 VSS.n16542 0.00197887
R74029 VSS.n15550 VSS.n15549 0.00197887
R74030 VSS.n15466 VSS.n15465 0.00197887
R74031 VSS.n15407 VSS.n15406 0.00197887
R74032 VSS.n15342 VSS.n15341 0.00197887
R74033 VSS.n8335 VSS.n8334 0.00197887
R74034 VSS.n19185 VSS.n19184 0.00197887
R74035 VSS.n19198 VSS.n19197 0.00197887
R74036 VSS.n19449 VSS.n19448 0.00197887
R74037 VSS.n19567 VSS.n19566 0.00197887
R74038 VSS.n19594 VSS.n19593 0.00197887
R74039 VSS.n19669 VSS.n19668 0.00197887
R74040 VSS.n19676 VSS.n19675 0.00197887
R74041 VSS.n19705 VSS.n19704 0.00197887
R74042 VSS.n19866 VSS.n19865 0.00197887
R74043 VSS.n19868 VSS.n19867 0.00197887
R74044 VSS.n19869 VSS.n19868 0.00197887
R74045 VSS.n19894 VSS.n19893 0.00197887
R74046 VSS.n19897 VSS.n19896 0.00197887
R74047 VSS.n19930 VSS.n19929 0.00197887
R74048 VSS.n19982 VSS.n19981 0.00197887
R74049 VSS.n19989 VSS.n19988 0.00197887
R74050 VSS.n20013 VSS.n20012 0.00197887
R74051 VSS.n758 VSS.n757 0.00197887
R74052 VSS.n795 VSS.n794 0.00197887
R74053 VSS.n1838 VSS.n1837 0.00197887
R74054 VSS.n1768 VSS.n1767 0.00197887
R74055 VSS.n1723 VSS.n1722 0.00197887
R74056 VSS.n1658 VSS.n1657 0.00197887
R74057 VSS.n8131 VSS.n8130 0.00197887
R74058 VSS.n2832 VSS.n2831 0.00197857
R74059 VSS.n2827 VSS.n2826 0.00197857
R74060 VSS.n2865 VSS.n2864 0.00197857
R74061 VSS.n5114 VSS.n5113 0.00197857
R74062 VSS.n5111 VSS.n5110 0.00197857
R74063 VSS.n5116 VSS.n5115 0.00197857
R74064 VSS.n5141 VSS.n5140 0.00197857
R74065 VSS.n7262 VSS.n7261 0.00197857
R74066 VSS.n7263 VSS.n7260 0.00197857
R74067 VSS.n7246 VSS.n7245 0.00197857
R74068 VSS.n4540 VSS.n4539 0.00197857
R74069 VSS.n4544 VSS.n4543 0.00197857
R74070 VSS.n4541 VSS.n4538 0.00197857
R74071 VSS.n4516 VSS.n4513 0.00197857
R74072 VSS.n18069 VSS.n18068 0.00197857
R74073 VSS.n18035 VSS.n18032 0.00197857
R74074 VSS.n18065 VSS.n18064 0.00197857
R74075 VSS.n17437 VSS.n17436 0.0019742
R74076 VSS.n11542 VSS.n11541 0.0019742
R74077 VSS.n11584 VSS.n11583 0.0019742
R74078 VSS.n5580 VSS.n5579 0.0019742
R74079 VSS.n9490 VSS.n9489 0.0019742
R74080 VSS.n9576 VSS.n9575 0.0019742
R74081 VSS.n9031 VSS.n9030 0.0019742
R74082 VSS.n9139 VSS.n9138 0.0019742
R74083 VSS.n9098 VSS.n9097 0.0019742
R74084 VSS.n11583 VSS.n11582 0.0019742
R74085 VSS.n11543 VSS.n11542 0.0019742
R74086 VSS.n13236 VSS.n13235 0.0019742
R74087 VSS.n12959 VSS.n12958 0.0019742
R74088 VSS.n12915 VSS.n12914 0.0019742
R74089 VSS.n12741 VSS.n12740 0.0019742
R74090 VSS.n12698 VSS.n12697 0.0019742
R74091 VSS.n11812 VSS.n11811 0.0019742
R74092 VSS.n11810 VSS.n11809 0.0019742
R74093 VSS.n12916 VSS.n12915 0.0019742
R74094 VSS.n12960 VSS.n12959 0.0019742
R74095 VSS.n13235 VSS.n13234 0.0019742
R74096 VSS.n17438 VSS.n17437 0.0019742
R74097 VSS.n2188 VSS.n2187 0.0019742
R74098 VSS.n15017 VSS.n15016 0.0019742
R74099 VSS.n15059 VSS.n15058 0.0019742
R74100 VSS.n16096 VSS.n16095 0.0019742
R74101 VSS.n9607 VSS.n9606 0.0019742
R74102 VSS.n9693 VSS.n9692 0.0019742
R74103 VSS.n9174 VSS.n9173 0.0019742
R74104 VSS.n9302 VSS.n9301 0.0019742
R74105 VSS.n9261 VSS.n9260 0.0019742
R74106 VSS.n2189 VSS.n2188 0.0019742
R74107 VSS.n15058 VSS.n15057 0.0019742
R74108 VSS.n15016 VSS.n15015 0.0019742
R74109 VSS.n13353 VSS.n13352 0.0019742
R74110 VSS.n20625 VSS.n20624 0.0019742
R74111 VSS.n20669 VSS.n20668 0.0019742
R74112 VSS.n21028 VSS.n21027 0.0019742
R74113 VSS.n6921 VSS.n6920 0.0019742
R74114 VSS.n6986 VSS.n6985 0.0019742
R74115 VSS.n6662 VSS.n6661 0.0019742
R74116 VSS.n6626 VSS.n6625 0.0019742
R74117 VSS.n6582 VSS.n6581 0.0019742
R74118 VSS.n13352 VSS.n13351 0.0019742
R74119 VSS.n20668 VSS.n20667 0.0019742
R74120 VSS.n20624 VSS.n20623 0.0019742
R74121 VSS.n13496 VSS.n13495 0.0019742
R74122 VSS.n20124 VSS.n20123 0.0019742
R74123 VSS.n20080 VSS.n20079 0.0019742
R74124 VSS.n1074 VSS.n1073 0.0019742
R74125 VSS.n6798 VSS.n6797 0.0019742
R74126 VSS.n6884 VSS.n6883 0.0019742
R74127 VSS.n6512 VSS.n6511 0.0019742
R74128 VSS.n6476 VSS.n6475 0.0019742
R74129 VSS.n6432 VSS.n6431 0.0019742
R74130 VSS.n20081 VSS.n20080 0.0019742
R74131 VSS.n20125 VSS.n20124 0.0019742
R74132 VSS.n13495 VSS.n13494 0.0019742
R74133 VSS.n21376 VSS.n21375 0.0019742
R74134 VSS.n21332 VSS.n21331 0.0019742
R74135 VSS.n7621 VSS.n7620 0.0019742
R74136 VSS.n7665 VSS.n7664 0.0019742
R74137 VSS.n7709 VSS.n7708 0.0019742
R74138 VSS.n7753 VSS.n7752 0.0019742
R74139 VSS.n7830 VSS.n7829 0.0019742
R74140 VSS.n7786 VSS.n7785 0.0019742
R74141 VSS.n21333 VSS.n21332 0.0019742
R74142 VSS.n21377 VSS.n21376 0.0019742
R74143 VSS.n9262 VSS.n9261 0.0019742
R74144 VSS.n11813 VSS.n11812 0.0019742
R74145 VSS.n11811 VSS.n11810 0.0019742
R74146 VSS.n7831 VSS.n7830 0.0019742
R74147 VSS.n11908 VSS.n11907 0.0019742
R74148 VSS.n6627 VSS.n6626 0.0019742
R74149 VSS.n6477 VSS.n6476 0.0019742
R74150 VSS.n9303 VSS.n9302 0.0019742
R74151 VSS.n9140 VSS.n9139 0.0019742
R74152 VSS.n7787 VSS.n7786 0.0019742
R74153 VSS.n6583 VSS.n6582 0.0019742
R74154 VSS.n6433 VSS.n6432 0.0019742
R74155 VSS.n9099 VSS.n9098 0.0019742
R74156 VSS.n9173 VSS.n9172 0.0019742
R74157 VSS.n7752 VSS.n7751 0.0019742
R74158 VSS.n9030 VSS.n9029 0.0019742
R74159 VSS.n7708 VSS.n7707 0.0019742
R74160 VSS.n6987 VSS.n6986 0.0019742
R74161 VSS.n6885 VSS.n6884 0.0019742
R74162 VSS.n9694 VSS.n9693 0.0019742
R74163 VSS.n9577 VSS.n9576 0.0019742
R74164 VSS.n6661 VSS.n6660 0.0019742
R74165 VSS.n6511 VSS.n6510 0.0019742
R74166 VSS.n9489 VSS.n9488 0.0019742
R74167 VSS.n9606 VSS.n9605 0.0019742
R74168 VSS.n6797 VSS.n6796 0.0019742
R74169 VSS.n6920 VSS.n6919 0.0019742
R74170 VSS.n12699 VSS.n12698 0.0019742
R74171 VSS.n7664 VSS.n7663 0.0019742
R74172 VSS.n7620 VSS.n7619 0.0019742
R74173 VSS.n12742 VSS.n12741 0.0019742
R74174 VSS.n21029 VSS.n21028 0.0019742
R74175 VSS.n1075 VSS.n1074 0.0019742
R74176 VSS.n16097 VSS.n16096 0.0019742
R74177 VSS.n5581 VSS.n5580 0.0019742
R74178 VSS.n11692 VSS.n11691 0.0019742
R74179 VSS.n11650 VSS.n11649 0.0019742
R74180 VSS.n6135 VSS.n6134 0.0019742
R74181 VSS.n6094 VSS.n6093 0.0019742
R74182 VSS.n6054 VSS.n6053 0.0019742
R74183 VSS.n6013 VSS.n6012 0.0019742
R74184 VSS.n5973 VSS.n5972 0.0019742
R74185 VSS.n5932 VSS.n5931 0.0019742
R74186 VSS.n11651 VSS.n11650 0.0019742
R74187 VSS.n6095 VSS.n6094 0.0019742
R74188 VSS.n6014 VSS.n6013 0.0019742
R74189 VSS.n5933 VSS.n5932 0.0019742
R74190 VSS.n6055 VSS.n6054 0.0019742
R74191 VSS.n5974 VSS.n5973 0.0019742
R74192 VSS.n6136 VSS.n6135 0.0019742
R74193 VSS.n11693 VSS.n11692 0.0019742
R74194 VSS.n649 VSS.n648 0.0019742
R74195 VSS.n608 VSS.n607 0.0019742
R74196 VSS.n10607 VSS.n10606 0.0019742
R74197 VSS.n10566 VSS.n10565 0.0019742
R74198 VSS.n9908 VSS.n9907 0.0019742
R74199 VSS.n8918 VSS.n8917 0.0019742
R74200 VSS.n8840 VSS.n8839 0.0019742
R74201 VSS.n10567 VSS.n10566 0.0019742
R74202 VSS.n9909 VSS.n9908 0.0019742
R74203 VSS.n10608 VSS.n10607 0.0019742
R74204 VSS.n609 VSS.n608 0.0019742
R74205 VSS.n650 VSS.n649 0.0019742
R74206 VSS.n7885 VSS.n7884 0.00197
R74207 VSS.n7978 VSS.n7977 0.00197
R74208 VSS.n11050 VSS.n11049 0.00197
R74209 VSS.n6320 VSS.n6319 0.00196667
R74210 VSS.n6345 VSS.n6344 0.00196667
R74211 VSS.n11114 VSS.n11113 0.00196667
R74212 VSS.n15492 VSS.n15489 0.00195724
R74213 VSS.n1793 VSS.n1792 0.00195724
R74214 VSS.n15489 VSS.n15488 0.00195724
R74215 VSS.n1794 VSS.n1793 0.00195724
R74216 VSS.n18182 VSS.n18181 0.00195058
R74217 VSS.n19674 VSS.n19673 0.00195058
R74218 VSS.n18798 VSS.n18797 0.0019505
R74219 VSS.n18838 VSS.n18837 0.0019505
R74220 VSS.n15369 VSS.n15368 0.0019505
R74221 VSS.n8571 VSS.n8570 0.0019505
R74222 VSS.n8426 VSS.n8425 0.0019505
R74223 VSS.n14897 VSS.n14896 0.0019505
R74224 VSS.n8427 VSS.n8426 0.0019505
R74225 VSS.n8572 VSS.n8571 0.0019505
R74226 VSS.n15370 VSS.n15369 0.0019505
R74227 VSS.n19510 VSS.n19509 0.0019505
R74228 VSS.n19968 VSS.n19967 0.0019505
R74229 VSS.n1686 VSS.n1685 0.0019505
R74230 VSS.n8722 VSS.n8721 0.0019505
R74231 VSS.n8234 VSS.n8233 0.0019505
R74232 VSS.n8723 VSS.n8722 0.0019505
R74233 VSS.n8235 VSS.n8234 0.0019505
R74234 VSS.n1685 VSS.n1684 0.0019505
R74235 VSS.n19470 VSS.n19469 0.0019505
R74236 VSS.n19511 VSS.n19510 0.0019505
R74237 VSS.n18839 VSS.n18838 0.0019505
R74238 VSS.n10652 VSS.n10651 0.00194
R74239 VSS.n9410 VSS.n9014 0.00194
R74240 VSS.n9802 VSS.n9476 0.00194
R74241 VSS.n10654 VSS.n10653 0.00194
R74242 VSS.n3962 VSS.n3961 0.00191732
R74243 VSS.n11540 VSS.n11539 0.00191732
R74244 VSS.n11586 VSS.n11585 0.00191732
R74245 VSS.n5743 VSS.n5742 0.00191732
R74246 VSS.n5627 VSS.n5626 0.00191732
R74247 VSS.n5610 VSS.n5609 0.00191732
R74248 VSS.n5583 VSS.n5582 0.00191732
R74249 VSS.n5559 VSS.n5558 0.00191732
R74250 VSS.n5555 VSS.n5554 0.00191732
R74251 VSS.n9492 VSS.n9491 0.00191732
R74252 VSS.n9541 VSS.n9540 0.00191732
R74253 VSS.n9579 VSS.n9578 0.00191732
R74254 VSS.n9033 VSS.n9032 0.00191732
R74255 VSS.n9142 VSS.n9141 0.00191732
R74256 VSS.n9096 VSS.n9095 0.00191732
R74257 VSS.n12962 VSS.n12961 0.00191732
R74258 VSS.n12913 VSS.n12912 0.00191732
R74259 VSS.n12744 VSS.n12743 0.00191732
R74260 VSS.n12696 VSS.n12695 0.00191732
R74261 VSS.n12689 VSS.n12688 0.00191732
R74262 VSS.n12560 VSS.n12559 0.00191732
R74263 VSS.n12529 VSS.n12528 0.00191732
R74264 VSS.n12322 VSS.n12321 0.00191732
R74265 VSS.n12277 VSS.n12276 0.00191732
R74266 VSS.n12256 VSS.n12255 0.00191732
R74267 VSS.n11967 VSS.n11966 0.00191732
R74268 VSS.n11932 VSS.n11931 0.00191732
R74269 VSS.n11914 VSS.n11913 0.00191732
R74270 VSS.n11805 VSS.n11804 0.00191732
R74271 VSS.n18963 VSS.n18962 0.00191732
R74272 VSS.n15014 VSS.n15013 0.00191732
R74273 VSS.n15061 VSS.n15060 0.00191732
R74274 VSS.n16191 VSS.n16190 0.00191732
R74275 VSS.n16149 VSS.n16148 0.00191732
R74276 VSS.n16126 VSS.n16125 0.00191732
R74277 VSS.n16099 VSS.n16098 0.00191732
R74278 VSS.n16069 VSS.n16068 0.00191732
R74279 VSS.n16065 VSS.n16064 0.00191732
R74280 VSS.n9609 VSS.n9608 0.00191732
R74281 VSS.n9658 VSS.n9657 0.00191732
R74282 VSS.n9696 VSS.n9695 0.00191732
R74283 VSS.n9176 VSS.n9175 0.00191732
R74284 VSS.n9305 VSS.n9304 0.00191732
R74285 VSS.n9259 VSS.n9258 0.00191732
R74286 VSS.n20622 VSS.n20621 0.00191732
R74287 VSS.n20671 VSS.n20670 0.00191732
R74288 VSS.n21133 VSS.n21132 0.00191732
R74289 VSS.n21077 VSS.n21076 0.00191732
R74290 VSS.n21060 VSS.n21059 0.00191732
R74291 VSS.n21031 VSS.n21030 0.00191732
R74292 VSS.n21008 VSS.n21007 0.00191732
R74293 VSS.n21004 VSS.n21003 0.00191732
R74294 VSS.n6923 VSS.n6922 0.00191732
R74295 VSS.n6947 VSS.n6946 0.00191732
R74296 VSS.n6989 VSS.n6988 0.00191732
R74297 VSS.n6664 VSS.n6663 0.00191732
R74298 VSS.n6629 VSS.n6628 0.00191732
R74299 VSS.n6580 VSS.n6579 0.00191732
R74300 VSS.n20127 VSS.n20126 0.00191732
R74301 VSS.n20078 VSS.n20077 0.00191732
R74302 VSS.n1183 VSS.n1182 0.00191732
R74303 VSS.n1129 VSS.n1128 0.00191732
R74304 VSS.n1106 VSS.n1105 0.00191732
R74305 VSS.n1077 VSS.n1076 0.00191732
R74306 VSS.n1054 VSS.n1053 0.00191732
R74307 VSS.n1050 VSS.n1049 0.00191732
R74308 VSS.n6800 VSS.n6799 0.00191732
R74309 VSS.n6845 VSS.n6844 0.00191732
R74310 VSS.n6887 VSS.n6886 0.00191732
R74311 VSS.n6514 VSS.n6513 0.00191732
R74312 VSS.n6479 VSS.n6478 0.00191732
R74313 VSS.n6430 VSS.n6429 0.00191732
R74314 VSS.n21644 VSS.n21643 0.00191732
R74315 VSS.n21647 VSS.n21646 0.00191732
R74316 VSS.n21648 VSS.n21647 0.00191732
R74317 VSS.n21656 VSS.n21655 0.00191732
R74318 VSS.n21658 VSS.n21657 0.00191732
R74319 VSS.n21379 VSS.n21378 0.00191732
R74320 VSS.n21330 VSS.n21329 0.00191732
R74321 VSS.n7618 VSS.n7617 0.00191732
R74322 VSS.n7667 VSS.n7666 0.00191732
R74323 VSS.n7706 VSS.n7705 0.00191732
R74324 VSS.n7755 VSS.n7754 0.00191732
R74325 VSS.n7833 VSS.n7832 0.00191732
R74326 VSS.n7784 VSS.n7783 0.00191732
R74327 VSS.n3873 VSS.n3872 0.00191732
R74328 VSS.n3876 VSS.n3875 0.00191732
R74329 VSS.n3877 VSS.n3876 0.00191732
R74330 VSS.n3885 VSS.n3884 0.00191732
R74331 VSS.n3887 VSS.n3886 0.00191732
R74332 VSS.n11695 VSS.n11694 0.00191732
R74333 VSS.n11648 VSS.n11647 0.00191732
R74334 VSS.n6138 VSS.n6137 0.00191732
R74335 VSS.n6092 VSS.n6091 0.00191732
R74336 VSS.n6057 VSS.n6056 0.00191732
R74337 VSS.n6011 VSS.n6010 0.00191732
R74338 VSS.n5976 VSS.n5975 0.00191732
R74339 VSS.n5930 VSS.n5929 0.00191732
R74340 VSS.n2596 VSS.n2595 0.00191732
R74341 VSS.n652 VSS.n651 0.00191732
R74342 VSS.n606 VSS.n605 0.00191732
R74343 VSS.n10610 VSS.n10609 0.00191732
R74344 VSS.n10564 VSS.n10563 0.00191732
R74345 VSS.n10557 VSS.n10556 0.00191732
R74346 VSS.n10504 VSS.n10503 0.00191732
R74347 VSS.n10474 VSS.n10473 0.00191732
R74348 VSS.n10268 VSS.n10267 0.00191732
R74349 VSS.n10226 VSS.n10225 0.00191732
R74350 VSS.n10204 VSS.n10203 0.00191732
R74351 VSS.n9970 VSS.n9969 0.00191732
R74352 VSS.n9933 VSS.n9932 0.00191732
R74353 VSS.n9915 VSS.n9914 0.00191732
R74354 VSS.n8967 VSS.n8966 0.00191732
R74355 VSS.n2681 VSS.n2678 0.00191429
R74356 VSS.n2726 VSS.n2722 0.00191429
R74357 VSS.n2786 VSS.n2782 0.00191429
R74358 VSS.n2853 VSS.n2852 0.00191429
R74359 VSS.n5130 VSS.n5129 0.00191429
R74360 VSS.n7169 VSS.n7168 0.00191429
R74361 VSS.n7166 VSS.n7165 0.00191429
R74362 VSS.n7110 VSS.n7109 0.00191429
R74363 VSS.n7107 VSS.n7106 0.00191429
R74364 VSS.n4525 VSS.n4524 0.00191429
R74365 VSS.n17547 VSS.n17546 0.00191429
R74366 VSS.n17489 VSS.n17488 0.00191429
R74367 VSS.n18045 VSS.n18044 0.00191429
R74368 VSS.n13659 VSS.n13658 0.00191342
R74369 VSS.n2925 VSS.n2924 0.0019116
R74370 VSS.n7945 DVSS 0.00191
R74371 VSS.n3220 VSS.n3219 0.00190845
R74372 VSS.n3424 VSS.n3423 0.00190845
R74373 VSS.n3482 VSS.n3481 0.00190845
R74374 VSS.n14153 VSS.n14152 0.00189982
R74375 VSS.n14203 VSS.n14202 0.00189982
R74376 VSS.n13672 VSS.n13671 0.00189982
R74377 VSS.n14204 VSS.n14203 0.00189982
R74378 VSS.n13673 VSS.n13672 0.00189982
R74379 VSS.n14122 VSS.n14121 0.00189982
R74380 VSS.n14123 VSS.n14122 0.00189982
R74381 VSS.n11557 VSS.n11556 0.00188565
R74382 VSS.n11569 VSS.n11568 0.00188565
R74383 VSS.n5540 VSS.n5539 0.00188565
R74384 VSS.n9562 VSS.n9561 0.00188565
R74385 VSS.n9017 VSS.n9016 0.00188565
R74386 VSS.n9125 VSS.n9124 0.00188565
R74387 VSS.n9112 VSS.n9111 0.00188565
R74388 VSS.n11570 VSS.n11569 0.00188565
R74389 VSS.n11556 VSS.n11555 0.00188565
R74390 VSS.n12945 VSS.n12944 0.00188565
R74391 VSS.n12929 VSS.n12928 0.00188565
R74392 VSS.n12728 VSS.n12727 0.00188565
R74393 VSS.n12712 VSS.n12711 0.00188565
R74394 VSS.n12521 VSS.n12520 0.00188565
R74395 VSS.n12311 VSS.n12310 0.00188565
R74396 VSS.n12281 VSS.n12280 0.00188565
R74397 VSS.n12278 VSS.n12277 0.00188565
R74398 VSS.n11906 VSS.n11905 0.00188565
R74399 VSS.n11846 VSS.n11845 0.00188565
R74400 VSS.n12946 VSS.n12945 0.00188565
R74401 VSS.n12930 VSS.n12929 0.00188565
R74402 VSS.n15031 VSS.n15030 0.00188565
R74403 VSS.n15045 VSS.n15044 0.00188565
R74404 VSS.n16050 VSS.n16049 0.00188565
R74405 VSS.n9679 VSS.n9678 0.00188565
R74406 VSS.n9160 VSS.n9159 0.00188565
R74407 VSS.n9288 VSS.n9287 0.00188565
R74408 VSS.n9275 VSS.n9274 0.00188565
R74409 VSS.n15030 VSS.n15029 0.00188565
R74410 VSS.n15044 VSS.n15043 0.00188565
R74411 VSS.n20639 VSS.n20638 0.00188565
R74412 VSS.n20655 VSS.n20654 0.00188565
R74413 VSS.n6907 VSS.n6906 0.00188565
R74414 VSS.n6972 VSS.n6971 0.00188565
R74415 VSS.n6648 VSS.n6647 0.00188565
R74416 VSS.n6612 VSS.n6611 0.00188565
R74417 VSS.n6596 VSS.n6595 0.00188565
R74418 VSS.n20638 VSS.n20637 0.00188565
R74419 VSS.n20654 VSS.n20653 0.00188565
R74420 VSS.n20110 VSS.n20109 0.00188565
R74421 VSS.n20094 VSS.n20093 0.00188565
R74422 VSS.n1024 VSS.n1023 0.00188565
R74423 VSS.n6870 VSS.n6869 0.00188565
R74424 VSS.n6498 VSS.n6497 0.00188565
R74425 VSS.n6462 VSS.n6461 0.00188565
R74426 VSS.n6446 VSS.n6445 0.00188565
R74427 VSS.n20111 VSS.n20110 0.00188565
R74428 VSS.n20095 VSS.n20094 0.00188565
R74429 VSS.n21650 VSS.n21649 0.00188565
R74430 VSS.n21526 VSS.n21525 0.00188565
R74431 VSS.n21476 VSS.n21475 0.00188565
R74432 VSS.n21362 VSS.n21361 0.00188565
R74433 VSS.n21346 VSS.n21345 0.00188565
R74434 VSS.n7634 VSS.n7633 0.00188565
R74435 VSS.n7651 VSS.n7650 0.00188565
R74436 VSS.n7723 VSS.n7722 0.00188565
R74437 VSS.n7739 VSS.n7738 0.00188565
R74438 VSS.n7816 VSS.n7815 0.00188565
R74439 VSS.n7800 VSS.n7799 0.00188565
R74440 VSS.n21363 VSS.n21362 0.00188565
R74441 VSS.n21347 VSS.n21346 0.00188565
R74442 VSS.n21525 VSS.n21524 0.00188565
R74443 VSS.n21477 VSS.n21476 0.00188565
R74444 VSS.n9289 VSS.n9288 0.00188565
R74445 VSS.n7817 VSS.n7816 0.00188565
R74446 VSS.n9126 VSS.n9125 0.00188565
R74447 VSS.n7801 VSS.n7800 0.00188565
R74448 VSS.n11847 VSS.n11846 0.00188565
R74449 VSS.n6597 VSS.n6596 0.00188565
R74450 VSS.n6447 VSS.n6446 0.00188565
R74451 VSS.n9276 VSS.n9275 0.00188565
R74452 VSS.n9113 VSS.n9112 0.00188565
R74453 VSS.n6613 VSS.n6612 0.00188565
R74454 VSS.n6463 VSS.n6462 0.00188565
R74455 VSS.n9680 VSS.n9679 0.00188565
R74456 VSS.n12522 VSS.n12521 0.00188565
R74457 VSS.n12312 VSS.n12311 0.00188565
R74458 VSS.n7722 VSS.n7721 0.00188565
R74459 VSS.n9563 VSS.n9562 0.00188565
R74460 VSS.n7738 VSS.n7737 0.00188565
R74461 VSS.n12279 VSS.n12278 0.00188565
R74462 VSS.n12280 VSS.n12279 0.00188565
R74463 VSS.n6647 VSS.n6646 0.00188565
R74464 VSS.n6497 VSS.n6496 0.00188565
R74465 VSS.n9159 VSS.n9158 0.00188565
R74466 VSS.n9016 VSS.n9015 0.00188565
R74467 VSS.n6973 VSS.n6972 0.00188565
R74468 VSS.n6871 VSS.n6870 0.00188565
R74469 VSS.n7650 VSS.n7649 0.00188565
R74470 VSS.n12713 VSS.n12712 0.00188565
R74471 VSS.n6906 VSS.n6905 0.00188565
R74472 VSS.n1025 VSS.n1024 0.00188565
R74473 VSS.n16051 VSS.n16050 0.00188565
R74474 VSS.n5541 VSS.n5540 0.00188565
R74475 VSS.n7635 VSS.n7634 0.00188565
R74476 VSS.n12727 VSS.n12726 0.00188565
R74477 VSS.n3879 VSS.n3878 0.00188565
R74478 VSS.n4142 VSS.n4141 0.00188565
R74479 VSS.n4761 VSS.n4760 0.00188565
R74480 VSS.n11678 VSS.n11677 0.00188565
R74481 VSS.n11664 VSS.n11663 0.00188565
R74482 VSS.n6121 VSS.n6120 0.00188565
R74483 VSS.n6108 VSS.n6107 0.00188565
R74484 VSS.n6040 VSS.n6039 0.00188565
R74485 VSS.n6027 VSS.n6026 0.00188565
R74486 VSS.n5959 VSS.n5958 0.00188565
R74487 VSS.n5946 VSS.n5945 0.00188565
R74488 VSS.n11679 VSS.n11678 0.00188565
R74489 VSS.n6122 VSS.n6121 0.00188565
R74490 VSS.n6041 VSS.n6040 0.00188565
R74491 VSS.n5960 VSS.n5959 0.00188565
R74492 VSS.n6028 VSS.n6027 0.00188565
R74493 VSS.n5947 VSS.n5946 0.00188565
R74494 VSS.n6109 VSS.n6108 0.00188565
R74495 VSS.n4760 VSS.n4759 0.00188565
R74496 VSS.n11665 VSS.n11664 0.00188565
R74497 VSS.n4143 VSS.n4142 0.00188565
R74498 VSS.n3878 VSS.n3877 0.00188565
R74499 VSS.n21649 VSS.n21648 0.00188565
R74500 VSS.n635 VSS.n634 0.00188565
R74501 VSS.n622 VSS.n621 0.00188565
R74502 VSS.n10594 VSS.n10593 0.00188565
R74503 VSS.n10580 VSS.n10579 0.00188565
R74504 VSS.n10466 VSS.n10465 0.00188565
R74505 VSS.n10229 VSS.n10228 0.00188565
R74506 VSS.n10227 VSS.n10226 0.00188565
R74507 VSS.n9906 VSS.n9905 0.00188565
R74508 VSS.n9004 VSS.n8999 0.00188565
R74509 VSS.n10467 VSS.n10466 0.00188565
R74510 VSS.n10259 VSS.n10258 0.00188565
R74511 VSS.n9907 VSS.n9906 0.00188565
R74512 VSS.n8999 VSS.n8998 0.00188565
R74513 VSS.n10581 VSS.n10580 0.00188565
R74514 VSS.n636 VSS.n635 0.00188565
R74515 VSS.n623 VSS.n622 0.00188565
R74516 VSS.n10593 VSS.n10592 0.00188565
R74517 VSS.n22254 VSS.n22177 0.00187029
R74518 VSS.n2685 VSS.n2684 0.00186769
R74519 VSS.n2686 VSS.n2685 0.00186769
R74520 VSS.n2691 VSS.n2690 0.00186769
R74521 VSS.n2694 VSS.n2693 0.00186769
R74522 VSS.n17588 VSS.n17587 0.00186769
R74523 VSS.n17540 VSS.n17539 0.00186769
R74524 VSS.n17539 VSS.n17538 0.00186769
R74525 VSS.n17534 VSS.n17533 0.00186769
R74526 VSS.n17533 VSS.n17532 0.00186769
R74527 VSS.n17483 VSS.n2278 0.00186769
R74528 VSS.n18104 VSS.n18103 0.00186769
R74529 VSS.n18100 VSS.n18099 0.00186769
R74530 VSS.n18098 VSS.n18097 0.00186769
R74531 VSS.n17976 VSS.n17975 0.00186769
R74532 VSS.n17967 VSS.n17873 0.00186769
R74533 VSS.n17822 VSS.n17821 0.00186769
R74534 VSS.n17814 VSS.n17813 0.00186769
R74535 VSS.n17535 VSS.n17534 0.00186769
R74536 VSS.n17538 VSS.n17537 0.00186769
R74537 VSS.n17532 VSS.n17531 0.00186769
R74538 VSS.n17541 VSS.n17540 0.00186769
R74539 VSS.n18105 VSS.n18104 0.00186769
R74540 VSS.n18101 VSS.n18100 0.00186769
R74541 VSS.n18105 VSS.n2278 0.00186769
R74542 VSS.n18099 VSS.n18098 0.00186769
R74543 VSS.n17823 VSS.n17822 0.00186769
R74544 VSS.n17815 VSS.n17814 0.00186769
R74545 VSS.n17873 VSS.n17872 0.00186769
R74546 VSS.n17977 VSS.n17976 0.00186769
R74547 VSS.n2692 VSS.n2691 0.00186769
R74548 VSS.n2684 VSS.n2683 0.00186769
R74549 VSS.n2693 VSS.n2692 0.00186769
R74550 VSS.n2687 VSS.n2686 0.00186769
R74551 VSS.n17589 VSS.n17588 0.00186769
R74552 VSS.n2730 VSS.n2729 0.00186769
R74553 VSS.n2732 VSS.n2731 0.00186769
R74554 VSS.n2736 VSS.n2735 0.00186769
R74555 VSS.n2738 VSS.n2737 0.00186769
R74556 VSS.n2790 VSS.n2789 0.00186769
R74557 VSS.n2792 VSS.n2791 0.00186769
R74558 VSS.n2796 VSS.n2795 0.00186769
R74559 VSS.n2798 VSS.n2797 0.00186769
R74560 VSS.n2934 VSS.n2933 0.00186769
R74561 VSS.n2936 VSS.n2935 0.00186769
R74562 VSS.n2990 VSS.n2989 0.00186769
R74563 VSS.n2998 VSS.n2997 0.00186769
R74564 VSS.n3000 VSS.n2999 0.00186769
R74565 VSS.n3038 VSS.n3037 0.00186769
R74566 VSS.n3046 VSS.n3045 0.00186769
R74567 VSS.n3048 VSS.n3047 0.00186769
R74568 VSS.n2729 VSS.n2728 0.00186769
R74569 VSS.n2735 VSS.n2734 0.00186769
R74570 VSS.n3045 VSS.n3044 0.00186769
R74571 VSS.n17584 VSS.n17583 0.00186769
R74572 VSS.n17578 VSS.n17577 0.00186769
R74573 VSS.n17968 VSS.n17967 0.00186769
R74574 VSS.n17812 VSS.n17811 0.00186769
R74575 VSS.n17778 VSS.n17777 0.00186769
R74576 VSS.n17769 VSS.n17768 0.00186769
R74577 VSS.n17767 VSS.n17766 0.00186769
R74578 VSS.n17777 VSS.n17776 0.00186769
R74579 VSS.n17768 VSS.n17767 0.00186769
R74580 VSS.n17770 VSS.n17769 0.00186769
R74581 VSS.n2795 VSS.n2794 0.00186769
R74582 VSS.n2789 VSS.n2788 0.00186769
R74583 VSS.n2997 VSS.n2996 0.00186769
R74584 VSS.n17813 VSS.n17812 0.00186769
R74585 VSS.n17969 VSS.n17968 0.00186769
R74586 VSS.n2933 VSS.n2932 0.00186769
R74587 VSS.n2791 VSS.n2790 0.00186769
R74588 VSS.n2935 VSS.n2934 0.00186769
R74589 VSS.n2797 VSS.n2796 0.00186769
R74590 VSS.n2999 VSS.n2998 0.00186769
R74591 VSS.n2989 VSS.n2988 0.00186769
R74592 VSS.n3047 VSS.n3046 0.00186769
R74593 VSS.n3037 VSS.n3036 0.00186769
R74594 VSS.n2737 VSS.n2736 0.00186769
R74595 VSS.n2731 VSS.n2730 0.00186769
R74596 VSS.n17587 VSS.n17584 0.00186769
R74597 VSS.n17579 VSS.n17578 0.00186769
R74598 VSS.n22177 VSS.n22176 0.0018651
R74599 VSS.n6270 VSS.n6269 0.00186
R74600 VSS.n6295 VSS.n6294 0.00186
R74601 VSS.n11139 VSS.n11138 0.00186
R74602 VSS.n11899 VSS.n11898 0.00185432
R74603 VSS.n14164 VSS.n14163 0.00185
R74604 VSS.n14191 VSS.n14190 0.00185
R74605 VSS.n19408 VSS.n19406 0.00185
R74606 VSS.n18258 VSS.n18257 0.00185
R74607 VSS.n16613 VSS.n16612 0.00185
R74608 VSS.n16516 VSS.n16514 0.00185
R74609 VSS.n2887 VSS.n2885 0.00185
R74610 VSS.n2849 VSS.n2848 0.00185
R74611 VSS.n2892 VSS.n2891 0.00185
R74612 VSS.n5127 VSS.n5126 0.00185
R74613 VSS.n5159 VSS.n5156 0.00185
R74614 VSS.n5162 VSS.n5161 0.00185
R74615 VSS.n7366 VSS.n7365 0.00185
R74616 VSS.n7363 VSS.n7362 0.00185
R74617 VSS.n7312 VSS.n7311 0.00185
R74618 VSS.n7309 VSS.n7308 0.00185
R74619 VSS.n7222 VSS.n7221 0.00185
R74620 VSS.n4528 VSS.n4527 0.00185
R74621 VSS.n4498 VSS.n4497 0.00185
R74622 VSS.n4493 VSS.n4492 0.00185
R74623 VSS.n18048 VSS.n18047 0.00185
R74624 VSS.n18009 VSS.n18008 0.00185
R74625 VSS.n18013 VSS.n18011 0.00185
R74626 VSS.n15698 VSS.n15697 0.00185
R74627 VSS.n7857 DVSS 0.00184667
R74628 VSS.n10321 VSS.n10316 0.00184615
R74629 VSS.n10439 VSS.n10434 0.00184615
R74630 VSS.n10347 VSS.n10342 0.00184615
R74631 VSS.n10154 VSS.n10149 0.00184615
R74632 VSS.n10062 VSS.n10057 0.00184615
R74633 VSS.n10023 VSS.n10022 0.00184615
R74634 VSS.n12375 VSS.n12370 0.00184615
R74635 VSS.n12493 VSS.n12488 0.00184615
R74636 VSS.n12401 VSS.n12396 0.00184615
R74637 VSS.n12205 VSS.n12200 0.00184615
R74638 VSS.n12113 VSS.n12108 0.00184615
R74639 VSS.n12074 VSS.n12073 0.00184615
R74640 VSS.n18805 VSS.n18804 0.00184491
R74641 VSS.n18452 VSS.n18451 0.00184491
R74642 VSS.n16589 VSS.n16588 0.00184491
R74643 VSS.n15536 VSS.n15535 0.00184491
R74644 VSS.n8514 VSS.n8513 0.00184491
R74645 VSS.n18453 VSS.n18452 0.00184491
R74646 VSS.n14890 VSS.n14889 0.00184491
R74647 VSS.n16638 VSS.n16637 0.00184491
R74648 VSS.n16590 VSS.n16589 0.00184491
R74649 VSS.n15537 VSS.n15536 0.00184491
R74650 VSS.n8513 VSS.n8512 0.00184491
R74651 VSS.n19587 VSS.n19586 0.00184491
R74652 VSS.n19961 VSS.n19960 0.00184491
R74653 VSS.n760 VSS.n759 0.00184491
R74654 VSS.n779 VSS.n778 0.00184491
R74655 VSS.n1824 VSS.n1823 0.00184491
R74656 VSS.n8665 VSS.n8664 0.00184491
R74657 VSS.n8664 VSS.n8663 0.00184491
R74658 VSS.n19586 VSS.n19585 0.00184491
R74659 VSS.n778 VSS.n777 0.00184491
R74660 VSS.n19477 VSS.n19476 0.00184491
R74661 VSS.n1825 VSS.n1824 0.00184491
R74662 VSS.n3446 VSS.n3445 0.00183803
R74663 VSS.n3461 VSS.n3460 0.00183803
R74664 VSS.n3465 VSS.n3464 0.00183803
R74665 VSS.n3674 VSS.n3673 0.00183803
R74666 VSS.n3671 VSS.n3670 0.00183803
R74667 VSS.n3008 VSS.n3007 0.00183556
R74668 VSS.n3056 VSS.n3055 0.00183556
R74669 VSS.n3057 VSS.n3056 0.00183556
R74670 VSS.n3009 VSS.n3008 0.00183556
R74671 VSS.n9780 VSS.n9779 0.00182
R74672 VSS.n9726 VSS.n9725 0.00182
R74673 VSS.n10681 VSS.n10680 0.00182
R74674 VSS.n10743 VSS.n10742 0.00182
R74675 DVSS VSS.n11079 0.00180667
R74676 VSS.n4072 VSS.n4071 0.0017971
R74677 VSS.n11529 VSS.n11528 0.0017971
R74678 VSS.n5594 VSS.n5593 0.0017971
R74679 VSS.n9590 VSS.n9589 0.0017971
R74680 VSS.n9153 VSS.n9152 0.0017971
R74681 VSS.n11528 VSS.n11527 0.0017971
R74682 VSS.n4071 VSS.n4070 0.0017971
R74683 VSS.n13099 VSS.n13098 0.0017971
R74684 VSS.n12975 VSS.n12974 0.0017971
R74685 VSS.n12757 VSS.n12756 0.0017971
R74686 VSS.n12556 VSS.n12555 0.0017971
R74687 VSS.n12243 VSS.n12242 0.0017971
R74688 VSS.n11939 VSS.n11938 0.0017971
R74689 VSS.n12976 VSS.n12975 0.0017971
R74690 VSS.n13098 VSS.n13097 0.0017971
R74691 VSS.n18943 VSS.n18942 0.0017971
R74692 VSS.n15003 VSS.n15002 0.0017971
R74693 VSS.n16110 VSS.n16109 0.0017971
R74694 VSS.n9707 VSS.n9706 0.0017971
R74695 VSS.n9316 VSS.n9315 0.0017971
R74696 VSS.n15002 VSS.n15001 0.0017971
R74697 VSS.n18942 VSS.n18941 0.0017971
R74698 VSS.n21872 VSS.n21871 0.0017971
R74699 VSS.n20609 VSS.n20608 0.0017971
R74700 VSS.n21044 VSS.n21043 0.0017971
R74701 VSS.n7002 VSS.n7001 0.0017971
R74702 VSS.n6642 VSS.n6641 0.0017971
R74703 VSS.n20608 VSS.n20607 0.0017971
R74704 VSS.n21871 VSS.n21870 0.0017971
R74705 VSS.n19157 VSS.n19156 0.0017971
R74706 VSS.n20140 VSS.n20139 0.0017971
R74707 VSS.n1090 VSS.n1089 0.0017971
R74708 VSS.n6900 VSS.n6899 0.0017971
R74709 VSS.n6492 VSS.n6491 0.0017971
R74710 VSS.n20141 VSS.n20140 0.0017971
R74711 VSS.n19156 VSS.n19155 0.0017971
R74712 VSS.n21462 VSS.n21461 0.0017971
R74713 VSS.n21392 VSS.n21391 0.0017971
R74714 VSS.n7605 VSS.n7604 0.0017971
R74715 VSS.n7693 VSS.n7692 0.0017971
R74716 VSS.n7846 VSS.n7845 0.0017971
R74717 VSS.n21393 VSS.n21392 0.0017971
R74718 VSS.n21463 VSS.n21462 0.0017971
R74719 VSS.n9317 VSS.n9316 0.0017971
R74720 VSS.n7847 VSS.n7846 0.0017971
R74721 VSS.n9154 VSS.n9153 0.0017971
R74722 VSS.n6643 VSS.n6642 0.0017971
R74723 VSS.n6493 VSS.n6492 0.0017971
R74724 VSS.n9708 VSS.n9707 0.0017971
R74725 VSS.n12557 VSS.n12556 0.0017971
R74726 VSS.n12242 VSS.n12241 0.0017971
R74727 VSS.n7692 VSS.n7691 0.0017971
R74728 VSS.n9591 VSS.n9590 0.0017971
R74729 VSS.n6901 VSS.n6900 0.0017971
R74730 VSS.n7003 VSS.n7002 0.0017971
R74731 VSS.n7604 VSS.n7603 0.0017971
R74732 VSS.n12758 VSS.n12757 0.0017971
R74733 VSS.n16111 VSS.n16110 0.0017971
R74734 VSS.n5595 VSS.n5594 0.0017971
R74735 VSS.n21045 VSS.n21044 0.0017971
R74736 VSS.n1091 VSS.n1090 0.0017971
R74737 VSS.n4773 VSS.n4772 0.0017971
R74738 VSS.n11706 VSS.n11705 0.0017971
R74739 VSS.n6149 VSS.n6148 0.0017971
R74740 VSS.n6068 VSS.n6067 0.0017971
R74741 VSS.n5987 VSS.n5986 0.0017971
R74742 VSS.n11707 VSS.n11706 0.0017971
R74743 VSS.n6150 VSS.n6149 0.0017971
R74744 VSS.n6069 VSS.n6068 0.0017971
R74745 VSS.n5988 VSS.n5987 0.0017971
R74746 VSS.n4772 VSS.n4771 0.0017971
R74747 VSS.n2616 VSS.n2615 0.0017971
R74748 VSS.n2617 VSS.n2616 0.0017971
R74749 VSS.n663 VSS.n662 0.0017971
R74750 VSS.n10621 VSS.n10620 0.0017971
R74751 VSS.n10192 VSS.n10191 0.0017971
R74752 VSS.n9940 VSS.n9939 0.0017971
R74753 VSS.n10501 VSS.n10500 0.0017971
R74754 VSS.n9941 VSS.n9940 0.0017971
R74755 VSS.n10191 VSS.n10190 0.0017971
R74756 VSS.n10622 VSS.n10621 0.0017971
R74757 VSS.n664 VSS.n663 0.0017971
R74758 VSS.n6767 VSS.n6766 0.00179
R74759 VSS.n6707 VSS.n6706 0.00179
R74760 VSS.n8083 VSS.n8082 0.00179
R74761 VSS.n8023 VSS.n8022 0.00179
R74762 VSS.n10930 VSS.n10929 0.00179
R74763 VSS.n10997 VSS.n10996 0.00179
R74764 VSS.n2577 VSS.n2576 0.00178571
R74765 VSS.n7267 VSS.n7266 0.00178571
R74766 VSS.n7248 VSS.n7247 0.00178571
R74767 VSS.n7235 VSS.n7234 0.00178571
R74768 VSS.n7216 VSS.n7215 0.00178571
R74769 VSS.n4683 VSS.n4682 0.00178571
R74770 VSS.n17601 VSS.n17600 0.00178571
R74771 VSS.n3536 VSS.n3535 0.00176761
R74772 VSS.n3595 VSS.n3594 0.00176761
R74773 VSS.n3638 VSS.n3637 0.00176761
R74774 VSS.n3202 VSS.n3201 0.00176761
R74775 VSS.n3442 VSS.n3441 0.00176761
R74776 VSS.n3452 VSS.n3448 0.00176761
R74777 VSS.n3538 VSS.n3537 0.00176761
R74778 VSS.n3597 VSS.n3596 0.00176761
R74779 VSS.n3640 VSS.n3639 0.00176761
R74780 VSS.n3656 VSS.n3655 0.00176761
R74781 VSS.n18692 VSS.n18691 0.00176761
R74782 VSS.n18411 VSS.n18410 0.00176761
R74783 VSS.n18192 VSS.n18191 0.00176761
R74784 VSS.n17130 VSS.n17129 0.00176761
R74785 VSS.n17119 VSS.n17118 0.00176761
R74786 VSS.n16921 VSS.n16920 0.00176761
R74787 VSS.n16581 VSS.n16580 0.00176761
R74788 VSS.n16526 VSS.n16525 0.00176761
R74789 VSS.n14986 VSS.n14985 0.00176761
R74790 VSS.n15532 VSS.n15531 0.00176761
R74791 VSS.n15469 VSS.n15468 0.00176761
R74792 VSS.n15459 VSS.n15458 0.00176761
R74793 VSS.n15334 VSS.n15333 0.00176761
R74794 VSS.n19174 VSS.n19173 0.00176761
R74795 VSS.n19611 VSS.n19610 0.00176761
R74796 VSS.n19664 VSS.n19663 0.00176761
R74797 VSS.n19865 VSS.n19864 0.00176761
R74798 VSS.n19876 VSS.n19875 0.00176761
R74799 VSS.n19995 VSS.n19994 0.00176761
R74800 VSS.n787 VSS.n786 0.00176761
R74801 VSS.n812 VSS.n811 0.00176761
R74802 VSS.n822 VSS.n821 0.00176761
R74803 VSS.n1820 VSS.n1819 0.00176761
R74804 VSS.n1771 VSS.n1770 0.00176761
R74805 VSS.n1761 VSS.n1760 0.00176761
R74806 VSS.n1650 VSS.n1649 0.00176761
R74807 VSS.n8086 VSS.n8085 0.00176
R74808 VSS.n8026 VSS.n8025 0.00176
R74809 VSS.n10925 VSS.n10924 0.00176
R74810 VSS.n10992 VSS.n10991 0.00176
R74811 VSS.n6205 VSS.n6204 0.00175333
R74812 VSS.n6245 VSS.n6244 0.00175333
R74813 VSS.n11164 VSS.n11163 0.00175333
R74814 VSS.n4003 VSS.n4002 0.00174016
R74815 VSS.n4035 VSS.n4034 0.00174016
R74816 VSS.n3954 VSS.n3953 0.00174016
R74817 VSS.n2364 VSS.n2363 0.00174016
R74818 VSS.n17322 VSS.n17321 0.00174016
R74819 VSS.n11333 VSS.n11332 0.00174016
R74820 VSS.n5864 VSS.n5863 0.00174016
R74821 VSS.n5741 VSS.n5740 0.00174016
R74822 VSS.n5630 VSS.n5629 0.00174016
R74823 VSS.n5568 VSS.n5567 0.00174016
R74824 VSS.n9540 VSS.n9539 0.00174016
R74825 VSS.n9042 VSS.n9041 0.00174016
R74826 VSS.n13028 VSS.n13027 0.00174016
R74827 VSS.n13064 VSS.n13063 0.00174016
R74828 VSS.n13126 VSS.n13125 0.00174016
R74829 VSS.n13174 VSS.n13173 0.00174016
R74830 VSS.n12990 VSS.n12989 0.00174016
R74831 VSS.n12878 VSS.n12877 0.00174016
R74832 VSS.n12815 VSS.n12814 0.00174016
R74833 VSS.n12772 VSS.n12771 0.00174016
R74834 VSS.n12692 VSS.n12691 0.00174016
R74835 VSS.n12690 VSS.n12689 0.00174016
R74836 VSS.n12676 VSS.n12675 0.00174016
R74837 VSS.n12510 VSS.n12509 0.00174016
R74838 VSS.n12325 VSS.n12324 0.00174016
R74839 VSS.n12323 VSS.n12322 0.00174016
R74840 VSS.n12285 VSS.n12284 0.00174016
R74841 VSS.n12233 VSS.n12232 0.00174016
R74842 VSS.n11942 VSS.n11941 0.00174016
R74843 VSS.n11938 VSS.n11937 0.00174016
R74844 VSS.n11909 VSS.n11908 0.00174016
R74845 VSS.n11905 VSS.n11904 0.00174016
R74846 VSS.n11890 VSS.n11889 0.00174016
R74847 VSS.n11856 VSS.n11855 0.00174016
R74848 VSS.n11835 VSS.n11834 0.00174016
R74849 VSS.n18874 VSS.n18873 0.00174016
R74850 VSS.n18906 VSS.n18905 0.00174016
R74851 VSS.n18971 VSS.n18970 0.00174016
R74852 VSS.n2263 VSS.n2262 0.00174016
R74853 VSS.n14414 VSS.n14413 0.00174016
R74854 VSS.n15134 VSS.n15133 0.00174016
R74855 VSS.n16225 VSS.n16224 0.00174016
R74856 VSS.n16189 VSS.n16188 0.00174016
R74857 VSS.n16152 VSS.n16151 0.00174016
R74858 VSS.n16084 VSS.n16083 0.00174016
R74859 VSS.n9657 VSS.n9656 0.00174016
R74860 VSS.n9185 VSS.n9184 0.00174016
R74861 VSS.n21801 VSS.n21800 0.00174016
R74862 VSS.n21837 VSS.n21836 0.00174016
R74863 VSS.n21752 VSS.n21751 0.00174016
R74864 VSS.n2314 VSS.n2313 0.00174016
R74865 VSS.n20594 VSS.n20593 0.00174016
R74866 VSS.n20782 VSS.n20781 0.00174016
R74867 VSS.n21169 VSS.n21168 0.00174016
R74868 VSS.n21131 VSS.n21130 0.00174016
R74869 VSS.n21080 VSS.n21079 0.00174016
R74870 VSS.n21017 VSS.n21016 0.00174016
R74871 VSS.n6675 VSS.n6674 0.00174016
R74872 VSS.n19086 VSS.n19085 0.00174016
R74873 VSS.n19122 VSS.n19121 0.00174016
R74874 VSS.n19037 VSS.n19036 0.00174016
R74875 VSS.n17922 VSS.n17921 0.00174016
R74876 VSS.n20156 VSS.n20155 0.00174016
R74877 VSS.n2037 VSS.n2036 0.00174016
R74878 VSS.n1298 VSS.n1297 0.00174016
R74879 VSS.n1181 VSS.n1180 0.00174016
R74880 VSS.n1132 VSS.n1131 0.00174016
R74881 VSS.n1063 VSS.n1062 0.00174016
R74882 VSS.n6525 VSS.n6524 0.00174016
R74883 VSS.n21572 VSS.n21571 0.00174016
R74884 VSS.n21608 VSS.n21607 0.00174016
R74885 VSS.n21666 VSS.n21665 0.00174016
R74886 VSS.n21499 VSS.n21498 0.00174016
R74887 VSS.n21407 VSS.n21406 0.00174016
R74888 VSS.n21299 VSS.n21298 0.00174016
R74889 VSS.n7547 VSS.n7546 0.00174016
R74890 VSS.n7590 VSS.n7589 0.00174016
R74891 VSS.n7678 VSS.n7677 0.00174016
R74892 VSS.n7766 VSS.n7765 0.00174016
R74893 VSS.n3790 VSS.n3789 0.00174016
R74894 VSS.n3805 VSS.n3804 0.00174016
R74895 VSS.n3837 VSS.n3836 0.00174016
R74896 VSS.n4127 VSS.n4126 0.00174016
R74897 VSS.n4717 VSS.n4716 0.00174016
R74898 VSS.n11732 VSS.n11731 0.00174016
R74899 VSS.n11455 VSS.n11454 0.00174016
R74900 VSS.n11234 VSS.n11233 0.00174016
R74901 VSS.n11195 VSS.n11194 0.00174016
R74902 VSS.n6083 VSS.n6082 0.00174016
R74903 VSS.n6002 VSS.n6001 0.00174016
R74904 VSS.n3283 VSS.n3282 0.00174016
R74905 VSS.n2652 VSS.n2651 0.00174016
R74906 VSS.n670 VSS.n669 0.00174016
R74907 VSS.n573 VSS.n572 0.00174016
R74908 VSS.n514 VSS.n513 0.00174016
R74909 VSS.n475 VSS.n474 0.00174016
R74910 VSS.n10560 VSS.n10559 0.00174016
R74911 VSS.n10558 VSS.n10557 0.00174016
R74912 VSS.n10544 VSS.n10543 0.00174016
R74913 VSS.n10456 VSS.n10455 0.00174016
R74914 VSS.n10271 VSS.n10270 0.00174016
R74915 VSS.n10269 VSS.n10268 0.00174016
R74916 VSS.n10233 VSS.n10232 0.00174016
R74917 VSS.n10181 VSS.n10180 0.00174016
R74918 VSS.n9944 VSS.n9943 0.00174016
R74919 VSS.n9939 VSS.n9938 0.00174016
R74920 VSS.n9910 VSS.n9909 0.00174016
R74921 VSS.n9905 VSS.n9904 0.00174016
R74922 VSS.n8981 VSS.n8980 0.00174016
R74923 VSS.n8794 VSS.n8793 0.00174016
R74924 VSS.n8908 VSS.n8907 0.00174016
R74925 VSS.n18714 VSS.n18713 0.00173932
R74926 VSS.n18398 VSS.n18397 0.00173932
R74927 VSS.n18183 VSS.n18182 0.00173932
R74928 VSS.n14856 VSS.n14834 0.00173932
R74929 VSS.n18713 VSS.n18712 0.00173932
R74930 VSS.n19196 VSS.n19195 0.00173932
R74931 VSS.n19624 VSS.n19623 0.00173932
R74932 VSS.n19927 VSS.n19926 0.00173932
R74933 VSS.n19673 VSS.n19672 0.00173932
R74934 VSS.n19195 VSS.n19194 0.00173932
R74935 VSS.n7953 DVSS 0.00173
R74936 DVSS VSS.n7944 0.00173
R74937 VSS.n14208 VSS.n13943 0.00172143
R74938 VSS.n3081 VSS.n3080 0.00172143
R74939 VSS.n4344 VSS.n4343 0.00172143
R74940 VSS.n4341 VSS.n4340 0.00172143
R74941 VSS.n17736 VSS.n17735 0.00172143
R74942 VSS.n17733 VSS.n17732 0.00172143
R74943 VSS.n14131 VSS.n14130 0.00172143
R74944 VSS.n4207 VSS.n4206 0.00170855
R74945 VSS.n11344 VSS.n11343 0.00170855
R74946 VSS.n5852 VSS.n5851 0.00170855
R74947 VSS.n4206 VSS.n4205 0.00170855
R74948 VSS.n11345 VSS.n11344 0.00170855
R74949 VSS.n5853 VSS.n5852 0.00170855
R74950 VSS.n3996 VSS.n3995 0.00170855
R74951 VSS.n2376 VSS.n2375 0.00170855
R74952 VSS.n9538 VSS.n9537 0.00170855
R74953 VSS.n3995 VSS.n3994 0.00170855
R74954 VSS.n13146 VSS.n13145 0.00170855
R74955 VSS.n13188 VSS.n13187 0.00170855
R74956 VSS.n12864 VSS.n12863 0.00170855
R74957 VSS.n12801 VSS.n12800 0.00170855
R74958 VSS.n12251 VSS.n12250 0.00170855
R74959 VSS.n11851 VSS.n11850 0.00170855
R74960 VSS.n13145 VSS.n13144 0.00170855
R74961 VSS.n12865 VSS.n12864 0.00170855
R74962 VSS.n13021 VSS.n13020 0.00170855
R74963 VSS.n12802 VSS.n12801 0.00170855
R74964 VSS.n13187 VSS.n13186 0.00170855
R74965 VSS.n2375 VSS.n2374 0.00170855
R74966 VSS.n18867 VSS.n18866 0.00170855
R74967 VSS.n2237 VSS.n2236 0.00170855
R74968 VSS.n2275 VSS.n2274 0.00170855
R74969 VSS.n15146 VSS.n15145 0.00170855
R74970 VSS.n16213 VSS.n16212 0.00170855
R74971 VSS.n9655 VSS.n9654 0.00170855
R74972 VSS.n2236 VSS.n2235 0.00170855
R74973 VSS.n15145 VSS.n15144 0.00170855
R74974 VSS.n2274 VSS.n2273 0.00170855
R74975 VSS.n18866 VSS.n18865 0.00170855
R74976 VSS.n16214 VSS.n16213 0.00170855
R74977 VSS.n2286 VSS.n2285 0.00170855
R74978 VSS.n2328 VSS.n2327 0.00170855
R74979 VSS.n20796 VSS.n20795 0.00170855
R74980 VSS.n21155 VSS.n21154 0.00170855
R74981 VSS.n6944 VSS.n6943 0.00170855
R74982 VSS.n2285 VSS.n2284 0.00170855
R74983 VSS.n20795 VSS.n20794 0.00170855
R74984 VSS.n2327 VSS.n2326 0.00170855
R74985 VSS.n21794 VSS.n21793 0.00170855
R74986 VSS.n21156 VSS.n21155 0.00170855
R74987 VSS.n17894 VSS.n17893 0.00170855
R74988 VSS.n17936 VSS.n17935 0.00170855
R74989 VSS.n2023 VSS.n2022 0.00170855
R74990 VSS.n1284 VSS.n1283 0.00170855
R74991 VSS.n6842 VSS.n6841 0.00170855
R74992 VSS.n17893 VSS.n17892 0.00170855
R74993 VSS.n2024 VSS.n2023 0.00170855
R74994 VSS.n17935 VSS.n17934 0.00170855
R74995 VSS.n19079 VSS.n19078 0.00170855
R74996 VSS.n1285 VSS.n1284 0.00170855
R74997 VSS.n21565 VSS.n21564 0.00170855
R74998 VSS.n21531 VSS.n21530 0.00170855
R74999 VSS.n21485 VSS.n21484 0.00170855
R75000 VSS.n21469 VSS.n21468 0.00170855
R75001 VSS.n21437 VSS.n21436 0.00170855
R75002 VSS.n21285 VSS.n21284 0.00170855
R75003 VSS.n7561 VSS.n7560 0.00170855
R75004 VSS.n21286 VSS.n21285 0.00170855
R75005 VSS.n21468 VSS.n21467 0.00170855
R75006 VSS.n21486 VSS.n21485 0.00170855
R75007 VSS.n21530 VSS.n21529 0.00170855
R75008 VSS.n21438 VSS.n21437 0.00170855
R75009 VSS.n7560 VSS.n7559 0.00170855
R75010 VSS.n9537 VSS.n9536 0.00170855
R75011 VSS.n9654 VSS.n9653 0.00170855
R75012 VSS.n12252 VSS.n12251 0.00170855
R75013 VSS.n6943 VSS.n6942 0.00170855
R75014 VSS.n6841 VSS.n6840 0.00170855
R75015 VSS.n3798 VSS.n3797 0.00170855
R75016 VSS.n4147 VSS.n4146 0.00170855
R75017 VSS.n4729 VSS.n4728 0.00170855
R75018 VSS.n4768 VSS.n4767 0.00170855
R75019 VSS.n17393 VSS.n17392 0.00170855
R75020 VSS.n11443 VSS.n11442 0.00170855
R75021 VSS.n11222 VSS.n11221 0.00170855
R75022 VSS.n4767 VSS.n4766 0.00170855
R75023 VSS.n11444 VSS.n11443 0.00170855
R75024 VSS.n3797 VSS.n3796 0.00170855
R75025 VSS.n4728 VSS.n4727 0.00170855
R75026 VSS.n11223 VSS.n11222 0.00170855
R75027 VSS.n17393 VSS.n4796 0.00170855
R75028 VSS.n3276 VSS.n3275 0.00170855
R75029 VSS.n3275 VSS.n3274 0.00170855
R75030 VSS.n561 VSS.n560 0.00170855
R75031 VSS.n502 VSS.n501 0.00170855
R75032 VSS.n10200 VSS.n10199 0.00170855
R75033 VSS.n8973 VSS.n8972 0.00170855
R75034 VSS.n8973 VSS.n8970 0.00170855
R75035 VSS.n562 VSS.n561 0.00170855
R75036 VSS.n503 VSS.n502 0.00170855
R75037 VSS.n10788 VSS.n10787 0.0017
R75038 VSS.n10782 VSS.n10772 0.0017
R75039 VSS.n10771 VSS.n10761 0.0017
R75040 VSS.n9386 VSS.n9385 0.0017
R75041 VSS.n9332 VSS.n9331 0.0017
R75042 VSS.n8453 VSS.n8101 0.0017
R75043 VSS.n8785 VSS.n8454 0.0017
R75044 VSS.n10687 VSS.n10685 0.0017
R75045 VSS.n10749 VSS.n10747 0.0017
R75046 VSS.n10790 VSS.n10789 0.0017
R75047 VSS.n3655 VSS.n3654 0.00169718
R75048 VSS.n13941 VSS.n13613 0.00165714
R75049 VSS.n13943 VSS.n13942 0.00165714
R75050 VSS.n2950 VSS.n2949 0.00165714
R75051 VSS.n3014 VSS.n3013 0.00165714
R75052 VSS.n3062 VSS.n3061 0.00165714
R75053 VSS.n2548 VSS.n2547 0.00165714
R75054 VSS.n2859 VSS.n2855 0.00165714
R75055 VSS.n2560 VSS.n2559 0.00165714
R75056 VSS.n5209 VSS.n5208 0.00165714
R75057 VSS.n5260 VSS.n5259 0.00165714
R75058 VSS.n5295 VSS.n5294 0.00165714
R75059 VSS.n4950 VSS.n4949 0.00165714
R75060 VSS.n5135 VSS.n5131 0.00165714
R75061 VSS.n5211 VSS.n5210 0.00165714
R75062 VSS.n5262 VSS.n5261 0.00165714
R75063 VSS.n5297 VSS.n5296 0.00165714
R75064 VSS.n4958 VSS.n4957 0.00165714
R75065 VSS.n7162 VSS.n7161 0.00165714
R75066 VSS.n7103 VSS.n7102 0.00165714
R75067 VSS.n7066 VSS.n7065 0.00165714
R75068 VSS.n7528 VSS.n7527 0.00165714
R75069 VSS.n7163 VSS.n7159 0.00165714
R75070 VSS.n7104 VSS.n7100 0.00165714
R75071 VSS.n7067 VSS.n7062 0.00165714
R75072 VSS.n7529 VSS.n7524 0.00165714
R75073 VSS.n4446 VSS.n4445 0.00165714
R75074 VSS.n4395 VSS.n4394 0.00165714
R75075 VSS.n4360 VSS.n4359 0.00165714
R75076 VSS.n4314 VSS.n4313 0.00165714
R75077 VSS.n4523 VSS.n4522 0.00165714
R75078 VSS.n4447 VSS.n4443 0.00165714
R75079 VSS.n4396 VSS.n4392 0.00165714
R75080 VSS.n4361 VSS.n4357 0.00165714
R75081 VSS.n4326 VSS.n4325 0.00165714
R75082 VSS.n18042 VSS.n18041 0.00165714
R75083 VSS.n17718 VSS.n17717 0.00165714
R75084 VSS.n17860 VSS.n17859 0.00165714
R75085 VSS.n17799 VSS.n17798 0.00165714
R75086 VSS.n17754 VSS.n17753 0.00165714
R75087 VSS.n17704 VSS.n17703 0.00165714
R75088 VSS.n14130 VSS.n14129 0.00165714
R75089 VSS.n14128 VSS.n13947 0.00165714
R75090 VSS.n18705 VSS.n18704 0.00163371
R75091 VSS.n15673 VSS.n15672 0.00163371
R75092 VSS.n18704 VSS.n18703 0.00163371
R75093 VSS.n19187 VSS.n19186 0.00163371
R75094 VSS.n1931 VSS.n1930 0.00163371
R75095 VSS.n1930 VSS.n1929 0.00163371
R75096 VSS.n19186 VSS.n19185 0.00163371
R75097 VSS.n15672 VSS.n15671 0.00163371
R75098 VSS.n3470 VSS.n3469 0.00162676
R75099 VSS.n3188 VSS.n3187 0.00162676
R75100 VSS.n3303 VSS.n3302 0.00162676
R75101 VSS.n3341 VSS.n3340 0.00162676
R75102 VSS.n3395 VSS.n3394 0.00162676
R75103 VSS.n3472 VSS.n3471 0.00162676
R75104 VSS.n3473 VSS.n3472 0.00162676
R75105 VSS.n3662 VSS.n3661 0.00162676
R75106 VSS.n3659 VSS.n3658 0.00162676
R75107 VSS.n17149 VSS.n17148 0.001625
R75108 VSS.n17003 VSS.n17002 0.001625
R75109 VSS.n16993 VSS.n16992 0.001625
R75110 VSS.n4001 VSS.n4000 0.00161999
R75111 VSS.n4000 VSS.n3999 0.00161999
R75112 VSS.n13026 VSS.n13025 0.00161999
R75113 VSS.n12681 VSS.n12680 0.00161999
R75114 VSS.n12289 VSS.n12288 0.00161999
R75115 VSS.n11840 VSS.n11839 0.00161999
R75116 VSS.n13025 VSS.n13024 0.00161999
R75117 VSS.n18872 VSS.n18871 0.00161999
R75118 VSS.n18871 VSS.n18870 0.00161999
R75119 VSS.n21799 VSS.n21798 0.00161999
R75120 VSS.n21798 VSS.n21797 0.00161999
R75121 VSS.n19084 VSS.n19083 0.00161999
R75122 VSS.n19083 VSS.n19082 0.00161999
R75123 VSS.n21557 VSS.n21556 0.00161999
R75124 VSS.n21570 VSS.n21569 0.00161999
R75125 VSS.n21628 VSS.n21627 0.00161999
R75126 VSS.n21442 VSS.n21441 0.00161999
R75127 VSS.n21443 VSS.n21442 0.00161999
R75128 VSS.n21569 VSS.n21568 0.00161999
R75129 VSS.n21627 VSS.n21626 0.00161999
R75130 VSS.n21558 VSS.n21557 0.00161999
R75131 VSS.n11839 VSS.n11838 0.00161999
R75132 VSS.n12290 VSS.n12289 0.00161999
R75133 VSS.n3803 VSS.n3802 0.00161999
R75134 VSS.n3856 VSS.n3855 0.00161999
R75135 VSS.n4793 VSS.n4792 0.00161999
R75136 VSS.n4792 VSS.n4791 0.00161999
R75137 VSS.n3802 VSS.n3801 0.00161999
R75138 VSS.n3855 VSS.n3854 0.00161999
R75139 VSS.n3281 VSS.n3280 0.00161999
R75140 VSS.n3280 VSS.n3279 0.00161999
R75141 VSS.n10549 VSS.n10548 0.00161999
R75142 VSS.n10237 VSS.n10236 0.00161999
R75143 VSS.n8912 VSS.n8911 0.00161999
R75144 VSS.n10238 VSS.n10237 0.00161999
R75145 VSS.n10548 VSS.n10547 0.00161999
R75146 VSS.n12680 VSS.n12679 0.00161999
R75147 VSS.n2511 VSS.n2510 0.00161111
R75148 VSS.n21698 VSS.n21697 0.00161111
R75149 VSS.n2425 VSS.n2424 0.00161111
R75150 VSS.n365 VSS.n364 0.00161111
R75151 VSS.n3937 VSS.n3936 0.00161111
R75152 VSS.n21918 VSS.n21917 0.00161111
R75153 VSS.n2834 VSS.n2833 0.00159286
R75154 VSS.n3018 VSS.n3017 0.00159286
R75155 VSS.n2559 VSS.n2558 0.00159286
R75156 VSS.n5212 VSS.n5211 0.00159286
R75157 VSS.n5263 VSS.n5262 0.00159286
R75158 VSS.n5298 VSS.n5297 0.00159286
R75159 VSS.n4957 VSS.n4956 0.00159286
R75160 VSS.n7062 VSS.n7061 0.00159286
R75161 VSS.n7524 VSS.n7523 0.00159286
R75162 VSS.n4443 VSS.n4442 0.00159286
R75163 VSS.n4392 VSS.n4391 0.00159286
R75164 VSS.n4357 VSS.n4356 0.00159286
R75165 VSS.n4325 VSS.n4324 0.00159286
R75166 VSS.n18066 VSS.n18062 0.00159286
R75167 VSS.n17856 VSS.n17855 0.00159286
R75168 VSS.n17795 VSS.n17794 0.00159286
R75169 VSS.n17750 VSS.n17749 0.00159286
R75170 VSS.n17717 VSS.n17716 0.00159286
R75171 VSS.n3981 VSS.n3980 0.00156299
R75172 VSS.n2353 VSS.n2352 0.00156299
R75173 VSS.n17455 VSS.n17454 0.00156299
R75174 VSS.n11359 VSS.n11358 0.00156299
R75175 VSS.n5848 VSS.n5847 0.00156299
R75176 VSS.n5734 VSS.n5733 0.00156299
R75177 VSS.n5561 VSS.n5560 0.00156299
R75178 VSS.n13005 VSS.n13004 0.00156299
R75179 VSS.n13161 VSS.n13160 0.00156299
R75180 VSS.n12850 VSS.n12849 0.00156299
R75181 VSS.n12787 VSS.n12786 0.00156299
R75182 VSS.n12558 VSS.n12557 0.00156299
R75183 VSS.n12215 VSS.n11972 0.00156299
R75184 VSS.n11878 VSS.n11877 0.00156299
R75185 VSS.n11816 VSS.n11815 0.00156299
R75186 VSS.n11814 VSS.n11813 0.00156299
R75187 VSS.n11806 VSS.n11805 0.00156299
R75188 VSS.n18852 VSS.n18851 0.00156299
R75189 VSS.n2252 VSS.n2251 0.00156299
R75190 VSS.n2206 VSS.n2205 0.00156299
R75191 VSS.n15160 VSS.n15159 0.00156299
R75192 VSS.n16209 VSS.n16208 0.00156299
R75193 VSS.n16182 VSS.n16181 0.00156299
R75194 VSS.n16071 VSS.n16070 0.00156299
R75195 VSS.n21778 VSS.n21777 0.00156299
R75196 VSS.n2301 VSS.n2300 0.00156299
R75197 VSS.n20810 VSS.n20809 0.00156299
R75198 VSS.n21151 VSS.n21150 0.00156299
R75199 VSS.n21124 VSS.n21123 0.00156299
R75200 VSS.n21010 VSS.n21009 0.00156299
R75201 VSS.n19063 VSS.n19062 0.00156299
R75202 VSS.n17909 VSS.n17908 0.00156299
R75203 VSS.n2009 VSS.n2008 0.00156299
R75204 VSS.n1280 VSS.n1279 0.00156299
R75205 VSS.n1174 VSS.n1173 0.00156299
R75206 VSS.n1056 VSS.n1055 0.00156299
R75207 VSS.n21546 VSS.n21545 0.00156299
R75208 VSS.n21559 VSS.n21558 0.00156299
R75209 VSS.n21665 VSS.n21664 0.00156299
R75210 VSS.n21512 VSS.n21511 0.00156299
R75211 VSS.n21452 VSS.n21451 0.00156299
R75212 VSS.n21271 VSS.n21270 0.00156299
R75213 VSS.n7575 VSS.n7574 0.00156299
R75214 VSS.n3781 VSS.n3780 0.00156299
R75215 VSS.n3791 VSS.n3790 0.00156299
R75216 VSS.n4126 VSS.n4125 0.00156299
R75217 VSS.n4706 VSS.n4705 0.00156299
R75218 VSS.n4783 VSS.n4782 0.00156299
R75219 VSS.n11429 VSS.n11428 0.00156299
R75220 VSS.n11208 VSS.n11207 0.00156299
R75221 VSS.n3261 VSS.n3260 0.00156299
R75222 VSS.n547 VSS.n546 0.00156299
R75223 VSS.n488 VSS.n487 0.00156299
R75224 VSS.n10502 VSS.n10501 0.00156299
R75225 VSS.n10164 VSS.n9975 0.00156299
R75226 VSS.n8940 VSS.n8939 0.00156299
R75227 VSS.n8833 VSS.n8832 0.00156299
R75228 VSS.n8839 VSS.n8838 0.00156299
R75229 VSS.n8966 VSS.n8965 0.00156299
R75230 VSS.n3192 VSS.n3189 0.00155634
R75231 VSS.n3193 VSS.n3188 0.00155634
R75232 VSS.n3196 VSS.n3195 0.00155634
R75233 VSS.n3778 VSS.n3777 0.00155634
R75234 VSS.n3240 VSS.n3236 0.00155634
R75235 VSS.n3323 VSS.n3319 0.00155634
R75236 VSS.n3377 VSS.n3373 0.00155634
R75237 VSS.n3512 VSS.n3511 0.00155634
R75238 VSS.n3515 VSS.n3514 0.00155634
R75239 VSS.n3571 VSS.n3570 0.00155634
R75240 VSS.n3574 VSS.n3573 0.00155634
R75241 VSS.n3614 VSS.n3613 0.00155634
R75242 VSS.n3617 VSS.n3616 0.00155634
R75243 VSS.n18735 VSS.n18734 0.00155634
R75244 VSS.n18739 VSS.n18738 0.00155634
R75245 VSS.n18744 VSS.n18743 0.00155634
R75246 VSS.n18794 VSS.n18793 0.00155634
R75247 VSS.n18442 VSS.n18441 0.00155634
R75248 VSS.n18395 VSS.n18394 0.00155634
R75249 VSS.n18393 VSS.n18392 0.00155634
R75250 VSS.n18204 VSS.n18203 0.00155634
R75251 VSS.n17124 VSS.n17123 0.00155634
R75252 VSS.n17031 VSS.n17030 0.00155634
R75253 VSS.n14861 VSS.n14860 0.00155634
R75254 VSS.n14873 VSS.n14872 0.00155634
R75255 VSS.n16918 VSS.n16917 0.00155634
R75256 VSS.n15405 VSS.n15404 0.00155634
R75257 VSS.n15391 VSS.n15388 0.00155634
R75258 VSS.n15329 VSS.n15328 0.00155634
R75259 VSS.n19217 VSS.n19216 0.00155634
R75260 VSS.n19221 VSS.n19220 0.00155634
R75261 VSS.n19226 VSS.n19225 0.00155634
R75262 VSS.n19466 VSS.n19465 0.00155634
R75263 VSS.n19597 VSS.n19596 0.00155634
R75264 VSS.n19627 VSS.n19626 0.00155634
R75265 VSS.n19629 VSS.n19628 0.00155634
R75266 VSS.n19652 VSS.n19651 0.00155634
R75267 VSS.n19871 VSS.n19870 0.00155634
R75268 VSS.n19904 VSS.n19903 0.00155634
R75269 VSS.n19932 VSS.n19931 0.00155634
R75270 VSS.n19944 VSS.n19943 0.00155634
R75271 VSS.n19998 VSS.n19997 0.00155634
R75272 VSS.n1721 VSS.n1720 0.00155634
R75273 VSS.n1707 VSS.n1704 0.00155634
R75274 VSS.n1645 VSS.n1644 0.00155634
R75275 VSS.n2954 VSS.n2953 0.00154636
R75276 VSS.n3066 VSS.n3065 0.00154636
R75277 VSS.n3067 VSS.n3066 0.00154636
R75278 VSS.n2955 VSS.n2954 0.00154636
R75279 VSS.n3210 DVSS 0.00153286
R75280 VSS.n5879 VSS.n5878 0.00153143
R75281 VSS.n3991 VSS.n3990 0.00153143
R75282 VSS.n12819 VSS.n12818 0.00153143
R75283 VSS.n12538 VSS.n12537 0.00153143
R75284 VSS.n11893 VSS.n11892 0.00153143
R75285 VSS.n11802 VSS.n11801 0.00153143
R75286 VSS.n13017 VSS.n13016 0.00153143
R75287 VSS.n16380 VSS.n16379 0.00153143
R75288 VSS.n18862 VSS.n18861 0.00153143
R75289 VSS.n21188 VSS.n21187 0.00153143
R75290 VSS.n21790 VSS.n21789 0.00153143
R75291 VSS.n1463 VSS.n1462 0.00153143
R75292 VSS.n19075 VSS.n19074 0.00153143
R75293 VSS.n1464 VSS.n1463 0.00153143
R75294 VSS.n12820 VSS.n12819 0.00153143
R75295 VSS.n21189 VSS.n21188 0.00153143
R75296 VSS.n21622 VSS.n21621 0.00153143
R75297 VSS.n21670 VSS.n21669 0.00153143
R75298 VSS.n21673 VSS.n21672 0.00153143
R75299 VSS.n7544 VSS.n7543 0.00153143
R75300 VSS.n21669 VSS.n21668 0.00153143
R75301 VSS.n21672 VSS.n21671 0.00153143
R75302 VSS.n11894 VSS.n11893 0.00153143
R75303 VSS.n11801 VSS.n11800 0.00153143
R75304 VSS.n12238 VSS.n12237 0.00153143
R75305 VSS.n12539 VSS.n12538 0.00153143
R75306 VSS.n16381 VSS.n16380 0.00153143
R75307 VSS.n5880 VSS.n5879 0.00153143
R75308 VSS.n3851 VSS.n3850 0.00153143
R75309 VSS.n4130 VSS.n4129 0.00153143
R75310 VSS.n4134 VSS.n4133 0.00153143
R75311 VSS.n4133 VSS.n4132 0.00153143
R75312 VSS.n11238 VSS.n11237 0.00153143
R75313 VSS.n4131 VSS.n4130 0.00153143
R75314 VSS.n3850 VSS.n3849 0.00153143
R75315 VSS.n21621 VSS.n21620 0.00153143
R75316 VSS.n3271 VSS.n3270 0.00153143
R75317 VSS.n518 VSS.n517 0.00153143
R75318 VSS.n10483 VSS.n10482 0.00153143
R75319 VSS.n10186 VSS.n10185 0.00153143
R75320 VSS.n8985 VSS.n8983 0.00153143
R75321 VSS.n10187 VSS.n10186 0.00153143
R75322 VSS.n8985 VSS.n8984 0.00153143
R75323 VSS.n10484 VSS.n10483 0.00153143
R75324 VSS.n519 VSS.n518 0.00153143
R75325 VSS.n8904 VSS.n8903 0.00153143
R75326 VSS.n2875 VSS.n2874 0.00152857
R75327 VSS.n2525 VSS.n2524 0.00152857
R75328 VSS.n2769 VSS.n2768 0.00152857
R75329 VSS.n2879 VSS.n2878 0.00152857
R75330 VSS.n2957 VSS.n2956 0.00152857
R75331 VSS.n3021 VSS.n3020 0.00152857
R75332 VSS.n3069 VSS.n3068 0.00152857
R75333 VSS.n2566 VSS.n2565 0.00152857
R75334 VSS.n2563 VSS.n2562 0.00152857
R75335 VSS.n5151 VSS.n5150 0.00152857
R75336 VSS.n4935 VSS.n4934 0.00152857
R75337 VSS.n4989 VSS.n4988 0.00152857
R75338 VSS.n5019 VSS.n5018 0.00152857
R75339 VSS.n5065 VSS.n5064 0.00152857
R75340 VSS.n5153 VSS.n5152 0.00152857
R75341 VSS.n5154 VSS.n5153 0.00152857
R75342 VSS.n7229 VSS.n7228 0.00152857
R75343 VSS.n5907 VSS.n5906 0.00152857
R75344 VSS.n7406 VSS.n7405 0.00152857
R75345 VSS.n7351 VSS.n7350 0.00152857
R75346 VSS.n7297 VSS.n7296 0.00152857
R75347 VSS.n7230 VSS.n7225 0.00152857
R75348 VSS.n7225 VSS.n7224 0.00152857
R75349 VSS.n4505 VSS.n4504 0.00152857
R75350 VSS.n2434 VSS.n2433 0.00152857
R75351 VSS.n4636 VSS.n4635 0.00152857
R75352 VSS.n4590 VSS.n4589 0.00152857
R75353 VSS.n4506 VSS.n4501 0.00152857
R75354 VSS.n4501 VSS.n4500 0.00152857
R75355 VSS.n4332 VSS.n4331 0.00152857
R75356 VSS.n4329 VSS.n4328 0.00152857
R75357 VSS.n4735 VSS.n4734 0.00152857
R75358 VSS.n17560 VSS.n17559 0.00152857
R75359 VSS.n17502 VSS.n17501 0.00152857
R75360 VSS.n18020 VSS.n18019 0.00152857
R75361 VSS.n17854 VSS.n17853 0.00152857
R75362 VSS.n17793 VSS.n17792 0.00152857
R75363 VSS.n17748 VSS.n17747 0.00152857
R75364 VSS.n17724 VSS.n17723 0.00152857
R75365 VSS.n17721 VSS.n17720 0.00152857
R75366 VSS.n18024 VSS.n18023 0.00152857
R75367 VSS.n17084 VSS.n17083 0.00152817
R75368 VSS.n19881 VSS.n19880 0.00152817
R75369 VSS.n18730 VSS.n18729 0.00152811
R75370 VSS.n18438 VSS.n18437 0.00152811
R75371 VSS.n18729 VSS.n18728 0.00152811
R75372 VSS.n19212 VSS.n19211 0.00152811
R75373 VSS.n19601 VSS.n19600 0.00152811
R75374 VSS.n19211 VSS.n19210 0.00152811
R75375 VSS.n2665 VSS.n2664 0.00151423
R75376 VSS.n2709 VSS.n2708 0.00151423
R75377 VSS.n2708 VSS.n2707 0.00151423
R75378 VSS.n2664 VSS.n2663 0.00151423
R75379 VSS.n146 VSS.n145 0.00150559
R75380 VSS.n133 VSS.n130 0.00150559
R75381 VSS.n115 VSS.n114 0.00150559
R75382 VSS.n102 VSS.n99 0.00150559
R75383 VSS.n83 VSS.n82 0.00150559
R75384 VSS.n70 VSS.n67 0.00150559
R75385 VSS.n235 VSS.n232 0.00150559
R75386 VSS.n248 VSS.n247 0.00150559
R75387 VSS.n267 VSS.n264 0.00150559
R75388 VSS.n280 VSS.n279 0.00150559
R75389 VSS.n299 VSS.n296 0.00150559
R75390 VSS.n312 VSS.n311 0.00150559
R75391 VSS.n3438 VSS.n3435 0.00148592
R75392 VSS.n3438 VSS.n3437 0.00148592
R75393 VSS.n3433 VSS.n3432 0.00148592
R75394 VSS.n3434 VSS.n3433 0.00148592
R75395 VSS.n3439 VSS.n3434 0.00148592
R75396 VSS.n3440 VSS.n3439 0.00148592
R75397 VSS.n5779 VSS.n5776 0.00147867
R75398 VSS.n5828 VSS.n5827 0.00147867
R75399 VSS.n5806 VSS.n5805 0.00147867
R75400 VSS.n1200 VSS.n1199 0.00147867
R75401 VSS.n1258 VSS.n1257 0.00147867
R75402 VSS.n5807 VSS.n5806 0.00147867
R75403 VSS.n5829 VSS.n5828 0.00147867
R75404 VSS.n5776 VSS.n5775 0.00147867
R75405 VSS.n1261 VSS.n1258 0.00147867
R75406 VSS.n1203 VSS.n1200 0.00147867
R75407 VSS.n2528 VSS.n2526 0.00146429
R75408 VSS.n2670 VSS.n2667 0.00146429
R75409 VSS.n2714 VSS.n2711 0.00146429
R75410 VSS.n2774 VSS.n2771 0.00146429
R75411 VSS.n2529 VSS.n2525 0.00146429
R75412 VSS.n2532 VSS.n2531 0.00146429
R75413 VSS.n2535 VSS.n2534 0.00146429
R75414 VSS.n2589 VSS.n2588 0.00146429
R75415 VSS.n2706 VSS.n2705 0.00146429
R75416 VSS.n2766 VSS.n2765 0.00146429
R75417 VSS.n2882 VSS.n2881 0.00146429
R75418 VSS.n4939 VSS.n4936 0.00146429
R75419 VSS.n4993 VSS.n4990 0.00146429
R75420 VSS.n5023 VSS.n5020 0.00146429
R75421 VSS.n5069 VSS.n5066 0.00146429
R75422 VSS.n4940 VSS.n4935 0.00146429
R75423 VSS.n4994 VSS.n4989 0.00146429
R75424 VSS.n5024 VSS.n5019 0.00146429
R75425 VSS.n5070 VSS.n5065 0.00146429
R75426 VSS.n5910 VSS.n5908 0.00146429
R75427 VSS.n7403 VSS.n7400 0.00146429
R75428 VSS.n7371 VSS.n7368 0.00146429
R75429 VSS.n7317 VSS.n7314 0.00146429
R75430 VSS.n5911 VSS.n5907 0.00146429
R75431 VSS.n7405 VSS.n7404 0.00146429
R75432 VSS.n7373 VSS.n7372 0.00146429
R75433 VSS.n7319 VSS.n7318 0.00146429
R75434 VSS.n7187 VSS.n7186 0.00146429
R75435 VSS.n7184 VSS.n7183 0.00146429
R75436 VSS.n7128 VSS.n7127 0.00146429
R75437 VSS.n7125 VSS.n7124 0.00146429
R75438 VSS.n2438 VSS.n2435 0.00146429
R75439 VSS.n4633 VSS.n4630 0.00146429
R75440 VSS.n4587 VSS.n4584 0.00146429
R75441 VSS.n2439 VSS.n2434 0.00146429
R75442 VSS.n2442 VSS.n2441 0.00146429
R75443 VSS.n4693 VSS.n4692 0.00146429
R75444 VSS.n4635 VSS.n4634 0.00146429
R75445 VSS.n4589 VSS.n4588 0.00146429
R75446 VSS.n4740 VSS.n4735 0.00146429
R75447 VSS.n4743 VSS.n4742 0.00146429
R75448 VSS.n4746 VSS.n4745 0.00146429
R75449 VSS.n17562 VSS.n17561 0.00146429
R75450 VSS.n17504 VSS.n17503 0.00146429
R75451 VSS.n18018 VSS.n18017 0.00146429
R75452 VSS.n4739 VSS.n4736 0.00146429
R75453 VSS.n17556 VSS.n17553 0.00146429
R75454 VSS.n17498 VSS.n17495 0.00146429
R75455 VSS.n10276 VSS.n10275 0.00146154
R75456 VSS.n10291 VSS.n10286 0.00146154
R75457 VSS.n10409 VSS.n10404 0.00146154
R75458 VSS.n10394 VSS.n10393 0.00146154
R75459 VSS.n10124 VSS.n10119 0.00146154
R75460 VSS.n10109 VSS.n10108 0.00146154
R75461 VSS.n8837 VSS.n8836 0.00146154
R75462 VSS.n8865 VSS.n8850 0.00146154
R75463 VSS.n12330 VSS.n12329 0.00146154
R75464 VSS.n12345 VSS.n12340 0.00146154
R75465 VSS.n12463 VSS.n12458 0.00146154
R75466 VSS.n12448 VSS.n12447 0.00146154
R75467 VSS.n12175 VSS.n12170 0.00146154
R75468 VSS.n12160 VSS.n12159 0.00146154
R75469 VSS.n12027 VSS.n12022 0.00146154
R75470 VSS.n12012 VSS.n12011 0.00146154
R75471 VSS.n9851 VSS.n9850 0.00146154
R75472 VSS.n12648 VSS.n12647 0.00146154
R75473 VSS.n10887 VSS.n10886 0.00146
R75474 VSS.n10905 VSS.n10904 0.00146
R75475 VSS.n5686 VSS.n5685 0.00145745
R75476 VSS.n5675 VSS.n5673 0.00145745
R75477 VSS.n16019 VSS.n16016 0.00145745
R75478 VSS.n16009 VSS.n16007 0.00145745
R75479 VSS.n1000 VSS.n997 0.00145745
R75480 VSS.n990 VSS.n988 0.00145745
R75481 VSS.n20944 VSS.n20942 0.00145745
R75482 VSS.n20955 VSS.n20954 0.00145745
R75483 VSS.n5795 VSS.n5794 0.00145745
R75484 VSS.n1239 VSS.n1238 0.00145745
R75485 VSS.n1228 VSS.n1226 0.00145745
R75486 VSS.n14138 VSS.n14137 0.00144995
R75487 VSS.n4013 VSS.n4012 0.00144287
R75488 VSS.n4012 VSS.n4011 0.00144287
R75489 VSS.n13038 VSS.n13037 0.00144287
R75490 VSS.n12591 VSS.n12590 0.00144287
R75491 VSS.n12220 VSS.n12219 0.00144287
R75492 VSS.n11866 VSS.n11865 0.00144287
R75493 VSS.n13037 VSS.n13036 0.00144287
R75494 VSS.n18884 VSS.n18883 0.00144287
R75495 VSS.n18883 VSS.n18882 0.00144287
R75496 VSS.n21811 VSS.n21810 0.00144287
R75497 VSS.n21810 VSS.n21809 0.00144287
R75498 VSS.n19096 VSS.n19095 0.00144287
R75499 VSS.n19095 VSS.n19094 0.00144287
R75500 VSS.n21582 VSS.n21581 0.00144287
R75501 VSS.n21581 VSS.n21580 0.00144287
R75502 VSS.n12219 VSS.n12218 0.00144287
R75503 VSS.n11867 VSS.n11866 0.00144287
R75504 VSS.n12590 VSS.n12589 0.00144287
R75505 VSS.n3815 VSS.n3814 0.00144287
R75506 VSS.n3814 VSS.n3813 0.00144287
R75507 VSS.n3256 VSS.n3255 0.00144287
R75508 VSS.n3257 VSS.n3256 0.00144287
R75509 VSS.n10525 VSS.n10524 0.00144287
R75510 VSS.n10168 VSS.n10167 0.00144287
R75511 VSS.n8914 VSS.n8913 0.00144287
R75512 VSS.n1769 VSS.n1768 0.0014225
R75513 VSS.n18439 VSS.n18438 0.0014225
R75514 VSS.n16539 VSS.n16538 0.0014225
R75515 VSS.n15336 VSS.n15335 0.0014225
R75516 VSS.n16932 VSS.n16931 0.0014225
R75517 VSS.n16540 VSS.n16539 0.0014225
R75518 VSS.n18780 VSS.n18779 0.0014225
R75519 VSS.n18440 VSS.n18439 0.0014225
R75520 VSS.n15467 VSS.n15466 0.0014225
R75521 VSS.n15337 VSS.n15336 0.0014225
R75522 VSS.n19600 VSS.n19599 0.0014225
R75523 VSS.n19984 VSS.n19983 0.0014225
R75524 VSS.n799 VSS.n798 0.0014225
R75525 VSS.n1652 VSS.n1651 0.0014225
R75526 VSS.n1653 VSS.n1652 0.0014225
R75527 VSS.n798 VSS.n797 0.0014225
R75528 VSS.n19452 VSS.n19451 0.0014225
R75529 VSS.n19599 VSS.n19598 0.0014225
R75530 VSS.n4110 VSS.n4109 0.00141663
R75531 VSS.n21906 VSS.n21905 0.00141663
R75532 VSS.n21909 VSS.n21906 0.00141663
R75533 VSS.n4113 VSS.n4110 0.00141663
R75534 VSS.n3192 VSS.n3191 0.00141549
R75535 VSS.n3239 VSS.n3238 0.00141549
R75536 VSS.n3322 VSS.n3321 0.00141549
R75537 VSS.n3376 VSS.n3375 0.00141549
R75538 VSS.n3194 VSS.n3193 0.00141549
R75539 VSS.n3241 VSS.n3240 0.00141549
R75540 VSS.n3324 VSS.n3323 0.00141549
R75541 VSS.n3378 VSS.n3377 0.00141549
R75542 DVSS VSS.n7516 0.00141429
R75543 VSS.n689 VSS.n688 0.00140496
R75544 VSS.n690 VSS.n689 0.00140496
R75545 VSS.n6776 VSS.n6775 0.00140496
R75546 VSS.n6716 VSS.n6715 0.00140496
R75547 VSS.n6717 VSS.n6716 0.00140496
R75548 VSS.n6777 VSS.n6776 0.00140496
R75549 VSS.n9334 VSS.n9333 0.00140496
R75550 VSS.n9388 VSS.n9387 0.00140496
R75551 VSS.n9383 VSS.n9382 0.00140496
R75552 VSS.n9329 VSS.n9328 0.00140496
R75553 VSS.n6769 VSS.n6768 0.00140496
R75554 VSS.n6709 VSS.n6708 0.00140496
R75555 VSS.n8092 VSS.n8091 0.00140496
R75556 VSS.n8032 VSS.n8031 0.00140496
R75557 VSS.n9720 VSS.n9719 0.00140496
R75558 VSS.n9778 VSS.n9777 0.00140496
R75559 VSS.n9773 VSS.n9772 0.00140496
R75560 VSS.n9724 VSS.n9723 0.00140496
R75561 VSS.n8093 VSS.n8092 0.00140496
R75562 VSS.n8033 VSS.n8032 0.00140496
R75563 VSS.n14176 VSS.n14175 0.0014
R75564 VSS.n19397 VSS.n19396 0.0014
R75565 VSS.n19387 VSS.n19385 0.0014
R75566 VSS.n19383 VSS.n19382 0.0014
R75567 VSS.n19380 VSS.n19379 0.0014
R75568 VSS.n18269 VSS.n18267 0.0014
R75569 VSS.n16655 VSS.n16654 0.0014
R75570 VSS.n16622 VSS.n16621 0.0014
R75571 VSS.n2844 VSS.n2841 0.0014
R75572 VSS.n2844 VSS.n2843 0.0014
R75573 VSS.n2838 VSS.n2837 0.0014
R75574 VSS.n2839 VSS.n2838 0.0014
R75575 VSS.n2846 VSS.n2845 0.0014
R75576 VSS.n5123 VSS.n5120 0.0014
R75577 VSS.n5123 VSS.n5122 0.0014
R75578 VSS.n5118 VSS.n5117 0.0014
R75579 VSS.n5119 VSS.n5118 0.0014
R75580 VSS.n5124 VSS.n5119 0.0014
R75581 VSS.n5125 VSS.n5124 0.0014
R75582 VSS.n7255 VSS.n7252 0.0014
R75583 VSS.n7255 VSS.n7254 0.0014
R75584 VSS.n7259 VSS.n7258 0.0014
R75585 VSS.n7258 VSS.n7257 0.0014
R75586 VSS.n7257 VSS.n7256 0.0014
R75587 VSS.n7256 VSS.n7251 0.0014
R75588 VSS.n4533 VSS.n4530 0.0014
R75589 VSS.n4533 VSS.n4532 0.0014
R75590 VSS.n4537 VSS.n4536 0.0014
R75591 VSS.n4536 VSS.n4535 0.0014
R75592 VSS.n4535 VSS.n4534 0.0014
R75593 VSS.n4534 VSS.n4529 0.0014
R75594 VSS.n18059 VSS.n18058 0.0014
R75595 VSS.n18058 VSS.n18057 0.0014
R75596 VSS.n18055 VSS.n18050 0.0014
R75597 VSS.n18054 VSS.n18051 0.0014
R75598 VSS.n18054 VSS.n18053 0.0014
R75599 VSS.n9776 VSS.n9774 0.0014
R75600 VSS.n10688 VSS.n10687 0.0014
R75601 VSS.n10750 VSS.n10749 0.0014
R75602 VSS.n4019 VSS.n4018 0.00138583
R75603 VSS.n5628 VSS.n5627 0.00138583
R75604 VSS.n5614 VSS.n5613 0.00138583
R75605 VSS.n5556 VSS.n5555 0.00138583
R75606 VSS.n13044 VSS.n13043 0.00138583
R75607 VSS.n12586 VSS.n12585 0.00138583
R75608 VSS.n12559 VSS.n12558 0.00138583
R75609 VSS.n12543 VSS.n12542 0.00138583
R75610 VSS.n12292 VSS.n12291 0.00138583
R75611 VSS.n12276 VSS.n12275 0.00138583
R75612 VSS.n12275 VSS.n12274 0.00138583
R75613 VSS.n11944 VSS.n11943 0.00138583
R75614 VSS.n11931 VSS.n11930 0.00138583
R75615 VSS.n11930 VSS.n11929 0.00138583
R75616 VSS.n11815 VSS.n11814 0.00138583
R75617 VSS.n11799 VSS.n11798 0.00138583
R75618 VSS.n11797 VSS.n11796 0.00138583
R75619 VSS.n11794 VSS.n11793 0.00138583
R75620 VSS.n18890 VSS.n18889 0.00138583
R75621 VSS.n16150 VSS.n16149 0.00138583
R75622 VSS.n16130 VSS.n16129 0.00138583
R75623 VSS.n16066 VSS.n16065 0.00138583
R75624 VSS.n21817 VSS.n21816 0.00138583
R75625 VSS.n21078 VSS.n21077 0.00138583
R75626 VSS.n21064 VSS.n21063 0.00138583
R75627 VSS.n21005 VSS.n21004 0.00138583
R75628 VSS.n19102 VSS.n19101 0.00138583
R75629 VSS.n1130 VSS.n1129 0.00138583
R75630 VSS.n1110 VSS.n1109 0.00138583
R75631 VSS.n1051 VSS.n1050 0.00138583
R75632 VSS.n21588 VSS.n21587 0.00138583
R75633 VSS.n21675 VSS.n21674 0.00138583
R75634 VSS.n21678 VSS.n21677 0.00138583
R75635 VSS.n3821 VSS.n3820 0.00138583
R75636 VSS.n4136 VSS.n4135 0.00138583
R75637 VSS.n4139 VSS.n4138 0.00138583
R75638 VSS.n3250 VSS.n3249 0.00138583
R75639 VSS.n10521 VSS.n10520 0.00138583
R75640 VSS.n10503 VSS.n10502 0.00138583
R75641 VSS.n10488 VSS.n10487 0.00138583
R75642 VSS.n10240 VSS.n10239 0.00138583
R75643 VSS.n10225 VSS.n10224 0.00138583
R75644 VSS.n10224 VSS.n10223 0.00138583
R75645 VSS.n9946 VSS.n9945 0.00138583
R75646 VSS.n9932 VSS.n9931 0.00138583
R75647 VSS.n9931 VSS.n9930 0.00138583
R75648 VSS.n8838 VSS.n8833 0.00138583
R75649 VSS.n8902 VSS.n8901 0.00138583
R75650 VSS.n8900 VSS.n8899 0.00138583
R75651 VSS.n8897 VSS.n8896 0.00138583
R75652 VSS.n2768 VSS.n2767 0.00138568
R75653 VSS.n2881 VSS.n2880 0.00138568
R75654 VSS.n2767 VSS.n2766 0.00138568
R75655 VSS.n2880 VSS.n2879 0.00138568
R75656 VSS.n5624 VSS.n5623 0.00135432
R75657 VSS.n16146 VSS.n16145 0.00135432
R75658 VSS.n21074 VSS.n21073 0.00135432
R75659 VSS.n1126 VSS.n1125 0.00135432
R75660 VSS.n2346 VSS.n2345 0.0013543
R75661 VSS.n11353 VSS.n11352 0.0013543
R75662 VSS.n5563 VSS.n5562 0.0013543
R75663 VSS.n2347 VSS.n2346 0.0013543
R75664 VSS.n11352 VSS.n11351 0.0013543
R75665 VSS.n13155 VSS.n13154 0.0013543
R75666 VSS.n12856 VSS.n12855 0.0013543
R75667 VSS.n12793 VSS.n12792 0.0013543
R75668 VSS.n12546 VSS.n12545 0.0013543
R75669 VSS.n12302 VSS.n12301 0.0013543
R75670 VSS.n12296 VSS.n12295 0.0013543
R75671 VSS.n11951 VSS.n11950 0.0013543
R75672 VSS.n11947 VSS.n11946 0.0013543
R75673 VSS.n12794 VSS.n12793 0.0013543
R75674 VSS.n12857 VSS.n12856 0.0013543
R75675 VSS.n13154 VSS.n13153 0.0013543
R75676 VSS.n5564 VSS.n5563 0.0013543
R75677 VSS.n2246 VSS.n2245 0.0013543
R75678 VSS.n15154 VSS.n15153 0.0013543
R75679 VSS.n16079 VSS.n16072 0.0013543
R75680 VSS.n16080 VSS.n16079 0.0013543
R75681 VSS.n15153 VSS.n15152 0.0013543
R75682 VSS.n2245 VSS.n2244 0.0013543
R75683 VSS.n2295 VSS.n2294 0.0013543
R75684 VSS.n20804 VSS.n20803 0.0013543
R75685 VSS.n21012 VSS.n21011 0.0013543
R75686 VSS.n21013 VSS.n21012 0.0013543
R75687 VSS.n20803 VSS.n20802 0.0013543
R75688 VSS.n2294 VSS.n2293 0.0013543
R75689 VSS.n17903 VSS.n17902 0.0013543
R75690 VSS.n2015 VSS.n2014 0.0013543
R75691 VSS.n1058 VSS.n1057 0.0013543
R75692 VSS.n1059 VSS.n1058 0.0013543
R75693 VSS.n2016 VSS.n2015 0.0013543
R75694 VSS.n17902 VSS.n17901 0.0013543
R75695 VSS.n21518 VSS.n21517 0.0013543
R75696 VSS.n21473 VSS.n21472 0.0013543
R75697 VSS.n21460 VSS.n21459 0.0013543
R75698 VSS.n21277 VSS.n21276 0.0013543
R75699 VSS.n7569 VSS.n7568 0.0013543
R75700 VSS.n7568 VSS.n7567 0.0013543
R75701 VSS.n21278 VSS.n21277 0.0013543
R75702 VSS.n21474 VSS.n21473 0.0013543
R75703 VSS.n21519 VSS.n21518 0.0013543
R75704 VSS.n21461 VSS.n21460 0.0013543
R75705 VSS.n11948 VSS.n11947 0.0013543
R75706 VSS.n11952 VSS.n11951 0.0013543
R75707 VSS.n12297 VSS.n12296 0.0013543
R75708 VSS.n12303 VSS.n12302 0.0013543
R75709 VSS.n12545 VSS.n12544 0.0013543
R75710 VSS.n4700 VSS.n4699 0.0013543
R75711 VSS.n4774 VSS.n4773 0.0013543
R75712 VSS.n11435 VSS.n11434 0.0013543
R75713 VSS.n11215 VSS.n11214 0.0013543
R75714 VSS.n4699 VSS.n4698 0.0013543
R75715 VSS.n4763 VSS.n4762 0.0013543
R75716 VSS.n11436 VSS.n11435 0.0013543
R75717 VSS.n11214 VSS.n11213 0.0013543
R75718 VSS.n4775 VSS.n4774 0.0013543
R75719 VSS.n553 VSS.n552 0.0013543
R75720 VSS.n495 VSS.n494 0.0013543
R75721 VSS.n10491 VSS.n10490 0.0013543
R75722 VSS.n10250 VSS.n10249 0.0013543
R75723 VSS.n10244 VSS.n10243 0.0013543
R75724 VSS.n9953 VSS.n9952 0.0013543
R75725 VSS.n9949 VSS.n9948 0.0013543
R75726 VSS.n10245 VSS.n10244 0.0013543
R75727 VSS.n9950 VSS.n9949 0.0013543
R75728 VSS.n10251 VSS.n10250 0.0013543
R75729 VSS.n9954 VSS.n9953 0.0013543
R75730 VSS.n10490 VSS.n10489 0.0013543
R75731 VSS.n554 VSS.n553 0.0013543
R75732 VSS.n494 VSS.n493 0.0013543
R75733 VSS.n3020 VSS.n3019 0.00135354
R75734 VSS.n3019 VSS.n3018 0.00135354
R75735 VSS.n3470 VSS.n3467 0.00134507
R75736 VSS.n3187 VSS.n3186 0.00134507
R75737 VSS.n3234 VSS.n3233 0.00134507
R75738 VSS.n3235 VSS.n3234 0.00134507
R75739 VSS.n3302 VSS.n3301 0.00134507
R75740 VSS.n3317 VSS.n3316 0.00134507
R75741 VSS.n3318 VSS.n3317 0.00134507
R75742 VSS.n3340 VSS.n3339 0.00134507
R75743 VSS.n3371 VSS.n3370 0.00134507
R75744 VSS.n3372 VSS.n3371 0.00134507
R75745 VSS.n3394 VSS.n3393 0.00134507
R75746 VSS.n3471 VSS.n3466 0.00134507
R75747 VSS.n3474 VSS.n3473 0.00134507
R75748 VSS.n3514 VSS.n3513 0.00134507
R75749 VSS.n3540 VSS.n3539 0.00134507
R75750 VSS.n3573 VSS.n3572 0.00134507
R75751 VSS.n3599 VSS.n3598 0.00134507
R75752 VSS.n3616 VSS.n3615 0.00134507
R75753 VSS.n3642 VSS.n3641 0.00134507
R75754 VSS.n18707 VSS.n18706 0.00134507
R75755 VSS.n18710 VSS.n18709 0.00134507
R75756 VSS.n18776 VSS.n18775 0.00134507
R75757 VSS.n18789 VSS.n18788 0.00134507
R75758 VSS.n18803 VSS.n18802 0.00134507
R75759 VSS.n18809 VSS.n18808 0.00134507
R75760 VSS.n18810 VSS.n18809 0.00134507
R75761 VSS.n18812 VSS.n18811 0.00134507
R75762 VSS.n18190 VSS.n18189 0.00134507
R75763 VSS.n18186 VSS.n18185 0.00134507
R75764 VSS.n17015 VSS.n17014 0.00134507
R75765 VSS.n17012 VSS.n17011 0.00134507
R75766 VSS.n17011 VSS.n17010 0.00134507
R75767 VSS.n16928 VSS.n16927 0.00134507
R75768 VSS.n16914 VSS.n16913 0.00134507
R75769 VSS.n16636 VSS.n16635 0.00134507
R75770 VSS.n16593 VSS.n16592 0.00134507
R75771 VSS.n15524 VSS.n15523 0.00134507
R75772 VSS.n15388 VSS.n15387 0.00134507
R75773 VSS.n15384 VSS.n15383 0.00134507
R75774 VSS.n15341 VSS.n15340 0.00134507
R75775 VSS.n15331 VSS.n15330 0.00134507
R75776 VSS.n8512 VSS.n8511 0.00134507
R75777 VSS.n19189 VSS.n19188 0.00134507
R75778 VSS.n19192 VSS.n19191 0.00134507
R75779 VSS.n19448 VSS.n19447 0.00134507
R75780 VSS.n19461 VSS.n19460 0.00134507
R75781 VSS.n19475 VSS.n19474 0.00134507
R75782 VSS.n19481 VSS.n19480 0.00134507
R75783 VSS.n19482 VSS.n19481 0.00134507
R75784 VSS.n19484 VSS.n19483 0.00134507
R75785 VSS.n19666 VSS.n19665 0.00134507
R75786 VSS.n19670 VSS.n19669 0.00134507
R75787 VSS.n19920 VSS.n19919 0.00134507
R75788 VSS.n19923 VSS.n19922 0.00134507
R75789 VSS.n19924 VSS.n19923 0.00134507
R75790 VSS.n19988 VSS.n19987 0.00134507
R75791 VSS.n20002 VSS.n20001 0.00134507
R75792 VSS.n762 VSS.n761 0.00134507
R75793 VSS.n775 VSS.n774 0.00134507
R75794 VSS.n1812 VSS.n1811 0.00134507
R75795 VSS.n1704 VSS.n1703 0.00134507
R75796 VSS.n1700 VSS.n1699 0.00134507
R75797 VSS.n1657 VSS.n1656 0.00134507
R75798 VSS.n1647 VSS.n1646 0.00134507
R75799 VSS.n8663 VSS.n8662 0.00134507
R75800 VSS.n20260 VSS.n20259 0.00134497
R75801 VSS.n20259 VSS.n20258 0.00134497
R75802 VSS.n20550 DVSS 0.00134
R75803 DVSS VSS.n20551 0.00134
R75804 DVSS VSS.n11076 0.00134
R75805 VSS.n11075 DVSS 0.00134
R75806 VSS.n2528 VSS.n2527 0.00133571
R75807 VSS.n2670 VSS.n2669 0.00133571
R75808 VSS.n2714 VSS.n2713 0.00133571
R75809 VSS.n2774 VSS.n2773 0.00133571
R75810 VSS.n2530 VSS.n2529 0.00133571
R75811 VSS.n2672 VSS.n2671 0.00133571
R75812 VSS.n2716 VSS.n2715 0.00133571
R75813 VSS.n2776 VSS.n2775 0.00133571
R75814 VSS.n2837 VSS.n2836 0.00133571
R75815 VSS.n2840 VSS.n2839 0.00133571
R75816 VSS.n2888 VSS.n2884 0.00133571
R75817 VSS.n4939 VSS.n4938 0.00133571
R75818 VSS.n4993 VSS.n4992 0.00133571
R75819 VSS.n5023 VSS.n5022 0.00133571
R75820 VSS.n5069 VSS.n5068 0.00133571
R75821 VSS.n4941 VSS.n4940 0.00133571
R75822 VSS.n4995 VSS.n4994 0.00133571
R75823 VSS.n5025 VSS.n5024 0.00133571
R75824 VSS.n5071 VSS.n5070 0.00133571
R75825 VSS.n5910 VSS.n5909 0.00133571
R75826 VSS.n7403 VSS.n7402 0.00133571
R75827 VSS.n7371 VSS.n7370 0.00133571
R75828 VSS.n7317 VSS.n7316 0.00133571
R75829 VSS.n5912 VSS.n5911 0.00133571
R75830 VSS.n7404 VSS.n7399 0.00133571
R75831 VSS.n7372 VSS.n7367 0.00133571
R75832 VSS.n7318 VSS.n7313 0.00133571
R75833 VSS.n2438 VSS.n2436 0.00133571
R75834 VSS.n4633 VSS.n4632 0.00133571
R75835 VSS.n4587 VSS.n4586 0.00133571
R75836 VSS.n2440 VSS.n2439 0.00133571
R75837 VSS.n4634 VSS.n4629 0.00133571
R75838 VSS.n4588 VSS.n4583 0.00133571
R75839 VSS.n4741 VSS.n4740 0.00133571
R75840 VSS.n17557 VSS.n17552 0.00133571
R75841 VSS.n17499 VSS.n17494 0.00133571
R75842 VSS.n18060 VSS.n18059 0.00133571
R75843 VSS.n18057 VSS.n18056 0.00133571
R75844 VSS.n18015 VSS.n18014 0.00133571
R75845 VSS.n4739 VSS.n4738 0.00133571
R75846 VSS.n17556 VSS.n17555 0.00133571
R75847 VSS.n17498 VSS.n17497 0.00133571
R75848 VSS.n4166 VSS.n4165 0.00133333
R75849 VSS.n21708 VSS.n21707 0.00133333
R75850 VSS.n17402 VSS.n17401 0.00133333
R75851 VSS.n13284 VSS.n375 0.00133333
R75852 VSS.n18807 VSS.n18806 0.00131688
R75853 VSS.n18167 VSS.n18166 0.00131688
R75854 VSS.n14988 VSS.n14987 0.00131688
R75855 VSS.n8524 VSS.n8523 0.00131688
R75856 VSS.n8342 VSS.n8341 0.00131688
R75857 VSS.n16898 VSS.n16897 0.00131688
R75858 VSS.n16591 VSS.n16590 0.00131688
R75859 VSS.n18806 VSS.n18805 0.00131688
R75860 VSS.n18168 VSS.n18167 0.00131688
R75861 VSS.n15394 VSS.n15393 0.00131688
R75862 VSS.n8341 VSS.n8340 0.00131688
R75863 VSS.n8523 VSS.n8522 0.00131688
R75864 VSS.n15387 VSS.n15386 0.00131688
R75865 VSS.n19479 VSS.n19478 0.00131688
R75866 VSS.n19689 VSS.n19688 0.00131688
R75867 VSS.n20018 VSS.n20017 0.00131688
R75868 VSS.n777 VSS.n776 0.00131688
R75869 VSS.n824 VSS.n823 0.00131688
R75870 VSS.n8675 VSS.n8674 0.00131688
R75871 VSS.n8138 VSS.n8137 0.00131688
R75872 VSS.n8137 VSS.n8136 0.00131688
R75873 VSS.n8674 VSS.n8673 0.00131688
R75874 VSS.n1703 VSS.n1702 0.00131688
R75875 VSS.n1710 VSS.n1709 0.00131688
R75876 VSS.n19688 VSS.n19687 0.00131688
R75877 VSS.n19478 VSS.n19477 0.00131688
R75878 VSS.n20204 VSS.n20203 0.00131498
R75879 VSS.n20205 VSS.n20204 0.00131498
R75880 VSS.n731 VSS.n730 0.00131
R75881 VSS.n20587 VSS.n20586 0.00131
R75882 VSS.n20505 VSS.n20504 0.00131
R75883 VSS.n20537 VSS.n20524 0.00131
R75884 VSS.n20175 VSS.n20174 0.00131
R75885 VSS.n732 VSS.n729 0.00131
R75886 VSS.n20588 VSS.n20585 0.00131
R75887 VSS.n20571 VSS.n20570 0.00131
R75888 VSS.n20565 VSS.n20564 0.00131
R75889 VSS.n20542 VSS.n20541 0.00131
R75890 VSS.n20536 VSS.n20535 0.00131
R75891 VSS.n10933 VSS.n10932 0.00131
R75892 VSS.n11000 VSS.n10999 0.00131
R75893 VSS.n11053 VSS.n11052 0.00131
R75894 VSS.n6367 VSS.n6361 0.00131
R75895 VSS.n8080 VSS.n8079 0.00131
R75896 VSS.n8020 VSS.n8019 0.00131
R75897 VSS.n7975 VSS.n7974 0.00131
R75898 VSS.n7938 VSS.n7932 0.00131
R75899 VSS.n6764 VSS.n6763 0.00131
R75900 VSS.n6704 VSS.n6703 0.00131
R75901 VSS.n7882 VSS.n7881 0.00131
R75902 VSS.n7043 VSS.n7040 0.00131
R75903 VSS.n9387 VSS.n9386 0.00131
R75904 VSS.n9382 VSS.n9381 0.00131
R75905 VSS.n9333 VSS.n9332 0.00131
R75906 VSS.n9328 VSS.n9327 0.00131
R75907 VSS.n6768 VSS.n6767 0.00131
R75908 VSS.n6708 VSS.n6707 0.00131
R75909 VSS.n7883 VSS.n7879 0.00131
R75910 VSS.n7025 VSS.n7024 0.00131
R75911 VSS.n7044 VSS.n7038 0.00131
R75912 VSS.n9779 VSS.n9778 0.00131
R75913 VSS.n9774 VSS.n9773 0.00131
R75914 VSS.n9725 VSS.n9724 0.00131
R75915 VSS.n9719 VSS.n9718 0.00131
R75916 VSS.n8085 VSS.n8084 0.00131
R75917 VSS.n8084 VSS.n8083 0.00131
R75918 VSS.n8025 VSS.n8024 0.00131
R75919 VSS.n8024 VSS.n8023 0.00131
R75920 VSS.n7976 VSS.n7972 0.00131
R75921 VSS.n7947 VSS.n7946 0.00131
R75922 VSS.n7937 VSS.n7936 0.00131
R75923 VSS.n11055 VSS.n11054 0.00131
R75924 VSS.n6373 VSS.n6372 0.00131
R75925 VSS.n6366 VSS.n6365 0.00131
R75926 VSS.n20172 VSS.n20169 0.00128
R75927 VSS.n686 VSS.n683 0.00128
R75928 VSS.n20501 VSS.n20499 0.00128
R75929 VSS.n20547 VSS.n20519 0.00128
R75930 VSS.n20174 VSS.n20173 0.00128
R75931 VSS.n729 VSS.n728 0.00128
R75932 VSS.n688 VSS.n687 0.00128
R75933 VSS.n20585 VSS.n20584 0.00128
R75934 VSS.n20570 VSS.n20569 0.00128
R75935 VSS.n20564 VSS.n20563 0.00128
R75936 VSS.n20546 VSS.n20542 0.00128
R75937 VSS.n20535 VSS.n20534 0.00128
R75938 VSS.n10922 VSS.n10920 0.00128
R75939 VSS.n10989 VSS.n10987 0.00128
R75940 VSS.n11044 VSS.n11042 0.00128
R75941 VSS.n6377 VSS.n6369 0.00128
R75942 VSS.n8089 VSS.n8087 0.00128
R75943 VSS.n8029 VSS.n8027 0.00128
R75944 VSS.n7984 VSS.n7982 0.00128
R75945 VSS.n7952 VSS.n7951 0.00128
R75946 VSS.n6773 VSS.n6771 0.00128
R75947 VSS.n6713 VSS.n6711 0.00128
R75948 VSS.n7891 VSS.n7889 0.00128
R75949 VSS.n7854 VSS.n7022 0.00128
R75950 VSS.n6779 VSS.n6778 0.00128
R75951 VSS.n6775 VSS.n6774 0.00128
R75952 VSS.n6765 VSS.n6761 0.00128
R75953 VSS.n6760 VSS.n6759 0.00128
R75954 VSS.n6719 VSS.n6718 0.00128
R75955 VSS.n6715 VSS.n6714 0.00128
R75956 VSS.n6705 VSS.n6701 0.00128
R75957 VSS.n6700 VSS.n6699 0.00128
R75958 VSS.n7893 VSS.n7892 0.00128
R75959 VSS.n7853 VSS.n7025 0.00128
R75960 VSS.n7038 VSS.n7037 0.00128
R75961 VSS.n8095 VSS.n8094 0.00128
R75962 VSS.n8091 VSS.n8090 0.00128
R75963 VSS.n8081 VSS.n8077 0.00128
R75964 VSS.n8076 VSS.n8075 0.00128
R75965 VSS.n8035 VSS.n8034 0.00128
R75966 VSS.n8031 VSS.n8030 0.00128
R75967 VSS.n8021 VSS.n8017 0.00128
R75968 VSS.n8016 VSS.n8015 0.00128
R75969 VSS.n7986 VSS.n7985 0.00128
R75970 VSS.n7950 VSS.n7947 0.00128
R75971 VSS.n7936 VSS.n7935 0.00128
R75972 VSS.n10923 VSS.n10919 0.00128
R75973 VSS.n10935 VSS.n10934 0.00128
R75974 VSS.n10990 VSS.n10986 0.00128
R75975 VSS.n11002 VSS.n11001 0.00128
R75976 VSS.n11045 VSS.n11041 0.00128
R75977 VSS.n6376 VSS.n6373 0.00128
R75978 VSS.n6365 VSS.n6364 0.00128
R75979 VSS.n3541 VSS.n3540 0.00127465
R75980 VSS.n3600 VSS.n3599 0.00127465
R75981 VSS.n3643 VSS.n3642 0.00127465
R75982 VSS.n3654 VSS.n3653 0.00127465
R75983 VSS.n2875 VSS.n2873 0.00127143
R75984 VSS.n2524 VSS.n2523 0.00127143
R75985 VSS.n2663 VSS.n2589 0.00127143
R75986 VSS.n2707 VSS.n2706 0.00127143
R75987 VSS.n2876 VSS.n2872 0.00127143
R75988 VSS.n5151 VSS.n5148 0.00127143
R75989 VSS.n4934 VSS.n4933 0.00127143
R75990 VSS.n4988 VSS.n4987 0.00127143
R75991 VSS.n5018 VSS.n5017 0.00127143
R75992 VSS.n5064 VSS.n5063 0.00127143
R75993 VSS.n5152 VSS.n5147 0.00127143
R75994 VSS.n5155 VSS.n5154 0.00127143
R75995 VSS.n7229 VSS.n7226 0.00127143
R75996 VSS.n5906 VSS.n5905 0.00127143
R75997 VSS.n7407 VSS.n7406 0.00127143
R75998 VSS.n7376 VSS.n7375 0.00127143
R75999 VSS.n7375 VSS.n7374 0.00127143
R76000 VSS.n7352 VSS.n7351 0.00127143
R76001 VSS.n7322 VSS.n7321 0.00127143
R76002 VSS.n7321 VSS.n7320 0.00127143
R76003 VSS.n7298 VSS.n7297 0.00127143
R76004 VSS.n7231 VSS.n7230 0.00127143
R76005 VSS.n7224 VSS.n7223 0.00127143
R76006 VSS.n7185 VSS.n7184 0.00127143
R76007 VSS.n7158 VSS.n7157 0.00127143
R76008 VSS.n7126 VSS.n7125 0.00127143
R76009 VSS.n7099 VSS.n7098 0.00127143
R76010 VSS.n4505 VSS.n4502 0.00127143
R76011 VSS.n2433 VSS.n2432 0.00127143
R76012 VSS.n4637 VSS.n4636 0.00127143
R76013 VSS.n4591 VSS.n4590 0.00127143
R76014 VSS.n4507 VSS.n4506 0.00127143
R76015 VSS.n4500 VSS.n4499 0.00127143
R76016 VSS.n4734 VSS.n4733 0.00127143
R76017 VSS.n17561 VSS.n17560 0.00127143
R76018 VSS.n17503 VSS.n17502 0.00127143
R76019 VSS.n18026 VSS.n18025 0.00127143
R76020 VSS.n18019 VSS.n18018 0.00127143
R76021 VSS.n18024 VSS.n18022 0.00127143
R76022 VSS.n6572 VSS.n6571 0.00126575
R76023 VSS.n6422 VSS.n6421 0.00126575
R76024 VSS.n4042 VSS.n4041 0.00126573
R76025 VSS.n17473 VSS.n17472 0.00126573
R76026 VSS.n17316 VSS.n17315 0.00126573
R76027 VSS.n5617 VSS.n5616 0.00126573
R76028 VSS.n9548 VSS.n9547 0.00126573
R76029 VSS.n9049 VSS.n9048 0.00126573
R76030 VSS.n17315 VSS.n17314 0.00126573
R76031 VSS.n4041 VSS.n4040 0.00126573
R76032 VSS.n13071 VSS.n13070 0.00126573
R76033 VSS.n13196 VSS.n13195 0.00126573
R76034 VSS.n13201 VSS.n13200 0.00126573
R76035 VSS.n12983 VSS.n12982 0.00126573
R76036 VSS.n12765 VSS.n12764 0.00126573
R76037 VSS.n12588 VSS.n12587 0.00126573
R76038 VSS.n12984 VSS.n12983 0.00126573
R76039 VSS.n13070 VSS.n13069 0.00126573
R76040 VSS.n13200 VSS.n13199 0.00126573
R76041 VSS.n17474 VSS.n17473 0.00126573
R76042 VSS.n13197 VSS.n13196 0.00126573
R76043 VSS.n18913 VSS.n18912 0.00126573
R76044 VSS.n2224 VSS.n2223 0.00126573
R76045 VSS.n14407 VSS.n14406 0.00126573
R76046 VSS.n16133 VSS.n16132 0.00126573
R76047 VSS.n9665 VSS.n9664 0.00126573
R76048 VSS.n9192 VSS.n9191 0.00126573
R76049 VSS.n2225 VSS.n2224 0.00126573
R76050 VSS.n14408 VSS.n14407 0.00126573
R76051 VSS.n18912 VSS.n18911 0.00126573
R76052 VSS.n5618 VSS.n5617 0.00126573
R76053 VSS.n16134 VSS.n16133 0.00126573
R76054 VSS.n21844 VSS.n21843 0.00126573
R76055 VSS.n2333 VSS.n2332 0.00126573
R76056 VSS.n13318 VSS.n13317 0.00126573
R76057 VSS.n20601 VSS.n20600 0.00126573
R76058 VSS.n21067 VSS.n21066 0.00126573
R76059 VSS.n6955 VSS.n6954 0.00126573
R76060 VSS.n6682 VSS.n6681 0.00126573
R76061 VSS.n21068 VSS.n21067 0.00126573
R76062 VSS.n20600 VSS.n20599 0.00126573
R76063 VSS.n2332 VSS.n2331 0.00126573
R76064 VSS.n21843 VSS.n21842 0.00126573
R76065 VSS.n13317 VSS.n13316 0.00126573
R76066 VSS.n19129 VSS.n19128 0.00126573
R76067 VSS.n17955 VSS.n17954 0.00126573
R76068 VSS.n17950 VSS.n17949 0.00126573
R76069 VSS.n20163 VSS.n20162 0.00126573
R76070 VSS.n1113 VSS.n1112 0.00126573
R76071 VSS.n6853 VSS.n6852 0.00126573
R76072 VSS.n6532 VSS.n6531 0.00126573
R76073 VSS.n1114 VSS.n1113 0.00126573
R76074 VSS.n20162 VSS.n20161 0.00126573
R76075 VSS.n17954 VSS.n17953 0.00126573
R76076 VSS.n19128 VSS.n19127 0.00126573
R76077 VSS.n17951 VSS.n17950 0.00126573
R76078 VSS.n21615 VSS.n21614 0.00126573
R76079 VSS.n21653 VSS.n21652 0.00126573
R76080 VSS.n21400 VSS.n21399 0.00126573
R76081 VSS.n7597 VSS.n7596 0.00126573
R76082 VSS.n7685 VSS.n7684 0.00126573
R76083 VSS.n7773 VSS.n7772 0.00126573
R76084 VSS.n21401 VSS.n21400 0.00126573
R76085 VSS.n21652 VSS.n21651 0.00126573
R76086 VSS.n21614 VSS.n21613 0.00126573
R76087 VSS.n7772 VSS.n7771 0.00126573
R76088 VSS.n11960 VSS.n11959 0.00126573
R76089 VSS.n6681 VSS.n6680 0.00126573
R76090 VSS.n6531 VSS.n6530 0.00126573
R76091 VSS.n9191 VSS.n9190 0.00126573
R76092 VSS.n9048 VSS.n9047 0.00126573
R76093 VSS.n7684 VSS.n7683 0.00126573
R76094 VSS.n6954 VSS.n6953 0.00126573
R76095 VSS.n6852 VSS.n6851 0.00126573
R76096 VSS.n9664 VSS.n9663 0.00126573
R76097 VSS.n9547 VSS.n9546 0.00126573
R76098 VSS.n12589 VSS.n12588 0.00126573
R76099 VSS.n7596 VSS.n7595 0.00126573
R76100 VSS.n12766 VSS.n12765 0.00126573
R76101 VSS.n3844 VSS.n3843 0.00126573
R76102 VSS.n3882 VSS.n3881 0.00126573
R76103 VSS.n11725 VSS.n11724 0.00126573
R76104 VSS.n11188 VSS.n11187 0.00126573
R76105 VSS.n6076 VSS.n6075 0.00126573
R76106 VSS.n5995 VSS.n5994 0.00126573
R76107 VSS.n5996 VSS.n5995 0.00126573
R76108 VSS.n6077 VSS.n6076 0.00126573
R76109 VSS.n11726 VSS.n11725 0.00126573
R76110 VSS.n3843 VSS.n3842 0.00126573
R76111 VSS.n11189 VSS.n11188 0.00126573
R76112 VSS.n3881 VSS.n3880 0.00126573
R76113 VSS.n2659 VSS.n2658 0.00126573
R76114 VSS.n2658 VSS.n2657 0.00126573
R76115 VSS.n677 VSS.n676 0.00126573
R76116 VSS.n468 VSS.n467 0.00126573
R76117 VSS.n9962 VSS.n9961 0.00126573
R76118 VSS.n10523 VSS.n10522 0.00126573
R76119 VSS.n9963 VSS.n9962 0.00126573
R76120 VSS.n676 VSS.n675 0.00126573
R76121 VSS.n469 VSS.n468 0.00126573
R76122 VSS.n6750 VSS.n6749 0.00125499
R76123 VSS.n6690 VSS.n6689 0.00125499
R76124 VSS.n7869 VSS.n7868 0.00125499
R76125 VSS.n7030 VSS.n7029 0.00125499
R76126 VSS.n7868 VSS.n7867 0.00125499
R76127 VSS.n7029 VSS.n7028 0.00125499
R76128 VSS.n6689 VSS.n6688 0.00125499
R76129 VSS.n6749 VSS.n6748 0.00125499
R76130 VSS.n8066 VSS.n8065 0.00125499
R76131 VSS.n8006 VSS.n8005 0.00125499
R76132 VSS.n7962 VSS.n7961 0.00125499
R76133 VSS.n7927 VSS.n7926 0.00125499
R76134 VSS.n7961 VSS.n7960 0.00125499
R76135 VSS.n7926 VSS.n7925 0.00125499
R76136 VSS.n8005 VSS.n8004 0.00125499
R76137 VSS.n8065 VSS.n8064 0.00125499
R76138 VSS.n6356 VSS.n6355 0.00125499
R76139 VSS.n6355 VSS.n6354 0.00125499
R76140 VSS.n20232 VSS.n20231 0.00125
R76141 VSS.n11720 VSS.n464 0.00125
R76142 VSS.n20374 VSS.n20373 0.00125
R76143 VSS.n20343 VSS.n20342 0.00125
R76144 VSS.n20297 VSS.n20296 0.00125
R76145 VSS.n10838 VSS.n10837 0.00125
R76146 VSS.n8745 VSS.n8744 0.00125
R76147 VSS.n8288 VSS.n8287 0.00125
R76148 VSS.n8809 VSS.n8808 0.00125
R76149 VSS.n9006 VSS.n9005 0.00125
R76150 VSS.n9396 VSS.n9395 0.00125
R76151 VSS.n9342 VSS.n9341 0.00125
R76152 VSS.n8281 VSS.n8280 0.00125
R76153 VSS.n6758 VSS.n6757 0.00125
R76154 VSS.n6698 VSS.n6697 0.00125
R76155 VSS.n9422 VSS.n9421 0.00125
R76156 VSS.n9468 VSS.n9467 0.00125
R76157 VSS.n9787 VSS.n9786 0.00125
R76158 VSS.n9733 VSS.n9732 0.00125
R76159 VSS.n8738 VSS.n8737 0.00125
R76160 VSS.n8074 VSS.n8073 0.00125
R76161 VSS.n8014 VSS.n8013 0.00125
R76162 VSS.n11183 VSS.n11182 0.00125
R76163 VSS.n10641 VSS.n10640 0.00125
R76164 VSS.n2891 VSS.n2890 0.00122499
R76165 VSS.n2890 VSS.n2889 0.00122499
R76166 VSS.n17191 VSS.n17190 0.00122499
R76167 VSS.n17197 VSS.n17196 0.00122499
R76168 VSS.n17205 VSS.n17204 0.00122499
R76169 VSS.n17211 VSS.n17210 0.00122499
R76170 VSS.n17217 VSS.n17216 0.00122499
R76171 VSS.n17202 VSS.n17201 0.00122499
R76172 VSS.n20400 VSS.n462 0.00122
R76173 VSS.n20371 VSS.n20368 0.00122
R76174 VSS.n20340 VSS.n20338 0.00122
R76175 VSS.n20294 VSS.n20292 0.00122
R76176 VSS.n20399 VSS.n464 0.00122
R76177 VSS.n20373 VSS.n20372 0.00122
R76178 VSS.n20342 VSS.n20341 0.00122
R76179 VSS.n20296 VSS.n20295 0.00122
R76180 VSS.n20225 VSS.n20224 0.00122
R76181 VSS.n20222 VSS.n20221 0.00122
R76182 VSS.n11180 VSS.n6164 0.00122
R76183 VSS.n10631 VSS.n10629 0.00122
R76184 VSS.n10678 VSS.n10676 0.00122
R76185 VSS.n10740 VSS.n10738 0.00122
R76186 VSS.n11026 VSS.n11025 0.00122
R76187 VSS.n9424 VSS.n9423 0.00122
R76188 VSS.n9458 VSS.n9456 0.00122
R76189 VSS.n9783 VSS.n9781 0.00122
R76190 VSS.n9729 VSS.n9727 0.00122
R76191 VSS.n8812 VSS.n8810 0.00122
R76192 VSS.n8924 VSS.n8922 0.00122
R76193 VSS.n9392 VSS.n9390 0.00122
R76194 VSS.n9338 VSS.n9336 0.00122
R76195 VSS.n11023 VSS.n11022 0.00122
R76196 VSS.n8813 VSS.n8809 0.00122
R76197 VSS.n8925 VSS.n8921 0.00122
R76198 VSS.n9398 VSS.n9397 0.00122
R76199 VSS.n9344 VSS.n9343 0.00122
R76200 VSS.n8279 VSS.n8278 0.00122
R76201 VSS.n7906 VSS.n7007 0.00122
R76202 VSS.n7897 VSS.n7896 0.00122
R76203 VSS.n7894 VSS.n7893 0.00122
R76204 VSS.n9425 VSS.n9422 0.00122
R76205 VSS.n9459 VSS.n9455 0.00122
R76206 VSS.n9789 VSS.n9788 0.00122
R76207 VSS.n9735 VSS.n9734 0.00122
R76208 VSS.n8736 VSS.n8735 0.00122
R76209 VSS.n8001 VSS.n7999 0.00122
R76210 VSS.n7990 VSS.n7989 0.00122
R76211 VSS.n7987 VSS.n7986 0.00122
R76212 VSS.n11182 VSS.n11181 0.00122
R76213 VSS.n10632 VSS.n10628 0.00122
R76214 VSS.n10684 VSS.n10683 0.00122
R76215 VSS.n10746 VSS.n10745 0.00122
R76216 VSS.n10927 VSS.n10926 0.00122
R76217 VSS.n10994 VSS.n10993 0.00122
R76218 VSS.n11028 VSS.n11027 0.00122
R76219 VSS.n11038 VSS.n11037 0.00122
R76220 VSS.n11041 VSS.n11040 0.00122
R76221 VSS.n18822 VSS.n18821 0.00121126
R76222 VSS.n18833 VSS.n18832 0.00121126
R76223 VSS.n18689 VSS.n18688 0.00121126
R76224 VSS.n18681 VSS.n18680 0.00121126
R76225 VSS.n18672 VSS.n18671 0.00121126
R76226 VSS.n18145 VSS.n18144 0.00121126
R76227 VSS.n14865 VSS.n14864 0.00121126
R76228 VSS.n16906 VSS.n16905 0.00121126
R76229 VSS.n15654 VSS.n15653 0.00121126
R76230 VSS.n15627 VSS.n15626 0.00121126
R76231 VSS.n15604 VSS.n15603 0.00121126
R76232 VSS.n15528 VSS.n15527 0.00121126
R76233 VSS.n15443 VSS.n15442 0.00121126
R76234 VSS.n15399 VSS.n15398 0.00121126
R76235 VSS.n15349 VSS.n15348 0.00121126
R76236 VSS.n8470 VSS.n8469 0.00121126
R76237 VSS.n8481 VSS.n8480 0.00121126
R76238 VSS.n8484 VSS.n8483 0.00121126
R76239 VSS.n8551 VSS.n8550 0.00121126
R76240 VSS.n8318 VSS.n8317 0.00121126
R76241 VSS.n8406 VSS.n8405 0.00121126
R76242 VSS.n8370 VSS.n8369 0.00121126
R76243 VSS.n8352 VSS.n8351 0.00121126
R76244 VSS.n15605 VSS.n15604 0.00121126
R76245 VSS.n15628 VSS.n15627 0.00121126
R76246 VSS.n15655 VSS.n15654 0.00121126
R76247 VSS.n16907 VSS.n16906 0.00121126
R76248 VSS.n14864 VSS.n14863 0.00121126
R76249 VSS.n17026 VSS.n17025 0.00121126
R76250 VSS.n16531 VSS.n16530 0.00121126
R76251 VSS.n18201 VSS.n18200 0.00121126
R76252 VSS.n18144 VSS.n18143 0.00121126
R76253 VSS.n15444 VSS.n15443 0.00121126
R76254 VSS.n15400 VSS.n15399 0.00121126
R76255 VSS.n15529 VSS.n15528 0.00121126
R76256 VSS.n8371 VSS.n8370 0.00121126
R76257 VSS.n8407 VSS.n8406 0.00121126
R76258 VSS.n8317 VSS.n8316 0.00121126
R76259 VSS.n8552 VSS.n8551 0.00121126
R76260 VSS.n8483 VSS.n8482 0.00121126
R76261 VSS.n8469 VSS.n8468 0.00121126
R76262 VSS.n15350 VSS.n15349 0.00121126
R76263 VSS.n19494 VSS.n19493 0.00121126
R76264 VSS.n19505 VSS.n19504 0.00121126
R76265 VSS.n19515 VSS.n19514 0.00121126
R76266 VSS.n19523 VSS.n19522 0.00121126
R76267 VSS.n19531 VSS.n19530 0.00121126
R76268 VSS.n19711 VSS.n19710 0.00121126
R76269 VSS.n19909 VSS.n19908 0.00121126
R76270 VSS.n19936 VSS.n19935 0.00121126
R76271 VSS.n20010 VSS.n20009 0.00121126
R76272 VSS.n807 VSS.n806 0.00121126
R76273 VSS.n1912 VSS.n1911 0.00121126
R76274 VSS.n1895 VSS.n1894 0.00121126
R76275 VSS.n1878 VSS.n1877 0.00121126
R76276 VSS.n1817 VSS.n1816 0.00121126
R76277 VSS.n1745 VSS.n1744 0.00121126
R76278 VSS.n1715 VSS.n1714 0.00121126
R76279 VSS.n1665 VSS.n1664 0.00121126
R76280 VSS.n8620 VSS.n8619 0.00121126
R76281 VSS.n8632 VSS.n8631 0.00121126
R76282 VSS.n8635 VSS.n8634 0.00121126
R76283 VSS.n8702 VSS.n8701 0.00121126
R76284 VSS.n8114 VSS.n8113 0.00121126
R76285 VSS.n8214 VSS.n8213 0.00121126
R76286 VSS.n8178 VSS.n8177 0.00121126
R76287 VSS.n8160 VSS.n8159 0.00121126
R76288 VSS.n8634 VSS.n8633 0.00121126
R76289 VSS.n8113 VSS.n8112 0.00121126
R76290 VSS.n8179 VSS.n8178 0.00121126
R76291 VSS.n8703 VSS.n8702 0.00121126
R76292 VSS.n8215 VSS.n8214 0.00121126
R76293 VSS.n8621 VSS.n8620 0.00121126
R76294 VSS.n1666 VSS.n1665 0.00121126
R76295 VSS.n20009 VSS.n20008 0.00121126
R76296 VSS.n19935 VSS.n19934 0.00121126
R76297 VSS.n1913 VSS.n1912 0.00121126
R76298 VSS.n1896 VSS.n1895 0.00121126
R76299 VSS.n1879 VSS.n1878 0.00121126
R76300 VSS.n19655 VSS.n19654 0.00121126
R76301 VSS.n19712 VSS.n19711 0.00121126
R76302 VSS.n1816 VSS.n1815 0.00121126
R76303 VSS.n1746 VSS.n1745 0.00121126
R76304 VSS.n1716 VSS.n1715 0.00121126
R76305 VSS.n18671 VSS.n18670 0.00121126
R76306 VSS.n19532 VSS.n19531 0.00121126
R76307 VSS.n18680 VSS.n18679 0.00121126
R76308 VSS.n18823 VSS.n18822 0.00121126
R76309 VSS.n19495 VSS.n19494 0.00121126
R76310 VSS.n18832 VSS.n18831 0.00121126
R76311 VSS.n19504 VSS.n19503 0.00121126
R76312 VSS.n19522 VSS.n19521 0.00121126
R76313 VSS.n8631 VSS.n8630 0.00121126
R76314 VSS.n8480 VSS.n8479 0.00121126
R76315 VSS.n8161 VSS.n8160 0.00121126
R76316 VSS.n8353 VSS.n8352 0.00121126
R76317 VSS.n19514 VSS.n19513 0.00121126
R76318 VSS.n18690 VSS.n18689 0.00121126
R76319 VSS.n20251 VSS.n20250 0.00120999
R76320 VSS.n20250 VSS.n20249 0.00120999
R76321 VSS.n10819 VSS.n10818 0.00120999
R76322 VSS.n10820 VSS.n10819 0.00120999
R76323 VSS.n3993 VSS.n3992 0.00120866
R76324 VSS.n3997 VSS.n3996 0.00120866
R76325 VSS.n4024 VSS.n4023 0.00120866
R76326 VSS.n5841 VSS.n5840 0.00120866
R76327 VSS.n5742 VSS.n5741 0.00120866
R76328 VSS.n5613 VSS.n5612 0.00120866
R76329 VSS.n5609 VSS.n5608 0.00120866
R76330 VSS.n5567 VSS.n5566 0.00120866
R76331 VSS.n5558 VSS.n5557 0.00120866
R76332 VSS.n9536 VSS.n9535 0.00120866
R76333 VSS.n13019 VSS.n13018 0.00120866
R76334 VSS.n13022 VSS.n13021 0.00120866
R76335 VSS.n13051 VSS.n13050 0.00120866
R76336 VSS.n12574 VSS.n12573 0.00120866
R76337 VSS.n12550 VSS.n12549 0.00120866
R76338 VSS.n12294 VSS.n12293 0.00120866
R76339 VSS.n11968 VSS.n11967 0.00120866
R76340 VSS.n11965 VSS.n11964 0.00120866
R76341 VSS.n11880 VSS.n11879 0.00120866
R76342 VSS.n11870 VSS.n11869 0.00120866
R76343 VSS.n18864 VSS.n18863 0.00120866
R76344 VSS.n18868 VSS.n18867 0.00120866
R76345 VSS.n18895 VSS.n18894 0.00120866
R76346 VSS.n16202 VSS.n16201 0.00120866
R76347 VSS.n16190 VSS.n16189 0.00120866
R76348 VSS.n16129 VSS.n16128 0.00120866
R76349 VSS.n16125 VSS.n16124 0.00120866
R76350 VSS.n16083 VSS.n16082 0.00120866
R76351 VSS.n16068 VSS.n16067 0.00120866
R76352 VSS.n9653 VSS.n9652 0.00120866
R76353 VSS.n21792 VSS.n21791 0.00120866
R76354 VSS.n21795 VSS.n21794 0.00120866
R76355 VSS.n21824 VSS.n21823 0.00120866
R76356 VSS.n21144 VSS.n21143 0.00120866
R76357 VSS.n21132 VSS.n21131 0.00120866
R76358 VSS.n21063 VSS.n21062 0.00120866
R76359 VSS.n21059 VSS.n21058 0.00120866
R76360 VSS.n21016 VSS.n21015 0.00120866
R76361 VSS.n21007 VSS.n21006 0.00120866
R76362 VSS.n6942 VSS.n6941 0.00120866
R76363 VSS.n19077 VSS.n19076 0.00120866
R76364 VSS.n19080 VSS.n19079 0.00120866
R76365 VSS.n19109 VSS.n19108 0.00120866
R76366 VSS.n1273 VSS.n1272 0.00120866
R76367 VSS.n1182 VSS.n1181 0.00120866
R76368 VSS.n1109 VSS.n1108 0.00120866
R76369 VSS.n1105 VSS.n1104 0.00120866
R76370 VSS.n1062 VSS.n1061 0.00120866
R76371 VSS.n1053 VSS.n1052 0.00120866
R76372 VSS.n6840 VSS.n6839 0.00120866
R76373 VSS.n21562 VSS.n21561 0.00120866
R76374 VSS.n21566 VSS.n21565 0.00120866
R76375 VSS.n21595 VSS.n21594 0.00120866
R76376 VSS.n21465 VSS.n21464 0.00120866
R76377 VSS.n3794 VSS.n3793 0.00120866
R76378 VSS.n3799 VSS.n3798 0.00120866
R76379 VSS.n3826 VSS.n3825 0.00120866
R76380 VSS.n4770 VSS.n4769 0.00120866
R76381 VSS.n3273 VSS.n3272 0.00120866
R76382 VSS.n3277 VSS.n3276 0.00120866
R76383 VSS.n3245 VSS.n3244 0.00120866
R76384 VSS.n10509 VSS.n10508 0.00120866
R76385 VSS.n10495 VSS.n10494 0.00120866
R76386 VSS.n10242 VSS.n10241 0.00120866
R76387 VSS.n9971 VSS.n9970 0.00120866
R76388 VSS.n9968 VSS.n9967 0.00120866
R76389 VSS.n8942 VSS.n8941 0.00120866
R76390 VSS.n8791 VSS.n8790 0.00120866
R76391 VSS.n2666 VSS.n2665 0.00120714
R76392 VSS.n2710 VSS.n2709 0.00120714
R76393 VSS.n2770 VSS.n2769 0.00120714
R76394 VSS.n2878 VSS.n2877 0.00120714
R76395 VSS.n2956 VSS.n2955 0.00120714
R76396 VSS.n3068 VSS.n3067 0.00120714
R76397 VSS.n2558 VSS.n2557 0.00120714
R76398 VSS.n5213 VSS.n5212 0.00120714
R76399 VSS.n5264 VSS.n5263 0.00120714
R76400 VSS.n5299 VSS.n5298 0.00120714
R76401 VSS.n4956 VSS.n4955 0.00120714
R76402 VSS.n7157 VSS.n7156 0.00120714
R76403 VSS.n7098 VSS.n7097 0.00120714
R76404 VSS.n7061 VSS.n7060 0.00120714
R76405 VSS.n7523 VSS.n7522 0.00120714
R76406 VSS.n4442 VSS.n4441 0.00120714
R76407 VSS.n4391 VSS.n4390 0.00120714
R76408 VSS.n4356 VSS.n4355 0.00120714
R76409 VSS.n4324 VSS.n4323 0.00120714
R76410 VSS.n17559 VSS.n17558 0.00120714
R76411 VSS.n17501 VSS.n17500 0.00120714
R76412 VSS.n18021 VSS.n18020 0.00120714
R76413 VSS.n17855 VSS.n17854 0.00120714
R76414 VSS.n17794 VSS.n17793 0.00120714
R76415 VSS.n17749 VSS.n17748 0.00120714
R76416 VSS.n17716 VSS.n17715 0.00120714
R76417 VSS.n3536 VSS.n3534 0.00120422
R76418 VSS.n3595 VSS.n3593 0.00120422
R76419 VSS.n3638 VSS.n3636 0.00120422
R76420 VSS.n3203 VSS.n3202 0.00120422
R76421 VSS.n3779 VSS.n3778 0.00120422
R76422 VSS.n3537 VSS.n3533 0.00120422
R76423 VSS.n3596 VSS.n3592 0.00120422
R76424 VSS.n3639 VSS.n3635 0.00120422
R76425 VSS.n3661 VSS.n3660 0.00120422
R76426 VSS.n3657 VSS.n3656 0.00120422
R76427 VSS.n20255 VSS.n20254 0.00119
R76428 VSS.n20235 VSS.n20230 0.00119
R76429 VSS.n20256 VSS.n20252 0.00119
R76430 VSS.n20227 VSS.n20226 0.00119
R76431 VSS.n10813 VSS.n10812 0.00119
R76432 VSS.n10841 VSS.n10836 0.00119
R76433 VSS.n8770 VSS.n8769 0.00119
R76434 VSS.n8748 VSS.n8743 0.00119
R76435 VSS.n8438 VSS.n8437 0.00119
R76436 VSS.n8291 VSS.n8286 0.00119
R76437 VSS.n8442 VSS.n8441 0.00119
R76438 VSS.n8295 VSS.n8294 0.00119
R76439 VSS.n8283 VSS.n8282 0.00119
R76440 VSS.n8774 VSS.n8773 0.00119
R76441 VSS.n8752 VSS.n8751 0.00119
R76442 VSS.n8740 VSS.n8739 0.00119
R76443 VSS.n10682 VSS.n10681 0.00119
R76444 VSS.n10744 VSS.n10743 0.00119
R76445 VSS.n10846 VSS.n10845 0.00119
R76446 VSS.n10929 VSS.n10928 0.00119
R76447 VSS.n10996 VSS.n10995 0.00119
R76448 VSS.n20352 VSS.n20351 0.00117999
R76449 VSS.n20213 VSS.n20212 0.00117999
R76450 VSS.n20353 VSS.n20352 0.00117999
R76451 VSS.n8830 VSS.n8829 0.00117999
R76452 VSS.n9443 VSS.n9442 0.00117999
R76453 VSS.n20214 VSS.n20213 0.00117999
R76454 VSS.n9444 VSS.n9443 0.00117999
R76455 VSS.n8841 VSS.n8830 0.00117999
R76456 VSS.n4054 VSS.n4053 0.00117716
R76457 VSS.n4065 VSS.n4064 0.00117716
R76458 VSS.n3978 VSS.n3977 0.00117716
R76459 VSS.n3968 VSS.n3967 0.00117716
R76460 VSS.n3957 VSS.n3956 0.00117716
R76461 VSS.n17446 VSS.n17445 0.00117716
R76462 VSS.n11546 VSS.n11545 0.00117716
R76463 VSS.n11580 VSS.n11579 0.00117716
R76464 VSS.n5721 VSS.n5720 0.00117716
R76465 VSS.n5576 VSS.n5575 0.00117716
R76466 VSS.n9486 VSS.n9485 0.00117716
R76467 VSS.n9497 VSS.n9496 0.00117716
R76468 VSS.n9500 VSS.n9499 0.00117716
R76469 VSS.n9572 VSS.n9571 0.00117716
R76470 VSS.n9027 VSS.n9026 0.00117716
R76471 VSS.n9135 VSS.n9134 0.00117716
R76472 VSS.n9102 VSS.n9101 0.00117716
R76473 VSS.n9083 VSS.n9082 0.00117716
R76474 VSS.n11579 VSS.n11578 0.00117716
R76475 VSS.n11547 VSS.n11546 0.00117716
R76476 VSS.n13083 VSS.n13082 0.00117716
R76477 VSS.n13093 VSS.n13092 0.00117716
R76478 VSS.n13103 VSS.n13102 0.00117716
R76479 VSS.n13112 VSS.n13111 0.00117716
R76480 VSS.n13123 VSS.n13122 0.00117716
R76481 VSS.n13228 VSS.n13227 0.00117716
R76482 VSS.n12955 VSS.n12954 0.00117716
R76483 VSS.n12919 VSS.n12918 0.00117716
R76484 VSS.n12737 VSS.n12736 0.00117716
R76485 VSS.n12702 VSS.n12701 0.00117716
R76486 VSS.n12530 VSS.n12529 0.00117716
R76487 VSS.n12512 VSS.n12511 0.00117716
R76488 VSS.n12309 VSS.n12308 0.00117716
R76489 VSS.n12253 VSS.n12252 0.00117716
R76490 VSS.n12244 VSS.n12243 0.00117716
R76491 VSS.n11898 VSS.n11897 0.00117716
R76492 VSS.n11822 VSS.n11821 0.00117716
R76493 VSS.n12920 VSS.n12919 0.00117716
R76494 VSS.n12956 VSS.n12955 0.00117716
R76495 VSS.n13227 VSS.n13226 0.00117716
R76496 VSS.n17447 VSS.n17446 0.00117716
R76497 VSS.n18925 VSS.n18924 0.00117716
R76498 VSS.n18936 VSS.n18935 0.00117716
R76499 VSS.n18947 VSS.n18946 0.00117716
R76500 VSS.n18957 VSS.n18956 0.00117716
R76501 VSS.n18968 VSS.n18967 0.00117716
R76502 VSS.n2198 VSS.n2197 0.00117716
R76503 VSS.n15021 VSS.n15020 0.00117716
R76504 VSS.n15055 VSS.n15054 0.00117716
R76505 VSS.n16362 VSS.n16361 0.00117716
R76506 VSS.n16317 VSS.n16316 0.00117716
R76507 VSS.n16282 VSS.n16281 0.00117716
R76508 VSS.n16168 VSS.n16167 0.00117716
R76509 VSS.n16092 VSS.n16091 0.00117716
R76510 VSS.n9603 VSS.n9602 0.00117716
R76511 VSS.n9614 VSS.n9613 0.00117716
R76512 VSS.n9617 VSS.n9616 0.00117716
R76513 VSS.n9689 VSS.n9688 0.00117716
R76514 VSS.n9170 VSS.n9169 0.00117716
R76515 VSS.n9298 VSS.n9297 0.00117716
R76516 VSS.n9265 VSS.n9264 0.00117716
R76517 VSS.n9247 VSS.n9246 0.00117716
R76518 VSS.n15054 VSS.n15053 0.00117716
R76519 VSS.n16363 VSS.n16362 0.00117716
R76520 VSS.n16318 VSS.n16317 0.00117716
R76521 VSS.n16283 VSS.n16282 0.00117716
R76522 VSS.n15020 VSS.n15019 0.00117716
R76523 VSS.n2197 VSS.n2196 0.00117716
R76524 VSS.n16169 VSS.n16168 0.00117716
R76525 VSS.n5720 VSS.n5719 0.00117716
R76526 VSS.n5623 VSS.n5622 0.00117716
R76527 VSS.n16145 VSS.n16138 0.00117716
R76528 VSS.n5845 VSS.n5844 0.00117716
R76529 VSS.n16206 VSS.n16205 0.00117716
R76530 VSS.n21856 VSS.n21855 0.00117716
R76531 VSS.n21866 VSS.n21865 0.00117716
R76532 VSS.n21775 VSS.n21774 0.00117716
R76533 VSS.n21766 VSS.n21765 0.00117716
R76534 VSS.n21755 VSS.n21754 0.00117716
R76535 VSS.n13344 VSS.n13343 0.00117716
R76536 VSS.n20629 VSS.n20628 0.00117716
R76537 VSS.n20665 VSS.n20664 0.00117716
R76538 VSS.n21109 VSS.n21108 0.00117716
R76539 VSS.n21024 VSS.n21023 0.00117716
R76540 VSS.n6917 VSS.n6916 0.00117716
R76541 VSS.n6928 VSS.n6927 0.00117716
R76542 VSS.n6931 VSS.n6930 0.00117716
R76543 VSS.n6982 VSS.n6981 0.00117716
R76544 VSS.n6658 VSS.n6657 0.00117716
R76545 VSS.n6622 VSS.n6621 0.00117716
R76546 VSS.n6586 VSS.n6585 0.00117716
R76547 VSS.n6567 VSS.n6566 0.00117716
R76548 VSS.n20664 VSS.n20663 0.00117716
R76549 VSS.n20628 VSS.n20627 0.00117716
R76550 VSS.n13345 VSS.n13344 0.00117716
R76551 VSS.n21148 VSS.n21147 0.00117716
R76552 VSS.n21108 VSS.n21107 0.00117716
R76553 VSS.n21073 VSS.n21072 0.00117716
R76554 VSS.n19141 VSS.n19140 0.00117716
R76555 VSS.n19151 VSS.n19150 0.00117716
R76556 VSS.n19060 VSS.n19059 0.00117716
R76557 VSS.n19051 VSS.n19050 0.00117716
R76558 VSS.n19040 VSS.n19039 0.00117716
R76559 VSS.n13487 VSS.n13486 0.00117716
R76560 VSS.n20120 VSS.n20119 0.00117716
R76561 VSS.n20084 VSS.n20083 0.00117716
R76562 VSS.n1443 VSS.n1442 0.00117716
R76563 VSS.n1398 VSS.n1397 0.00117716
R76564 VSS.n1363 VSS.n1362 0.00117716
R76565 VSS.n1158 VSS.n1157 0.00117716
R76566 VSS.n1070 VSS.n1069 0.00117716
R76567 VSS.n6794 VSS.n6793 0.00117716
R76568 VSS.n6805 VSS.n6804 0.00117716
R76569 VSS.n6808 VSS.n6807 0.00117716
R76570 VSS.n6880 VSS.n6879 0.00117716
R76571 VSS.n6508 VSS.n6507 0.00117716
R76572 VSS.n6472 VSS.n6471 0.00117716
R76573 VSS.n6436 VSS.n6435 0.00117716
R76574 VSS.n6417 VSS.n6416 0.00117716
R76575 VSS.n1159 VSS.n1158 0.00117716
R76576 VSS.n20085 VSS.n20084 0.00117716
R76577 VSS.n20121 VSS.n20120 0.00117716
R76578 VSS.n1364 VSS.n1363 0.00117716
R76579 VSS.n1399 VSS.n1398 0.00117716
R76580 VSS.n1444 VSS.n1443 0.00117716
R76581 VSS.n13488 VSS.n13487 0.00117716
R76582 VSS.n1277 VSS.n1276 0.00117716
R76583 VSS.n1125 VSS.n1118 0.00117716
R76584 VSS.n21629 VSS.n21628 0.00117716
R76585 VSS.n21640 VSS.n21639 0.00117716
R76586 VSS.n21535 VSS.n21534 0.00117716
R76587 VSS.n21372 VSS.n21371 0.00117716
R76588 VSS.n21336 VSS.n21335 0.00117716
R76589 VSS.n7625 VSS.n7624 0.00117716
R76590 VSS.n7661 VSS.n7660 0.00117716
R76591 VSS.n7713 VSS.n7712 0.00117716
R76592 VSS.n7749 VSS.n7748 0.00117716
R76593 VSS.n7826 VSS.n7825 0.00117716
R76594 VSS.n7790 VSS.n7789 0.00117716
R76595 VSS.n21337 VSS.n21336 0.00117716
R76596 VSS.n21373 VSS.n21372 0.00117716
R76597 VSS.n21630 VSS.n21629 0.00117716
R76598 VSS.n21536 VSS.n21535 0.00117716
R76599 VSS.n9266 VSS.n9265 0.00117716
R76600 VSS.n7827 VSS.n7826 0.00117716
R76601 VSS.n11900 VSS.n11899 0.00117716
R76602 VSS.n6623 VSS.n6622 0.00117716
R76603 VSS.n6473 VSS.n6472 0.00117716
R76604 VSS.n9299 VSS.n9298 0.00117716
R76605 VSS.n9136 VSS.n9135 0.00117716
R76606 VSS.n7791 VSS.n7790 0.00117716
R76607 VSS.n6587 VSS.n6586 0.00117716
R76608 VSS.n6437 VSS.n6436 0.00117716
R76609 VSS.n9103 VSS.n9102 0.00117716
R76610 VSS.n9169 VSS.n9168 0.00117716
R76611 VSS.n12531 VSS.n12530 0.00117716
R76612 VSS.n12254 VSS.n12253 0.00117716
R76613 VSS.n7748 VSS.n7747 0.00117716
R76614 VSS.n9026 VSS.n9025 0.00117716
R76615 VSS.n7712 VSS.n7711 0.00117716
R76616 VSS.n12513 VSS.n12512 0.00117716
R76617 VSS.n6983 VSS.n6982 0.00117716
R76618 VSS.n6881 VSS.n6880 0.00117716
R76619 VSS.n9690 VSS.n9689 0.00117716
R76620 VSS.n9573 VSS.n9572 0.00117716
R76621 VSS.n12310 VSS.n12309 0.00117716
R76622 VSS.n12245 VSS.n12244 0.00117716
R76623 VSS.n6657 VSS.n6656 0.00117716
R76624 VSS.n6507 VSS.n6506 0.00117716
R76625 VSS.n6930 VSS.n6929 0.00117716
R76626 VSS.n6807 VSS.n6806 0.00117716
R76627 VSS.n9616 VSS.n9615 0.00117716
R76628 VSS.n9499 VSS.n9498 0.00117716
R76629 VSS.n9485 VSS.n9484 0.00117716
R76630 VSS.n9602 VSS.n9601 0.00117716
R76631 VSS.n6916 VSS.n6915 0.00117716
R76632 VSS.n12703 VSS.n12702 0.00117716
R76633 VSS.n7660 VSS.n7659 0.00117716
R76634 VSS.n6793 VSS.n6792 0.00117716
R76635 VSS.n16093 VSS.n16092 0.00117716
R76636 VSS.n7624 VSS.n7623 0.00117716
R76637 VSS.n12738 VSS.n12737 0.00117716
R76638 VSS.n21025 VSS.n21024 0.00117716
R76639 VSS.n1071 VSS.n1070 0.00117716
R76640 VSS.n5577 VSS.n5576 0.00117716
R76641 VSS.n3857 VSS.n3856 0.00117716
R76642 VSS.n3869 VSS.n3868 0.00117716
R76643 VSS.n4151 VSS.n4150 0.00117716
R76644 VSS.n11688 VSS.n11687 0.00117716
R76645 VSS.n11654 VSS.n11653 0.00117716
R76646 VSS.n6131 VSS.n6130 0.00117716
R76647 VSS.n6098 VSS.n6097 0.00117716
R76648 VSS.n6050 VSS.n6049 0.00117716
R76649 VSS.n6017 VSS.n6016 0.00117716
R76650 VSS.n5969 VSS.n5968 0.00117716
R76651 VSS.n5936 VSS.n5935 0.00117716
R76652 VSS.n11655 VSS.n11654 0.00117716
R76653 VSS.n6099 VSS.n6098 0.00117716
R76654 VSS.n6018 VSS.n6017 0.00117716
R76655 VSS.n5937 VSS.n5936 0.00117716
R76656 VSS.n6051 VSS.n6050 0.00117716
R76657 VSS.n5970 VSS.n5969 0.00117716
R76658 VSS.n11689 VSS.n11688 0.00117716
R76659 VSS.n3858 VSS.n3857 0.00117716
R76660 VSS.n4152 VSS.n4151 0.00117716
R76661 VSS.n6132 VSS.n6131 0.00117716
R76662 VSS.n3958 VSS.n3957 0.00117716
R76663 VSS.n18967 VSS.n18966 0.00117716
R76664 VSS.n19041 VSS.n19040 0.00117716
R76665 VSS.n21756 VSS.n21755 0.00117716
R76666 VSS.n13122 VSS.n13121 0.00117716
R76667 VSS.n4053 VSS.n4052 0.00117716
R76668 VSS.n18924 VSS.n18923 0.00117716
R76669 VSS.n19140 VSS.n19139 0.00117716
R76670 VSS.n21855 VSS.n21854 0.00117716
R76671 VSS.n13082 VSS.n13081 0.00117716
R76672 VSS.n13092 VSS.n13091 0.00117716
R76673 VSS.n19052 VSS.n19051 0.00117716
R76674 VSS.n21767 VSS.n21766 0.00117716
R76675 VSS.n13111 VSS.n13110 0.00117716
R76676 VSS.n21639 VSS.n21638 0.00117716
R76677 VSS.n19150 VSS.n19149 0.00117716
R76678 VSS.n21865 VSS.n21864 0.00117716
R76679 VSS.n4064 VSS.n4063 0.00117716
R76680 VSS.n18935 VSS.n18934 0.00117716
R76681 VSS.n3969 VSS.n3968 0.00117716
R76682 VSS.n18956 VSS.n18955 0.00117716
R76683 VSS.n2634 VSS.n2633 0.00117716
R76684 VSS.n2624 VSS.n2623 0.00117716
R76685 VSS.n2612 VSS.n2611 0.00117716
R76686 VSS.n2603 VSS.n2602 0.00117716
R76687 VSS.n2591 VSS.n2590 0.00117716
R76688 VSS.n2592 VSS.n2591 0.00117716
R76689 VSS.n2635 VSS.n2634 0.00117716
R76690 VSS.n2623 VSS.n2622 0.00117716
R76691 VSS.n2602 VSS.n2601 0.00117716
R76692 VSS.n645 VSS.n644 0.00117716
R76693 VSS.n612 VSS.n611 0.00117716
R76694 VSS.n10603 VSS.n10602 0.00117716
R76695 VSS.n10570 VSS.n10569 0.00117716
R76696 VSS.n10475 VSS.n10474 0.00117716
R76697 VSS.n10458 VSS.n10457 0.00117716
R76698 VSS.n10257 VSS.n10256 0.00117716
R76699 VSS.n10193 VSS.n10192 0.00117716
R76700 VSS.n9899 VSS.n9898 0.00117716
R76701 VSS.n9897 VSS.n9896 0.00117716
R76702 VSS.n8933 VSS.n8932 0.00117716
R76703 VSS.n10476 VSS.n10475 0.00117716
R76704 VSS.n10202 VSS.n10201 0.00117716
R76705 VSS.n10571 VSS.n10570 0.00117716
R76706 VSS.n10194 VSS.n10193 0.00117716
R76707 VSS.n9898 VSS.n9897 0.00117716
R76708 VSS.n9900 VSS.n9899 0.00117716
R76709 VSS.n613 VSS.n612 0.00117716
R76710 VSS.n646 VSS.n645 0.00117716
R76711 VSS.n10604 VSS.n10603 0.00117716
R76712 VSS.n8932 VSS.n8931 0.00117716
R76713 VSS.n9496 VSS.n9495 0.00117716
R76714 VSS.n6804 VSS.n6803 0.00117716
R76715 VSS.n6927 VSS.n6926 0.00117716
R76716 VSS.n9613 VSS.n9612 0.00117716
R76717 VSS.n6418 VSS.n6417 0.00117716
R76718 VSS.n9084 VSS.n9083 0.00117716
R76719 VSS.n9248 VSS.n9247 0.00117716
R76720 VSS.n6568 VSS.n6567 0.00117716
R76721 VSS.n3979 VSS.n3978 0.00117716
R76722 VSS.n2613 VSS.n2612 0.00117716
R76723 VSS.n3868 VSS.n3867 0.00117716
R76724 VSS.n18946 VSS.n18945 0.00117716
R76725 VSS.n13102 VSS.n13101 0.00117716
R76726 VSS.n21776 VSS.n21775 0.00117716
R76727 VSS.n19061 VSS.n19060 0.00117716
R76728 VSS.n17110 VSS.n17109 0.001175
R76729 VSS.n17050 VSS.n17049 0.001175
R76730 VSS.n16952 VSS.n16951 0.001175
R76731 VSS.n14911 VSS.n14910 0.001175
R76732 VSS.n719 VSS.n718 0.00116499
R76733 VSS.n20557 VSS.n20556 0.00116499
R76734 VSS.n20528 VSS.n20527 0.00116499
R76735 VSS.n20558 VSS.n20557 0.00116499
R76736 VSS.n720 VSS.n719 0.00116499
R76737 VSS.n20529 VSS.n20528 0.00116499
R76738 VSS.n10952 VSS.n10951 0.00116499
R76739 VSS.n11069 VSS.n11068 0.00116499
R76740 VSS.n11068 VSS.n11067 0.00116499
R76741 VSS.n10951 VSS.n10950 0.00116499
R76742 VSS.n2829 VSS.n2828 0.00116071
R76743 VSS.n2851 VSS.n2850 0.00116071
R76744 VSS.n2828 VSS.n2827 0.00116071
R76745 VSS.n2850 VSS.n2849 0.00116071
R76746 VSS.n20239 VSS.n20238 0.00116
R76747 VSS.n9394 VSS.n9393 0.00116
R76748 VSS.n9340 VSS.n9339 0.00116
R76749 VSS.n8298 VSS.n8297 0.00116
R76750 VSS.n9785 VSS.n9784 0.00116
R76751 VSS.n9731 VSS.n9730 0.00116
R76752 VSS.n8755 VSS.n8754 0.00116
R76753 VSS.n10679 VSS.n10675 0.00116
R76754 VSS.n10741 VSS.n10737 0.00116
R76755 VSS.n10937 VSS.n10936 0.00116
R76756 VSS.n10940 VSS.n10939 0.00116
R76757 VSS.n11004 VSS.n11003 0.00116
R76758 VSS.n11008 VSS.n11007 0.00116
R76759 VSS.n13941 VSS.n13615 0.00114286
R76760 VSS.n13942 VSS.n13612 0.00114286
R76761 VSS.n2950 VSS.n2948 0.00114286
R76762 VSS.n2549 VSS.n2548 0.00114286
R76763 VSS.n2534 VSS.n2533 0.00114286
R76764 VSS.n2951 VSS.n2947 0.00114286
R76765 VSS.n2953 VSS.n2952 0.00114286
R76766 VSS.n3015 VSS.n3012 0.00114286
R76767 VSS.n3017 VSS.n3016 0.00114286
R76768 VSS.n3063 VSS.n3060 0.00114286
R76769 VSS.n3065 VSS.n3064 0.00114286
R76770 VSS.n2565 VSS.n2564 0.00114286
R76771 VSS.n2561 VSS.n2560 0.00114286
R76772 VSS.n5209 VSS.n5207 0.00114286
R76773 VSS.n5260 VSS.n5258 0.00114286
R76774 VSS.n5295 VSS.n5293 0.00114286
R76775 VSS.n4951 VSS.n4950 0.00114286
R76776 VSS.n5210 VSS.n5206 0.00114286
R76777 VSS.n5261 VSS.n5257 0.00114286
R76778 VSS.n5296 VSS.n5292 0.00114286
R76779 VSS.n4959 VSS.n4958 0.00114286
R76780 VSS.n7162 VSS.n7160 0.00114286
R76781 VSS.n7103 VSS.n7101 0.00114286
R76782 VSS.n7066 VSS.n7063 0.00114286
R76783 VSS.n7528 VSS.n7525 0.00114286
R76784 VSS.n7164 VSS.n7163 0.00114286
R76785 VSS.n7105 VSS.n7104 0.00114286
R76786 VSS.n7068 VSS.n7067 0.00114286
R76787 VSS.n7530 VSS.n7529 0.00114286
R76788 VSS.n4446 VSS.n4444 0.00114286
R76789 VSS.n4395 VSS.n4393 0.00114286
R76790 VSS.n4360 VSS.n4358 0.00114286
R76791 VSS.n4315 VSS.n4314 0.00114286
R76792 VSS.n4694 VSS.n4693 0.00114286
R76793 VSS.n4448 VSS.n4447 0.00114286
R76794 VSS.n4397 VSS.n4396 0.00114286
R76795 VSS.n4362 VSS.n4361 0.00114286
R76796 VSS.n4331 VSS.n4330 0.00114286
R76797 VSS.n4327 VSS.n4326 0.00114286
R76798 VSS.n4745 VSS.n4744 0.00114286
R76799 VSS.n17862 VSS.n17861 0.00114286
R76800 VSS.n17857 VSS.n17856 0.00114286
R76801 VSS.n17801 VSS.n17800 0.00114286
R76802 VSS.n17796 VSS.n17795 0.00114286
R76803 VSS.n17756 VSS.n17755 0.00114286
R76804 VSS.n17751 VSS.n17750 0.00114286
R76805 VSS.n17723 VSS.n17722 0.00114286
R76806 VSS.n17719 VSS.n17718 0.00114286
R76807 VSS.n17860 VSS.n17858 0.00114286
R76808 VSS.n17799 VSS.n17797 0.00114286
R76809 VSS.n17754 VSS.n17752 0.00114286
R76810 VSS.n17705 VSS.n17704 0.00114286
R76811 VSS.n14128 VSS.n14127 0.00114286
R76812 VSS.n6205 VSS.n6180 0.00114
R76813 VSS.n6245 VSS.n6220 0.00114
R76814 VSS.n11165 VSS.n11164 0.00114
R76815 VSS.n18699 VSS.n18698 0.0011338
R76816 VSS.n18747 VSS.n18746 0.0011338
R76817 VSS.n18753 VSS.n18752 0.0011338
R76818 VSS.n18403 VSS.n18402 0.0011338
R76819 VSS.n18170 VSS.n18169 0.0011338
R76820 VSS.n17080 VSS.n17079 0.0011338
R76821 VSS.n17017 VSS.n17016 0.0011338
R76822 VSS.n14868 VSS.n14867 0.0011338
R76823 VSS.n16920 VSS.n16919 0.0011338
R76824 VSS.n16915 VSS.n16914 0.0011338
R76825 VSS.n16910 VSS.n16909 0.0011338
R76826 VSS.n16901 VSS.n16900 0.0011338
R76827 VSS.n16634 VSS.n16633 0.0011338
R76828 VSS.n16631 VSS.n16630 0.0011338
R76829 VSS.n16587 VSS.n16586 0.0011338
R76830 VSS.n14983 VSS.n14982 0.0011338
R76831 VSS.n14991 VSS.n14990 0.0011338
R76832 VSS.n15452 VSS.n15451 0.0011338
R76833 VSS.n15376 VSS.n15375 0.0011338
R76834 VSS.n19181 VSS.n19180 0.0011338
R76835 VSS.n19229 VSS.n19228 0.0011338
R76836 VSS.n19235 VSS.n19234 0.0011338
R76837 VSS.n19619 VSS.n19618 0.0011338
R76838 VSS.n19686 VSS.n19685 0.0011338
R76839 VSS.n19885 VSS.n19884 0.0011338
R76840 VSS.n19918 VSS.n19917 0.0011338
R76841 VSS.n19939 VSS.n19938 0.0011338
R76842 VSS.n19996 VSS.n19995 0.0011338
R76843 VSS.n20001 VSS.n20000 0.0011338
R76844 VSS.n20006 VSS.n20005 0.0011338
R76845 VSS.n20015 VSS.n20014 0.0011338
R76846 VSS.n764 VSS.n763 0.0011338
R76847 VSS.n767 VSS.n766 0.0011338
R76848 VSS.n781 VSS.n780 0.0011338
R76849 VSS.n819 VSS.n818 0.0011338
R76850 VSS.n827 VSS.n826 0.0011338
R76851 VSS.n1754 VSS.n1753 0.0011338
R76852 VSS.n1692 VSS.n1691 0.0011338
R76853 VSS.n20209 VSS.n20207 0.00113
R76854 VSS.n20242 VSS.n20241 0.00113
R76855 VSS.n20211 VSS.n20210 0.00113
R76856 VSS.n10867 VSS.n10865 0.00113
R76857 VSS.n8601 VSS.n8599 0.00113
R76858 VSS.n8264 VSS.n8262 0.00113
R76859 VSS.n8992 VSS.n8927 0.00113
R76860 VSS.n8259 VSS.n8258 0.00113
R76861 VSS.n7886 VSS.n7885 0.00113
R76862 VSS.n9462 VSS.n9461 0.00113
R76863 VSS.n8596 VSS.n8595 0.00113
R76864 VSS.n7979 VSS.n7978 0.00113
R76865 VSS.n10635 VSS.n10634 0.00113
R76866 VSS.n10671 VSS.n10670 0.00113
R76867 VSS.n10674 VSS.n10673 0.00113
R76868 VSS.n10733 VSS.n10732 0.00113
R76869 VSS.n10736 VSS.n10735 0.00113
R76870 VSS.n11049 VSS.n11048 0.00113
R76871 VSS.n168 VSS.n167 0.00112569
R76872 VSS.n5902 VSS.n5901 0.00112569
R76873 VSS.n169 VSS.n168 0.00112569
R76874 VSS.n5901 VSS.n5900 0.00112569
R76875 VSS.n18719 VSS.n18718 0.00110563
R76876 VSS.n18750 VSS.n18749 0.00110563
R76877 VSS.n18817 VSS.n18816 0.00110563
R76878 VSS.n18153 VSS.n18152 0.00110563
R76879 VSS.n14881 VSS.n14880 0.00110563
R76880 VSS.n16922 VSS.n16921 0.00110563
R76881 VSS.n15634 VSS.n15633 0.00110563
R76882 VSS.n15611 VSS.n15610 0.00110563
R76883 VSS.n15588 VSS.n15587 0.00110563
R76884 VSS.n15471 VSS.n15470 0.00110563
R76885 VSS.n15413 VSS.n15412 0.00110563
R76886 VSS.n15379 VSS.n15378 0.00110563
R76887 VSS.n8464 VSS.n8463 0.00110563
R76888 VSS.n8545 VSS.n8544 0.00110563
R76889 VSS.n8312 VSS.n8311 0.00110563
R76890 VSS.n8400 VSS.n8399 0.00110563
R76891 VSS.n8376 VSS.n8375 0.00110563
R76892 VSS.n14880 VSS.n14879 0.00110563
R76893 VSS.n17085 VSS.n17084 0.00110563
R76894 VSS.n16923 VSS.n16922 0.00110563
R76895 VSS.n15635 VSS.n15634 0.00110563
R76896 VSS.n15612 VSS.n15611 0.00110563
R76897 VSS.n15589 VSS.n15588 0.00110563
R76898 VSS.n18816 VSS.n18815 0.00110563
R76899 VSS.n18718 VSS.n18717 0.00110563
R76900 VSS.n18154 VSS.n18153 0.00110563
R76901 VSS.n15414 VSS.n15413 0.00110563
R76902 VSS.n15380 VSS.n15379 0.00110563
R76903 VSS.n15470 VSS.n15469 0.00110563
R76904 VSS.n8401 VSS.n8400 0.00110563
R76905 VSS.n8377 VSS.n8376 0.00110563
R76906 VSS.n8546 VSS.n8545 0.00110563
R76907 VSS.n8311 VSS.n8310 0.00110563
R76908 VSS.n8463 VSS.n8462 0.00110563
R76909 VSS.n15343 VSS.n15342 0.00110563
R76910 VSS.n19201 VSS.n19200 0.00110563
R76911 VSS.n19488 VSS.n19487 0.00110563
R76912 VSS.n19703 VSS.n19702 0.00110563
R76913 VSS.n19952 VSS.n19951 0.00110563
R76914 VSS.n19994 VSS.n19993 0.00110563
R76915 VSS.n1902 VSS.n1901 0.00110563
R76916 VSS.n1885 VSS.n1884 0.00110563
R76917 VSS.n1868 VSS.n1867 0.00110563
R76918 VSS.n1772 VSS.n1771 0.00110563
R76919 VSS.n1729 VSS.n1728 0.00110563
R76920 VSS.n1696 VSS.n1695 0.00110563
R76921 VSS.n8615 VSS.n8614 0.00110563
R76922 VSS.n8696 VSS.n8695 0.00110563
R76923 VSS.n8108 VSS.n8107 0.00110563
R76924 VSS.n8208 VSS.n8207 0.00110563
R76925 VSS.n8184 VSS.n8183 0.00110563
R76926 VSS.n8697 VSS.n8696 0.00110563
R76927 VSS.n8209 VSS.n8208 0.00110563
R76928 VSS.n8107 VSS.n8106 0.00110563
R76929 VSS.n8185 VSS.n8184 0.00110563
R76930 VSS.n8614 VSS.n8613 0.00110563
R76931 VSS.n1773 VSS.n1772 0.00110563
R76932 VSS.n19993 VSS.n19992 0.00110563
R76933 VSS.n19951 VSS.n19950 0.00110563
R76934 VSS.n19880 VSS.n19879 0.00110563
R76935 VSS.n1903 VSS.n1902 0.00110563
R76936 VSS.n1886 VSS.n1885 0.00110563
R76937 VSS.n1869 VSS.n1868 0.00110563
R76938 VSS.n19232 VSS.n19231 0.00110563
R76939 VSS.n19200 VSS.n19199 0.00110563
R76940 VSS.n19489 VSS.n19488 0.00110563
R76941 VSS.n19702 VSS.n19701 0.00110563
R76942 VSS.n1730 VSS.n1729 0.00110563
R76943 VSS.n1695 VSS.n1694 0.00110563
R76944 VSS.n1659 VSS.n1658 0.00110563
R76945 VSS.n8261 VSS.n8260 0.001105
R76946 VSS.n8598 VSS.n8597 0.001105
R76947 VSS.n10871 VSS.n10870 0.001105
R76948 VSS.n8597 VSS.n8596 0.001105
R76949 VSS.n8260 VSS.n8259 0.001105
R76950 VSS.n10872 VSS.n10871 0.001105
R76951 VSS.n10808 VSS.n10807 0.0011
R76952 VSS.n10833 VSS.n10832 0.0011
R76953 VSS.n10849 VSS.n10848 0.0011
R76954 VSS.n10873 VSS.n10872 0.0011
R76955 VSS.n2676 VSS.n2675 0.00109643
R76956 VSS.n2719 VSS.n2718 0.00109643
R76957 VSS.n2780 VSS.n2779 0.00109643
R76958 VSS.n2870 VSS.n2869 0.00109643
R76959 VSS.n2720 VSS.n2719 0.00109643
R76960 VSS.n2779 VSS.n2778 0.00109643
R76961 VSS.n2869 VSS.n2868 0.00109643
R76962 VSS.n2675 VSS.n2674 0.00109643
R76963 VSS.n4005 VSS.n4004 0.00108858
R76964 VSS.n4058 VSS.n4057 0.00108858
R76965 VSS.n4068 VSS.n4067 0.00108858
R76966 VSS.n3974 VSS.n3973 0.00108858
R76967 VSS.n3964 VSS.n3963 0.00108858
R76968 VSS.n11553 VSS.n11552 0.00108858
R76969 VSS.n11573 VSS.n11572 0.00108858
R76970 VSS.n11574 VSS.n11573 0.00108858
R76971 VSS.n11552 VSS.n11551 0.00108858
R76972 VSS.n3963 VSS.n3962 0.00108858
R76973 VSS.n4069 VSS.n4068 0.00108858
R76974 VSS.n4057 VSS.n4056 0.00108858
R76975 VSS.n4006 VSS.n4005 0.00108858
R76976 VSS.n13217 VSS.n13216 0.00108858
R76977 VSS.n12731 VSS.n12730 0.00108858
R76978 VSS.n13216 VSS.n13215 0.00108858
R76979 VSS.n9254 VSS.n9253 0.00108858
R76980 VSS.n6573 VSS.n6572 0.00108858
R76981 VSS.n6423 VSS.n6422 0.00108858
R76982 VSS.n9253 VSS.n9252 0.00108858
R76983 VSS.n12732 VSS.n12731 0.00108858
R76984 VSS.n2608 VSS.n2607 0.00108858
R76985 VSS.n2597 VSS.n2596 0.00108858
R76986 VSS.n2598 VSS.n2597 0.00108858
R76987 VSS.n4048 VSS.n4047 0.00108858
R76988 VSS.n17475 VSS.n17474 0.00108858
R76989 VSS.n17466 VSS.n17465 0.00108858
R76990 VSS.n17457 VSS.n17456 0.00108858
R76991 VSS.n17453 VSS.n17452 0.00108858
R76992 VSS.n17443 VSS.n17442 0.00108858
R76993 VSS.n17434 VSS.n17433 0.00108858
R76994 VSS.n5636 VSS.n5635 0.00108858
R76995 VSS.n9480 VSS.n9479 0.00108858
R76996 VSS.n9566 VSS.n9565 0.00108858
R76997 VSS.n9021 VSS.n9020 0.00108858
R76998 VSS.n9129 VSS.n9128 0.00108858
R76999 VSS.n9108 VSS.n9107 0.00108858
R77000 VSS.n9089 VSS.n9088 0.00108858
R77001 VSS.n4047 VSS.n4046 0.00108858
R77002 VSS.n17458 VSS.n17457 0.00108858
R77003 VSS.n13031 VSS.n13030 0.00108858
R77004 VSS.n13077 VSS.n13076 0.00108858
R77005 VSS.n13107 VSS.n13106 0.00108858
R77006 VSS.n13230 VSS.n13229 0.00108858
R77007 VSS.n13238 VSS.n13237 0.00108858
R77008 VSS.n12949 VSS.n12948 0.00108858
R77009 VSS.n12925 VSS.n12924 0.00108858
R77010 VSS.n12708 VSS.n12707 0.00108858
R77011 VSS.n12523 VSS.n12522 0.00108858
R77012 VSS.n12320 VSS.n12319 0.00108858
R77013 VSS.n11921 VSS.n11920 0.00108858
R77014 VSS.n11885 VSS.n11884 0.00108858
R77015 VSS.n11837 VSS.n11836 0.00108858
R77016 VSS.n12950 VSS.n12949 0.00108858
R77017 VSS.n12926 VSS.n12925 0.00108858
R77018 VSS.n13086 VSS.n13085 0.00108858
R77019 VSS.n13096 VSS.n13095 0.00108858
R77020 VSS.n13076 VSS.n13075 0.00108858
R77021 VSS.n13030 VSS.n13029 0.00108858
R77022 VSS.n13116 VSS.n13115 0.00108858
R77023 VSS.n17435 VSS.n17434 0.00108858
R77024 VSS.n13208 VSS.n13207 0.00108858
R77025 VSS.n17476 VSS.n17475 0.00108858
R77026 VSS.n13199 VSS.n13198 0.00108858
R77027 VSS.n17467 VSS.n17466 0.00108858
R77028 VSS.n17454 VSS.n17453 0.00108858
R77029 VSS.n13221 VSS.n13220 0.00108858
R77030 VSS.n17444 VSS.n17443 0.00108858
R77031 VSS.n18877 VSS.n18876 0.00108858
R77032 VSS.n18919 VSS.n18918 0.00108858
R77033 VSS.n18929 VSS.n18928 0.00108858
R77034 VSS.n18940 VSS.n18939 0.00108858
R77035 VSS.n18952 VSS.n18951 0.00108858
R77036 VSS.n18962 VSS.n18961 0.00108858
R77037 VSS.n2226 VSS.n2225 0.00108858
R77038 VSS.n2217 VSS.n2216 0.00108858
R77039 VSS.n2208 VSS.n2207 0.00108858
R77040 VSS.n2204 VSS.n2203 0.00108858
R77041 VSS.n2194 VSS.n2193 0.00108858
R77042 VSS.n2185 VSS.n2184 0.00108858
R77043 VSS.n15027 VSS.n15026 0.00108858
R77044 VSS.n15049 VSS.n15048 0.00108858
R77045 VSS.n16324 VSS.n16323 0.00108858
R77046 VSS.n16289 VSS.n16288 0.00108858
R77047 VSS.n16253 VSS.n16252 0.00108858
R77048 VSS.n16158 VSS.n16157 0.00108858
R77049 VSS.n9597 VSS.n9596 0.00108858
R77050 VSS.n9683 VSS.n9682 0.00108858
R77051 VSS.n9164 VSS.n9163 0.00108858
R77052 VSS.n9292 VSS.n9291 0.00108858
R77053 VSS.n9271 VSS.n9270 0.00108858
R77054 VSS.n2186 VSS.n2185 0.00108858
R77055 VSS.n15026 VSS.n15025 0.00108858
R77056 VSS.n15048 VSS.n15047 0.00108858
R77057 VSS.n16325 VSS.n16324 0.00108858
R77058 VSS.n16290 VSS.n16289 0.00108858
R77059 VSS.n16254 VSS.n16253 0.00108858
R77060 VSS.n18961 VSS.n18960 0.00108858
R77061 VSS.n18951 VSS.n18950 0.00108858
R77062 VSS.n18939 VSS.n18938 0.00108858
R77063 VSS.n18918 VSS.n18917 0.00108858
R77064 VSS.n18876 VSS.n18875 0.00108858
R77065 VSS.n18928 VSS.n18927 0.00108858
R77066 VSS.n2227 VSS.n2226 0.00108858
R77067 VSS.n2218 VSS.n2217 0.00108858
R77068 VSS.n2209 VSS.n2208 0.00108858
R77069 VSS.n2205 VSS.n2204 0.00108858
R77070 VSS.n2195 VSS.n2194 0.00108858
R77071 VSS.n5637 VSS.n5636 0.00108858
R77072 VSS.n16159 VSS.n16158 0.00108858
R77073 VSS.n16121 VSS.n16120 0.00108858
R77074 VSS.n5605 VSS.n5604 0.00108858
R77075 VSS.n5745 VSS.n5744 0.00108858
R77076 VSS.n16193 VSS.n16192 0.00108858
R77077 VSS.n21804 VSS.n21803 0.00108858
R77078 VSS.n21850 VSS.n21849 0.00108858
R77079 VSS.n13334 VSS.n13333 0.00108858
R77080 VSS.n13347 VSS.n13346 0.00108858
R77081 VSS.n20635 VSS.n20634 0.00108858
R77082 VSS.n20659 VSS.n20658 0.00108858
R77083 VSS.n21135 VSS.n21134 0.00108858
R77084 VSS.n21086 VSS.n21085 0.00108858
R77085 VSS.n6911 VSS.n6910 0.00108858
R77086 VSS.n6976 VSS.n6975 0.00108858
R77087 VSS.n6652 VSS.n6651 0.00108858
R77088 VSS.n6616 VSS.n6615 0.00108858
R77089 VSS.n6592 VSS.n6591 0.00108858
R77090 VSS.n21055 VSS.n21054 0.00108858
R77091 VSS.n13355 VSS.n13354 0.00108858
R77092 VSS.n20634 VSS.n20633 0.00108858
R77093 VSS.n20658 VSS.n20657 0.00108858
R77094 VSS.n13333 VSS.n13332 0.00108858
R77095 VSS.n13325 VSS.n13324 0.00108858
R77096 VSS.n21869 VSS.n21868 0.00108858
R77097 VSS.n21849 VSS.n21848 0.00108858
R77098 VSS.n21803 VSS.n21802 0.00108858
R77099 VSS.n21762 VSS.n21761 0.00108858
R77100 VSS.n21859 VSS.n21858 0.00108858
R77101 VSS.n13316 VSS.n13315 0.00108858
R77102 VSS.n13338 VSS.n13337 0.00108858
R77103 VSS.n21087 VSS.n21086 0.00108858
R77104 VSS.n19089 VSS.n19088 0.00108858
R77105 VSS.n19135 VSS.n19134 0.00108858
R77106 VSS.n13477 VSS.n13476 0.00108858
R77107 VSS.n13490 VSS.n13489 0.00108858
R77108 VSS.n20114 VSS.n20113 0.00108858
R77109 VSS.n20090 VSS.n20089 0.00108858
R77110 VSS.n1405 VSS.n1404 0.00108858
R77111 VSS.n1370 VSS.n1369 0.00108858
R77112 VSS.n1334 VSS.n1333 0.00108858
R77113 VSS.n1138 VSS.n1137 0.00108858
R77114 VSS.n6788 VSS.n6787 0.00108858
R77115 VSS.n6874 VSS.n6873 0.00108858
R77116 VSS.n6502 VSS.n6501 0.00108858
R77117 VSS.n6466 VSS.n6465 0.00108858
R77118 VSS.n6442 VSS.n6441 0.00108858
R77119 VSS.n1185 VSS.n1184 0.00108858
R77120 VSS.n20115 VSS.n20114 0.00108858
R77121 VSS.n20091 VSS.n20090 0.00108858
R77122 VSS.n13498 VSS.n13497 0.00108858
R77123 VSS.n1406 VSS.n1405 0.00108858
R77124 VSS.n1371 VSS.n1370 0.00108858
R77125 VSS.n1335 VSS.n1334 0.00108858
R77126 VSS.n13476 VSS.n13475 0.00108858
R77127 VSS.n19088 VSS.n19087 0.00108858
R77128 VSS.n19134 VSS.n19133 0.00108858
R77129 VSS.n19144 VSS.n19143 0.00108858
R77130 VSS.n19154 VSS.n19153 0.00108858
R77131 VSS.n19047 VSS.n19046 0.00108858
R77132 VSS.n17952 VSS.n17951 0.00108858
R77133 VSS.n17943 VSS.n17942 0.00108858
R77134 VSS.n13481 VSS.n13480 0.00108858
R77135 VSS.n1139 VSS.n1138 0.00108858
R77136 VSS.n1101 VSS.n1100 0.00108858
R77137 VSS.n21575 VSS.n21574 0.00108858
R77138 VSS.n21540 VSS.n21539 0.00108858
R77139 VSS.n21532 VSS.n21531 0.00108858
R77140 VSS.n21454 VSS.n21453 0.00108858
R77141 VSS.n21451 VSS.n21450 0.00108858
R77142 VSS.n21366 VSS.n21365 0.00108858
R77143 VSS.n21342 VSS.n21341 0.00108858
R77144 VSS.n7631 VSS.n7630 0.00108858
R77145 VSS.n7655 VSS.n7654 0.00108858
R77146 VSS.n7719 VSS.n7718 0.00108858
R77147 VSS.n7743 VSS.n7742 0.00108858
R77148 VSS.n7820 VSS.n7819 0.00108858
R77149 VSS.n7796 VSS.n7795 0.00108858
R77150 VSS.n21367 VSS.n21366 0.00108858
R77151 VSS.n21343 VSS.n21342 0.00108858
R77152 VSS.n21450 VSS.n21449 0.00108858
R77153 VSS.n21541 VSS.n21540 0.00108858
R77154 VSS.n21574 VSS.n21573 0.00108858
R77155 VSS.n21634 VSS.n21633 0.00108858
R77156 VSS.n21533 VSS.n21532 0.00108858
R77157 VSS.n9090 VSS.n9089 0.00108858
R77158 VSS.n9293 VSS.n9292 0.00108858
R77159 VSS.n7821 VSS.n7820 0.00108858
R77160 VSS.n9130 VSS.n9129 0.00108858
R77161 VSS.n11920 VSS.n11919 0.00108858
R77162 VSS.n7797 VSS.n7796 0.00108858
R77163 VSS.n11838 VSS.n11837 0.00108858
R77164 VSS.n6593 VSS.n6592 0.00108858
R77165 VSS.n6617 VSS.n6616 0.00108858
R77166 VSS.n6443 VSS.n6442 0.00108858
R77167 VSS.n6467 VSS.n6466 0.00108858
R77168 VSS.n9272 VSS.n9271 0.00108858
R77169 VSS.n9109 VSS.n9108 0.00108858
R77170 VSS.n9684 VSS.n9683 0.00108858
R77171 VSS.n12321 VSS.n12320 0.00108858
R77172 VSS.n7718 VSS.n7717 0.00108858
R77173 VSS.n9567 VSS.n9566 0.00108858
R77174 VSS.n12524 VSS.n12523 0.00108858
R77175 VSS.n7742 VSS.n7741 0.00108858
R77176 VSS.n12269 VSS.n12268 0.00108858
R77177 VSS.n6651 VSS.n6650 0.00108858
R77178 VSS.n6501 VSS.n6500 0.00108858
R77179 VSS.n9163 VSS.n9162 0.00108858
R77180 VSS.n9020 VSS.n9019 0.00108858
R77181 VSS.n6977 VSS.n6976 0.00108858
R77182 VSS.n6875 VSS.n6874 0.00108858
R77183 VSS.n7654 VSS.n7653 0.00108858
R77184 VSS.n12709 VSS.n12708 0.00108858
R77185 VSS.n6910 VSS.n6909 0.00108858
R77186 VSS.n6787 VSS.n6786 0.00108858
R77187 VSS.n9596 VSS.n9595 0.00108858
R77188 VSS.n9479 VSS.n9478 0.00108858
R77189 VSS.n7630 VSS.n7629 0.00108858
R77190 VSS.n3808 VSS.n3807 0.00108858
R77191 VSS.n3863 VSS.n3862 0.00108858
R77192 VSS.n4156 VSS.n4155 0.00108858
R77193 VSS.n4149 VSS.n4148 0.00108858
R77194 VSS.n4785 VSS.n4784 0.00108858
R77195 VSS.n11682 VSS.n11681 0.00108858
R77196 VSS.n11660 VSS.n11659 0.00108858
R77197 VSS.n6125 VSS.n6124 0.00108858
R77198 VSS.n6104 VSS.n6103 0.00108858
R77199 VSS.n6044 VSS.n6043 0.00108858
R77200 VSS.n6023 VSS.n6022 0.00108858
R77201 VSS.n5963 VSS.n5962 0.00108858
R77202 VSS.n5942 VSS.n5941 0.00108858
R77203 VSS.n3862 VSS.n3861 0.00108858
R77204 VSS.n4157 VSS.n4156 0.00108858
R77205 VSS.n11683 VSS.n11682 0.00108858
R77206 VSS.n6126 VSS.n6125 0.00108858
R77207 VSS.n6045 VSS.n6044 0.00108858
R77208 VSS.n5964 VSS.n5963 0.00108858
R77209 VSS.n6024 VSS.n6023 0.00108858
R77210 VSS.n5943 VSS.n5942 0.00108858
R77211 VSS.n6105 VSS.n6104 0.00108858
R77212 VSS.n11661 VSS.n11660 0.00108858
R77213 VSS.n3807 VSS.n3806 0.00108858
R77214 VSS.n4781 VSS.n4780 0.00108858
R77215 VSS.n4784 VSS.n4783 0.00108858
R77216 VSS.n3286 VSS.n3285 0.00108858
R77217 VSS.n2640 VSS.n2639 0.00108858
R77218 VSS.n2630 VSS.n2629 0.00108858
R77219 VSS.n2619 VSS.n2618 0.00108858
R77220 VSS.n2620 VSS.n2619 0.00108858
R77221 VSS.n2641 VSS.n2640 0.00108858
R77222 VSS.n3285 VSS.n3284 0.00108858
R77223 VSS.n2631 VSS.n2630 0.00108858
R77224 VSS.n639 VSS.n638 0.00108858
R77225 VSS.n618 VSS.n617 0.00108858
R77226 VSS.n10597 VSS.n10596 0.00108858
R77227 VSS.n10576 VSS.n10575 0.00108858
R77228 VSS.n10468 VSS.n10467 0.00108858
R77229 VSS.n10217 VSS.n10216 0.00108858
R77230 VSS.n9922 VSS.n9921 0.00108858
R77231 VSS.n8947 VSS.n8946 0.00108858
R77232 VSS.n8910 VSS.n8909 0.00108858
R77233 VSS.n10267 VSS.n10266 0.00108858
R77234 VSS.n8948 VSS.n8947 0.00108858
R77235 VSS.n10469 VSS.n10468 0.00108858
R77236 VSS.n10218 VSS.n10217 0.00108858
R77237 VSS.n9921 VSS.n9920 0.00108858
R77238 VSS.n10577 VSS.n10576 0.00108858
R77239 VSS.n10598 VSS.n10597 0.00108858
R77240 VSS.n640 VSS.n639 0.00108858
R77241 VSS.n619 VSS.n618 0.00108858
R77242 VSS.n11080 DVSS 0.00108667
R77243 VSS.n14209 VSS.n14208 0.00107857
R77244 VSS.n14131 VSS.n13945 0.00107857
R77245 VSS.n10306 VSS.n10305 0.00107692
R77246 VSS.n10424 VSS.n10423 0.00107692
R77247 VSS.n10139 VSS.n10138 0.00107692
R77248 VSS.n10047 VSS.n10046 0.00107692
R77249 VSS.n10038 VSS.n10033 0.00107692
R77250 VSS.n12360 VSS.n12359 0.00107692
R77251 VSS.n12478 VSS.n12477 0.00107692
R77252 VSS.n12190 VSS.n12189 0.00107692
R77253 VSS.n12098 VSS.n12097 0.00107692
R77254 VSS.n12089 VSS.n12084 0.00107692
R77255 VSS.n8297 VSS.n8296 0.001075
R77256 VSS.n8296 VSS.n8295 0.001075
R77257 VSS.n8754 VSS.n8753 0.001075
R77258 VSS.n8753 VSS.n8752 0.001075
R77259 VSS.n10831 VSS.n10830 0.001075
R77260 VSS.n10832 VSS.n10831 0.001075
R77261 VSS.n8293 VSS.n8292 0.00107
R77262 VSS.n8750 VSS.n8749 0.00107
R77263 VSS.n10829 VSS.n10828 0.00107
R77264 VSS.n10842 VSS.n10835 0.00107
R77265 VSS.n10852 VSS.n10851 0.00107
R77266 VSS.n2512 VSS.n2511 0.00106944
R77267 VSS.n5476 VSS.n5475 0.00106944
R77268 VSS.n4921 VSS.n4920 0.00106944
R77269 VSS.n4857 VSS.n4856 0.00106944
R77270 VSS.n14292 VSS.n14291 0.00106944
R77271 VSS.n17309 VSS.n17308 0.00106944
R77272 VSS.n2427 VSS.n2426 0.00106944
R77273 VSS.n2426 VSS.n2425 0.00106944
R77274 VSS.n17308 VSS.n17307 0.00106944
R77275 VSS.n14293 VSS.n14292 0.00106944
R77276 VSS.n4856 VSS.n4855 0.00106944
R77277 VSS.n4920 VSS.n4919 0.00106944
R77278 VSS.n5475 VSS.n5474 0.00106944
R77279 VSS.n2513 VSS.n2512 0.00106944
R77280 VSS.n3939 VSS.n3938 0.00106944
R77281 VSS.n3938 VSS.n3937 0.00106944
R77282 VSS.n2945 VSS.n2944 0.00106429
R77283 VSS.n2944 VSS.n2943 0.00106429
R77284 VSS.n3219 VSS.n3218 0.00106338
R77285 VSS.n3672 VSS.n3671 0.00106338
R77286 DVSS VSS.n7856 0.00104667
R77287 VSS.n724 VSS.n723 0.00104
R77288 VSS.n20487 VSS.n20486 0.00104
R77289 VSS.n20509 VSS.n20508 0.00104
R77290 VSS.n20522 VSS.n20521 0.00104
R77291 VSS.n20237 VSS.n20236 0.00104
R77292 VSS.n725 VSS.n721 0.00104
R77293 VSS.n20581 VSS.n20580 0.00104
R77294 VSS.n20560 VSS.n20559 0.00104
R77295 VSS.n20531 VSS.n20530 0.00104
R77296 VSS.n10945 VSS.n10944 0.00104
R77297 VSS.n11013 VSS.n11012 0.00104
R77298 VSS.n11064 VSS.n11063 0.00104
R77299 VSS.n6358 VSS.n6351 0.00104
R77300 VSS.n8070 VSS.n8069 0.00104
R77301 VSS.n8010 VSS.n8009 0.00104
R77302 VSS.n7965 VSS.n7964 0.00104
R77303 VSS.n7929 VSS.n7922 0.00104
R77304 VSS.n6754 VSS.n6753 0.00104
R77305 VSS.n6694 VSS.n6693 0.00104
R77306 VSS.n7872 VSS.n7871 0.00104
R77307 VSS.n7033 VSS.n7032 0.00104
R77308 VSS.n7873 VSS.n7869 0.00104
R77309 VSS.n7034 VSS.n7030 0.00104
R77310 VSS.n7966 VSS.n7962 0.00104
R77311 VSS.n7928 VSS.n7927 0.00104
R77312 VSS.n11066 VSS.n11065 0.00104
R77313 VSS.n6357 VSS.n6356 0.00104
R77314 VSS.n11140 VSS.n11139 0.00103333
R77315 VSS.n2924 VSS.n2923 0.00103214
R77316 VSS.n2987 VSS.n2986 0.00103214
R77317 VSS.n3035 VSS.n3034 0.00103214
R77318 VSS.n3036 VSS.n3035 0.00103214
R77319 VSS.n2988 VSS.n2987 0.00103214
R77320 VSS.n2923 VSS.n2922 0.00103214
R77321 VSS.n3986 VSS.n3985 0.0010315
R77322 VSS.n2358 VSS.n2357 0.0010315
R77323 VSS.n17478 VSS.n17477 0.0010315
R77324 VSS.n11364 VSS.n11363 0.0010315
R77325 VSS.n5729 VSS.n5728 0.0010315
R77326 VSS.n5625 VSS.n5624 0.0010315
R77327 VSS.n5612 VSS.n5611 0.0010315
R77328 VSS.n5602 VSS.n5601 0.0010315
R77329 VSS.n13012 VSS.n13011 0.0010315
R77330 VSS.n13168 VSS.n13167 0.0010315
R77331 VSS.n12843 VSS.n12842 0.0010315
R77332 VSS.n12780 VSS.n12779 0.0010315
R77333 VSS.n12526 VSS.n12525 0.0010315
R77334 VSS.n12307 VSS.n12306 0.0010315
R77335 VSS.n11969 VSS.n11968 0.0010315
R77336 VSS.n11955 VSS.n11954 0.0010315
R77337 VSS.n11877 VSS.n11876 0.0010315
R77338 VSS.n11871 VSS.n11870 0.0010315
R77339 VSS.n18857 VSS.n18856 0.0010315
R77340 VSS.n2257 VSS.n2256 0.0010315
R77341 VSS.n2229 VSS.n2228 0.0010315
R77342 VSS.n15165 VSS.n15164 0.0010315
R77343 VSS.n16177 VSS.n16176 0.0010315
R77344 VSS.n16147 VSS.n16146 0.0010315
R77345 VSS.n16128 VSS.n16127 0.0010315
R77346 VSS.n16118 VSS.n16117 0.0010315
R77347 VSS.n21785 VSS.n21784 0.0010315
R77348 VSS.n2308 VSS.n2307 0.0010315
R77349 VSS.n20817 VSS.n20816 0.0010315
R77350 VSS.n21117 VSS.n21116 0.0010315
R77351 VSS.n21075 VSS.n21074 0.0010315
R77352 VSS.n21062 VSS.n21061 0.0010315
R77353 VSS.n21052 VSS.n21051 0.0010315
R77354 VSS.n19070 VSS.n19069 0.0010315
R77355 VSS.n17916 VSS.n17915 0.0010315
R77356 VSS.n2002 VSS.n2001 0.0010315
R77357 VSS.n1167 VSS.n1166 0.0010315
R77358 VSS.n1127 VSS.n1126 0.0010315
R77359 VSS.n1108 VSS.n1107 0.0010315
R77360 VSS.n1098 VSS.n1097 0.0010315
R77361 VSS.n21553 VSS.n21552 0.0010315
R77362 VSS.n21657 VSS.n21656 0.0010315
R77363 VSS.n21505 VSS.n21504 0.0010315
R77364 VSS.n21478 VSS.n21477 0.0010315
R77365 VSS.n21441 VSS.n21440 0.0010315
R77366 VSS.n21264 VSS.n21263 0.0010315
R77367 VSS.n7582 VSS.n7581 0.0010315
R77368 VSS.n3786 VSS.n3785 0.0010315
R77369 VSS.n3886 VSS.n3885 0.0010315
R77370 VSS.n4711 VSS.n4710 0.0010315
R77371 VSS.n4759 VSS.n4758 0.0010315
R77372 VSS.n4794 VSS.n4793 0.0010315
R77373 VSS.n11424 VSS.n11423 0.0010315
R77374 VSS.n11203 VSS.n11202 0.0010315
R77375 VSS.n3266 VSS.n3265 0.0010315
R77376 VSS.n542 VSS.n541 0.0010315
R77377 VSS.n483 VSS.n482 0.0010315
R77378 VSS.n10471 VSS.n10470 0.0010315
R77379 VSS.n10255 VSS.n10254 0.0010315
R77380 VSS.n9972 VSS.n9971 0.0010315
R77381 VSS.n9957 VSS.n9956 0.0010315
R77382 VSS.n8939 VSS.n8938 0.0010315
R77383 VSS.n8790 VSS.n8789 0.0010315
R77384 VSS.n11007 VSS.n11006 0.00103
R77385 VSS.n11059 VSS.n11058 0.00103
R77386 VSS.n11006 VSS.n11005 0.00103
R77387 VSS.n11058 VSS.n11057 0.00103
R77388 VSS.n2576 VSS.n2544 0.00101429
R77389 VSS.n2884 VSS.n2883 0.00101429
R77390 VSS.n2952 VSS.n2951 0.00101429
R77391 VSS.n3016 VSS.n3015 0.00101429
R77392 VSS.n3064 VSS.n3063 0.00101429
R77393 VSS.n3079 VSS.n3078 0.00101429
R77394 VSS.n4684 VSS.n4683 0.00101429
R77395 VSS.n4342 VSS.n4341 0.00101429
R77396 VSS.n17602 VSS.n17601 0.00101429
R77397 VSS.n18016 VSS.n18015 0.00101429
R77398 VSS.n17861 VSS.n17857 0.00101429
R77399 VSS.n17800 VSS.n17796 0.00101429
R77400 VSS.n17755 VSS.n17751 0.00101429
R77401 VSS.n17734 VSS.n17733 0.00101429
R77402 VSS.n22260 VSS 0.00101429
R77403 VSS.n721 VSS.n720 0.00101
R77404 VSS.n20580 VSS.n20579 0.00101
R77405 VSS.n20559 VSS.n20558 0.00101
R77406 VSS.n20530 VSS.n20529 0.00101
R77407 VSS.n8439 VSS.n8435 0.00101
R77408 VSS.n8771 VSS.n8767 0.00101
R77409 VSS.n10815 VSS.n10814 0.00101
R77410 VSS.n11067 VSS.n11066 0.00101
R77411 VSS.n3477 VSS.n3476 0.000992958
R77412 VSS.n3481 VSS.n3480 0.000992958
R77413 VSS.n20218 VSS.n20217 0.00098
R77414 VSS.n11712 VSS.n11711 0.00098
R77415 VSS.n20382 VSS.n20381 0.00098
R77416 VSS.n20351 VSS.n20350 0.00098
R77417 VSS.n20305 VSS.n20304 0.00098
R77418 VSS.n20219 VSS.n20215 0.00098
R77419 VSS.n20215 VSS.n20214 0.00098
R77420 VSS.n10856 VSS.n10855 0.00098
R77421 VSS.n8732 VSS.n8731 0.00098
R77422 VSS.n8275 VSS.n8274 0.00098
R77423 VSS.n8801 VSS.n8800 0.00098
R77424 VSS.n8842 VSS.n8841 0.00098
R77425 VSS.n9406 VSS.n9405 0.00098
R77426 VSS.n9352 VSS.n9351 0.00098
R77427 VSS.n8271 VSS.n8270 0.00098
R77428 VSS.n6747 VSS.n6746 0.00098
R77429 VSS.n6687 VSS.n6686 0.00098
R77430 VSS.n9414 VSS.n9413 0.00098
R77431 VSS.n9445 VSS.n9444 0.00098
R77432 VSS.n9797 VSS.n9796 0.00098
R77433 VSS.n9743 VSS.n9742 0.00098
R77434 VSS.n8728 VSS.n8727 0.00098
R77435 VSS.n8063 VSS.n8062 0.00098
R77436 VSS.n8003 VSS.n8002 0.00098
R77437 VSS.n6156 VSS.n6155 0.00098
R77438 VSS.n9819 VSS.n9818 0.00098
R77439 VSS.n10691 VSS.n10690 0.00098
R77440 VSS.n10753 VSS.n10752 0.00098
R77441 VSS.n10860 VSS.n10859 0.00098
R77442 VSS.n4322 DVSS 0.000957143
R77443 VSS.n18382 VSS.n18379 0.00095
R77444 VSS.n16561 VSS.n16560 0.00095
R77445 VSS.n2887 VSS.n2886 0.00095
R77446 VSS.n2889 VSS.n2888 0.00095
R77447 VSS.n11716 VSS.n11714 0.00095
R77448 VSS.n20379 VSS.n20377 0.00095
R77449 VSS.n20348 VSS.n20346 0.00095
R77450 VSS.n20302 VSS.n20300 0.00095
R77451 VSS.n11717 VSS.n11712 0.00095
R77452 VSS.n20381 VSS.n20380 0.00095
R77453 VSS.n20350 VSS.n20349 0.00095
R77454 VSS.n20304 VSS.n20303 0.00095
R77455 VSS.n5158 VSS.n5157 0.00095
R77456 VSS.n5160 VSS.n5159 0.00095
R77457 VSS.n5161 VSS.n5160 0.00095
R77458 VSS.n7220 VSS.n7219 0.00095
R77459 VSS.n7217 VSS.n7216 0.00095
R77460 VSS.n4496 VSS.n4495 0.00095
R77461 VSS.n4497 VSS.n4494 0.00095
R77462 VSS.n4494 VSS.n4493 0.00095
R77463 VSS.n18014 VSS.n18010 0.00095
R77464 VSS.n18010 VSS.n18009 0.00095
R77465 VSS.n18013 VSS.n18012 0.00095
R77466 VSS.n6159 VSS.n6157 0.00095
R77467 VSS.n9822 VSS.n9820 0.00095
R77468 VSS.n10666 VSS.n10664 0.00095
R77469 VSS.n10728 VSS.n10726 0.00095
R77470 VSS.n9417 VSS.n9415 0.00095
R77471 VSS.n9448 VSS.n9446 0.00095
R77472 VSS.n9793 VSS.n9791 0.00095
R77473 VSS.n9739 VSS.n9737 0.00095
R77474 VSS.n8804 VSS.n8802 0.00095
R77475 VSS.n8845 VSS.n8843 0.00095
R77476 VSS.n9402 VSS.n9400 0.00095
R77477 VSS.n9348 VSS.n9346 0.00095
R77478 VSS.n8805 VSS.n8801 0.00095
R77479 VSS.n8846 VSS.n8842 0.00095
R77480 VSS.n8920 VSS.n8919 0.00095
R77481 VSS.n9408 VSS.n9407 0.00095
R77482 VSS.n9354 VSS.n9353 0.00095
R77483 VSS.n8269 VSS.n8268 0.00095
R77484 VSS.n7878 VSS.n7877 0.00095
R77485 VSS.n9418 VSS.n9414 0.00095
R77486 VSS.n9449 VSS.n9445 0.00095
R77487 VSS.n9454 VSS.n9453 0.00095
R77488 VSS.n9799 VSS.n9798 0.00095
R77489 VSS.n9745 VSS.n9744 0.00095
R77490 VSS.n8606 VSS.n8605 0.00095
R77491 VSS.n7971 VSS.n7970 0.00095
R77492 VSS.n6160 VSS.n6156 0.00095
R77493 VSS.n9823 VSS.n9819 0.00095
R77494 VSS.n10627 VSS.n10626 0.00095
R77495 VSS.n10689 VSS.n10688 0.00095
R77496 VSS.n10751 VSS.n10750 0.00095
R77497 VSS.n10862 VSS.n10861 0.00095
R77498 VSS.n10916 VSS.n10915 0.00095
R77499 VSS.n10919 VSS.n10918 0.00095
R77500 VSS.n10983 VSS.n10982 0.00095
R77501 VSS.n10986 VSS.n10985 0.00095
R77502 VSS.n11057 VSS.n11056 0.00095
R77503 VSS.n11115 VSS.n11114 0.000926667
R77504 VSS.n3479 VSS.n3478 0.000922535
R77505 VSS.n18775 VSS.n18774 0.000922535
R77506 VSS.n18785 VSS.n18784 0.000922535
R77507 VSS.n18791 VSS.n18790 0.000922535
R77508 VSS.n18795 VSS.n18794 0.000922535
R77509 VSS.n18465 VSS.n18464 0.000922535
R77510 VSS.n18443 VSS.n18442 0.000922535
R77511 VSS.n18394 VSS.n18393 0.000922535
R77512 VSS.n18206 VSS.n18205 0.000922535
R77513 VSS.n18205 VSS.n18204 0.000922535
R77514 VSS.n18195 VSS.n18194 0.000922535
R77515 VSS.n18141 VSS.n18140 0.000922535
R77516 VSS.n17030 VSS.n17029 0.000922535
R77517 VSS.n14879 VSS.n14878 0.000922535
R77518 VSS.n16632 VSS.n16631 0.000922535
R77519 VSS.n16534 VSS.n16533 0.000922535
R77520 VSS.n16529 VSS.n16528 0.000922535
R77521 VSS.n15543 VSS.n15542 0.000922535
R77522 VSS.n15522 VSS.n15521 0.000922535
R77523 VSS.n8486 VSS.n8485 0.000922535
R77524 VSS.n8357 VSS.n8356 0.000922535
R77525 VSS.n19447 VSS.n19446 0.000922535
R77526 VSS.n19457 VSS.n19456 0.000922535
R77527 VSS.n19463 VSS.n19462 0.000922535
R77528 VSS.n19467 VSS.n19466 0.000922535
R77529 VSS.n19574 VSS.n19573 0.000922535
R77530 VSS.n19596 VSS.n19595 0.000922535
R77531 VSS.n19628 VSS.n19627 0.000922535
R77532 VSS.n19650 VSS.n19649 0.000922535
R77533 VSS.n19651 VSS.n19650 0.000922535
R77534 VSS.n19661 VSS.n19660 0.000922535
R77535 VSS.n19715 VSS.n19714 0.000922535
R77536 VSS.n19905 VSS.n19904 0.000922535
R77537 VSS.n19950 VSS.n19949 0.000922535
R77538 VSS.n766 VSS.n765 0.000922535
R77539 VSS.n804 VSS.n803 0.000922535
R77540 VSS.n809 VSS.n808 0.000922535
R77541 VSS.n1831 VSS.n1830 0.000922535
R77542 VSS.n1810 VSS.n1809 0.000922535
R77543 VSS.n8637 VSS.n8636 0.000922535
R77544 VSS.n8165 VSS.n8164 0.000922535
R77545 VSS.n20246 VSS.n20244 0.00092
R77546 VSS.n20246 VSS.n20245 0.00092
R77547 VSS.n20249 VSS.n20248 0.00092
R77548 VSS.n20248 VSS.n20247 0.00092
R77549 VSS.n20247 VSS.n20243 0.00092
R77550 VSS.n10825 VSS.n10823 0.00092
R77551 VSS.n10825 VSS.n10824 0.00092
R77552 VSS.n8759 VSS.n8757 0.00092
R77553 VSS.n8759 VSS.n8758 0.00092
R77554 VSS.n8302 VSS.n8300 0.00092
R77555 VSS.n8302 VSS.n8301 0.00092
R77556 VSS.n8432 VSS.n8431 0.00092
R77557 VSS.n8431 VSS.n8305 0.00092
R77558 VSS.n8303 VSS.n8299 0.00092
R77559 VSS.n8764 VSS.n8763 0.00092
R77560 VSS.n8763 VSS.n8762 0.00092
R77561 VSS.n8760 VSS.n8756 0.00092
R77562 VSS.n10821 VSS.n10820 0.00092
R77563 VSS.n10827 VSS.n10826 0.00092
R77564 VSS.n11716 VSS.n11715 0.00089
R77565 VSS.n20379 VSS.n20378 0.00089
R77566 VSS.n20348 VSS.n20347 0.00089
R77567 VSS.n20302 VSS.n20301 0.00089
R77568 VSS.n11718 VSS.n11717 0.00089
R77569 VSS.n20380 VSS.n20376 0.00089
R77570 VSS.n20349 VSS.n20345 0.00089
R77571 VSS.n20303 VSS.n20299 0.00089
R77572 VSS.n6159 VSS.n6158 0.00089
R77573 VSS.n9822 VSS.n9821 0.00089
R77574 VSS.n10666 VSS.n10665 0.00089
R77575 VSS.n10728 VSS.n10727 0.00089
R77576 VSS.n9417 VSS.n9416 0.00089
R77577 VSS.n9448 VSS.n9447 0.00089
R77578 VSS.n9793 VSS.n9792 0.00089
R77579 VSS.n9739 VSS.n9738 0.00089
R77580 VSS.n8804 VSS.n8803 0.00089
R77581 VSS.n8845 VSS.n8844 0.00089
R77582 VSS.n9402 VSS.n9401 0.00089
R77583 VSS.n9348 VSS.n9347 0.00089
R77584 VSS.n8806 VSS.n8805 0.00089
R77585 VSS.n8847 VSS.n8846 0.00089
R77586 VSS.n9403 VSS.n9399 0.00089
R77587 VSS.n9349 VSS.n9345 0.00089
R77588 VSS.n8433 VSS.n8432 0.00089
R77589 VSS.n8305 VSS.n8304 0.00089
R77590 VSS.n8266 VSS.n8265 0.00089
R77591 VSS.n9419 VSS.n9418 0.00089
R77592 VSS.n9450 VSS.n9449 0.00089
R77593 VSS.n9794 VSS.n9790 0.00089
R77594 VSS.n9740 VSS.n9736 0.00089
R77595 VSS.n8765 VSS.n8764 0.00089
R77596 VSS.n8762 VSS.n8761 0.00089
R77597 VSS.n8603 VSS.n8602 0.00089
R77598 VSS.n6161 VSS.n6160 0.00089
R77599 VSS.n9824 VSS.n9823 0.00089
R77600 VSS.n10668 VSS.n10667 0.00089
R77601 VSS.n10730 VSS.n10729 0.00089
R77602 VSS.n10818 VSS.n10817 0.00089
R77603 VSS.n10822 VSS.n10821 0.00089
R77604 VSS.n10868 VSS.n10864 0.00089
R77605 VSS.n2835 VSS.n2834 0.000885714
R77606 VSS.n2893 VSS.n2892 0.000885714
R77607 VSS.n7221 VSS.n7218 0.000885714
R77608 VSS.n18062 VSS.n18061 0.000885714
R77609 VSS.n18008 VSS.n18007 0.000885714
R77610 VSS.n20218 VSS.n20216 0.00086
R77611 VSS.n11711 VSS.n11710 0.00086
R77612 VSS.n20383 VSS.n20382 0.00086
R77613 VSS.n20306 VSS.n20305 0.00086
R77614 VSS.n20220 VSS.n20219 0.00086
R77615 VSS.n10856 VSS.n10854 0.00086
R77616 VSS.n8732 VSS.n8730 0.00086
R77617 VSS.n8275 VSS.n8273 0.00086
R77618 VSS.n8800 VSS.n8799 0.00086
R77619 VSS.n9407 VSS.n9406 0.00086
R77620 VSS.n9353 VSS.n9352 0.00086
R77621 VSS.n8277 VSS.n8276 0.00086
R77622 VSS.n8270 VSS.n8269 0.00086
R77623 VSS.n9413 VSS.n9412 0.00086
R77624 VSS.n9798 VSS.n9797 0.00086
R77625 VSS.n9744 VSS.n9743 0.00086
R77626 VSS.n8734 VSS.n8733 0.00086
R77627 VSS.n8727 VSS.n8606 0.00086
R77628 VSS.n6155 VSS.n6154 0.00086
R77629 VSS.n9818 VSS.n9817 0.00086
R77630 VSS.n10660 VSS.n10659 0.00086
R77631 VSS.n10661 VSS.n10660 0.00086
R77632 VSS.n10690 VSS.n10689 0.00086
R77633 VSS.n10722 VSS.n10721 0.00086
R77634 VSS.n10723 VSS.n10722 0.00086
R77635 VSS.n10752 VSS.n10751 0.00086
R77636 VSS.n10857 VSS.n10853 0.00086
R77637 VSS.n10861 VSS.n10860 0.00086
R77638 VSS.n10918 VSS.n10917 0.00086
R77639 VSS.n10950 VSS.n10949 0.00086
R77640 VSS.n10985 VSS.n10984 0.00086
R77641 VSS.n11018 VSS.n11017 0.00086
R77642 VSS.n4030 VSS.n4029 0.000854331
R77643 VSS.n3947 VSS.n3946 0.000854331
R77644 VSS.n2369 VSS.n2368 0.000854331
R77645 VSS.n17442 VSS.n17441 0.000854331
R77646 VSS.n11338 VSS.n11337 0.000854331
R77647 VSS.n5859 VSS.n5858 0.000854331
R77648 VSS.n5839 VSS.n5838 0.000854331
R77649 VSS.n9504 VSS.n9503 0.000854331
R77650 VSS.n13057 VSS.n13056 0.000854331
R77651 VSS.n13133 VSS.n13132 0.000854331
R77652 VSS.n13181 VSS.n13180 0.000854331
R77653 VSS.n13231 VSS.n13230 0.000854331
R77654 VSS.n12871 VSS.n12870 0.000854331
R77655 VSS.n12808 VSS.n12807 0.000854331
R77656 VSS.n12314 VSS.n12313 0.000854331
R77657 VSS.n12239 VSS.n12238 0.000854331
R77658 VSS.n12235 VSS.n12234 0.000854331
R77659 VSS.n11872 VSS.n11871 0.000854331
R77660 VSS.n11825 VSS.n11824 0.000854331
R77661 VSS.n11821 VSS.n11820 0.000854331
R77662 VSS.n18901 VSS.n18900 0.000854331
R77663 VSS.n18978 VSS.n18977 0.000854331
R77664 VSS.n2268 VSS.n2267 0.000854331
R77665 VSS.n2193 VSS.n2192 0.000854331
R77666 VSS.n15139 VSS.n15138 0.000854331
R77667 VSS.n16220 VSS.n16219 0.000854331
R77668 VSS.n16200 VSS.n16199 0.000854331
R77669 VSS.n9621 VSS.n9620 0.000854331
R77670 VSS.n21830 VSS.n21829 0.000854331
R77671 VSS.n21745 VSS.n21744 0.000854331
R77672 VSS.n2321 VSS.n2320 0.000854331
R77673 VSS.n13348 VSS.n13347 0.000854331
R77674 VSS.n20789 VSS.n20788 0.000854331
R77675 VSS.n21162 VSS.n21161 0.000854331
R77676 VSS.n21142 VSS.n21141 0.000854331
R77677 VSS.n6934 VSS.n6933 0.000854331
R77678 VSS.n19115 VSS.n19114 0.000854331
R77679 VSS.n19030 VSS.n19029 0.000854331
R77680 VSS.n17929 VSS.n17928 0.000854331
R77681 VSS.n13491 VSS.n13490 0.000854331
R77682 VSS.n2030 VSS.n2029 0.000854331
R77683 VSS.n1291 VSS.n1290 0.000854331
R77684 VSS.n1271 VSS.n1270 0.000854331
R77685 VSS.n6811 VSS.n6810 0.000854331
R77686 VSS.n21601 VSS.n21600 0.000854331
R77687 VSS.n21625 VSS.n21624 0.000854331
R77688 VSS.n21677 VSS.n21676 0.000854331
R77689 VSS.n21492 VSS.n21491 0.000854331
R77690 VSS.n21292 VSS.n21291 0.000854331
R77691 VSS.n7554 VSS.n7553 0.000854331
R77692 VSS.n3832 VSS.n3831 0.000854331
R77693 VSS.n3853 VSS.n3852 0.000854331
R77694 VSS.n4138 VSS.n4137 0.000854331
R77695 VSS.n4722 VSS.n4721 0.000854331
R77696 VSS.n11450 VSS.n11449 0.000854331
R77697 VSS.n11229 VSS.n11228 0.000854331
R77698 VSS.n2647 VSS.n2646 0.000854331
R77699 VSS.n568 VSS.n567 0.000854331
R77700 VSS.n509 VSS.n508 0.000854331
R77701 VSS.n10261 VSS.n10260 0.000854331
R77702 VSS.n10188 VSS.n10187 0.000854331
R77703 VSS.n10183 VSS.n10182 0.000854331
R77704 VSS.n8789 VSS.n8788 0.000854331
R77705 VSS.n8935 VSS.n8934 0.000854331
R77706 VSS.n8931 VSS.n8930 0.000854331
R77707 VSS.n3429 VSS.n3427 0.000852113
R77708 VSS.n3451 VSS.n3450 0.000852113
R77709 VSS.n3425 VSS.n3424 0.000852113
R77710 VSS.n3444 VSS.n3443 0.000852113
R77711 VSS.n3448 VSS.n3447 0.000852113
R77712 VSS.n3453 VSS.n3452 0.000852113
R77713 VSS.n3460 VSS.n3459 0.000852113
R77714 VSS.n3464 VSS.n3463 0.000852113
R77715 VSS.n3539 VSS.n3538 0.000852113
R77716 VSS.n3542 VSS.n3541 0.000852113
R77717 VSS.n3598 VSS.n3597 0.000852113
R77718 VSS.n3601 VSS.n3600 0.000852113
R77719 VSS.n3641 VSS.n3640 0.000852113
R77720 VSS.n3644 VSS.n3643 0.000852113
R77721 VSS.n20579 VSS.n20578 0.00083
R77722 VSS.n9405 VSS.n9404 0.00083
R77723 VSS.n9351 VSS.n9350 0.00083
R77724 VSS.n8272 VSS.n8271 0.00083
R77725 VSS.n6748 VSS.n6747 0.00083
R77726 VSS.n6688 VSS.n6687 0.00083
R77727 VSS.n7879 VSS.n7878 0.00083
R77728 VSS.n7876 VSS.n7875 0.00083
R77729 VSS.n7867 VSS.n7866 0.00083
R77730 VSS.n7028 VSS.n7027 0.00083
R77731 VSS.n9796 VSS.n9795 0.00083
R77732 VSS.n9742 VSS.n9741 0.00083
R77733 VSS.n8729 VSS.n8728 0.00083
R77734 VSS.n8064 VSS.n8063 0.00083
R77735 VSS.n8004 VSS.n8003 0.00083
R77736 VSS.n7972 VSS.n7971 0.00083
R77737 VSS.n7969 VSS.n7968 0.00083
R77738 VSS.n7960 VSS.n7959 0.00083
R77739 VSS.n7925 VSS.n7924 0.00083
R77740 VSS.n10658 VSS.n10657 0.00083
R77741 VSS.n10663 VSS.n10662 0.00083
R77742 VSS.n10692 VSS.n10691 0.00083
R77743 VSS.n10720 VSS.n10719 0.00083
R77744 VSS.n10725 VSS.n10724 0.00083
R77745 VSS.n10754 VSS.n10753 0.00083
R77746 VSS.n10859 VSS.n10858 0.00083
R77747 VSS.n10915 VSS.n10914 0.00083
R77748 VSS.n10954 VSS.n10953 0.00083
R77749 VSS.n10982 VSS.n10981 0.00083
R77750 VSS.n11019 VSS.n11018 0.00083
R77751 VSS.n11021 VSS.n11020 0.00083
R77752 VSS.n11056 VSS.n11055 0.00083
R77753 VSS.n11060 VSS.n11059 0.00083
R77754 VSS.n6354 VSS.n6353 0.00083
R77755 VSS.n2832 VSS.n2830 0.000821429
R77756 VSS.n2858 VSS.n2857 0.000821429
R77757 VSS.n2833 VSS.n2829 0.000821429
R77758 VSS.n2860 VSS.n2859 0.000821429
R77759 VSS.n2877 VSS.n2876 0.000821429
R77760 VSS.n5134 VSS.n5133 0.000821429
R77761 VSS.n5112 VSS.n5111 0.000821429
R77762 VSS.n5115 VSS.n5112 0.000821429
R77763 VSS.n5128 VSS.n5127 0.000821429
R77764 VSS.n5131 VSS.n5130 0.000821429
R77765 VSS.n5136 VSS.n5135 0.000821429
R77766 VSS.n7244 VSS.n7243 0.000821429
R77767 VSS.n7266 VSS.n7265 0.000821429
R77768 VSS.n7249 VSS.n7248 0.000821429
R77769 VSS.n7245 VSS.n7241 0.000821429
R77770 VSS.n7236 VSS.n7235 0.000821429
R77771 VSS.n7233 VSS.n7232 0.000821429
R77772 VSS.n7159 VSS.n7158 0.000821429
R77773 VSS.n7156 VSS.n7155 0.000821429
R77774 VSS.n7100 VSS.n7099 0.000821429
R77775 VSS.n7097 VSS.n7096 0.000821429
R77776 VSS.n4521 VSS.n4520 0.000821429
R77777 VSS.n4543 VSS.n4542 0.000821429
R77778 VSS.n4542 VSS.n4541 0.000821429
R77779 VSS.n4527 VSS.n4526 0.000821429
R77780 VSS.n4524 VSS.n4523 0.000821429
R77781 VSS.n4522 VSS.n4518 0.000821429
R77782 VSS.n18068 VSS.n18067 0.000821429
R77783 VSS.n18067 VSS.n18066 0.000821429
R77784 VSS.n18047 VSS.n18046 0.000821429
R77785 VSS.n18041 VSS.n18037 0.000821429
R77786 VSS.n18025 VSS.n18021 0.000821429
R77787 VSS.n18065 VSS.n18063 0.000821429
R77788 VSS.n18040 VSS.n18039 0.000821429
R77789 VSS.n11090 VSS.n11089 0.00082
R77790 VSS.n724 VSS.n722 0.0008
R77791 VSS.n20487 VSS.n20485 0.0008
R77792 VSS.n20509 VSS.n20507 0.0008
R77793 VSS.n20523 VSS.n20522 0.0008
R77794 VSS.n726 VSS.n725 0.0008
R77795 VSS.n20582 VSS.n20581 0.0008
R77796 VSS.n20561 VSS.n20560 0.0008
R77797 VSS.n20532 VSS.n20531 0.0008
R77798 VSS.n10945 VSS.n10943 0.0008
R77799 VSS.n11013 VSS.n11011 0.0008
R77800 VSS.n11064 VSS.n11062 0.0008
R77801 VSS.n6358 VSS.n6350 0.0008
R77802 VSS.n8070 VSS.n8068 0.0008
R77803 VSS.n8010 VSS.n8008 0.0008
R77804 VSS.n7965 VSS.n7963 0.0008
R77805 VSS.n7929 VSS.n7921 0.0008
R77806 VSS.n6754 VSS.n6752 0.0008
R77807 VSS.n6694 VSS.n6692 0.0008
R77808 VSS.n7872 VSS.n7870 0.0008
R77809 VSS.n7033 VSS.n7031 0.0008
R77810 VSS.n8849 VSS.n8848 0.0008
R77811 VSS.n8921 VSS.n8920 0.0008
R77812 VSS.n6756 VSS.n6755 0.0008
R77813 VSS.n6751 VSS.n6750 0.0008
R77814 VSS.n6696 VSS.n6695 0.0008
R77815 VSS.n6691 VSS.n6690 0.0008
R77816 VSS.n7874 VSS.n7873 0.0008
R77817 VSS.n7035 VSS.n7034 0.0008
R77818 VSS.n9452 VSS.n9451 0.0008
R77819 VSS.n9455 VSS.n9454 0.0008
R77820 VSS.n8072 VSS.n8071 0.0008
R77821 VSS.n8067 VSS.n8066 0.0008
R77822 VSS.n8012 VSS.n8011 0.0008
R77823 VSS.n8007 VSS.n8006 0.0008
R77824 VSS.n7967 VSS.n7966 0.0008
R77825 VSS.n7928 VSS.n7923 0.0008
R77826 VSS.n9826 VSS.n9825 0.0008
R77827 VSS.n10628 VSS.n10627 0.0008
R77828 VSS.n10946 VSS.n10942 0.0008
R77829 VSS.n10948 VSS.n10947 0.0008
R77830 VSS.n11014 VSS.n11010 0.0008
R77831 VSS.n11016 VSS.n11015 0.0008
R77832 VSS.n11065 VSS.n11061 0.0008
R77833 VSS.n6357 VSS.n6352 0.0008
R77834 VSS.n3775 VSS.n3199 0.00078169
R77835 VSS.n3293 VSS.n3292 0.00078169
R77836 VSS.n3331 VSS.n3330 0.00078169
R77837 VSS.n3385 VSS.n3384 0.00078169
R77838 VSS.n3776 VSS.n3197 0.00078169
R77839 VSS.n3233 VSS.n3232 0.00078169
R77840 VSS.n3236 VSS.n3235 0.00078169
R77841 VSS.n3290 VSS.n3289 0.00078169
R77842 VSS.n3295 VSS.n3294 0.00078169
R77843 VSS.n3297 VSS.n3296 0.00078169
R77844 VSS.n3316 VSS.n3315 0.00078169
R77845 VSS.n3319 VSS.n3318 0.00078169
R77846 VSS.n3328 VSS.n3327 0.00078169
R77847 VSS.n3333 VSS.n3332 0.00078169
R77848 VSS.n3335 VSS.n3334 0.00078169
R77849 VSS.n3370 VSS.n3369 0.00078169
R77850 VSS.n3373 VSS.n3372 0.00078169
R77851 VSS.n3382 VSS.n3381 0.00078169
R77852 VSS.n3387 VSS.n3386 0.00078169
R77853 VSS.n3389 VSS.n3388 0.00078169
R77854 VSS.n3522 VSS.n3521 0.00078169
R77855 VSS.n3530 VSS.n3529 0.00078169
R77856 VSS.n3581 VSS.n3580 0.00078169
R77857 VSS.n3589 VSS.n3588 0.00078169
R77858 VSS.n3624 VSS.n3623 0.00078169
R77859 VSS.n3632 VSS.n3631 0.00078169
R77860 VSS.n2540 VSS.n2537 0.000757143
R77861 VSS.n2680 VSS.n2679 0.000757143
R77862 VSS.n2725 VSS.n2724 0.000757143
R77863 VSS.n2785 VSS.n2784 0.000757143
R77864 VSS.n2542 VSS.n2541 0.000757143
R77865 VSS.n2671 VSS.n2666 0.000757143
R77866 VSS.n2682 VSS.n2681 0.000757143
R77867 VSS.n2715 VSS.n2710 0.000757143
R77868 VSS.n2727 VSS.n2726 0.000757143
R77869 VSS.n2775 VSS.n2770 0.000757143
R77870 VSS.n2787 VSS.n2786 0.000757143
R77871 VSS.n2826 VSS.n2825 0.000757143
R77872 VSS.n2854 VSS.n2853 0.000757143
R77873 VSS.n5410 VSS.n4946 0.000757143
R77874 VSS.n5000 VSS.n4999 0.000757143
R77875 VSS.n5030 VSS.n5029 0.000757143
R77876 VSS.n5076 VSS.n5075 0.000757143
R77877 VSS.n5411 VSS.n4943 0.000757143
R77878 VSS.n5002 VSS.n5001 0.000757143
R77879 VSS.n5032 VSS.n5031 0.000757143
R77880 VSS.n5078 VSS.n5077 0.000757143
R77881 VSS.n5920 VSS.n5919 0.000757143
R77882 VSS.n7394 VSS.n7393 0.000757143
R77883 VSS.n7360 VSS.n7359 0.000757143
R77884 VSS.n7306 VSS.n7305 0.000757143
R77885 VSS.n5922 VSS.n5921 0.000757143
R77886 VSS.n7395 VSS.n7392 0.000757143
R77887 VSS.n7377 VSS.n7376 0.000757143
R77888 VSS.n7374 VSS.n7373 0.000757143
R77889 VSS.n7364 VSS.n7363 0.000757143
R77890 VSS.n7361 VSS.n7358 0.000757143
R77891 VSS.n7357 VSS.n7356 0.000757143
R77892 VSS.n7323 VSS.n7322 0.000757143
R77893 VSS.n7320 VSS.n7319 0.000757143
R77894 VSS.n7310 VSS.n7309 0.000757143
R77895 VSS.n7307 VSS.n7304 0.000757143
R77896 VSS.n7303 VSS.n7302 0.000757143
R77897 VSS.n7176 VSS.n7175 0.000757143
R77898 VSS.n7168 VSS.n7167 0.000757143
R77899 VSS.n7117 VSS.n7116 0.000757143
R77900 VSS.n7109 VSS.n7108 0.000757143
R77901 VSS.n2445 VSS.n2444 0.000757143
R77902 VSS.n4624 VSS.n4623 0.000757143
R77903 VSS.n4578 VSS.n4577 0.000757143
R77904 VSS.n4691 VSS.n4690 0.000757143
R77905 VSS.n4625 VSS.n4622 0.000757143
R77906 VSS.n4579 VSS.n4576 0.000757143
R77907 VSS.n4752 VSS.n4751 0.000757143
R77908 VSS.n17558 VSS.n17557 0.000757143
R77909 VSS.n17546 VSS.n17542 0.000757143
R77910 VSS.n17500 VSS.n17499 0.000757143
R77911 VSS.n17488 VSS.n17484 0.000757143
R77912 VSS.n18070 VSS.n18069 0.000757143
R77913 VSS.n18044 VSS.n18043 0.000757143
R77914 VSS.n4750 VSS.n4748 0.000757143
R77915 VSS.n17545 VSS.n17544 0.000757143
R77916 VSS.n17487 VSS.n17486 0.000757143
R77917 VSS.n164 VSS.n163 0.000751397
R77918 VSS.n342 VSS.n339 0.000751397
R77919 VSS.n21240 VSS.n21237 0.000751397
R77920 VSS.n11253 VSS.n11251 0.000751397
R77921 VSS.n8267 VSS.n8266 0.00074
R77922 VSS.n6755 VSS.n6751 0.00074
R77923 VSS.n6695 VSS.n6691 0.00074
R77924 VSS.n8604 VSS.n8603 0.00074
R77925 VSS.n8071 VSS.n8067 0.00074
R77926 VSS.n8011 VSS.n8007 0.00074
R77927 VSS.n10864 VSS.n10863 0.00074
R77928 VSS.n10947 VSS.n10946 0.00074
R77929 VSS.n11015 VSS.n11014 0.00074
R77930 VSS.n19248 VSS.n19247 0.000725
R77931 VSS.n19271 VSS.n19268 0.000725
R77932 VSS.n16988 VSS.n16986 0.000725
R77933 VSS.n16972 VSS.n16971 0.000725
R77934 DVSS VSS.n16508 0.000725
R77935 VSS.n3779 VSS.n3196 0.000711268
R77936 VSS.n3289 VSS.n3243 0.000711268
R77937 VSS.n3327 VSS.n3326 0.000711268
R77938 VSS.n3381 VSS.n3380 0.000711268
R77939 VSS.n3423 VSS.n3422 0.000711268
R77940 VSS.n3426 VSS.n3425 0.000711268
R77941 VSS.n3443 VSS.n3442 0.000711268
R77942 VSS.n3447 VSS.n3446 0.000711268
R77943 VSS.n3457 VSS.n3454 0.000711268
R77944 VSS.n3463 VSS.n3462 0.000711268
R77945 VSS.n18728 VSS.n18727 0.000711268
R77946 VSS.n18733 VSS.n18732 0.000711268
R77947 VSS.n18754 VSS.n18753 0.000711268
R77948 VSS.n18412 VSS.n18411 0.000711268
R77949 VSS.n18409 VSS.n18408 0.000711268
R77950 VSS.n18198 VSS.n18197 0.000711268
R77951 VSS.n17082 VSS.n17081 0.000711268
R77952 VSS.n17066 VSS.n17065 0.000711268
R77953 VSS.n17021 VSS.n17020 0.000711268
R77954 VSS.n14876 VSS.n14875 0.000711268
R77955 VSS.n14878 VSS.n14877 0.000711268
R77956 VSS.n14885 VSS.n14884 0.000711268
R77957 VSS.n14899 VSS.n14898 0.000711268
R77958 VSS.n16886 VSS.n16885 0.000711268
R77959 VSS.n16577 VSS.n16546 0.000711268
R77960 VSS.n15401 VSS.n15400 0.000711268
R77961 VSS.n15363 VSS.n15362 0.000711268
R77962 VSS.n15330 VSS.n15329 0.000711268
R77963 VSS.n8565 VSS.n8564 0.000711268
R77964 VSS.n8331 VSS.n8330 0.000711268
R77965 VSS.n8420 VSS.n8419 0.000711268
R77966 VSS.n19210 VSS.n19209 0.000711268
R77967 VSS.n19215 VSS.n19214 0.000711268
R77968 VSS.n19236 VSS.n19235 0.000711268
R77969 VSS.n19610 VSS.n19609 0.000711268
R77970 VSS.n19613 VSS.n19612 0.000711268
R77971 VSS.n19658 VSS.n19657 0.000711268
R77972 VSS.n19883 VSS.n19882 0.000711268
R77973 VSS.n19899 VSS.n19898 0.000711268
R77974 VSS.n19914 VSS.n19913 0.000711268
R77975 VSS.n19947 VSS.n19946 0.000711268
R77976 VSS.n19949 VSS.n19948 0.000711268
R77977 VSS.n19956 VSS.n19955 0.000711268
R77978 VSS.n19970 VSS.n19969 0.000711268
R77979 VSS.n20030 VSS.n20029 0.000711268
R77980 VSS.n791 VSS.n790 0.000711268
R77981 VSS.n1717 VSS.n1716 0.000711268
R77982 VSS.n1679 VSS.n1678 0.000711268
R77983 VSS.n1646 VSS.n1645 0.000711268
R77984 VSS.n8716 VSS.n8715 0.000711268
R77985 VSS.n8127 VSS.n8126 0.000711268
R77986 VSS.n8228 VSS.n8227 0.000711268
R77987 VSS.n20209 VSS.n20208 0.00071
R77988 VSS.n20210 VSS.n20206 0.00071
R77989 VSS.n20206 VSS.n20205 0.00071
R77990 VSS.n10867 VSS.n10866 0.00071
R77991 VSS.n8601 VSS.n8600 0.00071
R77992 VSS.n8264 VSS.n8263 0.00071
R77993 VSS.n8993 VSS.n8992 0.00071
R77994 VSS.n8265 VSS.n8261 0.00071
R77995 VSS.n7887 VSS.n7886 0.00071
R77996 VSS.n9463 VSS.n9462 0.00071
R77997 VSS.n8602 VSS.n8598 0.00071
R77998 VSS.n7980 VSS.n7979 0.00071
R77999 VSS.n10636 VSS.n10635 0.00071
R78000 VSS.n11048 VSS.n11047 0.00071
R78001 VSS.n2533 VSS.n2532 0.000692857
R78002 VSS.n2864 VSS.n2861 0.000692857
R78003 VSS.n5413 VSS.n4942 0.000692857
R78004 VSS.n4997 VSS.n4996 0.000692857
R78005 VSS.n5027 VSS.n5026 0.000692857
R78006 VSS.n5073 VSS.n5072 0.000692857
R78007 VSS.n5140 VSS.n5137 0.000692857
R78008 VSS.n5145 VSS.n5144 0.000692857
R78009 VSS.n5914 VSS.n5913 0.000692857
R78010 VSS.n7398 VSS.n7397 0.000692857
R78011 VSS.n7365 VSS.n7364 0.000692857
R78012 VSS.n7311 VSS.n7310 0.000692857
R78013 VSS.n7268 VSS.n7267 0.000692857
R78014 VSS.n7265 VSS.n7264 0.000692857
R78015 VSS.n7250 VSS.n7249 0.000692857
R78016 VSS.n7247 VSS.n7246 0.000692857
R78017 VSS.n7240 VSS.n7239 0.000692857
R78018 VSS.n7234 VSS.n7233 0.000692857
R78019 VSS.n4694 VSS.n2442 0.000692857
R78020 VSS.n4628 VSS.n4627 0.000692857
R78021 VSS.n4582 VSS.n4581 0.000692857
R78022 VSS.n4517 VSS.n4516 0.000692857
R78023 VSS.n4510 VSS.n4509 0.000692857
R78024 VSS.n4744 VSS.n4743 0.000692857
R78025 VSS.n17550 VSS.n17549 0.000692857
R78026 VSS.n17492 VSS.n17491 0.000692857
R78027 VSS.n18036 VSS.n18035 0.000692857
R78028 VSS.n18029 VSS.n18028 0.000692857
R78029 VSS.n10534 VSS.n10529 0.000692308
R78030 VSS.n9893 VSS.n9892 0.000692308
R78031 VSS.n10385 VSS.n10380 0.000692308
R78032 VSS.n10362 VSS.n10361 0.000692308
R78033 VSS.n10100 VSS.n10095 0.000692308
R78034 VSS.n10077 VSS.n10076 0.000692308
R78035 VSS.n10008 VSS.n10003 0.000692308
R78036 VSS.n9985 VSS.n9984 0.000692308
R78037 VSS.n12600 VSS.n12595 0.000692308
R78038 VSS.n12572 VSS.n12571 0.000692308
R78039 VSS.n12439 VSS.n12434 0.000692308
R78040 VSS.n12416 VSS.n12415 0.000692308
R78041 VSS.n12151 VSS.n12146 0.000692308
R78042 VSS.n12128 VSS.n12127 0.000692308
R78043 VSS.n12059 VSS.n12054 0.000692308
R78044 VSS.n12036 VSS.n12035 0.000692308
R78045 VSS.n9844 VSS.n9843 0.000692308
R78046 VSS.n12636 VSS.n12635 0.000692308
R78047 VSS.n7859 DVSS 0.00068
R78048 VSS.n8435 VSS.n8434 0.00068
R78049 VSS.n8258 VSS.n8257 0.00068
R78050 DVSS VSS.n7860 0.00068
R78051 VSS.n8767 VSS.n8766 0.00068
R78052 VSS.n8595 VSS.n8594 0.00068
R78053 VSS.n10816 VSS.n10815 0.00068
R78054 VSS.n10869 VSS.n10868 0.00068
R78055 VSS.n10875 VSS.n10874 0.00068
R78056 VSS.n11535 VSS.n11534 0.000677165
R78057 VSS.n11591 VSS.n11590 0.000677165
R78058 VSS.n5588 VSS.n5587 0.000677165
R78059 VSS.n5569 VSS.n5568 0.000677165
R78060 VSS.n5557 VSS.n5556 0.000677165
R78061 VSS.n9503 VSS.n9502 0.000677165
R78062 VSS.n9584 VSS.n9583 0.000677165
R78063 VSS.n9038 VSS.n9037 0.000677165
R78064 VSS.n9147 VSS.n9146 0.000677165
R78065 VSS.n9088 VSS.n9087 0.000677165
R78066 VSS.n12969 VSS.n12968 0.000677165
R78067 VSS.n12906 VSS.n12905 0.000677165
R78068 VSS.n12751 VSS.n12750 0.000677165
R78069 VSS.n12688 VSS.n12687 0.000677165
R78070 VSS.n12678 VSS.n12677 0.000677165
R78071 VSS.n12675 VSS.n12674 0.000677165
R78072 VSS.n12593 VSS.n12592 0.000677165
R78073 VSS.n12573 VSS.n12563 0.000677165
R78074 VSS.n12540 VSS.n12539 0.000677165
R78075 VSS.n12519 VSS.n12518 0.000677165
R78076 VSS.n12504 VSS.n12503 0.000677165
R78077 VSS.n12271 VSS.n12270 0.000677165
R78078 VSS.n12270 VSS.n12269 0.000677165
R78079 VSS.n12266 VSS.n12265 0.000677165
R78080 VSS.n12249 VSS.n12248 0.000677165
R78081 VSS.n12227 VSS.n12226 0.000677165
R78082 VSS.n12216 VSS.n12215 0.000677165
R78083 VSS.n11926 VSS.n11925 0.000677165
R78084 VSS.n11925 VSS.n11924 0.000677165
R78085 VSS.n11924 VSS.n11923 0.000677165
R78086 VSS.n11917 VSS.n11916 0.000677165
R78087 VSS.n11903 VSS.n11902 0.000677165
R78088 VSS.n11876 VSS.n11875 0.000677165
R78089 VSS.n11854 VSS.n11853 0.000677165
R78090 VSS.n11850 VSS.n11849 0.000677165
R78091 VSS.n11842 VSS.n11841 0.000677165
R78092 VSS.n11820 VSS.n11819 0.000677165
R78093 VSS.n11795 VSS.n11794 0.000677165
R78094 VSS.n15009 VSS.n15008 0.000677165
R78095 VSS.n15066 VSS.n15065 0.000677165
R78096 VSS.n16104 VSS.n16103 0.000677165
R78097 VSS.n16085 VSS.n16084 0.000677165
R78098 VSS.n16067 VSS.n16066 0.000677165
R78099 VSS.n9620 VSS.n9619 0.000677165
R78100 VSS.n9701 VSS.n9700 0.000677165
R78101 VSS.n9181 VSS.n9180 0.000677165
R78102 VSS.n9310 VSS.n9309 0.000677165
R78103 VSS.n9252 VSS.n9251 0.000677165
R78104 VSS.n20615 VSS.n20614 0.000677165
R78105 VSS.n20678 VSS.n20677 0.000677165
R78106 VSS.n21038 VSS.n21037 0.000677165
R78107 VSS.n21006 VSS.n21005 0.000677165
R78108 VSS.n6996 VSS.n6995 0.000677165
R78109 VSS.n6671 VSS.n6670 0.000677165
R78110 VSS.n6636 VSS.n6635 0.000677165
R78111 VSS.n20134 VSS.n20133 0.000677165
R78112 VSS.n20071 VSS.n20070 0.000677165
R78113 VSS.n1084 VSS.n1083 0.000677165
R78114 VSS.n1052 VSS.n1051 0.000677165
R78115 VSS.n6894 VSS.n6893 0.000677165
R78116 VSS.n6521 VSS.n6520 0.000677165
R78117 VSS.n6486 VSS.n6485 0.000677165
R78118 VSS.n21645 VSS.n21644 0.000677165
R78119 VSS.n21528 VSS.n21527 0.000677165
R78120 VSS.n21386 VSS.n21385 0.000677165
R78121 VSS.n21323 VSS.n21322 0.000677165
R78122 VSS.n7611 VSS.n7610 0.000677165
R78123 VSS.n7674 VSS.n7673 0.000677165
R78124 VSS.n7699 VSS.n7698 0.000677165
R78125 VSS.n7762 VSS.n7761 0.000677165
R78126 VSS.n7840 VSS.n7839 0.000677165
R78127 VSS.n7777 VSS.n7776 0.000677165
R78128 VSS.n3874 VSS.n3873 0.000677165
R78129 VSS.n4145 VSS.n4144 0.000677165
R78130 VSS.n11700 VSS.n11699 0.000677165
R78131 VSS.n11643 VSS.n11642 0.000677165
R78132 VSS.n6143 VSS.n6142 0.000677165
R78133 VSS.n6087 VSS.n6086 0.000677165
R78134 VSS.n6062 VSS.n6061 0.000677165
R78135 VSS.n6006 VSS.n6005 0.000677165
R78136 VSS.n5981 VSS.n5980 0.000677165
R78137 VSS.n5925 VSS.n5924 0.000677165
R78138 VSS.n657 VSS.n656 0.000677165
R78139 VSS.n601 VSS.n600 0.000677165
R78140 VSS.n10615 VSS.n10614 0.000677165
R78141 VSS.n10556 VSS.n10555 0.000677165
R78142 VSS.n10546 VSS.n10545 0.000677165
R78143 VSS.n10543 VSS.n10542 0.000677165
R78144 VSS.n10527 VSS.n10526 0.000677165
R78145 VSS.n10508 VSS.n10507 0.000677165
R78146 VSS.n10485 VSS.n10484 0.000677165
R78147 VSS.n10464 VSS.n10463 0.000677165
R78148 VSS.n10450 VSS.n10449 0.000677165
R78149 VSS.n10220 VSS.n10219 0.000677165
R78150 VSS.n10219 VSS.n10218 0.000677165
R78151 VSS.n10214 VSS.n10213 0.000677165
R78152 VSS.n10198 VSS.n10197 0.000677165
R78153 VSS.n10175 VSS.n10174 0.000677165
R78154 VSS.n10165 VSS.n10164 0.000677165
R78155 VSS.n9927 VSS.n9926 0.000677165
R78156 VSS.n9926 VSS.n9925 0.000677165
R78157 VSS.n9925 VSS.n9924 0.000677165
R78158 VSS.n9918 VSS.n9917 0.000677165
R78159 VSS.n9903 VSS.n9902 0.000677165
R78160 VSS.n8938 VSS.n8937 0.000677165
R78161 VSS.n8796 VSS.n8795 0.000677165
R78162 VSS.n8972 VSS.n8971 0.000677165
R78163 VSS.n9001 VSS.n9000 0.000677165
R78164 VSS.n8930 VSS.n8929 0.000677165
R78165 VSS.n8898 VSS.n8897 0.000677165
R78166 VSS.n20255 VSS.n20253 0.00065
R78167 VSS.n20235 VSS.n20234 0.00065
R78168 VSS.n20258 VSS.n20257 0.00065
R78169 VSS.n20257 VSS.n20256 0.00065
R78170 VSS.n20241 VSS.n20240 0.00065
R78171 VSS.n20238 VSS.n20237 0.00065
R78172 VSS.n20236 VSS.n20229 0.00065
R78173 VSS.n10813 VSS.n10811 0.00065
R78174 VSS.n10841 VSS.n10840 0.00065
R78175 VSS.n8770 VSS.n8768 0.00065
R78176 VSS.n8748 VSS.n8747 0.00065
R78177 VSS.n8438 VSS.n8436 0.00065
R78178 VSS.n8291 VSS.n8290 0.00065
R78179 VSS.n8441 VSS.n8440 0.00065
R78180 VSS.n8440 VSS.n8439 0.00065
R78181 VSS.n8292 VSS.n8285 0.00065
R78182 VSS.n8276 VSS.n8272 0.00065
R78183 VSS.n8773 VSS.n8772 0.00065
R78184 VSS.n8772 VSS.n8771 0.00065
R78185 VSS.n8749 VSS.n8742 0.00065
R78186 VSS.n8733 VSS.n8729 0.00065
R78187 VSS.n10809 VSS.n10808 0.00065
R78188 VSS.n10843 VSS.n10842 0.00065
R78189 VSS.n10848 VSS.n10847 0.00065
R78190 VSS.n10851 VSS.n10850 0.00065
R78191 VSS.n10858 VSS.n10857 0.00065
R78192 VSS.n10949 VSS.n10948 0.00065
R78193 VSS.n10953 VSS.n10952 0.00065
R78194 VSS.n11017 VSS.n11016 0.00065
R78195 VSS.n11020 VSS.n11019 0.00065
R78196 VSS.n3517 VSS.n3516 0.000640845
R78197 VSS.n3576 VSS.n3575 0.000640845
R78198 VSS.n3619 VSS.n3618 0.000640845
R78199 VSS.n3211 VSS.n3207 0.000640845
R78200 VSS.n3215 VSS.n3214 0.000640845
R78201 VSS.n3430 VSS.n3426 0.000640845
R78202 VSS.n3459 VSS.n3458 0.000640845
R78203 VSS.n3519 VSS.n3518 0.000640845
R78204 VSS.n3531 VSS.n3530 0.000640845
R78205 VSS.n3578 VSS.n3577 0.000640845
R78206 VSS.n3590 VSS.n3589 0.000640845
R78207 VSS.n3621 VSS.n3620 0.000640845
R78208 VSS.n3633 VSS.n3632 0.000640845
R78209 VSS.n3669 VSS.n3668 0.000640845
R78210 VSS.n3667 VSS.n3666 0.000640845
R78211 VSS.n3660 VSS.n3659 0.000640845
R78212 VSS.n2518 VSS.n2516 0.000638889
R78213 VSS.n21692 VSS.n21689 0.000638889
R78214 VSS.n11416 VSS.n11415 0.000638889
R78215 VSS.n437 VSS.n434 0.000638889
R78216 VSS.n11468 VSS.n11466 0.000638889
R78217 VSS.n420 VSS.n417 0.000638889
R78218 VSS.n11639 VSS.n11638 0.000638889
R78219 VSS.n403 VSS.n400 0.000638889
R78220 VSS.n17238 VSS.n17237 0.000638889
R78221 VSS.n14288 VSS.n14287 0.000638889
R78222 VSS.n17385 VSS.n17384 0.000638889
R78223 VSS.n385 VSS.n382 0.000638889
R78224 VSS.n17396 VSS.n17394 0.000638889
R78225 VSS.n359 VSS.n356 0.000638889
R78226 VSS.n4119 VSS.n4118 0.000638889
R78227 VSS.n21930 VSS.n21927 0.000638889
R78228 VSS.n2929 VSS.n2928 0.000628571
R78229 VSS.n2993 VSS.n2992 0.000628571
R78230 VSS.n3041 VSS.n3040 0.000628571
R78231 VSS.n2574 VSS.n2555 0.000628571
R78232 VSS.n3184 VSS.n3183 0.000628571
R78233 VSS.n2678 VSS.n2677 0.000628571
R78234 VSS.n2722 VSS.n2721 0.000628571
R78235 VSS.n2782 VSS.n2781 0.000628571
R78236 VSS.n2866 VSS.n2865 0.000628571
R78237 VSS.n2931 VSS.n2930 0.000628571
R78238 VSS.n2995 VSS.n2994 0.000628571
R78239 VSS.n3010 VSS.n3009 0.000628571
R78240 VSS.n3043 VSS.n3042 0.000628571
R78241 VSS.n3058 VSS.n3057 0.000628571
R78242 VSS.n2573 VSS.n2572 0.000628571
R78243 VSS.n2571 VSS.n2570 0.000628571
R78244 VSS.n2564 VSS.n2563 0.000628571
R78245 VSS.n5195 VSS.n5194 0.000628571
R78246 VSS.n5246 VSS.n5245 0.000628571
R78247 VSS.n5280 VSS.n5279 0.000628571
R78248 VSS.n4972 VSS.n4966 0.000628571
R78249 VSS.n5142 VSS.n5141 0.000628571
R78250 VSS.n5197 VSS.n5196 0.000628571
R78251 VSS.n5205 VSS.n5204 0.000628571
R78252 VSS.n5248 VSS.n5247 0.000628571
R78253 VSS.n5256 VSS.n5255 0.000628571
R78254 VSS.n5282 VSS.n5281 0.000628571
R78255 VSS.n5291 VSS.n5290 0.000628571
R78256 VSS.n4971 VSS.n4970 0.000628571
R78257 VSS.n4961 VSS.n4960 0.000628571
R78258 VSS.n7181 VSS.n7180 0.000628571
R78259 VSS.n7122 VSS.n7121 0.000628571
R78260 VSS.n7080 VSS.n7079 0.000628571
R78261 VSS.n7519 VSS.n7048 0.000628571
R78262 VSS.n7264 VSS.n7263 0.000628571
R78263 VSS.n7182 VSS.n7178 0.000628571
R78264 VSS.n7167 VSS.n7166 0.000628571
R78265 VSS.n7123 VSS.n7119 0.000628571
R78266 VSS.n7108 VSS.n7107 0.000628571
R78267 VSS.n7081 VSS.n7077 0.000628571
R78268 VSS.n7070 VSS.n7069 0.000628571
R78269 VSS.n7521 VSS.n7520 0.000628571
R78270 VSS.n7532 VSS.n7531 0.000628571
R78271 VSS.n4460 VSS.n4459 0.000628571
R78272 VSS.n4409 VSS.n4408 0.000628571
R78273 VSS.n4374 VSS.n4373 0.000628571
R78274 VSS.n4320 VSS.n4319 0.000628571
R78275 VSS.n4688 VSS.n4687 0.000628571
R78276 VSS.n4513 VSS.n4512 0.000628571
R78277 VSS.n4461 VSS.n4457 0.000628571
R78278 VSS.n4450 VSS.n4449 0.000628571
R78279 VSS.n4410 VSS.n4406 0.000628571
R78280 VSS.n4399 VSS.n4398 0.000628571
R78281 VSS.n4375 VSS.n4371 0.000628571
R78282 VSS.n4364 VSS.n4363 0.000628571
R78283 VSS.n4339 VSS.n4338 0.000628571
R78284 VSS.n4337 VSS.n4336 0.000628571
R78285 VSS.n4330 VSS.n4329 0.000628571
R78286 VSS.n4754 VSS.n2338 0.000628571
R78287 VSS.n17548 VSS.n17547 0.000628571
R78288 VSS.n17490 VSS.n17489 0.000628571
R78289 VSS.n18032 VSS.n18031 0.000628571
R78290 VSS.n17974 VSS.n17970 0.000628571
R78291 VSS.n17865 VSS.n17864 0.000628571
R78292 VSS.n17820 VSS.n17816 0.000628571
R78293 VSS.n17804 VSS.n17803 0.000628571
R78294 VSS.n17775 VSS.n17771 0.000628571
R78295 VSS.n17759 VSS.n17758 0.000628571
R78296 VSS.n17731 VSS.n17730 0.000628571
R78297 VSS.n17729 VSS.n17728 0.000628571
R78298 VSS.n17722 VSS.n17721 0.000628571
R78299 VSS.n17973 VSS.n17972 0.000628571
R78300 VSS.n17819 VSS.n17818 0.000628571
R78301 VSS.n17774 VSS.n17773 0.000628571
R78302 VSS.n17713 VSS.n17709 0.000628571
R78303 VSS.n20400 VSS.n463 0.00062
R78304 VSS.n20371 VSS.n20370 0.00062
R78305 VSS.n20340 VSS.n20339 0.00062
R78306 VSS.n20294 VSS.n20293 0.00062
R78307 VSS.n20399 VSS.n20398 0.00062
R78308 VSS.n20372 VSS.n20367 0.00062
R78309 VSS.n20341 VSS.n20337 0.00062
R78310 VSS.n20295 VSS.n20291 0.00062
R78311 DVSS VSS.n7917 0.00062
R78312 VSS.n11180 VSS.n11179 0.00062
R78313 VSS.n10631 VSS.n10630 0.00062
R78314 VSS.n10678 VSS.n10677 0.00062
R78315 VSS.n10740 VSS.n10739 0.00062
R78316 VSS.n9458 VSS.n9457 0.00062
R78317 VSS.n9783 VSS.n9782 0.00062
R78318 VSS.n9729 VSS.n9728 0.00062
R78319 VSS.n8812 VSS.n8811 0.00062
R78320 VSS.n8924 VSS.n8923 0.00062
R78321 VSS.n9392 VSS.n9391 0.00062
R78322 VSS.n9338 VSS.n9337 0.00062
R78323 VSS.n8814 VSS.n8813 0.00062
R78324 VSS.n8926 VSS.n8925 0.00062
R78325 VSS.n9404 VSS.n9403 0.00062
R78326 VSS.n9393 VSS.n9389 0.00062
R78327 VSS.n9350 VSS.n9349 0.00062
R78328 VSS.n9339 VSS.n9335 0.00062
R78329 VSS.n8443 VSS.n8442 0.00062
R78330 VSS.n8294 VSS.n8293 0.00062
R78331 VSS.n9426 VSS.n9425 0.00062
R78332 VSS.n9460 VSS.n9459 0.00062
R78333 VSS.n9795 VSS.n9794 0.00062
R78334 VSS.n9784 VSS.n9780 0.00062
R78335 VSS.n9741 VSS.n9740 0.00062
R78336 VSS.n9730 VSS.n9726 0.00062
R78337 VSS.n8775 VSS.n8774 0.00062
R78338 VSS.n8751 VSS.n8750 0.00062
R78339 VSS.n11181 VSS.n6163 0.00062
R78340 VSS.n10633 VSS.n10632 0.00062
R78341 VSS.n10659 VSS.n10658 0.00062
R78342 VSS.n10662 VSS.n10661 0.00062
R78343 VSS.n10667 VSS.n10663 0.00062
R78344 VSS.n10673 VSS.n10672 0.00062
R78345 VSS.n10680 VSS.n10679 0.00062
R78346 VSS.n10683 VSS.n10682 0.00062
R78347 VSS.n10721 VSS.n10720 0.00062
R78348 VSS.n10724 VSS.n10723 0.00062
R78349 VSS.n10729 VSS.n10725 0.00062
R78350 VSS.n10735 VSS.n10734 0.00062
R78351 VSS.n10742 VSS.n10741 0.00062
R78352 VSS.n10745 VSS.n10744 0.00062
R78353 VSS.n10806 VSS.n10805 0.00062
R78354 VSS.n10835 VSS.n10834 0.00062
R78355 VSS.n10928 VSS.n10927 0.00062
R78356 VSS.n10938 VSS.n10937 0.00062
R78357 VSS.n10995 VSS.n10994 0.00062
R78358 VSS.n11005 VSS.n11004 0.00062
R78359 VSS.n20233 VSS.n20232 0.00059
R78360 VSS.n11720 VSS.n11719 0.00059
R78361 VSS.n20375 VSS.n20374 0.00059
R78362 VSS.n20344 VSS.n20343 0.00059
R78363 VSS.n20298 VSS.n20297 0.00059
R78364 VSS.n20228 VSS.n20227 0.00059
R78365 VSS.n20223 VSS.n20222 0.00059
R78366 VSS.n10839 VSS.n10838 0.00059
R78367 VSS.n8746 VSS.n8745 0.00059
R78368 VSS.n8289 VSS.n8288 0.00059
R78369 VSS.n8808 VSS.n8807 0.00059
R78370 VSS.n8919 VSS.n8849 0.00059
R78371 VSS.n9005 VSS.n8996 0.00059
R78372 VSS.n9397 VSS.n9396 0.00059
R78373 VSS.n9343 VSS.n9342 0.00059
R78374 VSS.n8284 VSS.n8283 0.00059
R78375 VSS.n8280 VSS.n8279 0.00059
R78376 VSS.n7895 VSS.n7894 0.00059
R78377 VSS.n9421 VSS.n9420 0.00059
R78378 VSS.n9453 VSS.n9452 0.00059
R78379 VSS.n9467 VSS.n9466 0.00059
R78380 VSS.n9788 VSS.n9787 0.00059
R78381 VSS.n9734 VSS.n9733 0.00059
R78382 VSS.n8741 VSS.n8740 0.00059
R78383 VSS.n8737 VSS.n8736 0.00059
R78384 VSS.n7988 VSS.n7987 0.00059
R78385 VSS.n11183 VSS.n6162 0.00059
R78386 VSS.n10626 VSS.n9826 0.00059
R78387 VSS.n10640 VSS.n10639 0.00059
R78388 VSS.n10670 VSS.n10669 0.00059
R78389 VSS.n10672 VSS.n10671 0.00059
R78390 VSS.n10685 VSS.n10684 0.00059
R78391 VSS.n10732 VSS.n10731 0.00059
R78392 VSS.n10734 VSS.n10733 0.00059
R78393 VSS.n10747 VSS.n10746 0.00059
R78394 VSS.n10807 VSS.n10806 0.00059
R78395 VSS.n10810 VSS.n10809 0.00059
R78396 VSS.n10830 VSS.n10829 0.00059
R78397 VSS.n10834 VSS.n10833 0.00059
R78398 VSS.n10845 VSS.n10844 0.00059
R78399 VSS.n10850 VSS.n10849 0.00059
R78400 VSS.n10926 VSS.n10925 0.00059
R78401 VSS.n10941 VSS.n10940 0.00059
R78402 VSS.n10993 VSS.n10992 0.00059
R78403 VSS.n11009 VSS.n11008 0.00059
R78404 VSS.n11040 VSS.n11039 0.00059
R78405 VSS.n4973 DVSS 0.000585714
R78406 VSS.n3526 VSS.n3524 0.000570422
R78407 VSS.n3585 VSS.n3583 0.000570422
R78408 VSS.n3628 VSS.n3626 0.000570422
R78409 VSS.n3206 VSS.n3205 0.000570422
R78410 VSS.n3445 VSS.n3444 0.000570422
R78411 VSS.n3462 VSS.n3461 0.000570422
R78412 VSS.n3480 VSS.n3479 0.000570422
R78413 VSS.n3483 VSS.n3482 0.000570422
R78414 VSS.n3513 VSS.n3512 0.000570422
R78415 VSS.n3527 VSS.n3523 0.000570422
R78416 VSS.n3572 VSS.n3571 0.000570422
R78417 VSS.n3586 VSS.n3582 0.000570422
R78418 VSS.n3615 VSS.n3614 0.000570422
R78419 VSS.n3629 VSS.n3625 0.000570422
R78420 VSS.n3673 VSS.n3672 0.000570422
R78421 VSS.n3664 VSS.n3663 0.000570422
R78422 VSS.n13675 VSS.n13674 0.000564286
R78423 VSS.n13677 VSS.n13676 0.000564286
R78424 VSS.n2554 VSS.n2553 0.000564286
R78425 VSS.n2845 VSS.n2840 0.000564286
R78426 VSS.n2848 VSS.n2847 0.000564286
R78427 VSS.n2852 VSS.n2851 0.000564286
R78428 VSS.n2855 VSS.n2854 0.000564286
R78429 VSS.n2868 VSS.n2867 0.000564286
R78430 VSS.n2940 VSS.n2937 0.000564286
R78431 VSS.n2942 VSS.n2941 0.000564286
R78432 VSS.n3005 VSS.n3001 0.000564286
R78433 VSS.n3007 VSS.n3006 0.000564286
R78434 VSS.n3053 VSS.n3049 0.000564286
R78435 VSS.n3055 VSS.n3054 0.000564286
R78436 VSS.n3080 VSS.n3079 0.000564286
R78437 VSS.n2568 VSS.n2567 0.000564286
R78438 VSS.n5287 VSS.n5285 0.000564286
R78439 VSS.n4965 VSS.n4964 0.000564286
R78440 VSS.n5129 VSS.n5128 0.000564286
R78441 VSS.n5144 VSS.n5143 0.000564286
R78442 VSS.n5191 VSS.n5190 0.000564286
R78443 VSS.n5202 VSS.n5199 0.000564286
R78444 VSS.n5242 VSS.n5241 0.000564286
R78445 VSS.n5253 VSS.n5250 0.000564286
R78446 VSS.n5277 VSS.n5276 0.000564286
R78447 VSS.n5288 VSS.n5284 0.000564286
R78448 VSS.n5309 VSS.n5308 0.000564286
R78449 VSS.n7172 VSS.n7170 0.000564286
R78450 VSS.n7113 VSS.n7111 0.000564286
R78451 VSS.n7538 VSS.n7534 0.000564286
R78452 VSS.n7218 VSS.n7217 0.000564286
R78453 VSS.n7215 VSS.n7214 0.000564286
R78454 VSS.n7186 VSS.n7185 0.000564286
R78455 VSS.n7174 VSS.n7173 0.000564286
R78456 VSS.n7127 VSS.n7126 0.000564286
R78457 VSS.n7115 VSS.n7114 0.000564286
R78458 VSS.n7084 VSS.n7083 0.000564286
R78459 VSS.n7075 VSS.n7074 0.000564286
R78460 VSS.n7052 VSS.n7051 0.000564286
R78461 VSS.n7540 VSS.n7539 0.000564286
R78462 VSS.n4318 VSS.n4317 0.000564286
R78463 VSS.n4526 VSS.n4525 0.000564286
R78464 VSS.n4511 VSS.n4510 0.000564286
R78465 VSS.n4464 VSS.n4463 0.000564286
R78466 VSS.n4455 VSS.n4454 0.000564286
R78467 VSS.n4413 VSS.n4412 0.000564286
R78468 VSS.n4404 VSS.n4403 0.000564286
R78469 VSS.n4378 VSS.n4377 0.000564286
R78470 VSS.n4369 VSS.n4368 0.000564286
R78471 VSS.n4343 VSS.n4342 0.000564286
R78472 VSS.n4334 VSS.n4333 0.000564286
R78473 VSS.n18056 VSS.n18055 0.000564286
R78474 VSS.n18049 VSS.n18048 0.000564286
R78475 VSS.n18046 VSS.n18045 0.000564286
R78476 VSS.n18043 VSS.n18042 0.000564286
R78477 VSS.n18030 VSS.n18029 0.000564286
R78478 VSS.n17978 VSS.n17977 0.000564286
R78479 VSS.n17871 VSS.n17870 0.000564286
R78480 VSS.n17867 VSS.n17866 0.000564286
R78481 VSS.n17824 VSS.n17823 0.000564286
R78482 VSS.n17810 VSS.n17809 0.000564286
R78483 VSS.n17806 VSS.n17805 0.000564286
R78484 VSS.n17779 VSS.n17778 0.000564286
R78485 VSS.n17765 VSS.n17764 0.000564286
R78486 VSS.n17761 VSS.n17760 0.000564286
R78487 VSS.n17735 VSS.n17734 0.000564286
R78488 VSS.n17726 VSS.n17725 0.000564286
R78489 VSS.n17708 VSS.n17707 0.000564286
R78490 VSS.n14125 VSS.n14119 0.000564286
R78491 VSS.n20172 VSS.n20171 0.00056
R78492 VSS.n686 VSS.n685 0.00056
R78493 VSS.n20501 VSS.n20500 0.00056
R78494 VSS.n20547 VSS.n20539 0.00056
R78495 VSS.n20226 VSS.n20225 0.00056
R78496 VSS.n20173 VSS.n20168 0.00056
R78497 VSS.n728 VSS.n727 0.00056
R78498 VSS.n687 VSS.n460 0.00056
R78499 VSS.n20584 VSS.n20583 0.00056
R78500 VSS.n20569 VSS.n20568 0.00056
R78501 VSS.n20563 VSS.n20562 0.00056
R78502 VSS.n20546 VSS.n20545 0.00056
R78503 VSS.n20534 VSS.n20533 0.00056
R78504 VSS.n10922 VSS.n10921 0.00056
R78505 VSS.n10989 VSS.n10988 0.00056
R78506 VSS.n11044 VSS.n11043 0.00056
R78507 VSS.n6377 VSS.n6370 0.00056
R78508 VSS.n8089 VSS.n8088 0.00056
R78509 VSS.n8029 VSS.n8028 0.00056
R78510 VSS.n7984 VSS.n7983 0.00056
R78511 VSS.n7951 VSS.n7941 0.00056
R78512 VSS.n6773 VSS.n6772 0.00056
R78513 VSS.n6713 VSS.n6712 0.00056
R78514 VSS.n7891 VSS.n7890 0.00056
R78515 VSS.n7854 VSS.n7023 0.00056
R78516 VSS.n9395 VSS.n9394 0.00056
R78517 VSS.n9341 VSS.n9340 0.00056
R78518 VSS.n8282 VSS.n8281 0.00056
R78519 VSS.n6774 VSS.n6770 0.00056
R78520 VSS.n6759 VSS.n6758 0.00056
R78521 VSS.n6714 VSS.n6710 0.00056
R78522 VSS.n6699 VSS.n6698 0.00056
R78523 VSS.n7892 VSS.n7888 0.00056
R78524 VSS.n7877 VSS.n7876 0.00056
R78525 VSS.n7853 VSS.n7852 0.00056
R78526 VSS.n7037 VSS.n7036 0.00056
R78527 VSS.n9786 VSS.n9785 0.00056
R78528 VSS.n9732 VSS.n9731 0.00056
R78529 VSS.n8739 VSS.n8738 0.00056
R78530 VSS.n8090 VSS.n8086 0.00056
R78531 VSS.n8075 VSS.n8074 0.00056
R78532 VSS.n8030 VSS.n8026 0.00056
R78533 VSS.n8015 VSS.n8014 0.00056
R78534 VSS.n7985 VSS.n7981 0.00056
R78535 VSS.n7970 VSS.n7969 0.00056
R78536 VSS.n7950 VSS.n7949 0.00056
R78537 VSS.n7935 VSS.n7934 0.00056
R78538 VSS.n10675 VSS.n10674 0.00056
R78539 VSS.n10737 VSS.n10736 0.00056
R78540 VSS.n10814 VSS.n10810 0.00056
R78541 VSS.n10847 VSS.n10846 0.00056
R78542 VSS.n10924 VSS.n10923 0.00056
R78543 VSS.n10939 VSS.n10938 0.00056
R78544 VSS.n10991 VSS.n10990 0.00056
R78545 VSS.n11046 VSS.n11045 0.00056
R78546 VSS.n6376 VSS.n6375 0.00056
R78547 VSS.n6364 VSS.n6363 0.00056
R78548 VSS.n13852 VSS 0.000557143
R78549 VSS.n20505 VSS.n20503 0.00053
R78550 VSS.n20538 VSS.n20537 0.00053
R78551 VSS.n20240 VSS.n20239 0.00053
R78552 VSS.n20224 VSS.n20223 0.00053
R78553 VSS.n20176 VSS.n20175 0.00053
R78554 VSS.n733 VSS.n732 0.00053
R78555 VSS.n691 VSS.n690 0.00053
R78556 VSS.n20589 VSS.n20588 0.00053
R78557 VSS.n20572 VSS.n20571 0.00053
R78558 VSS.n20566 VSS.n20565 0.00053
R78559 VSS.n20541 VSS.n20540 0.00053
R78560 VSS.n10933 VSS.n10931 0.00053
R78561 VSS.n11000 VSS.n10998 0.00053
R78562 VSS.n11053 VSS.n11051 0.00053
R78563 VSS.n6367 VSS.n6360 0.00053
R78564 VSS.n8080 VSS.n8078 0.00053
R78565 VSS.n8020 VSS.n8018 0.00053
R78566 VSS.n7975 VSS.n7973 0.00053
R78567 VSS.n7938 VSS.n7931 0.00053
R78568 VSS.n6764 VSS.n6762 0.00053
R78569 VSS.n6704 VSS.n6702 0.00053
R78570 VSS.n7882 VSS.n7880 0.00053
R78571 VSS.n7043 VSS.n7039 0.00053
R78572 VSS.n8304 VSS.n8303 0.00053
R78573 VSS.n6778 VSS.n6777 0.00053
R78574 VSS.n6766 VSS.n6765 0.00053
R78575 VSS.n6761 VSS.n6760 0.00053
R78576 VSS.n6718 VSS.n6717 0.00053
R78577 VSS.n6706 VSS.n6705 0.00053
R78578 VSS.n6701 VSS.n6700 0.00053
R78579 VSS.n7896 VSS.n7895 0.00053
R78580 VSS.n7884 VSS.n7883 0.00053
R78581 VSS.n7024 VSS.n7008 0.00053
R78582 VSS.n7045 VSS.n7044 0.00053
R78583 VSS.n8761 VSS.n8760 0.00053
R78584 VSS.n8094 VSS.n8093 0.00053
R78585 VSS.n8082 VSS.n8081 0.00053
R78586 VSS.n8077 VSS.n8076 0.00053
R78587 VSS.n8034 VSS.n8033 0.00053
R78588 VSS.n8022 VSS.n8021 0.00053
R78589 VSS.n8017 VSS.n8016 0.00053
R78590 VSS.n7989 VSS.n7988 0.00053
R78591 VSS.n7977 VSS.n7976 0.00053
R78592 VSS.n7946 VSS.n7945 0.00053
R78593 VSS.n7937 VSS.n7933 0.00053
R78594 VSS.n10826 VSS.n10822 0.00053
R78595 VSS.n10870 VSS.n10869 0.00053
R78596 VSS.n10874 VSS.n10873 0.00053
R78597 VSS.n10917 VSS.n10916 0.00053
R78598 VSS.n10934 VSS.n10930 0.00053
R78599 VSS.n10936 VSS.n10935 0.00053
R78600 VSS.n10984 VSS.n10983 0.00053
R78601 VSS.n11001 VSS.n10997 0.00053
R78602 VSS.n11003 VSS.n11002 0.00053
R78603 VSS.n11039 VSS.n11038 0.00053
R78604 VSS.n11054 VSS.n11050 0.00053
R78605 VSS.n6372 VSS.n6371 0.00053
R78606 VSS.n6366 VSS.n6362 0.00053
R78607 VSS.n20548 DVSS 0.000526667
C0 DVDD VDD 48.2f
C1 DVDD ASIG5V 0.626p
C2 DVSS VDD 51f
C3 DVSS ASIG5V 0.486p
C4 ASIG5V VDD 21.9f
C5 DVSS DVDD 1.56p
.ends


* NGSPICE file created from waffle_1984.ext - technology: gf180mcuD

.subckt waffle_1984
X0 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X2 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X3 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X4 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X5 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X6 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X7 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X8 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X9 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X10 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X11 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X12 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X13 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X14 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X15 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X16 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X17 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X18 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X19 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X20 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X21 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X22 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X23 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X24 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X25 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=2.56795p ps=9.38u w=4.38u l=0.5u
X26 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X27 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X28 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X29 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X30 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X31 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X32 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X33 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X34 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X35 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X36 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X37 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X38 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X39 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X40 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X41 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X42 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X43 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X44 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X45 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X46 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X47 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X48 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X49 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X50 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X51 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X52 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X53 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X54 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X55 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X56 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X57 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X58 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X59 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X60 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X61 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X62 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X63 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X64 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X65 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X66 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X67 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X68 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X69 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X70 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X71 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X72 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X73 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X74 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X75 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X76 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X77 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X78 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X79 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X80 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X81 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X82 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X83 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X84 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X85 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X86 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X87 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X88 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X89 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X90 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X91 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X92 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X93 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X94 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X95 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X96 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X97 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X98 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X99 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X100 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X101 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X102 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X103 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X104 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X105 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X106 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X107 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X108 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X109 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X110 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X111 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X112 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X113 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X114 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X115 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X116 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X117 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X118 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X119 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X120 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X121 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X122 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X123 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X124 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X125 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X126 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X127 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X128 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X129 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X130 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X131 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X132 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X133 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X134 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X135 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X136 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X137 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X138 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X139 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X140 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X141 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X142 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X143 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X144 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X145 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X146 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X147 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X148 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X149 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X150 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X151 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X152 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X153 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X154 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X155 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X156 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X157 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X158 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X159 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X160 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X161 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X162 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X163 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X164 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X165 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X166 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X167 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X168 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X169 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X170 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X171 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X172 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X173 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X174 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X175 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X176 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X177 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X178 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X179 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X180 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X181 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X182 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X183 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X184 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X185 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X186 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X187 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X188 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X189 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X190 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X191 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X192 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X193 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X194 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X195 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X196 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X197 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X198 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X199 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X200 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X201 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X202 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X203 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X204 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X205 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X206 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X207 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X208 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X209 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X210 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X211 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X212 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X213 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X214 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X215 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X216 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X217 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X218 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X219 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X220 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X221 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X222 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X223 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X224 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X225 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X226 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X227 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X228 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X229 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X230 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X231 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X232 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X233 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X234 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X235 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X236 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X237 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X238 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X239 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X240 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X241 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X242 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X243 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X244 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X245 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X246 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X247 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X248 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X249 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X250 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X251 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X252 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X253 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X254 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X255 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X256 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X257 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X258 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X259 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X260 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X261 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X262 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X263 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X264 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X265 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X266 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X267 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X268 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X269 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X270 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X271 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X272 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X273 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X274 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X275 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X276 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X277 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X278 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X279 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X280 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X281 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X282 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X283 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X284 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X285 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X286 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X287 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X288 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X289 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X290 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X291 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X292 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X293 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X294 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X295 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X296 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X297 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X298 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X299 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X300 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X301 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X302 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X303 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X304 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X305 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X306 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X307 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X308 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X309 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X310 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X311 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X312 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X313 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X314 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X315 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X316 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X317 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X318 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X319 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X320 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X321 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X322 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X323 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X324 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X325 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X326 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X327 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X328 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X329 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X330 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X331 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X332 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X333 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X334 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X335 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X336 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X337 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X338 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X339 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X340 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X341 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X342 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X343 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X344 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X345 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X346 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X347 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X348 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X349 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X350 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X351 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X352 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X353 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X354 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X355 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X356 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X357 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X358 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X359 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X360 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X361 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X362 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X363 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X364 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X365 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X366 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X367 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X368 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X369 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X370 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X371 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X372 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X373 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X374 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X375 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X376 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X377 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X378 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X379 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X380 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X381 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X382 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X383 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X384 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X385 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X386 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X387 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X388 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X389 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X390 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X391 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X392 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X393 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X394 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X395 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X396 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X397 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X398 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X399 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X400 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X401 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X402 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X403 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X404 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X405 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X406 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X407 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X408 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X409 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X410 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X411 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X412 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X413 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X414 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X415 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X416 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X417 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X418 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X419 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X420 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X421 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X422 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X423 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X424 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X425 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X426 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X427 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X428 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X429 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X430 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X431 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X432 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X433 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X434 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X435 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X436 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X437 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X438 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X439 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X440 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X441 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X442 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X443 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X444 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X445 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X446 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X447 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X448 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X449 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X450 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X451 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X452 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X453 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X454 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X455 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X456 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X457 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X458 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X459 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X460 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X461 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X462 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X463 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X464 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X465 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X466 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X467 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X468 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X469 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X470 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X471 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X472 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X473 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X474 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X475 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X476 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X477 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X478 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X479 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X480 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X481 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X482 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X483 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X484 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X485 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X486 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X487 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X488 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X489 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X490 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X491 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X492 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X493 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X494 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X495 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X496 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X497 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X498 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X499 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X500 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X501 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X502 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X503 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X504 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X505 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X506 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X507 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X508 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X509 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X510 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X511 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X512 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X513 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X514 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X515 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X516 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X517 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X518 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X519 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X520 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X521 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X522 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X523 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X524 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X525 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X526 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X527 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X528 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X529 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X530 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X531 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X532 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X533 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X534 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X535 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X536 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X537 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X538 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X539 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X540 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X541 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X542 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X543 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X544 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X545 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X546 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X547 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X548 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X549 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X550 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X551 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X552 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X553 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X554 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X555 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X556 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X557 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X558 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X559 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X560 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X561 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X562 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X563 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X564 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X565 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X566 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X567 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X568 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X569 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X570 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X571 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X572 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X573 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X574 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X575 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X576 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X577 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X578 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X579 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X580 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X581 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X582 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X583 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X584 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X585 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X586 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X587 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X588 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X589 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X590 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X591 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X592 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X593 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X594 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X595 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X596 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X597 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X598 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X599 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X600 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X601 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X602 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X603 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X604 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X605 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X606 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X607 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X608 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X609 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X610 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X611 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X612 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X613 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X614 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X615 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X616 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X617 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X618 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X619 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X620 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X621 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X622 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X623 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X624 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X625 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X626 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X627 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X628 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X629 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X630 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X631 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X632 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X633 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X634 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X635 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X636 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X637 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X638 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X639 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X640 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X641 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X642 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X643 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X644 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X645 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X646 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X647 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X648 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X649 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X650 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X651 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X652 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X653 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X654 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X655 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X656 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X657 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X658 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X659 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X660 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X661 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X662 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X663 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X664 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X665 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X666 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X667 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X668 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X669 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X670 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X671 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X672 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X673 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X674 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X675 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X676 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X677 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X678 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X679 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X680 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X681 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X682 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X683 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X684 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X685 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X686 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X687 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X688 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X689 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X690 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X691 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X692 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X693 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X694 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X695 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X696 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X697 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X698 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X699 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X700 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X701 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X702 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X703 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X704 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X705 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X706 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X707 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X708 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X709 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X710 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X711 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X712 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X713 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X714 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X715 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X716 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X717 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X718 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X719 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X720 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X721 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X722 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X723 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X724 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X725 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X726 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X727 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X728 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X729 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X730 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X731 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X732 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X733 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X734 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X735 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X736 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X737 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X738 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X739 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X740 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X741 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X742 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X743 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X744 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X745 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X746 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X747 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X748 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X749 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X750 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X751 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X752 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X753 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X754 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X755 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X756 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X757 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X758 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X759 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X760 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X761 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X762 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X763 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X764 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X765 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X766 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X767 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X768 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X769 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X770 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X771 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X772 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X773 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X774 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X775 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X776 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X777 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X778 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X779 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X780 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X781 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X782 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X783 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X784 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X785 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X786 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X787 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X788 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X789 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X790 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X791 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X792 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X793 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X794 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X795 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X796 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X797 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X798 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X799 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X800 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X801 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X802 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X803 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X804 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X805 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X806 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X807 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X808 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X809 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X810 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X811 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X812 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X813 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X814 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X815 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X816 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X817 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X818 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X819 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X820 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X821 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X822 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X823 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X824 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X825 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X826 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X827 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X828 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X829 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X830 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X831 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X832 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X833 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X834 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X835 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X836 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X837 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X838 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X839 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X840 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X841 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X842 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X843 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X844 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X845 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X846 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X847 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X848 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X849 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X850 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X851 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X852 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X853 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X854 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X855 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X856 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X857 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X858 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X859 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X860 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X861 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X862 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X863 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X864 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X865 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X866 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X867 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X868 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X869 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X870 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X871 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X872 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X873 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X874 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X875 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X876 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X877 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X878 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X879 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X880 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X881 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X882 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X883 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X884 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X885 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X886 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X887 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X888 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X889 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X890 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X891 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X892 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X893 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X894 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X895 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X896 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X897 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X898 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X899 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X900 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X901 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X902 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X903 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X904 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X905 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X906 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X907 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X908 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X909 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X910 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X911 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X912 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X913 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X914 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X915 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X916 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X917 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X918 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X919 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X920 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X921 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X922 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X923 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X924 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X925 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X926 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X927 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X928 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X929 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X930 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X931 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=2.56795p ps=9.38u w=4.38u l=0.5u
X932 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X933 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X934 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X935 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X936 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X937 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X938 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X939 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X940 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X941 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X942 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X943 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X944 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X945 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X946 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X947 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X948 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X949 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X950 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X951 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X952 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X953 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X954 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X955 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X956 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X957 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X958 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X959 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X960 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X961 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X962 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X963 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X964 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X965 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X966 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=2.56795p ps=9.38u w=4.38u l=0.5u
X967 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X968 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X969 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X970 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X971 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X972 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X973 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X974 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X975 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X976 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X977 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X978 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X979 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X980 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X981 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X982 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X983 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X984 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X985 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X986 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X987 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X988 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X989 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X990 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X991 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X992 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X993 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X994 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X995 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X996 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X997 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X998 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X999 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1000 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1001 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1002 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1003 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1004 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1005 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1006 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1007 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1008 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1009 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1010 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1011 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1012 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1013 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1014 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1015 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1016 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1017 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1018 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1019 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1020 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1021 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1022 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1023 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1024 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1025 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1026 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=2.56795p ps=9.38u w=4.38u l=0.5u
X1027 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1028 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1029 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1030 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1031 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1032 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1033 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1034 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1035 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1036 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1037 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1038 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1039 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1040 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1041 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1042 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1043 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1044 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1045 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1046 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1047 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1048 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1049 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1050 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1051 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1052 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1053 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1054 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1055 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1056 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1057 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1058 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1059 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1060 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1061 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1062 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1063 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1064 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1065 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1066 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1067 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=2.56795p pd=9.38u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1068 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1069 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1070 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1071 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1072 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1073 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1074 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1075 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1076 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1077 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1078 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1079 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1080 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1081 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1082 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1083 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1084 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1085 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1086 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1087 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1088 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1089 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1090 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1091 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1092 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1093 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1094 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1095 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1096 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1097 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1098 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1099 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1100 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1101 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1102 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1103 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1104 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1105 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1106 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1107 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1108 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1109 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1110 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1111 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1112 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1113 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1114 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1115 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1116 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1117 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1118 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1119 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1120 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1121 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1122 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1123 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1124 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1125 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1126 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1127 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1128 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1129 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1130 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1131 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1132 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1133 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1134 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1135 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1136 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1137 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1138 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1139 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1140 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1141 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1142 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1143 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1144 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1145 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1146 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1147 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1148 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=2.56795p pd=9.38u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1149 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1150 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1151 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1152 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1153 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1154 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1155 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1156 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1157 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1158 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1159 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1160 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1161 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1162 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1163 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1164 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1165 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1166 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1167 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1168 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1169 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1170 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1171 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1172 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1173 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1174 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1175 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1176 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1177 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1178 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1179 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1180 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1181 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1182 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1183 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1184 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1185 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1186 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1187 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1188 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1189 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1190 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1191 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1192 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1193 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1194 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1195 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1196 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1197 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1198 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1199 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1200 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1201 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1202 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1203 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1204 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1205 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1206 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1207 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1208 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1209 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1210 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1211 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1212 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1213 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1214 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1215 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1216 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1217 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1218 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1219 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1220 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1221 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1222 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1223 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1224 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1225 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1226 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1227 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1228 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1229 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1230 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1231 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1232 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1233 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1234 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1235 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1236 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1237 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1238 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1239 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1240 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1241 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1242 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1243 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1244 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1245 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1246 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1247 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1248 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1249 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1250 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1251 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1252 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1253 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1254 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1255 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1256 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1257 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1258 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1259 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1260 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1261 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1262 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1263 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1264 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1265 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1266 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1267 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1268 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1269 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1270 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1271 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1272 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1273 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1274 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1275 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1276 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1277 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1278 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1279 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1280 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1281 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1282 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1283 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1284 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1285 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1286 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1287 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1288 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1289 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1290 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1291 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1292 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1293 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1294 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1295 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1296 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1297 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1298 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1299 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1300 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1301 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1302 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1303 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1304 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1305 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1306 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1307 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1308 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1309 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1310 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1311 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1312 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1313 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1314 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1315 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1316 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1317 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1318 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1319 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1320 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1321 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1322 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1323 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1324 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1325 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1326 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1327 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1328 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1329 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1330 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1331 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1332 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1333 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1334 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1335 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1336 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1337 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1338 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1339 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1340 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1341 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1342 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1343 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1344 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1345 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1346 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1347 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1348 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1349 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1350 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1351 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1352 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1353 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1354 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1355 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1356 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1357 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1358 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1359 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1360 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1361 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1362 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1363 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=2.56795p pd=9.38u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1364 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1365 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1366 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1367 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1368 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1369 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1370 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1371 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1372 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1373 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1374 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1375 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1376 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1377 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1378 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1379 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1380 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1381 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1382 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1383 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1384 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1385 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1386 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1387 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1388 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1389 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1390 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1391 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1392 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1393 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1394 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1395 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1396 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1397 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1398 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1399 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1400 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1401 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1402 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1403 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1404 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1405 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1406 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1407 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1408 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1409 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1410 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1411 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1412 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1413 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1414 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1415 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1416 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1417 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1418 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1419 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1420 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1421 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1422 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1423 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1424 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1425 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1426 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1427 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1428 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1429 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1430 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1431 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1432 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1433 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1434 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1435 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1436 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1437 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1438 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1439 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1440 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1441 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1442 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1443 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1444 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1445 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1446 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1447 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1448 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1449 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1450 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1451 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1452 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1453 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1454 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1455 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1456 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1457 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1458 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1459 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1460 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1461 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1462 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1463 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1464 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1465 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1466 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1467 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1468 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1469 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1470 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1471 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1472 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1473 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1474 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1475 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1476 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1477 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1478 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1479 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1480 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1481 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1482 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1483 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1484 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1485 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1486 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1487 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1488 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1489 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1490 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1491 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1492 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1493 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1494 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1495 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1496 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1497 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1498 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1499 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1500 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1501 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1502 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1503 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1504 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1505 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1506 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1507 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1508 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1509 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1510 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1511 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1512 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1513 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1514 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1515 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1516 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1517 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1518 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1519 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1520 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1521 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1522 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1523 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1524 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1525 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1526 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1527 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1528 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1529 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1530 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1531 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1532 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1533 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1534 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1535 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1536 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1537 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1538 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1539 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1540 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1541 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1542 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1543 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1544 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1545 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1546 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1547 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1548 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1549 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1550 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1551 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1552 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1553 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1554 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1555 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1556 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1557 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1558 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1559 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1560 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1561 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1562 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1563 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1564 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1565 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1566 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1567 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1568 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1569 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1570 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1571 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1572 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1573 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1574 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1575 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1576 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1577 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1578 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1579 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1580 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1581 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1582 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1583 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1584 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1585 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1586 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1587 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1588 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1589 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1590 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1591 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1592 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1593 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1594 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1595 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1596 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1597 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1598 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1599 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1600 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1601 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1602 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1603 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1604 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1605 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1606 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1607 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1608 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1609 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1610 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1611 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1612 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1613 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1614 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1615 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1616 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1617 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1618 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1619 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1620 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1621 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1622 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1623 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1624 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1625 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1626 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1627 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1628 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1629 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1630 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1631 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1632 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1633 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1634 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1635 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1636 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1637 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1638 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1639 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1640 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1641 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1642 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1643 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1644 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1645 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1646 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1647 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1648 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1649 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1650 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1651 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1652 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1653 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1654 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1655 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1656 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1657 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1658 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1659 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1660 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1661 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1662 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1663 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1664 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1665 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1666 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1667 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1668 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1669 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1670 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1671 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1672 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1673 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1674 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1675 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1676 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1677 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1678 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1679 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1680 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1681 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1682 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1683 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1684 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1685 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1686 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1687 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1688 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1689 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1690 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1691 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1692 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1693 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1694 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1695 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1696 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1697 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1698 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1699 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1700 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1701 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1702 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1703 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1704 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1705 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1706 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1707 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1708 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1709 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1710 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1711 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1712 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1713 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1714 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1715 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1716 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1717 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1718 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1719 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1720 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1721 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1722 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1723 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1724 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1725 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1726 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1727 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1728 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1729 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1730 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1731 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1732 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1733 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1734 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1735 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1736 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1737 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1738 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1739 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1740 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1741 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1742 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1743 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1744 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1745 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1746 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1747 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1748 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1749 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1750 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1751 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1752 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1753 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1754 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1755 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1756 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1757 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1758 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1759 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1760 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1761 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1762 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1763 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1764 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1765 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1766 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1767 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1768 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1769 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1770 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1771 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1772 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1773 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1774 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1775 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1776 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1777 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1778 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1779 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1780 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1781 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1782 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1783 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1784 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1785 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1786 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1787 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1788 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1789 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1790 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1791 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1792 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1793 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1794 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1795 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1796 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1797 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1798 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1799 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1800 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1801 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1802 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1803 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1804 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1805 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1806 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1807 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1808 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=2.56795p pd=9.38u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1809 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1810 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1811 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1812 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1813 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1814 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1815 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1816 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1817 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1818 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1819 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1820 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1821 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1822 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1823 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1824 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1825 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1826 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1827 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1828 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1829 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1830 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1831 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1832 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1833 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1834 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1835 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1836 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1837 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1838 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1839 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1840 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1841 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1842 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1843 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1844 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1845 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1846 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1847 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1848 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1849 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1850 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1851 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1852 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1853 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1854 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1855 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1856 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1857 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1858 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1859 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1860 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1861 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1862 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1863 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1864 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1865 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1866 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1867 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1868 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1869 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1870 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1871 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1872 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1873 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1874 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1875 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1876 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1877 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1878 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1879 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1880 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1881 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1882 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1883 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1884 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1885 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1886 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1887 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1888 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1889 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1890 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1891 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1892 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1893 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1894 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1895 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1896 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1897 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1898 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1899 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1900 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1901 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1902 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1903 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1904 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1905 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1906 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1907 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1908 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1909 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1910 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1911 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1912 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1913 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1914 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1915 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1916 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1917 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1918 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1919 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1920 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1921 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1922 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1923 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1924 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1925 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1926 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1927 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1928 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1929 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1930 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1931 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1932 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1933 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1934 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1935 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1936 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1937 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1938 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1939 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1940 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1941 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1942 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1943 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1944 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1945 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1946 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1947 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1948 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1949 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1950 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1951 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1952 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1953 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1954 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1955 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1956 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1957 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1958 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1959 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1960 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1961 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1962 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1963 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1964 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1965 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1966 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1967 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1968 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1969 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1970 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1971 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1972 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1973 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1974 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1975 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1976 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1977 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1978 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1979 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1980 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1981 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
X1982 external-guardring-trck-3-5.5-10-216.0_0/S gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/D external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=3.8399p pd=13.78u as=3.8399p ps=13.78u w=4.38u l=0.5u
X1983 external-guardring-trck-3-5.5-10-216.0_0/D gate_mesh-5.5-0.5-2.25_0/G external-guardring-trck-3-5.5-10-216.0_0/S external-guardring-trck-3-5.5-10-216.0_0/S pfet_03v3 ad=5.0878p pd=17.599998u as=5.0878p ps=17.599998u w=4.38u l=0.5u
.ends


** sch_path: /home/tsuchiya/chipathon/chipathon2023/BGR/xschem/bgr_diode.sch
.subckt bgr_diode vss vdd vout
*.PININFO vdd:B vss:B vout:O
M5 net2 net1 net4 net4 nfet_03v3_dn L=1.12u W=11.2u nf=1 m=30
M6 net2 net2 vdd vdd pfet_03v3 L=1.12u W=11.2u nf=1 m=30
M7 net1 net1 net3 net3 nfet_03v3_dn L=1.12u W=11.2u nf=1 m=30
M8 net1 net2 vdd vdd pfet_03v3 L=1.12u W=11.2u nf=1 m=30
Q1 net5 net5 vss vss npn_10p00x10p00 m=1
Q20 net6 net6 vss vss npn_10p00x10p00 m=1
Q21 net6 net6 vss vss npn_10p00x10p00 m=1
Q22 net6 net6 vss vss npn_10p00x10p00 m=1
Q23 net6 net6 vss vss npn_10p00x10p00 m=1
Q24 net6 net6 vss vss npn_10p00x10p00 m=1
Q25 net6 net6 vss vss npn_10p00x10p00 m=1
Q26 net6 net6 vss vss npn_10p00x10p00 m=1
Q27 net6 net6 vss vss npn_10p00x10p00 m=1
Q28 net6 net6 vss vss npn_10p00x10p00 m=1
Q29 net6 net6 vss vss npn_10p00x10p00 m=1
Q2a net6 net6 vss vss npn_10p00x10p00 m=1
Q2b net6 net6 vss vss npn_10p00x10p00 m=1
Q2c net6 net6 vss vss npn_10p00x10p00 m=1
Q2d net6 net6 vss vss npn_10p00x10p00 m=1
Q2e net6 net6 vss vss npn_10p00x10p00 m=1
Q2f net6 net6 vss vss npn_10p00x10p00 m=1
M1 vout net2 vdd vdd pfet_03v3 L=1.12u W=11.2u nf=1 m=30
Q3 net7 net7 vss vss npn_10p00x10p00 m=1
R1 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R2 net6 net4 vss ppolyf_u W=1.6u L=0.8u m=1
R3 net7 vout vss ppolyf_u W=1.6u L=5.4u m=1
R4 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R5 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R6 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R7 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R8 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R9 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R10 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R11 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
R12 net5 net3 vss ppolyf_u W=1.6u L=0.8u m=1
.ends
.end

* Extracted by KLayout with GF180MCU LVS runset on : 03/02/2024 16:29

.SUBCKT resistor B OUT1 OUT2 IN2 IN1
R$1 B B B 3500 ppolyf_u r_length=20U r_width=2U
R$12 OUT2 IN2 B 42000 ppolyf_u r_length=120U r_width=1U
R$16 OUT1 IN1 B 70000 ppolyf_u r_length=200U r_width=1U
.ENDS resistor

* NGSPICE file created from sar.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_455_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_68# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X5 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6 VSS a_36_68# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 VDD a_36_68# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 VDD Q CLK VSS D VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1 Q a_2304_115# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X3 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X5 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X6 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X7 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X9 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X10 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X11 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X12 Q a_2304_115# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X13 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X14 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X15 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X17 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X18 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X19 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X20 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X21 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X22 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X23 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A2 VDD VNW pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VNW VPW
X0 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 Z VSS VDD I VNW VPW
X0 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X1 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X3 a_224_552# I VSS VPW nfet_06v0 ad=0.2662p pd=2.09u as=0.2662p ps=2.09u w=0.605u l=0.6u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X8 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.2002p ps=1.79u w=0.455u l=0.6u
X9 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X10 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 B1 C VDD VSS ZN A1 A2 B2 VNW VPW
X0 a_692_68# C a_36_68# VPW nfet_06v0 ad=0.246p pd=1.42u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 a_932_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.38575p ps=1.92u w=1.22u l=0.5u
X2 VSS B2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 ZN A2 a_692_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.246p ps=1.42u w=0.82u l=0.6u
X4 a_244_472# B2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.6588p ps=3.52u w=1.22u l=0.5u
X5 ZN A1 a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6 VDD C ZN VNW pfet_06v0 ad=0.38575p pd=1.92u as=0.3952p ps=1.94u w=0.945u l=0.5u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.3952p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 a_36_68# B1 VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_692_68# A1 ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D VDD VSS CLK Q VNW VPW
X0 VSS a_2304_115# Q VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS CLK a_36_151# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2 Q a_2304_115# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X4 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X8 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 VDD a_2304_115# Q VNW pfet_06v0 ad=0.854p pd=3.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X12 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 Q a_2304_115# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X15 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X16 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X17 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X18 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X19 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X21 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X22 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X23 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X24 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X25 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VNW VPW
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.234325p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VPW nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X1 a_428_148# A2 a_244_148# VPW nfet_06v0 ad=79.799995f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VPW nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VPW nfet_06v0 ad=0.2424p pd=1.635u as=79.799995f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VPW nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 Z VSS VDD I VNW VPW
X0 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3 a_224_552# I VDD VNW pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X4 VDD I a_224_552# VNW pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X7 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X10 VSS a_224_552# Z VPW nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X11 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X12 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X13 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X15 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X16 VDD I a_224_552# VNW pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X17 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X18 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X19 Z a_224_552# VSS VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X20 Z a_224_552# VDD VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X21 a_224_552# I VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X22 VSS a_224_552# Z VPW nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.4087p pd=1.89u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.3477p pd=1.79u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 VDD VSS Z I VNW VPW
X0 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X11 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X12 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X13 VDD a_224_552# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X15 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X16 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X17 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X18 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X19 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X20 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X21 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X22 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X23 VSS I a_224_552# VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X24 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X25 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X26 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X27 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X28 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X29 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X30 a_224_552# I VSS VPW nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X31 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X32 VSS a_224_552# Z VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X33 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X34 VSS a_224_552# Z VPW nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X35 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X36 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X37 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X38 Z a_224_552# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X39 a_224_552# I VDD VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X40 a_224_552# I VSS VPW nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X41 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X42 VDD I a_224_552# VNW pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X43 VDD a_224_552# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X44 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X45 Z a_224_552# VSS VPW nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VNW VPW
X0 VSS B a_36_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VNW VPW
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5 VSS B ZN VPW nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_728_472# a_56_604# VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X1 Z A1 a_728_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2 VSS A1 a_56_604# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3 a_728_472# A2 Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4 Z a_56_604# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X5 VSS A2 a_952_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6 a_244_604# A2 a_56_604# VNW pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X7 a_56_604# A2 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X8 a_952_68# A1 Z VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 VDD A1 a_244_604# VNW pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 Z I VDD VSS VNW VPW
X0 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2 VDD a_224_472# Z VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3 a_224_472# I VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 VDD I a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_472# Z VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7 VSS a_224_472# Z VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8 VSS a_224_472# Z VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X9 a_224_472# I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X10 VSS I a_224_472# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 Z a_224_472# VSS VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VPW nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VPW nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VPW nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3 VSS I a_36_113# VPW nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VPW nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VPW nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VPW nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VPW nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 B C VDD VSS ZN A1 A2 VNW VPW
X0 a_692_68# B a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X3 VDD B ZN VNW pfet_06v0 ad=0.2561p pd=1.505u as=0.4016p ps=1.94u w=0.985u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4016p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.44325p pd=2.87u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6 VSS C a_692_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VPW nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 VDD VSS ZN A1 A2 VNW VPW
X0 a_1140_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2 ZN A1 a_1140_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X4 a_1588_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X5 VDD A2 a_1588_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6 ZN A1 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7 a_244_472# A2 VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X8 ZN A1 a_244_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X9 a_692_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X11 VDD A2 a_692_472# VNW pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X12 VSS A1 ZN VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X13 VSS A2 ZN VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X14 VSS A1 ZN VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X15 ZN A2 VSS VPW nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 a_224_604# A1 a_36_88# VNW pfet_06v0 ad=0.1736p pd=1.18u as=0.2464p ps=2u w=0.56u l=0.5u
X1 a_36_88# A2 VSS VPW nfet_06v0 ad=0.14p pd=1.1u as=0.104p ps=0.92u w=0.4u l=0.6u
X2 Z a_36_88# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.389p ps=2.02u w=1.22u l=0.5u
X3 VSS A1 a_36_88# VPW nfet_06v0 ad=0.104p pd=0.92u as=0.176p ps=1.68u w=0.4u l=0.6u
X4 a_448_604# A2 a_224_604# VNW pfet_06v0 ad=0.224p pd=1.36u as=0.1736p ps=1.18u w=0.56u l=0.5u
X5 VSS A3 a_36_88# VPW nfet_06v0 ad=0.224p pd=1.52u as=0.14p ps=1.1u w=0.4u l=0.6u
X6 VDD A3 a_448_604# VNW pfet_06v0 ad=0.389p pd=2.02u as=0.224p ps=1.36u w=0.56u l=0.5u
X7 Z a_36_88# VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.224p ps=1.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A4 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X1 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4 a_275_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5 a_673_68# A2 a_469_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X6 a_469_68# A3 a_275_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X7 ZN A1 a_673_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VNW VPW
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VPW nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2384p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1617p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VPW nfet_06v0 ad=0.2384p pd=1.51u as=0.1232p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VPW nfet_06v0 ad=0.2541p pd=1.605u as=0.1196p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.4514p pd=1.96u as=0.3172p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.3782p pd=1.84u as=0.4514p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VPW nfet_06v0 ad=0.1617p pd=1.19u as=0.4466p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VPW nfet_06v0 ad=0.2002p pd=1.29u as=0.1232p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3172p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VPW nfet_06v0 ad=0.264p pd=1.66u as=0.1196p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.2541p ps=1.605u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VPW nfet_06v0 ad=0.1196p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.7076p pd=2.38u as=0.3782p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VPW nfet_06v0 ad=0.2024p pd=1.8u as=0.1196p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VPW nfet_06v0 ad=0.1232p pd=1.09u as=0.2002p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.7076p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 a_1458_68# A3 a_1254_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VPW nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VPW nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VPW nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VPW nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
.ends

.subckt sar_logic VDD VSS clk comp current_state[0] current_state[1] dbot[0] dbot[10] dbot[11]
+ dbot[1] dbot[2] dbot[3] dbot[4] dbot[5] dbot[6] dbot[7] dbot[8] dbot[9] dtop[0]
+ dtop[10] dtop[11] dtop[1] dtop[2] dtop[3] dtop[4] dtop[5] dtop[6] dtop[7] dtop[8]
+ dtop[9] rst
X_200_ _062_ VDD VSS _065_ net33 _034_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_131_ VDD VSS net13 _098_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput20 VSS dtop[1] net20 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput7 VSS dbot[11] net7 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_142 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_130_ VDD VSS net12 _097_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_259_ VDD net12 clknet_2_1_0_clk VSS _021_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput21 VSS dtop[2] net21 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput10 VSS dbot[3] net10 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput8 VSS dbot[1] net8 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_258_ VDD net11 clknet_2_0_0_clk VSS _020_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_189_ VDD VSS _057_ _104_ _052_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_97 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput11 VSS dbot[4] net11 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput22 VSS dtop[3] net22 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput9 dbot[2] VSS VDD net9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_1_133 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_257_ VDD net10 clknet_2_3_0_clk VSS _019_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_188_ VDD VSS _056_ _105_ _050_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput23 VSS dtop[4] net23 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput12 dbot[5] VSS VDD net12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_256_ VDD net9 clknet_2_3_0_clk VSS _018_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_187_ _055_ net29 VDD VSS _009_ _093_ _054_ _115_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_21_44 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_239_ _001_ VDD VSS clknet_2_1_0_clk current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_21_146 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 VSS dtop[5] net24 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput13 dbot[6] VSS VDD net13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_255_ VDD net8 clknet_2_3_0_clk VSS _017_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_186_ VDD VSS _055_ _102_ _052_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_238_ _000_ VDD VSS clknet_2_0_0_clk current_bit\[0\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_21_89 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_169_ _039_ VDD VSS _041_ net34 _032_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_114 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput14 VSS dbot[7] net14 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput25 dtop[6] VSS VDD net25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_254_ VDD net5 clknet_2_0_0_clk VSS _016_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_185_ VDD VSS _054_ _103_ _050_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_142 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_237_ VDD VSS _029_ _100_ net29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_168_ VDD VSS _040_ _089_ _104_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_34 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_79 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput26 VSS dtop[7] net26 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput15 VSS dbot[8] net15 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_115 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_3_0_clk clknet_2_3_0_clk VSS VDD clknet_1_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_19_57 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_253_ VDD net19 clknet_2_3_0_clk VSS _015_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_184_ _053_ net29 VDD VSS _008_ _092_ _051_ _115_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_21_36 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_167_ VDD VSS _039_ net32 _105_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_236_ _117_ VDD VSS _028_ net3 net2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_21_138 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_219_ _106_ VDD VSS _077_ net32 net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput27 dtop[8] VSS VDD net27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput16 VSS dbot[9] net16 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_0_clk VDD VSS clknet_0_clk clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_2_2_0_clk clknet_2_2_0_clk VSS VDD clknet_1_1_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_252_ VDD net18 clknet_2_2_0_clk VSS _014_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_183_ VDD VSS _053_ _106_ _052_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_59 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_235_ VDD net31 _085_ _027_ _072_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_166_ VDD net30 _038_ _005_ _036_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_128 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_218_ VDD net31 _076_ _019_ _049_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_149_ VDD VSS _112_ net3 _087_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput28 VSS dtop[9] net28 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput17 dtop[0] VSS VDD net17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_17_80 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_251_ VDD net28 clknet_2_2_0_clk VSS _013_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout30 net30 VSS VDD net31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_182_ VDD VSS _052_ _089_ net33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_165_ net20 VDD VSS _038_ _032_ _034_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_234_ net7 VDD VSS _085_ _045_ _062_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_2_1_0_clk clknet_2_1_0_clk VSS VDD clknet_1_0_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_217_ net10 VDD VSS _076_ _032_ _045_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_148_ VDD VSS _003_ _101_ _110_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput18 VSS dtop[10] net18 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_21_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_37 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_250_ VDD net27 clknet_2_2_0_clk VSS _012_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout31 VSS net31 _112_ VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_181_ _050_ VDD VSS _051_ current_bit\[1\] current_bit\[0\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_164_ _034_ VDD VSS _037_ net33 _032_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_233_ _084_ VDD VSS _026_ net31 _068_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_18_8 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_147_ VDD VSS _111_ current_bit\[3\] _107_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_216_ _075_ VDD VSS _018_ net30 _042_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput19 VSS dtop[11] net19 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_2_0_0_clk clknet_2_0_0_clk VSS VDD clknet_1_0_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout32 net32 current_bit\[2\] VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_180_ net32 VDD VSS _050_ _087_ _088_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_3_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_163_ _034_ VDD VSS _036_ net34 _032_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_232_ VDD net6 _063_ _084_ _040_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_18 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_215_ VDD net9 _040_ _075_ _033_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_146_ VDD VSS _110_ _088_ _107_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_129_ VDD VSS net11 _096_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout33 net33 VSS VDD net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_231_ _083_ VDD VSS _025_ net31 _065_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_162_ VDD VSS _035_ _089_ _102_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput1 VSS net1 comp VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_214_ _074_ VDD VSS _017_ net30 _037_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_145_ VDD VSS _109_ current_bit\[3\] _107_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_128_ VDD VSS net26 _095_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout34 VSS net34 net1 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_230_ VDD net16 _063_ _083_ _035_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_161_ VDD VSS _034_ net32 _103_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput2 VSS net2 rst VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_213_ VDD net8 _035_ _074_ _033_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_144_ VDD VSS _002_ _101_ _108_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_122 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_127_ VDD VSS net25 _094_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_160_ VDD VSS _033_ _111_ _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_212_ _073_ VDD VSS _016_ net29 _116_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_143_ VDD VSS _108_ _089_ _106_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_126_ VDD VSS net24 _093_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_142_ current_bit\[0\] VDD VSS _107_ net32 current_bit\[1\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_211_ VDD VSS _073_ net5 _117_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_125_ VDD VSS net23 _092_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_10 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_146 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_100 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_210_ _071_ net30 VDD VSS _015_ net34 _070_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_141_ VDD VSS _106_ current_bit\[1\] current_bit\[0\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_124_ VDD VSS current_bit\[0\] _091_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_88 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_115 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_126 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_140_ _105_ VDD VSS _001_ _101_ _103_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_123_ VDD VSS current_bit\[1\] _090_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_45 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_104 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_199_ _062_ VDD VSS _064_ net34 _034_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_1_1_0_clk clknet_1_1_0_clk VSS VDD clknet_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_122_ VDD VSS net32 _089_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_0_138 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout29 VSS net29 net31 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_198_ VDD VSS _063_ _110_ _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_267_ _029_ VDD VSS clknet_2_0_0_clk net4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_121_ VDD VSS current_bit\[3\] _088_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xclkbuf_1_0_0_clk clknet_1_0_0_clk VSS VDD clknet_0_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_91 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_197_ VDD VSS _062_ _110_ _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_266_ _028_ VDD VSS clknet_2_0_0_clk net3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_120_ VSS _087_ net4 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_249_ VDD net26 clknet_2_1_0_clk VSS _011_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_16 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_37 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_265_ VDD net7 clknet_2_3_0_clk VSS _027_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_196_ _061_ VDD VSS _012_ net30 _060_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_248_ VDD net25 clknet_2_1_0_clk VSS _010_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_179_ _048_ net30 VDD VSS _007_ net33 _047_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_0_119 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_70 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_195_ VDD net27 _031_ _061_ _109_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_264_ VDD net6 clknet_2_3_0_clk VSS _026_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_247_ VDD net24 clknet_2_3_0_clk VSS _009_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_178_ _046_ VDD VSS _049_ net33 _033_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_20_83 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_93 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_194_ _031_ VDD VSS _060_ net34 _109_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_263_ VDD net16 clknet_2_3_0_clk VSS _025_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_246_ VDD net23 clknet_2_0_0_clk VSS _008_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_177_ VDD net22 _046_ _048_ _033_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_229_ _082_ VDD VSS _024_ net30 _081_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_193_ _059_ net29 VDD VSS _011_ _095_ _058_ _115_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_262_ VDD net15 clknet_2_2_0_clk VSS _024_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_245_ VDD net22 clknet_2_3_0_clk VSS _007_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_176_ VDD VSS _047_ _032_ _045_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_159_ VDD VSS _032_ _111_ _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_228_ _106_ _113_ VDD VSS _082_ current_bit\[3\] net34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_261_ VDD net14 clknet_2_1_0_clk VSS _023_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_192_ _052_ VDD VSS _059_ current_bit\[1\] current_bit\[0\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_244_ VDD net21 clknet_2_2_0_clk VSS _006_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_175_ VSS _046_ _045_ VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_227_ VDD net15 _031_ _081_ _109_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_158_ _087_ _113_ _114_ VDD VSS _031_ net3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_20_53 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_260_ VDD net13 clknet_2_1_0_clk VSS _022_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_191_ VDD VSS _058_ _044_ _050_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_243_ VDD net20 clknet_2_2_0_clk VSS _005_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_174_ VDD VSS _045_ net32 _044_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_157_ VDD VSS _004_ net29 _030_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_226_ _080_ net31 VDD VSS _023_ _099_ _058_ _115_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_209_ _063_ VDD VSS _072_ net1 _046_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_15_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_190_ _057_ net29 VDD VSS _010_ _094_ _056_ _115_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_4_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_173_ VDD VSS _044_ current_bit\[1\] current_bit\[0\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_242_ VDD net17 clknet_2_0_0_clk VSS _004_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_156_ VDD _116_ _118_ _030_ net17 VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_225_ current_bit\[0\] net33 VDD VSS _080_ current_bit\[2\] current_bit\[1\] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_208_ VDD net19 _063_ _071_ _046_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_139_ VDD VSS _105_ current_bit\[1\] _091_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_142 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_172_ VDD net30 _043_ _006_ _041_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_241_ _003_ VDD VSS clknet_2_2_0_clk current_bit\[3\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_155_ VDD VSS _117_ _118_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_224_ _079_ net29 VDD VSS _022_ _098_ _056_ _115_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_207_ VDD VSS _070_ _045_ _062_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_138_ VDD VSS _104_ _090_ current_bit\[0\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_171_ net21 VDD VSS _043_ _032_ _039_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_240_ VDD current_bit\[2\] clknet_2_2_0_clk VSS _002_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_146 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _104_ VDD VSS _079_ net32 net33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_154_ VDD VSS _117_ _107_ _114_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_206_ VDD net30 _069_ _014_ _067_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_137_ VDD VSS _103_ _090_ current_bit\[0\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_78 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_136 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_170_ _039_ VDD VSS _042_ net33 _032_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_222_ _078_ net29 VDD VSS _021_ _097_ _054_ _115_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_153_ net34 _107_ VDD VSS _116_ _087_ _088_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_205_ net18 VDD VSS _069_ _039_ _062_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_136_ VDD VSS _102_ current_bit\[1\] _091_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_142 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_119_ VDD VSS net3 _086_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_101 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_221_ _102_ VDD VSS _078_ net32 net33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_152_ VDD VSS _115_ _113_ _114_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_204_ _062_ VDD VSS _068_ net33 _039_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_36 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_37 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_135_ current_bit\[0\] VDD VSS _000_ _086_ net4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput3 VSS current_state[0] net3 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_151_ VDD VSS _114_ net4 current_bit\[3\] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_220_ _077_ net29 VDD VSS _020_ _096_ _051_ _031_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_134_ VDD VSS _101_ _086_ net4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_203_ _062_ VDD VSS _067_ net34 _039_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_70 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput4 VSS current_state[1] net4 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_150_ VDD VSS _113_ net4 net32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_0_2 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_202_ VDD net30 _066_ _013_ _064_ VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_133_ VDD VSS net2 _100_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput5 VSS dbot[0] net5 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_132_ VDD VSS net14 _099_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_201_ net28 VDD VSS _066_ _034_ _062_ VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_135 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_18 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_82 VDD VSS VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 VSS dbot[10] net6 VDD VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
.ends


* NGSPICE file created from resistor-pex.ext - technology: gf180mcuD

.subckt resistor-pex B OUT1 OUT2 VDD VSS
X0 OUT2.t0 a_4000_1800.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X1 a_n132_5400.t0 a_4000_4800.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X2 a_n132_7800.t0 a_4000_9000.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X3 a_n132_1200.t1 a_4000_2400.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X4 a_n132_6000.t0 a_4000_4200.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X5 VDD.t0 a_4000_9000.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X6 a_n132_3000.t1 a_4000_2400.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X7 B.t3 B.t4 B.t0 ppolyf_u r_width=1u r_length=20u
X8 a_n132_6000.t1 a_4000_6600.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X9 OUT1.t0 a_4000_600.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X10 a_n132_3600.t1 a_4000_1800.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X11 a_n132_5400.t1 a_4000_7200.t1 B.t0 ppolyf_u r_width=1u r_length=20u
X12 a_n132_3600.t0 a_4000_4200.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X13 a_n132_7800.t1 a_4000_7200.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X14 a_n132_1200.t0 a_4000_600.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X15 a_n132_3000.t0 a_4000_4800.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X16 VSS.t0 a_4000_6600.t0 B.t0 ppolyf_u r_width=1u r_length=20u
X17 B.t1 B.t2 B.t0 ppolyf_u r_width=1u r_length=20u
R0 OUT2 OUT2.t0 19.8748
R1 a_4000_1800.t0 a_4000_1800.t1 40.1685
R2 B.n3 B.t0 679.019
R3 B.n2 B.t1 12.4939
R4 B.n0 B.t3 12.4939
R5 B.n0 B.t4 10.4095
R6 B.n2 B.t2 10.4095
R7 B.n3 B.n1 5.05707
R8 B B.n4 2.66425
R9 B.n4 B.n2 2.36639
R10 B B.n1 0.6382
R11 B.n1 B.n0 0.412158
R12 B.n4 B.n3 0.0879041
R13 a_n132_5400.t0 a_n132_5400.t1 40.1685
R14 a_4000_4800.t0 a_4000_4800.t1 39.9885
R15 a_n132_7800.t0 a_n132_7800.t1 39.8985
R16 a_4000_9000.t0 a_4000_9000.t1 39.9885
R17 a_n132_1200.t0 a_n132_1200.t1 39.8985
R18 a_4000_2400.t0 a_4000_2400.t1 39.9885
R19 a_n132_6000.t0 a_n132_6000.t1 39.9885
R20 a_4000_4200.t0 a_4000_4200.t1 40.1685
R21 VDD VDD.t0 19.8653
R22 a_n132_3000.t0 a_n132_3000.t1 40.1685
R23 a_4000_6600.t0 a_4000_6600.t1 40.1685
R24 OUT1 OUT1.t0 19.8788
R25 a_4000_600.t0 a_4000_600.t1 39.9885
R26 a_n132_3600.t0 a_n132_3600.t1 39.9885
R27 a_4000_7200.t0 a_4000_7200.t1 39.9885
R28 VSS VSS.t0 19.8671
C0 OUT1 m1_n1166_0# 0.041547f
C1 m1_n1166_9000# VSS 0.041547f
C2 m1_4966_6600# m1_4966_6000# 0.041547f
C3 m1_4566_0# m1_4966_0# 0.080033f
C4 VDD m1_n1166_10200# 0.041547f
C5 VDD m1_n766_10200# 0.023331f
C6 m1_n1166_4800# m1_n1166_5400# 0.041547f
C7 m1_n1166_3000# m1_n1166_2400# 0.041547f
C8 m1_n1166_7200# m1_n1166_7800# 0.041547f
C9 m1_4966_10200# m1_4566_10200# 0.080033f
C10 VDD VSS 0.008902f
C11 OUT2 OUT1 0.025988f
C12 m1_n1166_7800# VSS 0.041547f
C13 m1_n766_0# m1_n1166_0# 0.080033f
C14 m1_n766_10200# m1_n1166_10200# 0.080033f
C15 VDD m1_n1166_9000# 0.041547f
C16 m1_n766_0# OUT1 0.023331f
C17 OUT2 m1_n1166_2400# 0.041547f
C18 m1_4966_4200# m1_4966_3600# 0.041547f
C19 OUT1 B 1.02531f
C20 OUT2 B 0.86077f
C21 VSS B 0.841918f
C22 VDD B 1.00646f
C23 m1_4966_0# B 0.227912f $ **FLOATING
C24 m1_4566_0# B 0.248546f $ **FLOATING
C25 m1_n766_0# B 0.260418f $ **FLOATING
C26 m1_n1166_0# B 0.227912f $ **FLOATING
C27 m1_4966_1800# B 0.187856f $ **FLOATING
C28 m1_4966_3600# B 0.187856f $ **FLOATING
C29 m1_n1166_2400# B 0.187856f $ **FLOATING
C30 m1_4966_4200# B 0.187856f $ **FLOATING
C31 m1_4966_6000# B 0.187856f $ **FLOATING
C32 m1_n1166_3000# B 0.187856f $ **FLOATING
C33 m1_n1166_4800# B 0.187856f $ **FLOATING
C34 m1_4966_6600# B 0.187856f $ **FLOATING
C35 m1_4966_8400# B 0.187856f $ **FLOATING
C36 m1_n1166_5400# B 0.187856f $ **FLOATING
C37 m1_n1166_7200# B 0.187856f $ **FLOATING
C38 m1_n1166_7800# B 0.187856f $ **FLOATING
C39 m1_n1166_9000# B 0.187856f $ **FLOATING
C40 m1_4966_10200# B 0.227912f $ **FLOATING
C41 m1_4566_10200# B 0.248546f $ **FLOATING
C42 m1_n766_10200# B 0.260418f $ **FLOATING
C43 m1_n1166_10200# B 0.227912f $ **FLOATING
.ends


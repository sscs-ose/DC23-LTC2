* Extracted by KLayout with GF180MCU LVS runset on : 18/01/2024 00:22

.SUBCKT waffle_1984 G
M$1 \$4 G \$8 \$4 pfet_03v3 L=0.5U W=8689.92U AS=5051.0418P AD=5049.1178P
+ PS=17554.32U PD=17507.92U
.ENDS waffle_1984

* 10-bit Counter
.SUBCKT 10bit_Counter OUT0 OUT1 OUT2 OUT3 OUT4 OUT5 OUT6 OUT7 OUT8 OUT9
* Output configuration
VPULSE_0 OUT0 0 PULSE(0V 3.3V 10n 2n 2n 23n 50n) 
VPULSE_1 OUT1 0 PULSE(0V 3.3V 35n 2n 2n 48n 100n) 
VPULSE_2 OUT2 0 PULSE(0V 3.3V 85n 2n 2n 98n 200n) 
VPULSE_3 OUT3 0 PULSE(0V 3.3V 185n 2n 2n 198n 400n) 
VPULSE_4 OUT4 0 PULSE(0V 3.3V 385n 2n 2n 398n 800n) 
VPULSE_5 OUT5 0 PULSE(0V 3.3V 785n 2n 2n 798n 1600n) 
VPULSE_6 OUT6 0 PULSE(0V 3.3V 1585n 2n 2n 1598n 3200n) 
VPULSE_7 OUT7 0 PULSE(0V 3.3V 3185n 2n 2n 3198n 6400n) 
VPULSE_8 OUT8 0 PULSE(0V 3.3V 6385n 2n 2n 6398n 12800n) 
VPULSE_9 OUT9 0 PULSE(0V 3.3V 12785n 2n 2n 12798n 25600n) 
.ENDS
